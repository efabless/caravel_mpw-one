magic
tech sky130A
magscale 1 2
timestamp 1625155807
<< metal1 >>
rect 585042 996344 585048 996396
rect 585100 996384 585106 996396
rect 674742 996384 674748 996396
rect 585100 996356 674748 996384
rect 585100 996344 585106 996356
rect 674742 996344 674748 996356
rect 674800 996344 674806 996396
rect 342162 990836 342168 990888
rect 342220 990876 342226 990888
rect 673546 990876 673552 990888
rect 342220 990848 673552 990876
rect 342220 990836 342226 990848
rect 673546 990836 673552 990848
rect 673604 990836 673610 990888
rect 42242 990156 42248 990208
rect 42300 990196 42306 990208
rect 342254 990196 342260 990208
rect 42300 990168 342260 990196
rect 42300 990156 42306 990168
rect 342254 990156 342260 990168
rect 342312 990156 342318 990208
rect 44910 990088 44916 990140
rect 44968 990128 44974 990140
rect 673454 990128 673460 990140
rect 44968 990100 673460 990128
rect 44968 990088 44974 990100
rect 673454 990088 673460 990100
rect 673512 990088 673518 990140
rect 42334 990020 42340 990072
rect 42392 990060 42398 990072
rect 673638 990060 673644 990072
rect 42392 990032 673644 990060
rect 42392 990020 42398 990032
rect 673638 990020 673644 990032
rect 673696 990020 673702 990072
rect 673638 875780 673644 875832
rect 673696 875820 673702 875832
rect 675386 875820 675392 875832
rect 673696 875792 675392 875820
rect 673696 875780 673702 875792
rect 675386 875780 675392 875792
rect 675444 875780 675450 875832
rect 673546 874488 673552 874540
rect 673604 874528 673610 874540
rect 675386 874528 675392 874540
rect 673604 874500 675392 874528
rect 673604 874488 673610 874500
rect 675386 874488 675392 874500
rect 675444 874488 675450 874540
rect 673454 872380 673460 872432
rect 673512 872420 673518 872432
rect 674006 872420 674012 872432
rect 673512 872392 674012 872420
rect 673512 872380 673518 872392
rect 674006 872380 674012 872392
rect 674064 872420 674070 872432
rect 675386 872420 675392 872432
rect 674064 872392 675392 872420
rect 674064 872380 674070 872392
rect 675386 872380 675392 872392
rect 675444 872380 675450 872432
rect 673730 871292 673736 871344
rect 673788 871332 673794 871344
rect 675294 871332 675300 871344
rect 673788 871304 675300 871332
rect 673788 871292 673794 871304
rect 675294 871292 675300 871304
rect 675352 871292 675358 871344
rect 673914 870136 673920 870188
rect 673972 870176 673978 870188
rect 675386 870176 675392 870188
rect 673972 870148 675392 870176
rect 673972 870136 673978 870148
rect 675386 870136 675392 870148
rect 675444 870136 675450 870188
rect 673822 864220 673828 864272
rect 673880 864260 673886 864272
rect 675386 864260 675392 864272
rect 673880 864232 675392 864260
rect 673880 864220 673886 864232
rect 675386 864220 675392 864232
rect 675444 864220 675450 864272
rect 673914 863200 673920 863252
rect 673972 863240 673978 863252
rect 675386 863240 675392 863252
rect 673972 863212 675392 863240
rect 673972 863200 673978 863212
rect 675386 863200 675392 863212
rect 675444 863200 675450 863252
rect 675294 818320 675300 818372
rect 675352 818360 675358 818372
rect 677594 818360 677600 818372
rect 675352 818332 677600 818360
rect 675352 818320 675358 818332
rect 677594 818320 677600 818332
rect 677652 818320 677658 818372
rect 41782 797716 41788 797768
rect 41840 797756 41846 797768
rect 42610 797756 42616 797768
rect 41840 797728 42616 797756
rect 41840 797716 41846 797728
rect 42610 797716 42616 797728
rect 42668 797716 42674 797768
rect 41782 791936 41788 791988
rect 41840 791976 41846 791988
rect 42426 791976 42432 791988
rect 41840 791948 42432 791976
rect 41840 791936 41846 791948
rect 42426 791936 42432 791948
rect 42484 791936 42490 791988
rect 41782 791324 41788 791376
rect 41840 791364 41846 791376
rect 42518 791364 42524 791376
rect 41840 791336 42524 791364
rect 41840 791324 41846 791336
rect 42518 791324 42524 791336
rect 42576 791324 42582 791376
rect 41782 786972 41788 787024
rect 41840 787012 41846 787024
rect 42426 787012 42432 787024
rect 41840 786984 42432 787012
rect 41840 786972 41846 786984
rect 42426 786972 42432 786984
rect 42484 786972 42490 787024
rect 673730 785952 673736 786004
rect 673788 785992 673794 786004
rect 675202 785992 675208 786004
rect 673788 785964 675208 785992
rect 673788 785952 673794 785964
rect 675202 785952 675208 785964
rect 675260 785992 675266 786004
rect 675386 785992 675392 786004
rect 675260 785964 675392 785992
rect 675260 785952 675266 785964
rect 675386 785952 675392 785964
rect 675444 785952 675450 786004
rect 673454 785680 673460 785732
rect 673512 785720 673518 785732
rect 675386 785720 675392 785732
rect 673512 785692 675392 785720
rect 673512 785680 673518 785692
rect 675386 785680 675392 785692
rect 675444 785680 675450 785732
rect 673638 782280 673644 782332
rect 673696 782320 673702 782332
rect 674006 782320 674012 782332
rect 673696 782292 674012 782320
rect 673696 782280 673702 782292
rect 674006 782280 674012 782292
rect 674064 782320 674070 782332
rect 675386 782320 675392 782332
rect 674064 782292 675392 782320
rect 674064 782280 674070 782292
rect 675386 782280 675392 782292
rect 675444 782280 675450 782332
rect 673730 781600 673736 781652
rect 673788 781640 673794 781652
rect 675202 781640 675208 781652
rect 673788 781612 675208 781640
rect 673788 781600 673794 781612
rect 675202 781600 675208 781612
rect 675260 781640 675266 781652
rect 675386 781640 675392 781652
rect 675260 781612 675392 781640
rect 675260 781600 675266 781612
rect 675386 781600 675392 781612
rect 675444 781600 675450 781652
rect 675202 780988 675208 781040
rect 675260 781028 675266 781040
rect 675386 781028 675392 781040
rect 675260 781000 675392 781028
rect 675260 780988 675266 781000
rect 675386 780988 675392 781000
rect 675444 780988 675450 781040
rect 673822 775820 673828 775872
rect 673880 775860 673886 775872
rect 675386 775860 675392 775872
rect 673880 775832 675392 775860
rect 673880 775820 673886 775832
rect 675386 775820 675392 775832
rect 675444 775820 675450 775872
rect 42242 762220 42248 762272
rect 42300 762260 42306 762272
rect 42518 762260 42524 762272
rect 42300 762232 42524 762260
rect 42300 762220 42306 762232
rect 42518 762220 42524 762232
rect 42576 762220 42582 762272
rect 41782 755420 41788 755472
rect 41840 755460 41846 755472
rect 42610 755460 42616 755472
rect 41840 755432 42616 755460
rect 41840 755420 41846 755432
rect 42610 755420 42616 755432
rect 42668 755420 42674 755472
rect 41782 747668 41788 747720
rect 41840 747708 41846 747720
rect 42426 747708 42432 747720
rect 41840 747680 42432 747708
rect 41840 747668 41846 747680
rect 42426 747668 42432 747680
rect 42484 747668 42490 747720
rect 41782 743996 41788 744048
rect 41840 744036 41846 744048
rect 42518 744036 42524 744048
rect 41840 744008 42524 744036
rect 41840 743996 41846 744008
rect 42518 743996 42524 744008
rect 42576 743996 42582 744048
rect 673730 740936 673736 740988
rect 673788 740976 673794 740988
rect 675202 740976 675208 740988
rect 673788 740948 675208 740976
rect 673788 740936 673794 740948
rect 675202 740936 675208 740948
rect 675260 740976 675266 740988
rect 675386 740976 675392 740988
rect 675260 740948 675392 740976
rect 675260 740936 675266 740948
rect 675386 740936 675392 740948
rect 675444 740936 675450 740988
rect 673454 740324 673460 740376
rect 673512 740364 673518 740376
rect 675386 740364 675392 740376
rect 673512 740336 675392 740364
rect 673512 740324 673518 740336
rect 675386 740324 675392 740336
rect 675444 740324 675450 740376
rect 673638 738080 673644 738132
rect 673696 738120 673702 738132
rect 675386 738120 675392 738132
rect 673696 738092 675392 738120
rect 673696 738080 673702 738092
rect 675386 738080 675392 738092
rect 675444 738080 675450 738132
rect 673730 736992 673736 737044
rect 673788 737032 673794 737044
rect 675202 737032 675208 737044
rect 673788 737004 675208 737032
rect 673788 736992 673794 737004
rect 675202 736992 675208 737004
rect 675260 737032 675266 737044
rect 675386 737032 675392 737044
rect 675260 737004 675392 737032
rect 675260 736992 675266 737004
rect 675386 736992 675392 737004
rect 675444 736992 675450 737044
rect 673546 730872 673552 730924
rect 673604 730912 673610 730924
rect 673914 730912 673920 730924
rect 673604 730884 673920 730912
rect 673604 730872 673610 730884
rect 673914 730872 673920 730884
rect 673972 730912 673978 730924
rect 675386 730912 675392 730924
rect 673972 730884 675392 730912
rect 673972 730872 673978 730884
rect 675386 730872 675392 730884
rect 675444 730872 675450 730924
rect 41782 712240 41788 712292
rect 41840 712280 41846 712292
rect 42610 712280 42616 712292
rect 41840 712252 42616 712280
rect 41840 712240 41846 712252
rect 42610 712240 42616 712252
rect 42668 712240 42674 712292
rect 41782 703944 41788 703996
rect 41840 703984 41846 703996
rect 42426 703984 42432 703996
rect 41840 703956 42432 703984
rect 41840 703944 41846 703956
rect 42426 703944 42432 703956
rect 42484 703944 42490 703996
rect 41782 700816 41788 700868
rect 41840 700856 41846 700868
rect 42518 700856 42524 700868
rect 41840 700828 42524 700856
rect 41840 700816 41846 700828
rect 42518 700816 42524 700828
rect 42576 700816 42582 700868
rect 673730 695920 673736 695972
rect 673788 695960 673794 695972
rect 675202 695960 675208 695972
rect 673788 695932 675208 695960
rect 673788 695920 673794 695932
rect 675202 695920 675208 695932
rect 675260 695960 675266 695972
rect 675386 695960 675392 695972
rect 675260 695932 675392 695960
rect 675260 695920 675266 695932
rect 675386 695920 675392 695932
rect 675444 695920 675450 695972
rect 673454 695308 673460 695360
rect 673512 695348 673518 695360
rect 675386 695348 675392 695360
rect 673512 695320 675392 695348
rect 673512 695308 673518 695320
rect 675386 695308 675392 695320
rect 675444 695308 675450 695360
rect 673914 692248 673920 692300
rect 673972 692288 673978 692300
rect 675386 692288 675392 692300
rect 673972 692260 675392 692288
rect 673972 692248 673978 692260
rect 675386 692248 675392 692260
rect 675444 692248 675450 692300
rect 673730 692044 673736 692096
rect 673788 692084 673794 692096
rect 675202 692084 675208 692096
rect 673788 692056 675208 692084
rect 673788 692044 673794 692056
rect 675202 692044 675208 692056
rect 675260 692084 675266 692096
rect 675386 692084 675392 692096
rect 675260 692056 675392 692084
rect 675260 692044 675266 692056
rect 675386 692044 675392 692056
rect 675444 692044 675450 692096
rect 673546 685176 673552 685228
rect 673604 685216 673610 685228
rect 675386 685216 675392 685228
rect 673604 685188 675392 685216
rect 673604 685176 673610 685188
rect 675386 685176 675392 685188
rect 675444 685176 675450 685228
rect 41782 668108 41788 668160
rect 41840 668148 41846 668160
rect 42702 668148 42708 668160
rect 41840 668120 42708 668148
rect 41840 668108 41846 668120
rect 42702 668108 42708 668120
rect 42760 668108 42766 668160
rect 41782 661036 41788 661088
rect 41840 661076 41846 661088
rect 42426 661076 42432 661088
rect 41840 661048 42432 661076
rect 41840 661036 41846 661048
rect 42426 661036 42432 661048
rect 42484 661036 42490 661088
rect 41782 658656 41788 658708
rect 41840 658696 41846 658708
rect 42518 658696 42524 658708
rect 41840 658668 42524 658696
rect 41840 658656 41846 658668
rect 42518 658656 42524 658668
rect 42576 658656 42582 658708
rect 673730 651108 673736 651160
rect 673788 651148 673794 651160
rect 675386 651148 675392 651160
rect 673788 651120 675392 651148
rect 673788 651108 673794 651120
rect 675386 651108 675392 651120
rect 675444 651108 675450 651160
rect 673454 650496 673460 650548
rect 673512 650536 673518 650548
rect 675386 650536 675392 650548
rect 673512 650508 675392 650536
rect 673512 650496 673518 650508
rect 675386 650496 675392 650508
rect 675444 650496 675450 650548
rect 673454 647164 673460 647216
rect 673512 647204 673518 647216
rect 673638 647204 673644 647216
rect 673512 647176 673644 647204
rect 673512 647164 673518 647176
rect 673638 647164 673644 647176
rect 673696 647164 673702 647216
rect 673454 647028 673460 647080
rect 673512 647068 673518 647080
rect 673914 647068 673920 647080
rect 673512 647040 673920 647068
rect 673512 647028 673518 647040
rect 673914 647028 673920 647040
rect 673972 647068 673978 647080
rect 675386 647068 675392 647080
rect 673972 647040 675392 647068
rect 673972 647028 673978 647040
rect 675386 647028 675392 647040
rect 675444 647028 675450 647080
rect 673730 646416 673736 646468
rect 673788 646456 673794 646468
rect 675386 646456 675392 646468
rect 673788 646428 675392 646456
rect 673788 646416 673794 646428
rect 675386 646416 675392 646428
rect 675444 646416 675450 646468
rect 675202 645736 675208 645788
rect 675260 645776 675266 645788
rect 675386 645776 675392 645788
rect 675260 645748 675392 645776
rect 675260 645736 675266 645748
rect 675386 645736 675392 645748
rect 675444 645736 675450 645788
rect 673546 640636 673552 640688
rect 673604 640676 673610 640688
rect 675386 640676 675392 640688
rect 673604 640648 675392 640676
rect 673604 640636 673610 640648
rect 675386 640636 675392 640648
rect 675444 640636 675450 640688
rect 41782 624928 41788 624980
rect 41840 624968 41846 624980
rect 42518 624968 42524 624980
rect 41840 624940 42524 624968
rect 41840 624928 41846 624940
rect 42518 624928 42524 624940
rect 42576 624968 42582 624980
rect 42702 624968 42708 624980
rect 42576 624940 42708 624968
rect 42576 624928 42582 624940
rect 42702 624928 42708 624940
rect 42760 624928 42766 624980
rect 41782 618468 41788 618520
rect 41840 618508 41846 618520
rect 42426 618508 42432 618520
rect 41840 618480 42432 618508
rect 41840 618468 41846 618480
rect 42426 618468 42432 618480
rect 42484 618468 42490 618520
rect 41782 615476 41788 615528
rect 41840 615516 41846 615528
rect 42610 615516 42616 615528
rect 41840 615488 42616 615516
rect 41840 615476 41846 615488
rect 42610 615476 42616 615488
rect 42668 615476 42674 615528
rect 673730 605752 673736 605804
rect 673788 605792 673794 605804
rect 675202 605792 675208 605804
rect 673788 605764 675208 605792
rect 673788 605752 673794 605764
rect 675202 605752 675208 605764
rect 675260 605792 675266 605804
rect 675386 605792 675392 605804
rect 675260 605764 675392 605792
rect 675260 605752 675266 605764
rect 675386 605752 675392 605764
rect 675444 605752 675450 605804
rect 673638 605072 673644 605124
rect 673696 605112 673702 605124
rect 675386 605112 675392 605124
rect 673696 605084 675392 605112
rect 673696 605072 673702 605084
rect 675386 605072 675392 605084
rect 675444 605072 675450 605124
rect 673454 602896 673460 602948
rect 673512 602936 673518 602948
rect 675386 602936 675392 602948
rect 673512 602908 675392 602936
rect 673512 602896 673518 602908
rect 675386 602896 675392 602908
rect 675444 602896 675450 602948
rect 673730 601808 673736 601860
rect 673788 601848 673794 601860
rect 675202 601848 675208 601860
rect 673788 601820 675208 601848
rect 673788 601808 673794 601820
rect 675202 601808 675208 601820
rect 675260 601848 675266 601860
rect 675386 601848 675392 601860
rect 675260 601820 675392 601848
rect 675260 601808 675266 601820
rect 675386 601808 675392 601820
rect 675444 601808 675450 601860
rect 673546 595008 673552 595060
rect 673604 595048 673610 595060
rect 675386 595048 675392 595060
rect 673604 595020 675392 595048
rect 673604 595008 673610 595020
rect 675386 595008 675392 595020
rect 675444 595008 675450 595060
rect 41782 582632 41788 582684
rect 41840 582672 41846 582684
rect 42518 582672 42524 582684
rect 41840 582644 42524 582672
rect 41840 582632 41846 582644
rect 42518 582632 42524 582644
rect 42576 582632 42582 582684
rect 41782 574676 41788 574728
rect 41840 574716 41846 574728
rect 42426 574716 42432 574728
rect 41840 574688 42432 574716
rect 41840 574676 41846 574688
rect 42426 574676 42432 574688
rect 42484 574676 42490 574728
rect 41782 571208 41788 571260
rect 41840 571248 41846 571260
rect 42518 571248 42524 571260
rect 41840 571220 42524 571248
rect 41840 571208 41846 571220
rect 42518 571208 42524 571220
rect 42576 571248 42582 571260
rect 42702 571248 42708 571260
rect 42576 571220 42708 571248
rect 42576 571208 42582 571220
rect 42702 571208 42708 571220
rect 42760 571208 42766 571260
rect 673730 561212 673736 561264
rect 673788 561252 673794 561264
rect 675202 561252 675208 561264
rect 673788 561224 675208 561252
rect 673788 561212 673794 561224
rect 675202 561212 675208 561224
rect 675260 561252 675266 561264
rect 675386 561252 675392 561264
rect 675260 561224 675392 561252
rect 675260 561212 675266 561224
rect 675386 561212 675392 561224
rect 675444 561212 675450 561264
rect 673638 560940 673644 560992
rect 673696 560980 673702 560992
rect 675386 560980 675392 560992
rect 673696 560952 675392 560980
rect 673696 560940 673702 560952
rect 675386 560940 675392 560952
rect 675444 560940 675450 560992
rect 673454 557812 673460 557864
rect 673512 557852 673518 557864
rect 675386 557852 675392 557864
rect 673512 557824 675392 557852
rect 673512 557812 673518 557824
rect 675386 557812 675392 557824
rect 675444 557812 675450 557864
rect 675202 557268 675208 557320
rect 675260 557308 675266 557320
rect 675386 557308 675392 557320
rect 675260 557280 675392 557308
rect 675260 557268 675266 557280
rect 675386 557268 675392 557280
rect 675444 557268 675450 557320
rect 675202 555568 675208 555620
rect 675260 555608 675266 555620
rect 675386 555608 675392 555620
rect 675260 555580 675392 555608
rect 675260 555568 675266 555580
rect 675386 555568 675392 555580
rect 675444 555568 675450 555620
rect 673546 550468 673552 550520
rect 673604 550508 673610 550520
rect 675386 550508 675392 550520
rect 673604 550480 675392 550508
rect 673604 550468 673610 550480
rect 675386 550468 675392 550480
rect 675444 550468 675450 550520
rect 42334 545232 42340 545284
rect 42392 545232 42398 545284
rect 42352 545080 42380 545232
rect 42334 545028 42340 545080
rect 42392 545028 42398 545080
rect 41782 539452 41788 539504
rect 41840 539492 41846 539504
rect 42610 539492 42616 539504
rect 41840 539464 42616 539492
rect 41840 539452 41846 539464
rect 42610 539452 42616 539464
rect 42668 539452 42674 539504
rect 42242 532108 42248 532160
rect 42300 532148 42306 532160
rect 42426 532148 42432 532160
rect 42300 532120 42432 532148
rect 42300 532108 42306 532120
rect 42426 532108 42432 532120
rect 42484 532108 42490 532160
rect 41782 531156 41788 531208
rect 41840 531196 41846 531208
rect 42426 531196 42432 531208
rect 41840 531168 42432 531196
rect 41840 531156 41846 531168
rect 42426 531156 42432 531168
rect 42484 531156 42490 531208
rect 41782 528028 41788 528080
rect 41840 528068 41846 528080
rect 42518 528068 42524 528080
rect 41840 528040 42524 528068
rect 41840 528028 41846 528040
rect 42518 528028 42524 528040
rect 42576 528068 42582 528080
rect 42702 528068 42708 528080
rect 42576 528040 42708 528068
rect 42576 528028 42582 528040
rect 42702 528028 42708 528040
rect 42760 528028 42766 528080
rect 675294 513748 675300 513800
rect 675352 513788 675358 513800
rect 677686 513788 677692 513800
rect 675352 513760 677692 513788
rect 675352 513748 675358 513760
rect 677686 513748 677692 513760
rect 677744 513748 677750 513800
rect 674742 427796 674748 427848
rect 674800 427836 674806 427848
rect 677502 427836 677508 427848
rect 674800 427808 677508 427836
rect 674800 427796 674806 427808
rect 677502 427796 677508 427808
rect 677560 427796 677566 427848
rect 41782 410932 41788 410984
rect 41840 410972 41846 410984
rect 42518 410972 42524 410984
rect 41840 410944 42524 410972
rect 41840 410932 41846 410944
rect 42518 410932 42524 410944
rect 42576 410932 42582 410984
rect 41782 404472 41788 404524
rect 41840 404512 41846 404524
rect 42426 404512 42432 404524
rect 41840 404484 42432 404512
rect 41840 404472 41846 404484
rect 42426 404472 42432 404484
rect 42484 404512 42490 404524
rect 42610 404512 42616 404524
rect 42484 404484 42616 404512
rect 42484 404472 42490 404484
rect 42610 404472 42616 404484
rect 42668 404472 42674 404524
rect 41782 400800 41788 400852
rect 41840 400840 41846 400852
rect 42702 400840 42708 400852
rect 41840 400812 42708 400840
rect 41840 400800 41846 400812
rect 42702 400800 42708 400812
rect 42760 400800 42766 400852
rect 673546 382712 673552 382764
rect 673604 382752 673610 382764
rect 675386 382752 675392 382764
rect 673604 382724 675392 382752
rect 673604 382712 673610 382724
rect 675386 382712 675392 382724
rect 675444 382712 675450 382764
rect 673730 379652 673736 379704
rect 673788 379692 673794 379704
rect 675386 379692 675392 379704
rect 673788 379664 675392 379692
rect 673788 379652 673794 379664
rect 675386 379652 675392 379664
rect 675444 379652 675450 379704
rect 673638 379040 673644 379092
rect 673696 379080 673702 379092
rect 675386 379080 675392 379092
rect 673696 379052 675392 379080
rect 673696 379040 673702 379052
rect 675386 379040 675392 379052
rect 675444 379040 675450 379092
rect 673454 372308 673460 372360
rect 673512 372348 673518 372360
rect 675386 372348 675392 372360
rect 673512 372320 675392 372348
rect 673512 372308 673518 372320
rect 675386 372308 675392 372320
rect 675444 372308 675450 372360
rect 41782 368636 41788 368688
rect 41840 368676 41846 368688
rect 42334 368676 42340 368688
rect 41840 368648 42340 368676
rect 41840 368636 41846 368648
rect 42334 368636 42340 368648
rect 42392 368676 42398 368688
rect 42518 368676 42524 368688
rect 42392 368648 42524 368676
rect 42392 368636 42398 368648
rect 42518 368636 42524 368648
rect 42576 368636 42582 368688
rect 41782 361292 41788 361344
rect 41840 361332 41846 361344
rect 42334 361332 42340 361344
rect 41840 361304 42340 361332
rect 41840 361292 41846 361304
rect 42334 361292 42340 361304
rect 42392 361292 42398 361344
rect 41782 360680 41788 360732
rect 41840 360720 41846 360732
rect 42610 360720 42616 360732
rect 41840 360692 42616 360720
rect 41840 360680 41846 360692
rect 42610 360680 42616 360692
rect 42668 360680 42674 360732
rect 41782 357212 41788 357264
rect 41840 357252 41846 357264
rect 42518 357252 42524 357264
rect 41840 357224 42524 357252
rect 41840 357212 41846 357224
rect 42518 357212 42524 357224
rect 42576 357252 42582 357264
rect 42702 357252 42708 357264
rect 42576 357224 42708 357252
rect 42576 357212 42582 357224
rect 42702 357212 42708 357224
rect 42760 357212 42766 357264
rect 41782 356668 41788 356720
rect 41840 356708 41846 356720
rect 42334 356708 42340 356720
rect 41840 356680 42340 356708
rect 41840 356668 41846 356680
rect 42334 356668 42340 356680
rect 42392 356668 42398 356720
rect 673546 337492 673552 337544
rect 673604 337532 673610 337544
rect 675386 337532 675392 337544
rect 673604 337504 675392 337532
rect 673604 337492 673610 337504
rect 675386 337492 675392 337504
rect 675444 337492 675450 337544
rect 673914 334432 673920 334484
rect 673972 334472 673978 334484
rect 675386 334472 675392 334484
rect 673972 334444 675392 334472
rect 673972 334432 673978 334444
rect 675386 334432 675392 334444
rect 675444 334432 675450 334484
rect 673638 334228 673644 334280
rect 673696 334268 673702 334280
rect 675386 334268 675392 334280
rect 673696 334240 675392 334268
rect 673696 334228 673702 334240
rect 675386 334228 675392 334240
rect 675444 334228 675450 334280
rect 42242 330012 42248 330064
rect 42300 330052 42306 330064
rect 42426 330052 42432 330064
rect 42300 330024 42432 330052
rect 42300 330012 42306 330024
rect 42426 330012 42432 330024
rect 42484 330012 42490 330064
rect 673454 328040 673460 328092
rect 673512 328080 673518 328092
rect 675386 328080 675392 328092
rect 673512 328052 675392 328080
rect 673512 328040 673518 328052
rect 675386 328040 675392 328052
rect 675444 328040 675450 328092
rect 41782 325456 41788 325508
rect 41840 325496 41846 325508
rect 42426 325496 42432 325508
rect 41840 325468 42432 325496
rect 41840 325456 41846 325468
rect 42426 325456 42432 325468
rect 42484 325496 42490 325508
rect 42794 325496 42800 325508
rect 42484 325468 42800 325496
rect 42484 325456 42490 325468
rect 42794 325456 42800 325468
rect 42852 325456 42858 325508
rect 41782 317160 41788 317212
rect 41840 317200 41846 317212
rect 42610 317200 42616 317212
rect 41840 317172 42616 317200
rect 41840 317160 41846 317172
rect 42610 317160 42616 317172
rect 42668 317160 42674 317212
rect 41782 314032 41788 314084
rect 41840 314072 41846 314084
rect 42518 314072 42524 314084
rect 41840 314044 42524 314072
rect 41840 314032 41846 314044
rect 42518 314032 42524 314044
rect 42576 314072 42582 314084
rect 42702 314072 42708 314084
rect 42576 314044 42708 314072
rect 42576 314032 42582 314044
rect 42702 314032 42708 314044
rect 42760 314032 42766 314084
rect 673638 293768 673644 293820
rect 673696 293808 673702 293820
rect 675386 293808 675392 293820
rect 673696 293780 675392 293808
rect 673696 293768 673702 293780
rect 675386 293768 675392 293780
rect 675444 293768 675450 293820
rect 673546 293564 673552 293616
rect 673604 293604 673610 293616
rect 675386 293604 675392 293616
rect 673604 293576 675392 293604
rect 673604 293564 673610 293576
rect 675386 293564 675392 293576
rect 675444 293564 675450 293616
rect 673914 289824 673920 289876
rect 673972 289864 673978 289876
rect 675386 289864 675392 289876
rect 673972 289836 675392 289864
rect 673972 289824 673978 289836
rect 675386 289824 675392 289836
rect 675444 289824 675450 289876
rect 673454 282072 673460 282124
rect 673512 282112 673518 282124
rect 673730 282112 673736 282124
rect 673512 282084 673736 282112
rect 673512 282072 673518 282084
rect 673730 282072 673736 282084
rect 673788 282112 673794 282124
rect 675386 282112 675392 282124
rect 673788 282084 675392 282112
rect 673788 282072 673794 282084
rect 675386 282072 675392 282084
rect 675444 282072 675450 282124
rect 41782 281324 41788 281376
rect 41840 281364 41846 281376
rect 42426 281364 42432 281376
rect 41840 281336 42432 281364
rect 41840 281324 41846 281336
rect 42426 281324 42432 281336
rect 42484 281364 42490 281376
rect 42794 281364 42800 281376
rect 42484 281336 42800 281364
rect 42484 281324 42490 281336
rect 42794 281324 42800 281336
rect 42852 281324 42858 281376
rect 41782 274524 41788 274576
rect 41840 274564 41846 274576
rect 42610 274564 42616 274576
rect 41840 274536 42616 274564
rect 41840 274524 41846 274536
rect 42610 274524 42616 274536
rect 42668 274524 42674 274576
rect 41782 271872 41788 271924
rect 41840 271912 41846 271924
rect 42702 271912 42708 271924
rect 41840 271884 42708 271912
rect 41840 271872 41846 271884
rect 42702 271872 42708 271884
rect 42760 271872 42766 271924
rect 673638 249092 673644 249144
rect 673696 249132 673702 249144
rect 675386 249132 675392 249144
rect 673696 249104 675392 249132
rect 673696 249092 673702 249104
rect 675386 249092 675392 249104
rect 675444 249092 675450 249144
rect 673546 248548 673552 248600
rect 673604 248588 673610 248600
rect 675386 248588 675392 248600
rect 673604 248560 675392 248588
rect 673604 248548 673610 248560
rect 675386 248548 675392 248560
rect 675444 248548 675450 248600
rect 673914 244876 673920 244928
rect 673972 244916 673978 244928
rect 675386 244916 675392 244928
rect 673972 244888 675392 244916
rect 673972 244876 673978 244888
rect 675386 244876 675392 244888
rect 675444 244876 675450 244928
rect 673638 243992 673644 244044
rect 673696 244032 673702 244044
rect 673914 244032 673920 244044
rect 673696 244004 673920 244032
rect 673696 243992 673702 244004
rect 673914 243992 673920 244004
rect 673972 243992 673978 244044
rect 673822 243788 673828 243840
rect 673880 243828 673886 243840
rect 675386 243828 675392 243840
rect 673880 243800 675392 243828
rect 673880 243788 673886 243800
rect 675386 243788 675392 243800
rect 675444 243788 675450 243840
rect 41782 238076 41788 238128
rect 41840 238116 41846 238128
rect 42426 238116 42432 238128
rect 41840 238088 42432 238116
rect 41840 238076 41846 238088
rect 42426 238076 42432 238088
rect 42484 238076 42490 238128
rect 673914 237668 673920 237720
rect 673972 237708 673978 237720
rect 675386 237708 675392 237720
rect 673972 237680 675392 237708
rect 673972 237668 673978 237680
rect 675386 237668 675392 237680
rect 675444 237668 675450 237720
rect 41782 231684 41788 231736
rect 41840 231724 41846 231736
rect 42518 231724 42524 231736
rect 41840 231696 42524 231724
rect 41840 231684 41846 231696
rect 42518 231684 42524 231696
rect 42576 231684 42582 231736
rect 41782 228624 41788 228676
rect 41840 228664 41846 228676
rect 42610 228664 42616 228676
rect 41840 228636 42616 228664
rect 41840 228624 41846 228636
rect 42610 228624 42616 228636
rect 42668 228624 42674 228676
rect 42242 227468 42248 227520
rect 42300 227508 42306 227520
rect 42518 227508 42524 227520
rect 42300 227480 42524 227508
rect 42300 227468 42306 227480
rect 42518 227468 42524 227480
rect 42576 227468 42582 227520
rect 673822 203464 673828 203516
rect 673880 203504 673886 203516
rect 675294 203504 675300 203516
rect 673880 203476 675300 203504
rect 673880 203464 673886 203476
rect 675294 203464 675300 203476
rect 675352 203464 675358 203516
rect 673546 202308 673552 202360
rect 673604 202348 673610 202360
rect 675386 202348 675392 202360
rect 673604 202320 675392 202348
rect 673604 202308 673610 202320
rect 675386 202308 675392 202320
rect 675444 202308 675450 202360
rect 673638 199248 673644 199300
rect 673696 199288 673702 199300
rect 675386 199288 675392 199300
rect 673696 199260 675392 199288
rect 673696 199248 673702 199260
rect 675386 199248 675392 199260
rect 675444 199248 675450 199300
rect 673730 199044 673736 199096
rect 673788 199084 673794 199096
rect 675386 199084 675392 199096
rect 673788 199056 675392 199084
rect 673788 199044 673794 199056
rect 675386 199044 675392 199056
rect 675444 199044 675450 199096
rect 41782 195848 41788 195900
rect 41840 195888 41846 195900
rect 42518 195888 42524 195900
rect 41840 195860 42524 195888
rect 41840 195848 41846 195860
rect 42518 195848 42524 195860
rect 42576 195848 42582 195900
rect 673914 191904 673920 191956
rect 673972 191944 673978 191956
rect 675386 191944 675392 191956
rect 673972 191916 675392 191944
rect 673972 191904 673978 191916
rect 675386 191904 675392 191916
rect 675444 191904 675450 191956
rect 41782 189116 41788 189168
rect 41840 189156 41846 189168
rect 42426 189156 42432 189168
rect 41840 189128 42432 189156
rect 41840 189116 41846 189128
rect 42426 189116 42432 189128
rect 42484 189116 42490 189168
rect 41966 187552 41972 187604
rect 42024 187592 42030 187604
rect 42518 187592 42524 187604
rect 42024 187564 42524 187592
rect 42024 187552 42030 187564
rect 42518 187552 42524 187564
rect 42576 187552 42582 187604
rect 41782 184424 41788 184476
rect 41840 184464 41846 184476
rect 42610 184464 42616 184476
rect 41840 184436 42616 184464
rect 41840 184424 41846 184436
rect 42260 184204 42288 184436
rect 42610 184424 42616 184436
rect 42668 184424 42674 184476
rect 42242 184152 42248 184204
rect 42300 184152 42306 184204
rect 673730 158584 673736 158636
rect 673788 158624 673794 158636
rect 675386 158624 675392 158636
rect 673788 158596 675392 158624
rect 673788 158584 673794 158596
rect 675386 158584 675392 158596
rect 675444 158584 675450 158636
rect 673546 158312 673552 158364
rect 673604 158352 673610 158364
rect 675386 158352 675392 158364
rect 673604 158324 675392 158352
rect 673604 158312 673610 158324
rect 675386 158312 675392 158324
rect 675444 158312 675450 158364
rect 673638 155184 673644 155236
rect 673696 155224 673702 155236
rect 675386 155224 675392 155236
rect 673696 155196 675392 155224
rect 673696 155184 673702 155196
rect 675386 155184 675392 155196
rect 675444 155184 675450 155236
rect 673730 154096 673736 154148
rect 673788 154136 673794 154148
rect 675294 154136 675300 154148
rect 673788 154108 675300 154136
rect 673788 154096 673794 154108
rect 675294 154096 675300 154108
rect 675352 154096 675358 154148
rect 673822 146888 673828 146940
rect 673880 146928 673886 146940
rect 675386 146928 675392 146940
rect 673880 146900 675392 146928
rect 673880 146888 673886 146900
rect 675386 146888 675392 146900
rect 675444 146888 675450 146940
rect 42518 121456 42524 121508
rect 42576 121496 42582 121508
rect 44174 121496 44180 121508
rect 42576 121468 44180 121496
rect 42576 121456 42582 121468
rect 44174 121456 44180 121468
rect 44232 121456 44238 121508
rect 673638 113704 673644 113756
rect 673696 113744 673702 113756
rect 675386 113744 675392 113756
rect 673696 113716 675392 113744
rect 673696 113704 673702 113716
rect 675386 113704 675392 113716
rect 675444 113704 675450 113756
rect 673454 113160 673460 113212
rect 673512 113200 673518 113212
rect 675386 113200 675392 113212
rect 673512 113172 675392 113200
rect 673512 113160 673518 113172
rect 675386 113160 675392 113172
rect 675444 113160 675450 113212
rect 673546 109488 673552 109540
rect 673604 109528 673610 109540
rect 675386 109528 675392 109540
rect 673604 109500 675392 109528
rect 673604 109488 673610 109500
rect 675386 109488 675392 109500
rect 675444 109488 675450 109540
rect 673638 108400 673644 108452
rect 673696 108440 673702 108452
rect 675386 108440 675392 108452
rect 673696 108412 675392 108440
rect 673696 108400 673702 108412
rect 675386 108400 675392 108412
rect 675444 108400 675450 108452
rect 673730 101668 673736 101720
rect 673788 101708 673794 101720
rect 675386 101708 675392 101720
rect 673788 101680 675392 101708
rect 673788 101668 673794 101680
rect 675386 101668 675392 101680
rect 675444 101668 675450 101720
rect 42426 82832 42432 82884
rect 42484 82872 42490 82884
rect 44174 82872 44180 82884
rect 42484 82844 44180 82872
rect 42484 82832 42490 82844
rect 44174 82832 44180 82844
rect 44232 82832 44238 82884
rect 44818 46928 44824 46980
rect 44876 46928 44882 46980
rect 673638 46968 673644 46980
rect 200868 46940 297772 46968
rect 44836 46900 44864 46928
rect 200868 46912 200896 46940
rect 143534 46900 143540 46912
rect 44836 46872 143540 46900
rect 143534 46860 143540 46872
rect 143592 46860 143598 46912
rect 200850 46860 200856 46912
rect 200908 46860 200914 46912
rect 240888 46900 240916 46940
rect 297744 46912 297772 46940
rect 309428 46940 352604 46968
rect 309428 46912 309456 46940
rect 352576 46912 352604 46940
rect 364260 46940 407436 46968
rect 364260 46912 364288 46940
rect 407408 46912 407436 46940
rect 419092 46940 462176 46968
rect 419092 46912 419120 46940
rect 462148 46912 462176 46940
rect 473832 46940 517008 46968
rect 473832 46912 473860 46940
rect 516980 46912 517008 46940
rect 527468 46940 673644 46968
rect 527468 46912 527496 46940
rect 673638 46928 673644 46940
rect 673696 46928 673702 46980
rect 256234 46900 256240 46912
rect 240888 46872 256240 46900
rect 256234 46860 256240 46872
rect 256292 46860 256298 46912
rect 297726 46860 297732 46912
rect 297784 46860 297790 46912
rect 309410 46860 309416 46912
rect 309468 46860 309474 46912
rect 352558 46860 352564 46912
rect 352616 46860 352622 46912
rect 364242 46860 364248 46912
rect 364300 46860 364306 46912
rect 407390 46860 407396 46912
rect 407448 46860 407454 46912
rect 419074 46860 419080 46912
rect 419132 46860 419138 46912
rect 462130 46860 462136 46912
rect 462188 46860 462194 46912
rect 473814 46860 473820 46912
rect 473872 46860 473878 46912
rect 516962 46860 516968 46912
rect 517020 46860 517026 46912
rect 527450 46860 527456 46912
rect 527508 46860 527514 46912
rect 42242 45636 42248 45688
rect 42300 45676 42306 45688
rect 140958 45676 140964 45688
rect 42300 45648 140964 45676
rect 42300 45636 42306 45648
rect 140958 45636 140964 45648
rect 141016 45636 141022 45688
rect 42334 45568 42340 45620
rect 42392 45608 42398 45620
rect 143626 45608 143632 45620
rect 42392 45580 143632 45608
rect 42392 45568 42398 45580
rect 143626 45568 143632 45580
rect 143684 45568 143690 45620
rect 186682 45568 186688 45620
rect 186740 45608 186746 45620
rect 194686 45608 194692 45620
rect 186740 45580 194692 45608
rect 186740 45568 186746 45580
rect 194686 45568 194692 45580
rect 194744 45568 194750 45620
rect 523770 45568 523776 45620
rect 523828 45608 523834 45620
rect 673546 45608 673552 45620
rect 523828 45580 673552 45608
rect 523828 45568 523834 45580
rect 673546 45568 673552 45580
rect 673604 45568 673610 45620
rect 44910 45500 44916 45552
rect 44968 45540 44974 45552
rect 195974 45540 195980 45552
rect 44968 45512 195980 45540
rect 44968 45500 44974 45512
rect 195974 45500 195980 45512
rect 196032 45500 196038 45552
rect 518710 45500 518716 45552
rect 518768 45540 518774 45552
rect 673730 45540 673736 45552
rect 518768 45512 673736 45540
rect 518768 45500 518774 45512
rect 673730 45500 673736 45512
rect 673788 45500 673794 45552
rect 349982 44412 349988 44464
rect 350040 44452 350046 44464
rect 359366 44452 359372 44464
rect 350040 44424 359372 44452
rect 350040 44412 350046 44424
rect 359366 44412 359372 44424
rect 359424 44452 359430 44464
rect 414198 44452 414204 44464
rect 359424 44424 414204 44452
rect 359424 44412 359430 44424
rect 414198 44412 414204 44424
rect 414256 44412 414262 44464
rect 188522 44344 188528 44396
rect 188580 44384 188586 44396
rect 192846 44384 192852 44396
rect 188580 44356 192852 44384
rect 188580 44344 188586 44356
rect 192846 44344 192852 44356
rect 192904 44384 192910 44396
rect 297082 44384 297088 44396
rect 192904 44356 201540 44384
rect 192904 44344 192910 44356
rect 201512 44328 201540 44356
rect 284266 44356 297088 44384
rect 195974 44276 195980 44328
rect 196032 44316 196038 44328
rect 196032 44288 199792 44316
rect 196032 44276 196038 44288
rect 143626 44140 143632 44192
rect 143684 44180 143690 44192
rect 145098 44180 145104 44192
rect 143684 44152 145104 44180
rect 143684 44140 143690 44152
rect 145098 44140 145104 44152
rect 145156 44180 145162 44192
rect 195330 44180 195336 44192
rect 145156 44152 195336 44180
rect 145156 44140 145162 44152
rect 195330 44140 195336 44152
rect 195388 44180 195394 44192
rect 199654 44180 199660 44192
rect 195388 44152 199660 44180
rect 195388 44140 195394 44152
rect 199654 44140 199660 44152
rect 199712 44140 199718 44192
rect 199764 44180 199792 44288
rect 201494 44276 201500 44328
rect 201552 44316 201558 44328
rect 284266 44316 284294 44356
rect 297082 44344 297088 44356
rect 297140 44384 297146 44396
rect 299566 44384 299572 44396
rect 297140 44356 299572 44384
rect 297140 44344 297146 44356
rect 299566 44344 299572 44356
rect 299624 44384 299630 44396
rect 305730 44384 305736 44396
rect 299624 44356 305736 44384
rect 299624 44344 299630 44356
rect 305730 44344 305736 44356
rect 305788 44384 305794 44396
rect 305788 44356 322934 44384
rect 305788 44344 305794 44356
rect 201552 44288 284294 44316
rect 201552 44276 201558 44288
rect 295242 44276 295248 44328
rect 295300 44316 295306 44328
rect 303246 44316 303252 44328
rect 295300 44288 303252 44316
rect 295300 44276 295306 44288
rect 303246 44276 303252 44288
rect 303304 44276 303310 44328
rect 322906 44316 322934 44356
rect 468938 44344 468944 44396
rect 468996 44384 469002 44396
rect 523770 44384 523776 44396
rect 468996 44356 523776 44384
rect 468996 44344 469002 44356
rect 523770 44344 523776 44356
rect 523828 44344 523834 44396
rect 351914 44316 351920 44328
rect 303586 44288 303936 44316
rect 322906 44288 351920 44316
rect 199838 44208 199844 44260
rect 199896 44248 199902 44260
rect 303586 44248 303614 44288
rect 303908 44260 303936 44288
rect 351914 44276 351920 44288
rect 351972 44316 351978 44328
rect 354398 44316 354404 44328
rect 351972 44288 354404 44316
rect 351972 44276 351978 44288
rect 354398 44276 354404 44288
rect 354456 44316 354462 44328
rect 360562 44316 360568 44328
rect 354456 44288 360568 44316
rect 354456 44276 354462 44288
rect 360562 44276 360568 44288
rect 360620 44276 360626 44328
rect 363046 44316 363052 44328
rect 361546 44288 363052 44316
rect 199896 44220 303614 44248
rect 199896 44208 199902 44220
rect 303890 44208 303896 44260
rect 303948 44248 303954 44260
rect 308214 44248 308220 44260
rect 303948 44220 308220 44248
rect 303948 44208 303954 44220
rect 308214 44208 308220 44220
rect 308272 44248 308278 44260
rect 358722 44248 358728 44260
rect 308272 44220 358728 44248
rect 308272 44208 308278 44220
rect 358722 44208 358728 44220
rect 358780 44248 358786 44260
rect 361546 44248 361574 44288
rect 363046 44276 363052 44288
rect 363104 44316 363110 44328
rect 413554 44316 413560 44328
rect 363104 44288 413560 44316
rect 363104 44276 363110 44288
rect 413554 44276 413560 44288
rect 413612 44316 413618 44328
rect 417878 44316 417884 44328
rect 413612 44288 417884 44316
rect 413612 44276 413618 44288
rect 417878 44276 417884 44288
rect 417936 44316 417942 44328
rect 468294 44316 468300 44328
rect 417936 44288 468300 44316
rect 417936 44276 417942 44288
rect 468294 44276 468300 44288
rect 468352 44316 468358 44328
rect 472618 44316 472624 44328
rect 468352 44288 472624 44316
rect 468352 44276 468358 44288
rect 472618 44276 472624 44288
rect 472676 44316 472682 44328
rect 472676 44288 523172 44316
rect 472676 44276 472682 44288
rect 406746 44248 406752 44260
rect 358780 44220 361574 44248
rect 380866 44220 406752 44248
rect 358780 44208 358786 44220
rect 304534 44180 304540 44192
rect 199764 44152 304540 44180
rect 304534 44140 304540 44152
rect 304592 44180 304598 44192
rect 349982 44180 349988 44192
rect 304592 44152 349988 44180
rect 304592 44140 304598 44152
rect 349982 44140 349988 44152
rect 350040 44140 350046 44192
rect 350074 44140 350080 44192
rect 350132 44180 350138 44192
rect 358078 44180 358084 44192
rect 350132 44152 358084 44180
rect 350132 44140 350138 44152
rect 358078 44140 358084 44152
rect 358136 44140 358142 44192
rect 360562 44140 360568 44192
rect 360620 44180 360626 44192
rect 380866 44180 380894 44220
rect 406746 44208 406752 44220
rect 406804 44248 406810 44260
rect 461486 44248 461492 44260
rect 406804 44220 461492 44248
rect 406804 44208 406810 44220
rect 461486 44208 461492 44220
rect 461544 44248 461550 44260
rect 516318 44248 516324 44260
rect 461544 44220 516324 44248
rect 461544 44208 461550 44220
rect 516318 44208 516324 44220
rect 516376 44248 516382 44260
rect 518710 44248 518716 44260
rect 516376 44220 518716 44248
rect 516376 44208 516382 44220
rect 518710 44208 518716 44220
rect 518768 44208 518774 44260
rect 523144 44192 523172 44288
rect 360620 44152 380894 44180
rect 360620 44140 360626 44152
rect 414198 44140 414204 44192
rect 414256 44180 414262 44192
rect 468938 44180 468944 44192
rect 414256 44152 468944 44180
rect 414256 44140 414262 44152
rect 468938 44140 468944 44152
rect 468996 44140 469002 44192
rect 523126 44140 523132 44192
rect 523184 44180 523190 44192
rect 527450 44180 527456 44192
rect 523184 44152 527456 44180
rect 523184 44140 523190 44152
rect 527450 44140 527456 44152
rect 527508 44140 527514 44192
rect 579890 42712 579896 42764
rect 579948 42752 579954 42764
rect 673454 42752 673460 42764
rect 579948 42724 673460 42752
rect 579948 42712 579954 42724
rect 673454 42712 673460 42724
rect 673512 42712 673518 42764
rect 189258 41896 189264 41948
rect 189316 41936 189322 41948
rect 191098 41936 191104 41948
rect 189316 41908 191104 41936
rect 189316 41896 189322 41908
rect 191098 41896 191104 41908
rect 191156 41936 191162 41948
rect 192294 41936 192300 41948
rect 191156 41908 192300 41936
rect 191156 41896 191162 41908
rect 192294 41896 192300 41908
rect 192352 41936 192358 41948
rect 193582 41936 193588 41948
rect 192352 41908 193588 41936
rect 192352 41896 192358 41908
rect 193582 41896 193588 41908
rect 193640 41936 193646 41948
rect 196434 41936 196440 41948
rect 193640 41908 196440 41936
rect 193640 41896 193646 41908
rect 196434 41896 196440 41908
rect 196492 41896 196498 41948
rect 198458 41896 198464 41948
rect 198516 41936 198522 41948
rect 200114 41936 200120 41948
rect 198516 41908 200120 41936
rect 198516 41896 198522 41908
rect 200114 41896 200120 41908
rect 200172 41896 200178 41948
rect 297910 41896 297916 41948
rect 297968 41936 297974 41948
rect 300670 41936 300676 41948
rect 297968 41908 300676 41936
rect 297968 41896 297974 41908
rect 300670 41896 300676 41908
rect 300728 41896 300734 41948
rect 302234 41896 302240 41948
rect 302292 41936 302298 41948
rect 305270 41936 305276 41948
rect 302292 41908 305276 41936
rect 302292 41896 302298 41908
rect 305270 41896 305276 41908
rect 305328 41936 305334 41948
rect 306558 41936 306564 41948
rect 305328 41908 306564 41936
rect 305328 41896 305334 41908
rect 306558 41896 306564 41908
rect 306616 41936 306622 41948
rect 308674 41936 308680 41948
rect 306616 41908 308680 41936
rect 306616 41896 306622 41908
rect 308674 41896 308680 41908
rect 308732 41896 308738 41948
rect 352650 41896 352656 41948
rect 352708 41936 352714 41948
rect 355502 41936 355508 41948
rect 352708 41908 355508 41936
rect 352708 41896 352714 41908
rect 355502 41896 355508 41908
rect 355560 41896 355566 41948
rect 356974 41896 356980 41948
rect 357032 41936 357038 41948
rect 359826 41936 359832 41948
rect 357032 41908 359832 41936
rect 357032 41896 357038 41908
rect 359826 41896 359832 41908
rect 359884 41936 359890 41948
rect 361114 41936 361120 41948
rect 359884 41908 361120 41936
rect 359884 41896 359890 41908
rect 361114 41896 361120 41908
rect 361172 41936 361178 41948
rect 363506 41936 363512 41948
rect 361172 41908 363512 41936
rect 361172 41896 361178 41908
rect 363506 41896 363512 41908
rect 363564 41896 363570 41948
rect 407482 41896 407488 41948
rect 407540 41936 407546 41948
rect 410242 41936 410248 41948
rect 407540 41908 410248 41936
rect 407540 41896 407546 41908
rect 410242 41896 410248 41908
rect 410300 41936 410306 41948
rect 411530 41936 411536 41948
rect 410300 41908 411536 41936
rect 410300 41896 410306 41908
rect 411530 41896 411536 41908
rect 411588 41936 411594 41948
rect 414566 41936 414572 41948
rect 411588 41908 414572 41936
rect 411588 41896 411594 41908
rect 414566 41896 414572 41908
rect 414624 41936 414630 41948
rect 415854 41936 415860 41948
rect 414624 41908 415860 41936
rect 414624 41896 414630 41908
rect 415854 41896 415860 41908
rect 415912 41936 415918 41948
rect 418246 41936 418252 41948
rect 415912 41908 418252 41936
rect 415912 41896 415918 41908
rect 418246 41896 418252 41908
rect 418304 41896 418310 41948
rect 462314 41896 462320 41948
rect 462372 41936 462378 41948
rect 465074 41936 465080 41948
rect 462372 41908 465080 41936
rect 462372 41896 462378 41908
rect 465074 41896 465080 41908
rect 465132 41936 465138 41948
rect 466362 41936 466368 41948
rect 465132 41908 466368 41936
rect 465132 41896 465138 41908
rect 466362 41896 466368 41908
rect 466420 41936 466426 41948
rect 469398 41936 469404 41948
rect 466420 41908 469404 41936
rect 466420 41896 466426 41908
rect 469398 41896 469404 41908
rect 469456 41936 469462 41948
rect 470686 41936 470692 41948
rect 469456 41908 470692 41936
rect 469456 41896 469462 41908
rect 470686 41896 470692 41908
rect 470744 41936 470750 41948
rect 473078 41936 473084 41948
rect 470744 41908 473084 41936
rect 470744 41896 470750 41908
rect 473078 41896 473084 41908
rect 473136 41896 473142 41948
rect 517054 41896 517060 41948
rect 517112 41936 517118 41948
rect 519906 41936 519912 41948
rect 517112 41908 519912 41936
rect 517112 41896 517118 41908
rect 519906 41896 519912 41908
rect 519964 41936 519970 41948
rect 521194 41936 521200 41948
rect 519964 41908 521200 41936
rect 519964 41896 519970 41908
rect 521194 41896 521200 41908
rect 521252 41936 521258 41948
rect 524230 41936 524236 41948
rect 521252 41908 524236 41936
rect 521252 41896 521258 41908
rect 524230 41896 524236 41908
rect 524288 41936 524294 41948
rect 525518 41936 525524 41948
rect 524288 41908 525524 41936
rect 524288 41896 524294 41908
rect 525518 41896 525524 41908
rect 525576 41936 525582 41948
rect 527910 41936 527916 41948
rect 525576 41908 527916 41936
rect 525576 41896 525582 41908
rect 527910 41896 527916 41908
rect 527968 41896 527974 41948
rect 146294 41828 146300 41880
rect 146352 41868 146358 41880
rect 568850 41868 568856 41880
rect 146352 41840 568856 41868
rect 146352 41828 146358 41840
rect 568850 41828 568856 41840
rect 568908 41868 568914 41880
rect 579890 41868 579896 41880
rect 568908 41840 579896 41868
rect 568908 41828 568914 41840
rect 579890 41828 579896 41840
rect 579948 41828 579954 41880
rect 198918 41800 198924 41812
rect 168346 41772 198924 41800
rect 93762 41488 93768 41540
rect 93820 41528 93826 41540
rect 168346 41528 168374 41772
rect 198918 41760 198924 41772
rect 198976 41800 198982 41812
rect 307754 41800 307760 41812
rect 198976 41772 307760 41800
rect 198976 41760 198982 41772
rect 307754 41760 307760 41772
rect 307812 41800 307818 41812
rect 362494 41800 362500 41812
rect 307812 41772 362500 41800
rect 307812 41760 307818 41772
rect 362494 41760 362500 41772
rect 362552 41800 362558 41812
rect 362552 41772 380894 41800
rect 362552 41760 362558 41772
rect 93820 41500 168374 41528
rect 380866 41528 380894 41772
rect 409322 41760 409328 41812
rect 409380 41800 409386 41812
rect 412358 41800 412364 41812
rect 409380 41772 412364 41800
rect 409380 41760 409386 41772
rect 412358 41760 412364 41772
rect 412416 41800 412422 41812
rect 415210 41800 415216 41812
rect 412416 41772 415216 41800
rect 412416 41760 412422 41772
rect 415210 41760 415216 41772
rect 415268 41760 415274 41812
rect 417326 41800 417332 41812
rect 417252 41772 417332 41800
rect 417252 41528 417280 41772
rect 417326 41760 417332 41772
rect 417384 41760 417390 41812
rect 464154 41760 464160 41812
rect 464212 41800 464218 41812
rect 467190 41800 467196 41812
rect 464212 41772 467196 41800
rect 464212 41760 464218 41772
rect 467190 41760 467196 41772
rect 467248 41800 467254 41812
rect 470042 41800 470048 41812
rect 467248 41772 470048 41800
rect 467248 41760 467254 41772
rect 470042 41760 470048 41772
rect 470100 41760 470106 41812
rect 472158 41800 472164 41812
rect 472084 41772 472164 41800
rect 472084 41528 472112 41772
rect 472158 41760 472164 41772
rect 472216 41760 472222 41812
rect 526714 41800 526720 41812
rect 516106 41772 526720 41800
rect 516106 41528 516134 41772
rect 526714 41760 526720 41772
rect 526772 41760 526778 41812
rect 380866 41500 516134 41528
rect 93820 41488 93826 41500
rect 135162 40196 135168 40248
rect 135220 40236 135226 40248
rect 143534 40236 143540 40248
rect 135220 40208 143540 40236
rect 135220 40196 135226 40208
rect 143534 40196 143540 40208
rect 143592 40196 143598 40248
rect 140990 40060 140996 40112
rect 141048 40100 141054 40112
rect 143066 40100 143072 40112
rect 141048 40072 143072 40100
rect 141048 40060 141054 40072
rect 142586 39950 142614 40072
rect 143066 40060 143072 40072
rect 143124 40100 143130 40112
rect 144546 40100 144552 40112
rect 143124 40072 144552 40100
rect 143124 40060 143130 40072
rect 144546 40060 144552 40072
rect 144604 40100 144610 40112
rect 146294 40100 146300 40112
rect 144604 40072 146300 40100
rect 144604 40060 144610 40072
rect 146294 40060 146300 40072
rect 146352 40060 146358 40112
<< via1 >>
rect 585048 996344 585100 996396
rect 674748 996344 674800 996396
rect 342168 990836 342220 990888
rect 673552 990836 673604 990888
rect 42248 990156 42300 990208
rect 342260 990156 342312 990208
rect 44916 990088 44968 990140
rect 673460 990088 673512 990140
rect 42340 990020 42392 990072
rect 673644 990020 673696 990072
rect 673644 875780 673696 875832
rect 675392 875780 675444 875832
rect 673552 874488 673604 874540
rect 675392 874488 675444 874540
rect 673460 872380 673512 872432
rect 674012 872380 674064 872432
rect 675392 872380 675444 872432
rect 673736 871292 673788 871344
rect 675300 871292 675352 871344
rect 673920 870136 673972 870188
rect 675392 870136 675444 870188
rect 673828 864220 673880 864272
rect 675392 864220 675444 864272
rect 673920 863200 673972 863252
rect 675392 863200 675444 863252
rect 675300 818320 675352 818372
rect 677600 818320 677652 818372
rect 41788 797716 41840 797768
rect 42616 797716 42668 797768
rect 41788 791936 41840 791988
rect 42432 791936 42484 791988
rect 41788 791324 41840 791376
rect 42524 791324 42576 791376
rect 41788 786972 41840 787024
rect 42432 786972 42484 787024
rect 673736 785952 673788 786004
rect 675208 785952 675260 786004
rect 675392 785952 675444 786004
rect 673460 785680 673512 785732
rect 675392 785680 675444 785732
rect 673644 782280 673696 782332
rect 674012 782280 674064 782332
rect 675392 782280 675444 782332
rect 673736 781600 673788 781652
rect 675208 781600 675260 781652
rect 675392 781600 675444 781652
rect 675208 780988 675260 781040
rect 675392 780988 675444 781040
rect 673828 775820 673880 775872
rect 675392 775820 675444 775872
rect 42248 762220 42300 762272
rect 42524 762220 42576 762272
rect 41788 755420 41840 755472
rect 42616 755420 42668 755472
rect 41788 747668 41840 747720
rect 42432 747668 42484 747720
rect 41788 743996 41840 744048
rect 42524 743996 42576 744048
rect 673736 740936 673788 740988
rect 675208 740936 675260 740988
rect 675392 740936 675444 740988
rect 673460 740324 673512 740376
rect 675392 740324 675444 740376
rect 673644 738080 673696 738132
rect 675392 738080 675444 738132
rect 673736 736992 673788 737044
rect 675208 736992 675260 737044
rect 675392 736992 675444 737044
rect 673552 730872 673604 730924
rect 673920 730872 673972 730924
rect 675392 730872 675444 730924
rect 41788 712240 41840 712292
rect 42616 712240 42668 712292
rect 41788 703944 41840 703996
rect 42432 703944 42484 703996
rect 41788 700816 41840 700868
rect 42524 700816 42576 700868
rect 673736 695920 673788 695972
rect 675208 695920 675260 695972
rect 675392 695920 675444 695972
rect 673460 695308 673512 695360
rect 675392 695308 675444 695360
rect 673920 692248 673972 692300
rect 675392 692248 675444 692300
rect 673736 692044 673788 692096
rect 675208 692044 675260 692096
rect 675392 692044 675444 692096
rect 673552 685176 673604 685228
rect 675392 685176 675444 685228
rect 41788 668108 41840 668160
rect 42708 668108 42760 668160
rect 41788 661036 41840 661088
rect 42432 661036 42484 661088
rect 41788 658656 41840 658708
rect 42524 658656 42576 658708
rect 673736 651108 673788 651160
rect 675392 651108 675444 651160
rect 673460 650496 673512 650548
rect 675392 650496 675444 650548
rect 673460 647164 673512 647216
rect 673644 647164 673696 647216
rect 673460 647028 673512 647080
rect 673920 647028 673972 647080
rect 675392 647028 675444 647080
rect 673736 646416 673788 646468
rect 675392 646416 675444 646468
rect 675208 645736 675260 645788
rect 675392 645736 675444 645788
rect 673552 640636 673604 640688
rect 675392 640636 675444 640688
rect 41788 624928 41840 624980
rect 42524 624928 42576 624980
rect 42708 624928 42760 624980
rect 41788 618468 41840 618520
rect 42432 618468 42484 618520
rect 41788 615476 41840 615528
rect 42616 615476 42668 615528
rect 673736 605752 673788 605804
rect 675208 605752 675260 605804
rect 675392 605752 675444 605804
rect 673644 605072 673696 605124
rect 675392 605072 675444 605124
rect 673460 602896 673512 602948
rect 675392 602896 675444 602948
rect 673736 601808 673788 601860
rect 675208 601808 675260 601860
rect 675392 601808 675444 601860
rect 673552 595008 673604 595060
rect 675392 595008 675444 595060
rect 41788 582632 41840 582684
rect 42524 582632 42576 582684
rect 41788 574676 41840 574728
rect 42432 574676 42484 574728
rect 41788 571208 41840 571260
rect 42524 571208 42576 571260
rect 42708 571208 42760 571260
rect 673736 561212 673788 561264
rect 675208 561212 675260 561264
rect 675392 561212 675444 561264
rect 673644 560940 673696 560992
rect 675392 560940 675444 560992
rect 673460 557812 673512 557864
rect 675392 557812 675444 557864
rect 675208 557268 675260 557320
rect 675392 557268 675444 557320
rect 675208 555568 675260 555620
rect 675392 555568 675444 555620
rect 673552 550468 673604 550520
rect 675392 550468 675444 550520
rect 42340 545232 42392 545284
rect 42340 545028 42392 545080
rect 41788 539452 41840 539504
rect 42616 539452 42668 539504
rect 42248 532108 42300 532160
rect 42432 532108 42484 532160
rect 41788 531156 41840 531208
rect 42432 531156 42484 531208
rect 41788 528028 41840 528080
rect 42524 528028 42576 528080
rect 42708 528028 42760 528080
rect 675300 513748 675352 513800
rect 677692 513748 677744 513800
rect 674748 427796 674800 427848
rect 677508 427796 677560 427848
rect 41788 410932 41840 410984
rect 42524 410932 42576 410984
rect 41788 404472 41840 404524
rect 42432 404472 42484 404524
rect 42616 404472 42668 404524
rect 41788 400800 41840 400852
rect 42708 400800 42760 400852
rect 673552 382712 673604 382764
rect 675392 382712 675444 382764
rect 673736 379652 673788 379704
rect 675392 379652 675444 379704
rect 673644 379040 673696 379092
rect 675392 379040 675444 379092
rect 673460 372308 673512 372360
rect 675392 372308 675444 372360
rect 41788 368636 41840 368688
rect 42340 368636 42392 368688
rect 42524 368636 42576 368688
rect 41788 361292 41840 361344
rect 42340 361292 42392 361344
rect 41788 360680 41840 360732
rect 42616 360680 42668 360732
rect 41788 357212 41840 357264
rect 42524 357212 42576 357264
rect 42708 357212 42760 357264
rect 41788 356668 41840 356720
rect 42340 356668 42392 356720
rect 673552 337492 673604 337544
rect 675392 337492 675444 337544
rect 673920 334432 673972 334484
rect 675392 334432 675444 334484
rect 673644 334228 673696 334280
rect 675392 334228 675444 334280
rect 42248 330012 42300 330064
rect 42432 330012 42484 330064
rect 673460 328040 673512 328092
rect 675392 328040 675444 328092
rect 41788 325456 41840 325508
rect 42432 325456 42484 325508
rect 42800 325456 42852 325508
rect 41788 317160 41840 317212
rect 42616 317160 42668 317212
rect 41788 314032 41840 314084
rect 42524 314032 42576 314084
rect 42708 314032 42760 314084
rect 673644 293768 673696 293820
rect 675392 293768 675444 293820
rect 673552 293564 673604 293616
rect 675392 293564 675444 293616
rect 673920 289824 673972 289876
rect 675392 289824 675444 289876
rect 673460 282072 673512 282124
rect 673736 282072 673788 282124
rect 675392 282072 675444 282124
rect 41788 281324 41840 281376
rect 42432 281324 42484 281376
rect 42800 281324 42852 281376
rect 41788 274524 41840 274576
rect 42616 274524 42668 274576
rect 41788 271872 41840 271924
rect 42708 271872 42760 271924
rect 673644 249092 673696 249144
rect 675392 249092 675444 249144
rect 673552 248548 673604 248600
rect 675392 248548 675444 248600
rect 673920 244876 673972 244928
rect 675392 244876 675444 244928
rect 673644 243992 673696 244044
rect 673920 243992 673972 244044
rect 673828 243788 673880 243840
rect 675392 243788 675444 243840
rect 41788 238076 41840 238128
rect 42432 238076 42484 238128
rect 673920 237668 673972 237720
rect 675392 237668 675444 237720
rect 41788 231684 41840 231736
rect 42524 231684 42576 231736
rect 41788 228624 41840 228676
rect 42616 228624 42668 228676
rect 42248 227468 42300 227520
rect 42524 227468 42576 227520
rect 673828 203464 673880 203516
rect 675300 203464 675352 203516
rect 673552 202308 673604 202360
rect 675392 202308 675444 202360
rect 673644 199248 673696 199300
rect 675392 199248 675444 199300
rect 673736 199044 673788 199096
rect 675392 199044 675444 199096
rect 41788 195848 41840 195900
rect 42524 195848 42576 195900
rect 673920 191904 673972 191956
rect 675392 191904 675444 191956
rect 41788 189116 41840 189168
rect 42432 189116 42484 189168
rect 41972 187552 42024 187604
rect 42524 187552 42576 187604
rect 41788 184424 41840 184476
rect 42616 184424 42668 184476
rect 42248 184152 42300 184204
rect 673736 158584 673788 158636
rect 675392 158584 675444 158636
rect 673552 158312 673604 158364
rect 675392 158312 675444 158364
rect 673644 155184 673696 155236
rect 675392 155184 675444 155236
rect 673736 154096 673788 154148
rect 675300 154096 675352 154148
rect 673828 146888 673880 146940
rect 675392 146888 675444 146940
rect 42524 121456 42576 121508
rect 44180 121456 44232 121508
rect 673644 113704 673696 113756
rect 675392 113704 675444 113756
rect 673460 113160 673512 113212
rect 675392 113160 675444 113212
rect 673552 109488 673604 109540
rect 675392 109488 675444 109540
rect 673644 108400 673696 108452
rect 675392 108400 675444 108452
rect 673736 101668 673788 101720
rect 675392 101668 675444 101720
rect 42432 82832 42484 82884
rect 44180 82832 44232 82884
rect 44824 46928 44876 46980
rect 143540 46860 143592 46912
rect 200856 46860 200908 46912
rect 673644 46928 673696 46980
rect 256240 46860 256292 46912
rect 297732 46860 297784 46912
rect 309416 46860 309468 46912
rect 352564 46860 352616 46912
rect 364248 46860 364300 46912
rect 407396 46860 407448 46912
rect 419080 46860 419132 46912
rect 462136 46860 462188 46912
rect 473820 46860 473872 46912
rect 516968 46860 517020 46912
rect 527456 46860 527508 46912
rect 42248 45636 42300 45688
rect 140964 45636 141016 45688
rect 42340 45568 42392 45620
rect 143632 45568 143684 45620
rect 186688 45568 186740 45620
rect 194692 45568 194744 45620
rect 523776 45568 523828 45620
rect 673552 45568 673604 45620
rect 44916 45500 44968 45552
rect 195980 45500 196032 45552
rect 518716 45500 518768 45552
rect 673736 45500 673788 45552
rect 349988 44412 350040 44464
rect 359372 44412 359424 44464
rect 414204 44412 414256 44464
rect 188528 44344 188580 44396
rect 192852 44344 192904 44396
rect 195980 44276 196032 44328
rect 143632 44140 143684 44192
rect 145104 44140 145156 44192
rect 195336 44140 195388 44192
rect 199660 44140 199712 44192
rect 201500 44276 201552 44328
rect 297088 44344 297140 44396
rect 299572 44344 299624 44396
rect 305736 44344 305788 44396
rect 295248 44276 295300 44328
rect 303252 44276 303304 44328
rect 468944 44344 468996 44396
rect 523776 44344 523828 44396
rect 199844 44208 199896 44260
rect 351920 44276 351972 44328
rect 354404 44276 354456 44328
rect 360568 44276 360620 44328
rect 303896 44208 303948 44260
rect 308220 44208 308272 44260
rect 358728 44208 358780 44260
rect 363052 44276 363104 44328
rect 413560 44276 413612 44328
rect 417884 44276 417936 44328
rect 468300 44276 468352 44328
rect 472624 44276 472676 44328
rect 304540 44140 304592 44192
rect 349988 44140 350040 44192
rect 350080 44140 350132 44192
rect 358084 44140 358136 44192
rect 360568 44140 360620 44192
rect 406752 44208 406804 44260
rect 461492 44208 461544 44260
rect 516324 44208 516376 44260
rect 518716 44208 518768 44260
rect 414204 44140 414256 44192
rect 468944 44140 468996 44192
rect 523132 44140 523184 44192
rect 527456 44140 527508 44192
rect 579896 42712 579948 42764
rect 673460 42712 673512 42764
rect 189264 41896 189316 41948
rect 191104 41896 191156 41948
rect 192300 41896 192352 41948
rect 193588 41896 193640 41948
rect 196440 41896 196492 41948
rect 198464 41896 198516 41948
rect 200120 41896 200172 41948
rect 297916 41896 297968 41948
rect 300676 41896 300728 41948
rect 302240 41896 302292 41948
rect 305276 41896 305328 41948
rect 306564 41896 306616 41948
rect 308680 41896 308732 41948
rect 352656 41896 352708 41948
rect 355508 41896 355560 41948
rect 356980 41896 357032 41948
rect 359832 41896 359884 41948
rect 361120 41896 361172 41948
rect 363512 41896 363564 41948
rect 407488 41896 407540 41948
rect 410248 41896 410300 41948
rect 411536 41896 411588 41948
rect 414572 41896 414624 41948
rect 415860 41896 415912 41948
rect 418252 41896 418304 41948
rect 462320 41896 462372 41948
rect 465080 41896 465132 41948
rect 466368 41896 466420 41948
rect 469404 41896 469456 41948
rect 470692 41896 470744 41948
rect 473084 41896 473136 41948
rect 517060 41896 517112 41948
rect 519912 41896 519964 41948
rect 521200 41896 521252 41948
rect 524236 41896 524288 41948
rect 525524 41896 525576 41948
rect 527916 41896 527968 41948
rect 146300 41828 146352 41880
rect 568856 41828 568908 41880
rect 579896 41828 579948 41880
rect 93768 41488 93820 41540
rect 198924 41760 198976 41812
rect 307760 41760 307812 41812
rect 362500 41760 362552 41812
rect 409328 41760 409380 41812
rect 412364 41760 412416 41812
rect 415216 41760 415268 41812
rect 417332 41760 417384 41812
rect 464160 41760 464212 41812
rect 467196 41760 467248 41812
rect 470048 41760 470100 41812
rect 472164 41760 472216 41812
rect 526720 41760 526772 41812
rect 135168 40196 135220 40248
rect 143540 40196 143592 40248
rect 140996 40060 141048 40112
rect 143072 40060 143124 40112
rect 144552 40060 144604 40112
rect 146300 40060 146352 40112
<< metal2 >>
rect 230499 997600 235279 998010
rect 240478 997600 245258 1002732
rect 282099 997600 286879 998010
rect 292078 997600 296858 1002732
rect 383899 997600 388679 998010
rect 393878 997600 398658 1002732
rect 342166 997520 342222 997529
rect 342166 997455 342222 997464
rect 585046 997520 585102 997529
rect 585046 997455 585102 997464
rect 342180 990894 342208 997455
rect 585060 996402 585088 997455
rect 585048 996396 585100 996402
rect 585048 996338 585100 996344
rect 674748 996396 674800 996402
rect 674748 996338 674800 996344
rect 342168 990888 342220 990894
rect 673552 990888 673604 990894
rect 342220 990836 342300 990842
rect 342168 990830 342300 990836
rect 673552 990830 673604 990836
rect 342180 990814 342300 990830
rect 342180 990765 342208 990814
rect 342272 990214 342300 990814
rect 42248 990208 42300 990214
rect 42248 990150 42300 990156
rect 342260 990208 342312 990214
rect 342260 990150 342312 990156
rect 42260 800170 42288 990150
rect 44916 990140 44968 990146
rect 44916 990082 44968 990088
rect 673460 990140 673512 990146
rect 673460 990082 673512 990088
rect 42340 990072 42392 990078
rect 42340 990014 42392 990020
rect 42352 800306 42380 990014
rect 44928 888734 44956 990082
rect 44836 888706 44956 888734
rect 44836 870097 44864 888706
rect 673472 872438 673500 990082
rect 673564 874546 673592 990830
rect 673644 990072 673696 990078
rect 673644 990014 673696 990020
rect 673656 875838 673684 990014
rect 673644 875832 673696 875838
rect 673644 875774 673696 875780
rect 673552 874540 673604 874546
rect 673552 874482 673604 874488
rect 673460 872432 673512 872438
rect 673460 872374 673512 872380
rect 42430 870088 42486 870097
rect 42430 870023 42486 870032
rect 44822 870088 44878 870097
rect 44822 870023 44878 870032
rect 42444 805934 42472 870023
rect 42444 805906 42564 805934
rect 42352 800278 42472 800306
rect 42260 800142 42380 800170
rect 41722 800075 42288 800103
rect 41713 799417 42193 799473
rect 41722 798238 41828 798266
rect 41800 797774 41828 798238
rect 41788 797768 41840 797774
rect 41788 797710 41840 797716
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 795093 42193 795149
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 42260 792282 42288 800075
rect 41892 792254 42288 792282
rect 41892 792099 41920 792254
rect 41722 792071 41920 792099
rect 41788 791988 41840 791994
rect 41788 791930 41840 791936
rect 41800 791466 41828 791930
rect 41722 791438 41828 791466
rect 41788 791376 41840 791382
rect 41788 791318 41840 791324
rect 41800 790786 41828 791318
rect 41722 790758 41828 790786
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 42352 787930 42380 800142
rect 42444 791994 42472 800278
rect 42432 791988 42484 791994
rect 42432 791930 42484 791936
rect 41800 787902 42380 787930
rect 41800 787794 41828 787902
rect 41722 787766 41828 787794
rect 41722 787086 41828 787114
rect 41800 787030 41828 787086
rect 41788 787024 41840 787030
rect 41788 786966 41840 786972
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 41713 784697 42193 784753
rect 42260 762278 42288 787902
rect 42444 787030 42472 791930
rect 42536 791382 42564 805906
rect 42616 797768 42668 797774
rect 42616 797710 42668 797716
rect 42524 791376 42576 791382
rect 42524 791318 42576 791324
rect 42432 787024 42484 787030
rect 42432 786966 42484 786972
rect 42444 786706 42472 786966
rect 42352 786678 42472 786706
rect 42248 762272 42300 762278
rect 42248 762214 42300 762220
rect 41722 756894 42288 756922
rect 41713 756217 42193 756273
rect 41788 755472 41840 755478
rect 41788 755414 41840 755420
rect 41800 755063 41828 755414
rect 41722 755035 41828 755063
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751893 42193 751949
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 42260 749034 42288 756894
rect 41800 749006 42288 749034
rect 41800 748898 41828 749006
rect 41722 748870 41828 748898
rect 42352 748255 42380 786678
rect 42536 786614 42564 791318
rect 41722 748227 42380 748255
rect 42352 747974 42380 748227
rect 42260 747946 42380 747974
rect 42444 786586 42564 786614
rect 41788 747720 41840 747726
rect 41788 747662 41840 747668
rect 41800 747611 41828 747662
rect 41722 747583 41828 747611
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 41722 744547 41828 744575
rect 41800 744054 41828 744547
rect 41788 744048 41840 744054
rect 41788 743990 41840 743996
rect 42260 743931 42288 747946
rect 42444 747726 42472 786586
rect 42524 762272 42576 762278
rect 42524 762214 42576 762220
rect 42432 747720 42484 747726
rect 42432 747662 42484 747668
rect 41722 743903 42288 743931
rect 41713 743337 42193 743393
rect 41713 742693 42193 742749
rect 41713 742049 42193 742105
rect 41713 741497 42193 741553
rect 42260 728654 42288 743903
rect 42260 728626 42380 728654
rect 41722 713675 42288 713703
rect 41713 713017 42193 713073
rect 41788 712292 41840 712298
rect 41788 712234 41840 712240
rect 41800 711863 41828 712234
rect 41722 711835 41828 711863
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708693 42193 708749
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 42260 706194 42288 713675
rect 41800 706166 42288 706194
rect 41800 705699 41828 706166
rect 41722 705671 41828 705699
rect 41722 705027 41920 705055
rect 41892 704970 41920 705027
rect 42352 704970 42380 728626
rect 41892 704942 42380 704970
rect 41722 704398 41828 704426
rect 41800 704002 41828 704398
rect 41788 703996 41840 704002
rect 41788 703938 41840 703944
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 41722 701347 41828 701375
rect 41800 700874 41828 701347
rect 41788 700868 41840 700874
rect 41788 700810 41840 700816
rect 41722 700726 41920 700754
rect 41892 700618 41920 700726
rect 42260 700618 42288 704942
rect 42444 704002 42472 747662
rect 42536 744054 42564 762214
rect 42628 755478 42656 797710
rect 673564 786614 673592 874482
rect 674012 872432 674064 872438
rect 674012 872374 674064 872380
rect 673736 871344 673788 871350
rect 673736 871286 673788 871292
rect 673472 786586 673592 786614
rect 673472 785738 673500 786586
rect 673748 786010 673776 871286
rect 673920 870188 673972 870194
rect 673920 870130 673972 870136
rect 673828 864272 673880 864278
rect 673828 864214 673880 864220
rect 673736 786004 673788 786010
rect 673736 785946 673788 785952
rect 673460 785732 673512 785738
rect 673460 785674 673512 785680
rect 42616 755472 42668 755478
rect 42616 755414 42668 755420
rect 42524 744048 42576 744054
rect 42524 743990 42576 743996
rect 42432 703996 42484 704002
rect 42432 703938 42484 703944
rect 41892 700590 42288 700618
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 41713 698297 42193 698353
rect 42260 690014 42288 700590
rect 42260 689986 42380 690014
rect 41722 670475 42288 670503
rect 41713 669817 42193 669873
rect 41722 668630 41828 668658
rect 41800 668166 41828 668630
rect 41788 668160 41840 668166
rect 41788 668102 41840 668108
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 665493 42193 665549
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 42260 662538 42288 670475
rect 41708 662510 42288 662538
rect 41708 662485 41736 662510
rect 42352 661994 42380 689986
rect 41800 661966 42380 661994
rect 41800 661858 41828 661966
rect 41722 661830 41828 661858
rect 41722 661183 41828 661211
rect 41800 661094 41828 661183
rect 41788 661088 41840 661094
rect 41788 661030 41840 661036
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 41788 658708 41840 658714
rect 41788 658650 41840 658656
rect 41800 658186 41828 658650
rect 41722 658158 41828 658186
rect 42260 657642 42288 661966
rect 42444 661094 42472 703938
rect 42536 700874 42564 743990
rect 42628 712298 42656 755414
rect 673472 740382 673500 785674
rect 673644 782332 673696 782338
rect 673644 782274 673696 782280
rect 673460 740376 673512 740382
rect 673460 740318 673512 740324
rect 42616 712292 42668 712298
rect 42616 712234 42668 712240
rect 42524 700868 42576 700874
rect 42524 700810 42576 700816
rect 42432 661088 42484 661094
rect 42432 661030 42484 661036
rect 41892 657614 42288 657642
rect 41892 657506 41920 657614
rect 41722 657478 41920 657506
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 41713 655097 42193 655153
rect 42260 651374 42288 657614
rect 42260 651346 42380 651374
rect 41722 627286 42288 627314
rect 41713 626617 42193 626673
rect 41722 625435 41828 625463
rect 41800 624986 41828 625435
rect 41788 624980 41840 624986
rect 41788 624922 41840 624928
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 622293 42193 622349
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 42260 619426 42288 627286
rect 41800 619398 42288 619426
rect 41800 619290 41828 619398
rect 41722 619262 41828 619290
rect 42352 618746 42380 651346
rect 41800 618718 42380 618746
rect 41800 618655 41828 618718
rect 41722 618627 41828 618655
rect 41788 618520 41840 618526
rect 41788 618462 41840 618468
rect 41800 618011 41828 618462
rect 41722 617983 41828 618011
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41788 615528 41840 615534
rect 41788 615470 41840 615476
rect 41800 614975 41828 615470
rect 41722 614947 41828 614975
rect 42260 614331 42288 618718
rect 42444 618526 42472 661030
rect 42536 658714 42564 700810
rect 42628 690014 42656 712234
rect 673472 695366 673500 740318
rect 673656 738138 673684 782274
rect 673736 781652 673788 781658
rect 673736 781594 673788 781600
rect 673748 740994 673776 781594
rect 673840 775878 673868 864214
rect 673932 863258 673960 870130
rect 673920 863252 673972 863258
rect 673920 863194 673972 863200
rect 674024 782338 674052 872374
rect 674012 782332 674064 782338
rect 674012 782274 674064 782280
rect 673828 775872 673880 775878
rect 673828 775814 673880 775820
rect 673840 767294 673868 775814
rect 673840 767266 673960 767294
rect 673736 740988 673788 740994
rect 673736 740930 673788 740936
rect 673644 738132 673696 738138
rect 673644 738074 673696 738080
rect 673552 730924 673604 730930
rect 673552 730866 673604 730872
rect 673460 695360 673512 695366
rect 673460 695302 673512 695308
rect 42628 689986 42748 690014
rect 42720 668166 42748 689986
rect 42708 668160 42760 668166
rect 42708 668102 42760 668108
rect 42524 658708 42576 658714
rect 42524 658650 42576 658656
rect 42536 651374 42564 658650
rect 42536 651346 42656 651374
rect 42524 624980 42576 624986
rect 42524 624922 42576 624928
rect 42432 618520 42484 618526
rect 42432 618462 42484 618468
rect 41722 614303 42288 614331
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 41713 611897 42193 611953
rect 42260 584202 42288 614303
rect 42260 584174 42380 584202
rect 41722 584075 42288 584103
rect 41713 583417 42193 583473
rect 41788 582684 41840 582690
rect 41788 582626 41840 582632
rect 41800 582263 41828 582626
rect 41722 582235 41828 582263
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 579093 42193 579149
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 42260 576178 42288 584075
rect 41800 576150 42288 576178
rect 41800 576099 41828 576150
rect 41722 576071 41828 576099
rect 42352 575455 42380 584174
rect 41722 575427 42380 575455
rect 41722 574790 41828 574818
rect 41800 574734 41828 574790
rect 41788 574728 41840 574734
rect 41788 574670 41840 574676
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 41722 571747 41828 571775
rect 41800 571266 41828 571747
rect 41788 571260 41840 571266
rect 41788 571202 41840 571208
rect 41722 571118 41920 571146
rect 41892 570738 41920 571118
rect 42260 570738 42288 575427
rect 42444 574734 42472 618462
rect 42536 582690 42564 624922
rect 42628 615534 42656 651346
rect 42720 624986 42748 668102
rect 673472 650554 673500 695302
rect 673564 685234 673592 730866
rect 673656 692322 673684 738074
rect 673736 737044 673788 737050
rect 673736 736986 673788 736992
rect 673748 695978 673776 736986
rect 673932 730930 673960 767266
rect 673920 730924 673972 730930
rect 673920 730866 673972 730872
rect 673736 695972 673788 695978
rect 673736 695914 673788 695920
rect 673656 692306 673960 692322
rect 673656 692300 673972 692306
rect 673656 692294 673920 692300
rect 673920 692242 673972 692248
rect 673736 692096 673788 692102
rect 673736 692038 673788 692044
rect 673552 685228 673604 685234
rect 673552 685170 673604 685176
rect 673460 650548 673512 650554
rect 673460 650490 673512 650496
rect 673472 647222 673500 650490
rect 673460 647216 673512 647222
rect 673460 647158 673512 647164
rect 673460 647080 673512 647086
rect 673460 647022 673512 647028
rect 42708 624980 42760 624986
rect 42708 624922 42760 624928
rect 42616 615528 42668 615534
rect 42616 615470 42668 615476
rect 42628 612734 42656 615470
rect 42628 612706 42748 612734
rect 42524 582684 42576 582690
rect 42524 582626 42576 582632
rect 42432 574728 42484 574734
rect 42432 574670 42484 574676
rect 41892 570710 42288 570738
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 41713 568697 42193 568753
rect 42260 545170 42288 570710
rect 42444 554774 42472 574670
rect 42536 574094 42564 582626
rect 42536 574066 42656 574094
rect 42524 571260 42576 571266
rect 42524 571202 42576 571208
rect 42352 554746 42472 554774
rect 42352 545290 42380 554746
rect 42340 545284 42392 545290
rect 42340 545226 42392 545232
rect 42260 545142 42472 545170
rect 42340 545080 42392 545086
rect 42340 545022 42392 545028
rect 41722 540875 42288 540903
rect 41713 540217 42193 540273
rect 41788 539504 41840 539510
rect 41788 539446 41840 539452
rect 41800 539050 41828 539446
rect 41722 539022 41828 539050
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535893 42193 535949
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 42260 533066 42288 540875
rect 41800 533038 42288 533066
rect 41800 532899 41828 533038
rect 41722 532871 41828 532899
rect 41722 532222 41920 532250
rect 41892 532114 41920 532222
rect 42260 532166 42288 532197
rect 42248 532160 42300 532166
rect 41892 532108 42248 532114
rect 41892 532102 42300 532108
rect 41892 532086 42288 532102
rect 41722 531583 41828 531611
rect 41800 531214 41828 531583
rect 41788 531208 41840 531214
rect 41788 531150 41840 531156
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 41722 528550 41828 528578
rect 41800 528086 41828 528550
rect 41788 528080 41840 528086
rect 41788 528022 41840 528028
rect 41708 527898 41736 527917
rect 42260 527898 42288 532086
rect 42352 531298 42380 545022
rect 42444 532166 42472 545142
rect 42432 532160 42484 532166
rect 42432 532102 42484 532108
rect 42352 531270 42472 531298
rect 42444 531214 42472 531270
rect 42432 531208 42484 531214
rect 42432 531150 42484 531156
rect 41708 527870 42288 527898
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 41713 525497 42193 525553
rect 42260 419534 42288 527870
rect 42260 419506 42380 419534
rect 41722 413275 42288 413303
rect 41713 412617 42193 412673
rect 41722 411454 41828 411482
rect 41800 410990 41828 411454
rect 41788 410984 41840 410990
rect 41788 410926 41840 410932
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 408293 42193 408349
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 42260 405498 42288 413275
rect 41800 405470 42288 405498
rect 41800 405299 41828 405470
rect 41722 405271 41828 405299
rect 42352 405226 42380 419506
rect 41800 405198 42380 405226
rect 41800 404682 41828 405198
rect 41722 404654 41828 404682
rect 41788 404524 41840 404530
rect 41788 404466 41840 404472
rect 41800 404002 41828 404466
rect 41722 403974 41828 404002
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41722 400947 41828 400975
rect 41800 400858 41828 400947
rect 41788 400852 41840 400858
rect 41788 400794 41840 400800
rect 42352 400330 42380 405198
rect 42444 404530 42472 531150
rect 42536 528086 42564 571202
rect 42628 539510 42656 574066
rect 42720 571266 42748 612706
rect 673472 602954 673500 647022
rect 673564 640694 673592 685170
rect 673748 651166 673776 692038
rect 673736 651160 673788 651166
rect 673736 651102 673788 651108
rect 673644 647216 673696 647222
rect 673644 647158 673696 647164
rect 673552 640688 673604 640694
rect 673552 640630 673604 640636
rect 673460 602948 673512 602954
rect 673460 602890 673512 602896
rect 42708 571260 42760 571266
rect 42708 571202 42760 571208
rect 673472 557870 673500 602890
rect 673564 595066 673592 640630
rect 673656 605130 673684 647158
rect 673748 646474 673776 651102
rect 673932 647086 673960 692242
rect 673920 647080 673972 647086
rect 673920 647022 673972 647028
rect 673736 646468 673788 646474
rect 673736 646410 673788 646416
rect 673748 605810 673776 646410
rect 673736 605804 673788 605810
rect 673736 605746 673788 605752
rect 673644 605124 673696 605130
rect 673644 605066 673696 605072
rect 673552 595060 673604 595066
rect 673552 595002 673604 595008
rect 673460 557864 673512 557870
rect 673460 557806 673512 557812
rect 673564 550526 673592 595002
rect 673656 560998 673684 605066
rect 673736 601860 673788 601866
rect 673736 601802 673788 601808
rect 673748 561270 673776 601802
rect 673736 561264 673788 561270
rect 673736 561206 673788 561212
rect 673644 560992 673696 560998
rect 673644 560934 673696 560940
rect 673552 550520 673604 550526
rect 673552 550462 673604 550468
rect 673564 546494 673592 550462
rect 673472 546466 673592 546494
rect 42616 539504 42668 539510
rect 42616 539446 42668 539452
rect 42524 528080 42576 528086
rect 42524 528022 42576 528028
rect 42628 419534 42656 539446
rect 42708 528080 42760 528086
rect 42708 528022 42760 528028
rect 42536 419506 42656 419534
rect 42536 410990 42564 419506
rect 42524 410984 42576 410990
rect 42524 410926 42576 410932
rect 42432 404524 42484 404530
rect 42432 404466 42484 404472
rect 41722 400302 42380 400330
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 41713 397897 42193 397953
rect 42352 380894 42380 400302
rect 42352 380866 42472 380894
rect 41722 370075 42288 370103
rect 41713 369417 42193 369473
rect 41788 368688 41840 368694
rect 41788 368630 41840 368636
rect 41800 368263 41828 368630
rect 41722 368235 41828 368263
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 365093 42193 365149
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 42260 362250 42288 370075
rect 42340 368688 42392 368694
rect 42340 368630 42392 368636
rect 41892 362222 42288 362250
rect 41892 362114 41920 362222
rect 42352 362114 42380 368630
rect 41722 362086 41920 362114
rect 42260 362086 42380 362114
rect 41722 361406 41828 361434
rect 41800 361350 41828 361406
rect 41788 361344 41840 361350
rect 41788 361286 41840 361292
rect 41722 360783 41828 360811
rect 41800 360738 41828 360783
rect 41788 360732 41840 360738
rect 41788 360674 41840 360680
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41722 357734 41828 357762
rect 41800 357270 41828 357734
rect 41788 357264 41840 357270
rect 41788 357206 41840 357212
rect 41722 357103 41828 357131
rect 41800 356726 41828 357103
rect 41788 356720 41840 356726
rect 41788 356662 41840 356668
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 41713 354697 42193 354753
rect 42260 330070 42288 362086
rect 42444 361574 42472 380866
rect 42536 368694 42564 410926
rect 42616 404524 42668 404530
rect 42616 404466 42668 404472
rect 42524 368688 42576 368694
rect 42524 368630 42576 368636
rect 42352 361546 42472 361574
rect 42352 361350 42380 361546
rect 42340 361344 42392 361350
rect 42340 361286 42392 361292
rect 42352 356726 42380 361286
rect 42628 360738 42656 404466
rect 42720 400858 42748 528022
rect 42708 400852 42760 400858
rect 42708 400794 42760 400800
rect 42616 360732 42668 360738
rect 42616 360674 42668 360680
rect 42524 357264 42576 357270
rect 42524 357206 42576 357212
rect 42340 356720 42392 356726
rect 42340 356662 42392 356668
rect 42248 330064 42300 330070
rect 42248 330006 42300 330012
rect 41722 326862 41828 326890
rect 41800 326754 41828 326862
rect 41800 326726 42288 326754
rect 41713 326217 42193 326273
rect 41788 325508 41840 325514
rect 41788 325450 41840 325456
rect 41800 325063 41828 325450
rect 41722 325035 41828 325063
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321893 42193 321949
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 42260 318899 42288 326726
rect 41722 318871 42288 318899
rect 42352 318255 42380 356662
rect 42432 330064 42484 330070
rect 42432 330006 42484 330012
rect 42444 325514 42472 330006
rect 42432 325508 42484 325514
rect 42432 325450 42484 325456
rect 41722 318227 42380 318255
rect 41722 317583 41828 317611
rect 41800 317218 41828 317583
rect 41788 317212 41840 317218
rect 41788 317154 41840 317160
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 41722 314547 41828 314575
rect 41800 314090 41828 314547
rect 41788 314084 41840 314090
rect 41788 314026 41840 314032
rect 41722 313903 41828 313931
rect 41800 313834 41828 313903
rect 42260 313834 42288 318227
rect 42536 314090 42564 357206
rect 42628 317218 42656 360674
rect 42720 357270 42748 400794
rect 673472 372366 673500 546466
rect 674760 427854 674788 996338
rect 675407 878047 675887 878103
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675392 875832 675444 875838
rect 675392 875774 675444 875780
rect 675404 875697 675432 875774
rect 675312 875683 675432 875697
rect 675312 875669 675418 875683
rect 675312 871373 675340 875669
rect 675404 874546 675432 875039
rect 675392 874540 675444 874546
rect 675392 874482 675444 874488
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675392 872432 675444 872438
rect 675392 872374 675444 872380
rect 675404 872003 675432 872374
rect 675312 871350 675418 871373
rect 675300 871345 675418 871350
rect 675300 871344 675352 871345
rect 675300 871286 675352 871292
rect 675404 870194 675432 870740
rect 675392 870188 675444 870194
rect 675392 870130 675444 870136
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867651 675887 867707
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675404 864278 675432 864551
rect 675392 864272 675444 864278
rect 675392 864214 675444 864220
rect 675407 863327 675887 863383
rect 675392 863252 675444 863258
rect 675392 863194 675444 863200
rect 675404 862716 675432 863194
rect 677598 818408 677654 818417
rect 675300 818372 675352 818378
rect 677598 818343 677600 818352
rect 675300 818314 675352 818320
rect 677652 818343 677654 818352
rect 677600 818314 677652 818320
rect 675312 786614 675340 818314
rect 675407 788847 675887 788903
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 675128 786586 675340 786614
rect 675128 728906 675156 786586
rect 675404 786010 675432 786483
rect 675208 786004 675260 786010
rect 675208 785946 675260 785952
rect 675392 786004 675444 786010
rect 675392 785946 675444 785952
rect 675220 781658 675248 785946
rect 675404 785738 675432 785839
rect 675392 785732 675444 785738
rect 675392 785674 675444 785680
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675404 782338 675432 782803
rect 675392 782332 675444 782338
rect 675392 782274 675444 782280
rect 675404 781658 675432 782159
rect 675208 781652 675260 781658
rect 675208 781594 675260 781600
rect 675392 781652 675444 781658
rect 675392 781594 675444 781600
rect 675404 781046 675432 781524
rect 675208 781040 675260 781046
rect 675208 780982 675260 780988
rect 675392 781040 675444 781046
rect 675392 780982 675444 780988
rect 675220 773514 675248 780982
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 778451 675887 778507
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675392 775872 675444 775878
rect 675392 775814 675444 775820
rect 675404 775351 675432 775814
rect 675407 774127 675887 774183
rect 675220 773486 675418 773514
rect 675407 743847 675887 743903
rect 675407 743295 675887 743351
rect 675407 742651 675887 742707
rect 675407 742007 675887 742063
rect 675404 740994 675432 741483
rect 675208 740988 675260 740994
rect 675208 740930 675260 740936
rect 675392 740988 675444 740994
rect 675392 740930 675444 740936
rect 675220 737050 675248 740930
rect 675404 740382 675432 740860
rect 675392 740376 675444 740382
rect 675392 740318 675444 740324
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675392 738132 675444 738138
rect 675392 738074 675444 738080
rect 675404 737803 675432 738074
rect 675404 737050 675432 737159
rect 675208 737044 675260 737050
rect 675208 736986 675260 736992
rect 675392 737044 675444 737050
rect 675392 736986 675444 736992
rect 675312 736494 675418 736522
rect 675312 729042 675340 736494
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 733451 675887 733507
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675392 730924 675444 730930
rect 675392 730866 675444 730872
rect 675404 730351 675432 730866
rect 675407 729127 675887 729183
rect 675312 729014 675432 729042
rect 675128 728878 675340 728906
rect 675312 701054 675340 728878
rect 675404 728484 675432 729014
rect 675128 701026 675340 701054
rect 675128 681734 675156 701026
rect 675407 698847 675887 698903
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675404 695978 675432 696483
rect 675208 695972 675260 695978
rect 675208 695914 675260 695920
rect 675392 695972 675444 695978
rect 675392 695914 675444 695920
rect 675220 692102 675248 695914
rect 675404 695366 675432 695844
rect 675392 695360 675444 695366
rect 675392 695302 675444 695308
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675404 692306 675432 692803
rect 675392 692300 675444 692306
rect 675392 692242 675444 692248
rect 675404 692102 675432 692172
rect 675208 692096 675260 692102
rect 675208 692038 675260 692044
rect 675392 692096 675444 692102
rect 675392 692038 675444 692044
rect 675312 691614 675432 691642
rect 675312 683525 675340 691614
rect 675404 691492 675432 691614
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 688451 675887 688507
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675404 685234 675432 685372
rect 675392 685228 675444 685234
rect 675392 685170 675444 685176
rect 675407 684127 675887 684183
rect 675312 683497 675418 683525
rect 675128 681706 675340 681734
rect 675312 651374 675340 681706
rect 675407 653647 675887 653703
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 675128 651346 675340 651374
rect 675128 632054 675156 651346
rect 675404 651166 675432 651283
rect 675392 651160 675444 651166
rect 675392 651102 675444 651108
rect 675404 650554 675432 650639
rect 675392 650548 675444 650554
rect 675392 650490 675444 650496
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675404 647086 675432 647603
rect 675392 647080 675444 647086
rect 675392 647022 675444 647028
rect 675404 646474 675432 646959
rect 675392 646468 675444 646474
rect 675392 646410 675444 646416
rect 675404 645794 675432 646340
rect 675208 645788 675260 645794
rect 675208 645730 675260 645736
rect 675392 645788 675444 645794
rect 675392 645730 675444 645736
rect 675220 638330 675248 645730
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 643251 675887 643307
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675392 640688 675444 640694
rect 675392 640630 675444 640636
rect 675404 640151 675432 640630
rect 675407 638927 675887 638983
rect 675220 638302 675418 638330
rect 675128 632026 675340 632054
rect 675312 612734 675340 632026
rect 675128 612706 675340 612734
rect 675128 593722 675156 612706
rect 675407 608647 675887 608703
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 675404 605810 675432 606283
rect 675208 605804 675260 605810
rect 675208 605746 675260 605752
rect 675392 605804 675444 605810
rect 675392 605746 675444 605752
rect 675220 601866 675248 605746
rect 675404 605130 675432 605639
rect 675392 605124 675444 605130
rect 675392 605066 675444 605072
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675392 602948 675444 602954
rect 675392 602890 675444 602896
rect 675404 602603 675432 602890
rect 675404 601866 675432 601959
rect 675208 601860 675260 601866
rect 675208 601802 675260 601808
rect 675392 601860 675444 601866
rect 675392 601802 675444 601808
rect 675312 601310 675418 601338
rect 675312 593858 675340 601310
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 598251 675887 598307
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675404 595066 675432 595151
rect 675392 595060 675444 595066
rect 675392 595002 675444 595008
rect 675407 593927 675887 593983
rect 675312 593830 675432 593858
rect 675128 593694 675340 593722
rect 675312 574094 675340 593694
rect 675404 593300 675432 593830
rect 675128 574066 675340 574094
rect 675128 546494 675156 574066
rect 675407 563447 675887 563503
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 675208 561264 675260 561270
rect 675208 561206 675260 561212
rect 675392 561264 675444 561270
rect 675392 561206 675444 561212
rect 675220 557326 675248 561206
rect 675404 561068 675432 561206
rect 675392 560992 675444 560998
rect 675392 560934 675444 560940
rect 675404 560439 675432 560934
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675392 557864 675444 557870
rect 675392 557806 675444 557812
rect 675404 557396 675432 557806
rect 675208 557320 675260 557326
rect 675208 557262 675260 557268
rect 675392 557320 675444 557326
rect 675392 557262 675444 557268
rect 675404 556759 675432 557262
rect 675404 555626 675432 556115
rect 675208 555620 675260 555626
rect 675208 555562 675260 555568
rect 675392 555620 675444 555626
rect 675392 555562 675444 555568
rect 675220 548125 675248 555562
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 553051 675887 553107
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675392 550520 675444 550526
rect 675392 550462 675444 550468
rect 675404 549951 675432 550462
rect 675407 548727 675887 548783
rect 675220 548097 675418 548125
rect 675128 546466 675340 546494
rect 675312 513806 675340 546466
rect 675300 513800 675352 513806
rect 677692 513800 677744 513806
rect 675300 513742 675352 513748
rect 677690 513768 677692 513777
rect 677744 513768 677746 513777
rect 677690 513703 677746 513712
rect 674748 427848 674800 427854
rect 674748 427790 674800 427796
rect 677508 427848 677560 427854
rect 677508 427790 677560 427796
rect 677520 425649 677548 427790
rect 677506 425640 677562 425649
rect 677506 425575 677562 425584
rect 675407 386247 675887 386303
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 675312 383982 675432 384010
rect 673552 382764 673604 382770
rect 673552 382706 673604 382712
rect 673460 372360 673512 372366
rect 673460 372302 673512 372308
rect 42708 357264 42760 357270
rect 42708 357206 42760 357212
rect 673472 328098 673500 372302
rect 673564 337550 673592 382706
rect 673736 379704 673788 379710
rect 673736 379646 673788 379652
rect 673644 379092 673696 379098
rect 673644 379034 673696 379040
rect 673552 337544 673604 337550
rect 673552 337486 673604 337492
rect 673460 328092 673512 328098
rect 673460 328034 673512 328040
rect 42800 325508 42852 325514
rect 42800 325450 42852 325456
rect 42616 317212 42668 317218
rect 42616 317154 42668 317160
rect 42524 314084 42576 314090
rect 42524 314026 42576 314032
rect 41800 313806 42288 313834
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 41713 311497 42193 311553
rect 42260 303614 42288 313806
rect 42260 303586 42380 303614
rect 41722 283675 42288 283703
rect 41713 283017 42193 283073
rect 41722 281846 41828 281874
rect 41800 281382 41828 281846
rect 41788 281376 41840 281382
rect 41788 281318 41840 281324
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278693 42193 278749
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 42260 275699 42288 283675
rect 41722 275671 42288 275699
rect 42352 275210 42380 303586
rect 42432 281376 42484 281382
rect 42432 281318 42484 281324
rect 41800 275182 42380 275210
rect 41800 275074 41828 275182
rect 41722 275046 41828 275074
rect 41788 274576 41840 274582
rect 41788 274518 41840 274524
rect 41800 274394 41828 274518
rect 41722 274366 41828 274394
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 41788 271924 41840 271930
rect 41788 271866 41840 271872
rect 41800 271402 41828 271866
rect 41722 271374 41828 271402
rect 42260 270858 42288 275182
rect 41892 270830 42288 270858
rect 41892 270722 41920 270830
rect 41722 270694 41920 270722
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 41713 268297 42193 268353
rect 42260 264974 42288 270830
rect 42260 264946 42380 264974
rect 41722 240502 42288 240530
rect 41713 239817 42193 239873
rect 41722 238635 41828 238663
rect 41800 238134 41828 238635
rect 41788 238128 41840 238134
rect 41788 238070 41840 238076
rect 41713 237977 42193 238033
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 42260 232642 42288 240502
rect 41800 232614 42288 232642
rect 41800 232506 41828 232614
rect 41722 232478 41828 232506
rect 42352 231855 42380 264946
rect 42444 238134 42472 281318
rect 42628 274582 42656 317154
rect 42708 314084 42760 314090
rect 42708 314026 42760 314032
rect 42616 274576 42668 274582
rect 42536 274524 42616 274530
rect 42536 274518 42668 274524
rect 42536 274502 42656 274518
rect 42432 238128 42484 238134
rect 42432 238070 42484 238076
rect 41722 231827 42380 231855
rect 41788 231736 41840 231742
rect 41788 231678 41840 231684
rect 41800 231211 41828 231678
rect 41722 231183 41828 231211
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 41788 228676 41840 228682
rect 41788 228618 41840 228624
rect 41800 228154 41828 228618
rect 41722 228126 41828 228154
rect 42260 227610 42288 231827
rect 41800 227582 42380 227610
rect 41800 227531 41828 227582
rect 41722 227503 41828 227531
rect 42248 227520 42300 227526
rect 42248 227462 42300 227468
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 41713 225097 42193 225153
rect 42260 197418 42288 227462
rect 42352 197554 42380 227582
rect 42444 226334 42472 238070
rect 42536 231742 42564 274502
rect 42720 271930 42748 314026
rect 42812 281382 42840 325450
rect 673472 282130 673500 328034
rect 673564 293622 673592 337486
rect 673656 334286 673684 379034
rect 673748 342254 673776 379646
rect 675312 379573 675340 383982
rect 675404 383860 675432 383982
rect 675404 382770 675432 383239
rect 675392 382764 675444 382770
rect 675392 382706 675444 382712
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675404 379710 675432 380188
rect 675392 379704 675444 379710
rect 675392 379646 675444 379652
rect 675312 379559 675418 379573
rect 675312 379545 675432 379559
rect 675404 379098 675432 379545
rect 675392 379092 675444 379098
rect 675392 379034 675444 379040
rect 675312 378901 675418 378929
rect 675312 370925 675340 378901
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675404 372366 675432 372751
rect 675392 372360 675444 372366
rect 675392 372302 675444 372308
rect 675407 371527 675887 371583
rect 675312 370897 675418 370925
rect 673748 342226 673960 342254
rect 673932 334490 673960 342226
rect 675407 341047 675887 341103
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675404 338178 675432 338708
rect 675312 338150 675432 338178
rect 673920 334484 673972 334490
rect 673920 334426 673972 334432
rect 673644 334280 673696 334286
rect 673644 334222 673696 334228
rect 673656 293826 673684 334222
rect 673644 293820 673696 293826
rect 673644 293762 673696 293768
rect 673552 293616 673604 293622
rect 673552 293558 673604 293564
rect 673460 282124 673512 282130
rect 673460 282066 673512 282072
rect 42800 281376 42852 281382
rect 42800 281318 42852 281324
rect 42708 271924 42760 271930
rect 42708 271866 42760 271872
rect 42720 245654 42748 271866
rect 673564 248606 673592 293558
rect 673656 249150 673684 293762
rect 673932 289882 673960 334426
rect 675312 334370 675340 338150
rect 675404 337550 675432 338028
rect 675392 337544 675444 337550
rect 675392 337486 675444 337492
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675404 334490 675432 335003
rect 675392 334484 675444 334490
rect 675392 334426 675444 334432
rect 675312 334356 675418 334370
rect 675312 334342 675432 334356
rect 675404 334286 675432 334342
rect 675392 334280 675444 334286
rect 675392 334222 675444 334228
rect 675312 333701 675418 333729
rect 675312 325725 675340 333701
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675392 328092 675444 328098
rect 675392 328034 675444 328040
rect 675404 327556 675432 328034
rect 675407 326327 675887 326383
rect 675312 325697 675418 325725
rect 675407 296047 675887 296103
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 675392 293820 675444 293826
rect 675392 293762 675444 293768
rect 675404 293706 675432 293762
rect 675312 293692 675432 293706
rect 675312 293678 675418 293692
rect 673920 289876 673972 289882
rect 673920 289818 673972 289824
rect 673736 282124 673788 282130
rect 673736 282066 673788 282072
rect 673748 264974 673776 282066
rect 673748 264946 673868 264974
rect 673644 249144 673696 249150
rect 673644 249086 673696 249092
rect 673552 248600 673604 248606
rect 673552 248542 673604 248548
rect 42628 245626 42748 245654
rect 42524 231736 42576 231742
rect 42524 231678 42576 231684
rect 42536 227526 42564 231678
rect 42628 228682 42656 245626
rect 42616 228676 42668 228682
rect 42616 228618 42668 228624
rect 42524 227520 42576 227526
rect 42524 227462 42576 227468
rect 42444 226306 42564 226334
rect 42352 197526 42472 197554
rect 42260 197390 42380 197418
rect 41722 197254 42288 197282
rect 41713 196617 42193 196673
rect 41788 195900 41840 195906
rect 41788 195842 41840 195848
rect 41800 195463 41828 195842
rect 41722 195435 41828 195463
rect 41713 194777 42193 194833
rect 41713 192937 42193 192993
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 42260 189394 42288 197254
rect 41892 189366 42288 189394
rect 41892 189299 41920 189366
rect 41722 189271 41920 189299
rect 41788 189168 41840 189174
rect 41788 189110 41840 189116
rect 41800 188655 41828 189110
rect 41722 188627 41828 188655
rect 42352 188170 42380 197390
rect 42444 189174 42472 197526
rect 42536 195906 42564 226306
rect 42524 195900 42576 195906
rect 42524 195842 42576 195848
rect 42432 189168 42484 189174
rect 42432 189110 42484 189116
rect 41892 188142 42380 188170
rect 41892 188034 41920 188142
rect 41722 188006 41920 188034
rect 41984 187610 42012 188142
rect 42444 188034 42472 189110
rect 42260 188006 42472 188034
rect 41972 187604 42024 187610
rect 41972 187546 42024 187552
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 41722 184947 41828 184975
rect 41800 184482 41828 184947
rect 41788 184476 41840 184482
rect 41788 184418 41840 184424
rect 42260 184331 42288 188006
rect 42536 187694 42564 195842
rect 42444 187666 42564 187694
rect 41722 184303 42380 184331
rect 42248 184204 42300 184210
rect 42248 184146 42300 184152
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 41713 181897 42193 181953
rect 42260 45694 42288 184146
rect 42248 45688 42300 45694
rect 42248 45630 42300 45636
rect 42352 45626 42380 184303
rect 42444 82890 42472 187666
rect 42524 187604 42576 187610
rect 42524 187546 42576 187552
rect 42536 121514 42564 187546
rect 42628 184482 42656 228618
rect 673564 202366 673592 248542
rect 673644 244044 673696 244050
rect 673644 243986 673696 243992
rect 673552 202360 673604 202366
rect 673552 202302 673604 202308
rect 42616 184476 42668 184482
rect 42616 184418 42668 184424
rect 673564 158370 673592 202302
rect 673656 199306 673684 243986
rect 673840 243930 673868 264946
rect 673932 244934 673960 289818
rect 675312 289762 675340 293678
rect 675392 293616 675444 293622
rect 675392 293558 675444 293564
rect 675404 293012 675432 293558
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675404 289882 675432 290020
rect 675392 289876 675444 289882
rect 675392 289818 675444 289824
rect 675312 289734 675432 289762
rect 675404 289340 675432 289734
rect 675312 288701 675418 288729
rect 675312 280725 675340 288701
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 675404 282130 675432 282540
rect 675392 282124 675444 282130
rect 675392 282066 675444 282072
rect 675407 281327 675887 281383
rect 675312 280697 675418 280725
rect 675407 251047 675887 251103
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675392 249144 675444 249150
rect 675392 249086 675444 249092
rect 675404 248690 675432 249086
rect 675312 248676 675432 248690
rect 675312 248662 675418 248676
rect 673920 244928 673972 244934
rect 673920 244870 673972 244876
rect 673932 244050 673960 244870
rect 675312 244373 675340 248662
rect 675392 248600 675444 248606
rect 675392 248542 675444 248548
rect 675404 248039 675432 248542
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675404 244934 675432 245004
rect 675392 244928 675444 244934
rect 675392 244870 675444 244876
rect 675312 244359 675418 244373
rect 675312 244345 675432 244359
rect 673920 244044 673972 244050
rect 673920 243986 673972 243992
rect 673840 243902 673960 243930
rect 673828 243840 673880 243846
rect 673828 243782 673880 243788
rect 673840 203522 673868 243782
rect 673932 237726 673960 243902
rect 675404 243846 675432 244345
rect 675392 243840 675444 243846
rect 675392 243782 675444 243788
rect 675312 243701 675418 243729
rect 673920 237720 673972 237726
rect 673920 237662 673972 237668
rect 673828 203516 673880 203522
rect 673828 203458 673880 203464
rect 673644 199300 673696 199306
rect 673644 199242 673696 199248
rect 673552 158364 673604 158370
rect 673552 158306 673604 158312
rect 673564 158250 673592 158306
rect 673472 158222 673592 158250
rect 42524 121508 42576 121514
rect 42524 121450 42576 121456
rect 44180 121508 44232 121514
rect 44180 121450 44232 121456
rect 44192 110537 44220 121450
rect 673472 113218 673500 158222
rect 673656 155242 673684 199242
rect 673736 199096 673788 199102
rect 673736 199038 673788 199044
rect 673748 158642 673776 199038
rect 673932 191962 673960 237662
rect 675312 235725 675340 243701
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 675407 238167 675887 238223
rect 675392 237720 675444 237726
rect 675392 237662 675444 237668
rect 675404 237524 675432 237662
rect 675407 236327 675887 236383
rect 675312 235697 675418 235725
rect 675407 205847 675887 205903
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 675312 203522 675340 203580
rect 675300 203516 675352 203522
rect 675352 203469 675418 203497
rect 675300 203458 675352 203464
rect 675312 199186 675340 203458
rect 675404 202366 675432 202844
rect 675392 202360 675444 202366
rect 675392 202302 675444 202308
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675404 199306 675432 199803
rect 675392 199300 675444 199306
rect 675392 199242 675444 199248
rect 675312 199172 675418 199186
rect 675312 199158 675432 199172
rect 675404 199102 675432 199158
rect 675392 199096 675444 199102
rect 675392 199038 675444 199044
rect 675312 198614 675432 198642
rect 673920 191956 673972 191962
rect 673920 191898 673972 191904
rect 673736 158636 673788 158642
rect 673736 158578 673788 158584
rect 673644 155236 673696 155242
rect 673644 155178 673696 155184
rect 673656 149054 673684 155178
rect 673736 154148 673788 154154
rect 673736 154090 673788 154096
rect 673564 149026 673684 149054
rect 673460 113212 673512 113218
rect 673460 113154 673512 113160
rect 44178 110528 44234 110537
rect 44178 110463 44234 110472
rect 44822 110528 44878 110537
rect 44822 110463 44878 110472
rect 44836 110414 44864 110463
rect 44836 110386 44956 110414
rect 42432 82884 42484 82890
rect 42432 82826 42484 82832
rect 44180 82884 44232 82890
rect 44180 82826 44232 82832
rect 44192 71913 44220 82826
rect 44178 71904 44234 71913
rect 44178 71839 44234 71848
rect 44822 71904 44878 71913
rect 44822 71839 44878 71848
rect 44836 46986 44864 71839
rect 44824 46980 44876 46986
rect 44824 46922 44876 46928
rect 42340 45620 42392 45626
rect 42340 45562 42392 45568
rect 44928 45558 44956 110386
rect 143540 46912 143592 46918
rect 200856 46912 200908 46918
rect 143540 46854 143592 46860
rect 151726 46880 151782 46889
rect 140964 45688 141016 45694
rect 140964 45630 141016 45636
rect 44916 45552 44968 45558
rect 44916 45494 44968 45500
rect 93768 41540 93820 41546
rect 93768 41482 93820 41488
rect 93780 40225 93808 41482
rect 135168 40248 135220 40254
rect 93766 40216 93822 40225
rect 93766 40151 93822 40160
rect 135166 40216 135168 40225
rect 135220 40216 135222 40225
rect 140976 40202 141004 45630
rect 143552 40497 143580 46854
rect 151726 46815 151782 46824
rect 188526 46880 188582 46889
rect 200856 46854 200908 46860
rect 256240 46912 256292 46918
rect 256240 46854 256292 46860
rect 297732 46912 297784 46918
rect 297732 46854 297784 46860
rect 309416 46912 309468 46918
rect 309416 46854 309468 46860
rect 352564 46912 352616 46918
rect 352564 46854 352616 46860
rect 364248 46912 364300 46918
rect 364248 46854 364300 46860
rect 407396 46912 407448 46918
rect 407396 46854 407448 46860
rect 419080 46912 419132 46918
rect 419080 46854 419132 46860
rect 462136 46912 462188 46918
rect 462136 46854 462188 46860
rect 473820 46912 473872 46918
rect 473820 46854 473872 46860
rect 516968 46912 517020 46918
rect 516968 46854 517020 46860
rect 527456 46912 527508 46918
rect 527456 46854 527508 46860
rect 188526 46815 188582 46824
rect 143632 45620 143684 45626
rect 143632 45562 143684 45568
rect 143644 44198 143672 45562
rect 143632 44192 143684 44198
rect 143632 44134 143684 44140
rect 145104 44192 145156 44198
rect 145104 44134 145156 44140
rect 143538 40488 143594 40497
rect 143538 40423 143594 40432
rect 143540 40248 143592 40254
rect 143078 40216 143134 40225
rect 140976 40174 141036 40202
rect 135166 40151 135222 40160
rect 141008 40118 141036 40174
rect 143078 40151 143134 40160
rect 143538 40216 143540 40225
rect 143592 40216 143594 40225
rect 145116 40202 145144 44134
rect 146300 41880 146352 41886
rect 146300 41822 146352 41828
rect 143538 40151 143594 40160
rect 145103 40174 145144 40202
rect 143084 40118 143112 40151
rect 140996 40112 141048 40118
rect 140996 40054 141048 40060
rect 143072 40112 143124 40118
rect 143072 40054 143124 40060
rect 144552 40112 144604 40118
rect 144552 40054 144604 40060
rect 141008 39984 141036 40054
rect 143084 39916 143112 40054
rect 144564 39916 144592 40054
rect 145103 40000 145131 40174
rect 146312 40118 146340 41822
rect 151740 40497 151768 46815
rect 186688 45620 186740 45626
rect 186688 45562 186740 45568
rect 186700 41820 186728 45562
rect 188540 44402 188568 46815
rect 194692 45620 194744 45626
rect 194692 45562 194744 45568
rect 188528 44396 188580 44402
rect 188528 44338 188580 44344
rect 192852 44396 192904 44402
rect 192852 44338 192904 44344
rect 187327 41713 187383 42193
rect 188540 41820 188568 44338
rect 189264 41948 189316 41954
rect 189264 41890 189316 41896
rect 191104 41948 191156 41954
rect 191104 41890 191156 41896
rect 192300 41948 192352 41954
rect 192300 41890 192352 41896
rect 189276 41834 189304 41890
rect 191116 41834 191144 41890
rect 192312 41834 192340 41890
rect 189198 41806 189304 41834
rect 191038 41806 191144 41834
rect 192234 41806 192340 41834
rect 192864 41820 192892 44338
rect 193588 41948 193640 41954
rect 193588 41890 193640 41896
rect 193600 41834 193628 41890
rect 193522 41806 193628 41834
rect 194043 41713 194099 42193
rect 194704 41820 194732 45562
rect 195980 45552 196032 45558
rect 195980 45494 196032 45500
rect 195992 44334 196020 45494
rect 195980 44328 196032 44334
rect 195980 44270 196032 44276
rect 195336 44192 195388 44198
rect 195336 44134 195388 44140
rect 195348 41820 195376 44134
rect 195992 41820 196020 44270
rect 199844 44260 199896 44266
rect 199844 44202 199896 44208
rect 199660 44192 199712 44198
rect 199856 44146 199884 44202
rect 199712 44140 199884 44146
rect 199660 44134 199884 44140
rect 199672 44118 199884 44134
rect 196440 41948 196492 41954
rect 196440 41890 196492 41896
rect 198464 41948 198516 41954
rect 198464 41890 198516 41896
rect 196452 41834 196480 41890
rect 198476 41834 198504 41890
rect 196452 41806 198504 41834
rect 198936 41818 199042 41834
rect 199672 41820 199700 44118
rect 200120 41948 200172 41954
rect 200120 41890 200172 41896
rect 200132 41834 200160 41890
rect 200868 41834 200896 46854
rect 201500 44328 201552 44334
rect 201500 44270 201552 44276
rect 200132 41820 200896 41834
rect 201512 41820 201540 44270
rect 198924 41812 199042 41818
rect 198976 41806 199042 41812
rect 200132 41806 200882 41820
rect 198924 41754 198976 41760
rect 151726 40488 151782 40497
rect 151726 40423 151782 40432
rect 146300 40112 146352 40118
rect 146300 40054 146352 40060
rect 145091 39706 145143 40000
rect 256252 39545 256280 46854
rect 297088 44396 297140 44402
rect 297088 44338 297140 44344
rect 295248 44328 295300 44334
rect 295248 44270 295300 44276
rect 295260 41834 295288 44270
rect 297100 41834 297128 44338
rect 297744 41834 297772 46854
rect 299572 44396 299624 44402
rect 299572 44338 299624 44344
rect 305736 44396 305788 44402
rect 305736 44338 305788 44344
rect 297916 41948 297968 41954
rect 297916 41890 297968 41896
rect 297928 41834 297956 41890
rect 295260 41806 295311 41834
rect 297100 41806 297151 41834
rect 297744 41806 297956 41834
rect 299584 41834 299612 44338
rect 303252 44328 303304 44334
rect 303252 44270 303304 44276
rect 300676 41948 300728 41954
rect 300676 41890 300728 41896
rect 302240 41948 302292 41954
rect 302240 41890 302292 41896
rect 300688 41834 300716 41890
rect 302252 41834 302280 41890
rect 299584 41806 299635 41834
rect 300688 41806 302280 41834
rect 302643 41713 302699 42193
rect 303264 41834 303292 44270
rect 303896 44260 303948 44266
rect 303896 44202 303948 44208
rect 303908 41834 303936 44202
rect 304540 44192 304592 44198
rect 304540 44134 304592 44140
rect 304552 41834 304580 44134
rect 305276 41948 305328 41954
rect 305276 41890 305328 41896
rect 305288 41834 305316 41890
rect 303264 41806 303315 41834
rect 303908 41806 303959 41834
rect 304552 41806 304603 41834
rect 305155 41806 305316 41834
rect 305748 41834 305776 44338
rect 308220 44260 308272 44266
rect 308220 44202 308272 44208
rect 306564 41948 306616 41954
rect 306564 41890 306616 41896
rect 306576 41834 306604 41890
rect 305748 41806 305799 41834
rect 306443 41806 306604 41834
rect 306967 41713 307023 42193
rect 308232 41834 308260 44202
rect 308680 41948 308732 41954
rect 308680 41890 308732 41896
rect 308692 41834 308720 41890
rect 309428 41834 309456 46854
rect 349988 44464 350040 44470
rect 349988 44406 350040 44412
rect 350000 44198 350028 44406
rect 351920 44328 351972 44334
rect 351920 44270 351972 44276
rect 349988 44192 350040 44198
rect 349988 44134 350040 44140
rect 350080 44192 350132 44198
rect 350080 44134 350132 44140
rect 307639 41818 307800 41834
rect 307639 41812 307812 41818
rect 307639 41806 307760 41812
rect 308232 41806 308283 41834
rect 308692 41806 309479 41834
rect 307760 41754 307812 41760
rect 310095 41713 310151 42193
rect 350092 41820 350120 44134
rect 351932 41820 351960 44270
rect 352576 41970 352604 46854
rect 359372 44464 359424 44470
rect 359372 44406 359424 44412
rect 354404 44328 354456 44334
rect 354404 44270 354456 44276
rect 352576 41954 352696 41970
rect 352576 41948 352708 41954
rect 352576 41942 352656 41948
rect 352576 41820 352604 41942
rect 352656 41890 352708 41896
rect 354416 41820 354444 44270
rect 358728 44260 358780 44266
rect 358728 44202 358780 44208
rect 358084 44192 358136 44198
rect 358084 44134 358136 44140
rect 355508 41948 355560 41954
rect 355508 41890 355560 41896
rect 356980 41948 357032 41954
rect 356980 41890 357032 41896
rect 355520 41834 355548 41890
rect 356992 41834 357020 41890
rect 355520 41806 357020 41834
rect 357443 41713 357499 42193
rect 358096 41820 358124 44134
rect 358740 41820 358768 44202
rect 359384 41820 359412 44406
rect 360568 44328 360620 44334
rect 360568 44270 360620 44276
rect 363052 44328 363104 44334
rect 363052 44270 363104 44276
rect 360580 44198 360608 44270
rect 360568 44192 360620 44198
rect 360568 44134 360620 44140
rect 359832 41948 359884 41954
rect 359832 41890 359884 41896
rect 359844 41834 359872 41890
rect 359844 41806 359950 41834
rect 360580 41820 360608 44134
rect 361120 41948 361172 41954
rect 361120 41890 361172 41896
rect 361132 41834 361160 41890
rect 361132 41806 361238 41834
rect 361767 41713 361823 42193
rect 362434 41818 362540 41834
rect 363064 41820 363092 44270
rect 363512 41948 363564 41954
rect 363512 41890 363564 41896
rect 363524 41834 363552 41890
rect 364260 41834 364288 46854
rect 404910 44296 404966 44305
rect 404910 44231 404966 44240
rect 406752 44260 406804 44266
rect 363524 41820 364288 41834
rect 362434 41812 362552 41818
rect 362434 41806 362500 41812
rect 363524 41806 364274 41820
rect 362500 41754 362552 41760
rect 364895 41713 364951 42193
rect 404924 41820 404952 44231
rect 406752 44202 406804 44208
rect 405527 41713 405583 42193
rect 406764 41820 406792 44202
rect 407408 41970 407436 46854
rect 414204 44464 414256 44470
rect 411074 44432 411130 44441
rect 414204 44406 414256 44412
rect 411074 44367 411130 44376
rect 407408 41954 407528 41970
rect 407408 41948 407540 41954
rect 407408 41942 407488 41948
rect 407408 41820 407436 41942
rect 407488 41890 407540 41896
rect 410248 41948 410300 41954
rect 410248 41890 410300 41896
rect 410260 41834 410288 41890
rect 409262 41818 409368 41834
rect 409262 41812 409380 41818
rect 409262 41806 409328 41812
rect 410260 41806 410458 41834
rect 411088 41820 411116 44367
rect 413560 44328 413612 44334
rect 412914 44296 412970 44305
rect 413560 44270 413612 44276
rect 412914 44231 412970 44240
rect 411536 41948 411588 41954
rect 411536 41890 411588 41896
rect 411548 41834 411576 41890
rect 412243 41834 412299 42193
rect 411548 41806 411746 41834
rect 412243 41818 412404 41834
rect 412928 41820 412956 44231
rect 413572 41820 413600 44270
rect 414216 44198 414244 44406
rect 417884 44328 417936 44334
rect 417884 44270 417936 44276
rect 414204 44192 414256 44198
rect 414204 44134 414256 44140
rect 414216 41820 414244 44134
rect 414572 41948 414624 41954
rect 414572 41890 414624 41896
rect 415860 41948 415912 41954
rect 415860 41890 415912 41896
rect 414584 41834 414612 41890
rect 415872 41834 415900 41890
rect 412243 41812 412416 41818
rect 412243 41806 412364 41812
rect 409328 41754 409380 41760
rect 412243 41713 412299 41806
rect 414584 41806 414782 41834
rect 415228 41818 415426 41834
rect 415216 41812 415426 41818
rect 412364 41754 412416 41760
rect 415268 41806 415426 41812
rect 415872 41806 416070 41834
rect 415216 41754 415268 41760
rect 416567 41713 416623 42193
rect 417266 41818 417372 41834
rect 417896 41820 417924 44270
rect 418252 41948 418304 41954
rect 418252 41890 418304 41896
rect 418264 41834 418292 41890
rect 419092 41834 419120 46854
rect 419722 44296 419778 44305
rect 419722 44231 419778 44240
rect 459650 44296 459706 44305
rect 459650 44231 459706 44240
rect 461492 44260 461544 44266
rect 419736 42193 419764 44231
rect 418264 41820 419120 41834
rect 419695 41820 419764 42193
rect 459664 41834 459692 44231
rect 461492 44202 461544 44208
rect 417266 41812 417384 41818
rect 417266 41806 417332 41812
rect 418264 41806 419106 41820
rect 417332 41754 417384 41760
rect 419695 41713 419751 41820
rect 459664 41806 459711 41834
rect 460327 41713 460383 42193
rect 461504 41834 461532 44202
rect 462148 41834 462176 46854
rect 465814 44432 465870 44441
rect 465814 44367 465870 44376
rect 468944 44396 468996 44402
rect 462320 41948 462372 41954
rect 462320 41890 462372 41896
rect 465080 41948 465132 41954
rect 465080 41890 465132 41896
rect 462332 41834 462360 41890
rect 465092 41834 465120 41890
rect 465828 41834 465856 44367
rect 468944 44338 468996 44344
rect 468300 44328 468352 44334
rect 467654 44296 467710 44305
rect 468300 44270 468352 44276
rect 467654 44231 467710 44240
rect 466368 41948 466420 41954
rect 466368 41890 466420 41896
rect 466380 41834 466408 41890
rect 467043 41834 467099 42193
rect 467668 41834 467696 44231
rect 468312 41834 468340 44270
rect 468956 44198 468984 44338
rect 472624 44328 472676 44334
rect 472624 44270 472676 44276
rect 468944 44192 468996 44198
rect 468944 44134 468996 44140
rect 468956 41834 468984 44134
rect 469404 41948 469456 41954
rect 469404 41890 469456 41896
rect 470692 41948 470744 41954
rect 470692 41890 470744 41896
rect 469416 41834 469444 41890
rect 470704 41834 470732 41890
rect 461504 41806 461551 41834
rect 462148 41806 462360 41834
rect 464035 41818 464200 41834
rect 464035 41812 464212 41818
rect 464035 41806 464160 41812
rect 465092 41806 465231 41834
rect 465828 41806 465875 41834
rect 466380 41806 466519 41834
rect 467043 41818 467236 41834
rect 467043 41812 467248 41818
rect 467043 41806 467196 41812
rect 464160 41754 464212 41760
rect 467043 41713 467099 41806
rect 467668 41806 467715 41834
rect 468312 41806 468359 41834
rect 468956 41806 469003 41834
rect 469416 41806 469555 41834
rect 470060 41818 470199 41834
rect 470048 41812 470199 41818
rect 467196 41754 467248 41760
rect 470100 41806 470199 41812
rect 470704 41806 470843 41834
rect 470048 41754 470100 41760
rect 471367 41713 471423 42193
rect 472636 41834 472664 44270
rect 473084 41948 473136 41954
rect 473084 41890 473136 41896
rect 473096 41834 473124 41890
rect 473832 41834 473860 46854
rect 474462 44432 474518 44441
rect 474462 44367 474518 44376
rect 474476 42193 474504 44367
rect 514482 44296 514538 44305
rect 514482 44231 514538 44240
rect 516324 44260 516376 44266
rect 472039 41818 472204 41834
rect 472039 41812 472216 41818
rect 472039 41806 472164 41812
rect 472636 41806 472683 41834
rect 473096 41806 473879 41834
rect 474476 41806 474551 42193
rect 514496 41820 514524 44231
rect 516324 44202 516376 44208
rect 472164 41754 472216 41760
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 516336 41820 516364 44202
rect 516980 41970 517008 46854
rect 523776 45620 523828 45626
rect 523776 45562 523828 45568
rect 518716 45552 518768 45558
rect 518716 45494 518768 45500
rect 518728 44266 518756 45494
rect 522486 44432 522542 44441
rect 523788 44402 523816 45562
rect 522486 44367 522542 44376
rect 523776 44396 523828 44402
rect 518806 44296 518862 44305
rect 518716 44260 518768 44266
rect 518806 44231 518862 44240
rect 518716 44202 518768 44208
rect 516980 41954 517100 41970
rect 516980 41948 517112 41954
rect 516980 41942 517060 41948
rect 516980 41820 517008 41942
rect 517060 41890 517112 41896
rect 518820 41820 518848 44231
rect 519912 41948 519964 41954
rect 519912 41890 519964 41896
rect 519924 41834 519952 41890
rect 519924 41806 520030 41834
rect 520647 41713 520703 42193
rect 521200 41948 521252 41954
rect 521200 41890 521252 41896
rect 521212 41834 521240 41890
rect 521212 41806 521318 41834
rect 521843 41713 521899 42193
rect 522500 41820 522528 44367
rect 523776 44338 523828 44344
rect 523132 44192 523184 44198
rect 523132 44134 523184 44140
rect 523144 41820 523172 44134
rect 523788 41820 523816 44338
rect 524970 44296 525026 44305
rect 524970 44231 525026 44240
rect 524984 42193 525012 44231
rect 527468 44198 527496 46854
rect 527456 44192 527508 44198
rect 527456 44134 527508 44140
rect 524236 41948 524288 41954
rect 524236 41890 524288 41896
rect 524248 41834 524276 41890
rect 524248 41806 524354 41834
rect 524971 41713 525027 42193
rect 525524 41948 525576 41954
rect 525524 41890 525576 41896
rect 525536 41834 525564 41890
rect 525536 41806 525642 41834
rect 526167 41713 526223 42193
rect 526732 41818 526838 41834
rect 527468 41820 527496 44134
rect 673472 42770 673500 113154
rect 673564 109546 673592 149026
rect 673748 139346 673776 154090
rect 673932 149054 673960 191898
rect 675312 190525 675340 198614
rect 675404 198492 675432 198614
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 675407 194807 675887 194863
rect 675407 192967 675887 193023
rect 675404 191962 675432 192372
rect 675392 191956 675444 191962
rect 675392 191898 675444 191904
rect 675407 191127 675887 191183
rect 675312 190497 675418 190525
rect 675407 160847 675887 160903
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675392 158636 675444 158642
rect 675392 158578 675444 158584
rect 675404 158522 675432 158578
rect 675312 158508 675432 158522
rect 675312 158494 675418 158508
rect 675312 154170 675340 158494
rect 675392 158364 675444 158370
rect 675392 158306 675444 158312
rect 675404 157828 675432 158306
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675392 155236 675444 155242
rect 675392 155178 675444 155184
rect 675404 154803 675432 155178
rect 675312 154154 675418 154170
rect 675300 154148 675418 154154
rect 675352 154142 675418 154148
rect 675300 154090 675352 154096
rect 675312 154059 675340 154090
rect 673840 149026 673960 149054
rect 675312 153501 675418 153529
rect 673840 146946 673868 149026
rect 673828 146940 673880 146946
rect 673828 146882 673880 146888
rect 673656 139318 673776 139346
rect 673656 113762 673684 139318
rect 673840 129734 673868 146882
rect 675312 145525 675340 153501
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675404 146946 675432 147356
rect 675392 146940 675444 146946
rect 675392 146882 675444 146888
rect 675407 146127 675887 146183
rect 675312 145497 675418 145525
rect 673748 129706 673868 129734
rect 673644 113756 673696 113762
rect 673644 113698 673696 113704
rect 673552 109540 673604 109546
rect 673552 109482 673604 109488
rect 673564 45626 673592 109482
rect 673644 108452 673696 108458
rect 673644 108394 673696 108400
rect 673656 46986 673684 108394
rect 673748 101726 673776 129706
rect 675407 115647 675887 115703
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675392 113756 675444 113762
rect 675392 113698 675444 113704
rect 675404 113297 675432 113698
rect 675312 113283 675432 113297
rect 675312 113269 675418 113283
rect 675312 108973 675340 113269
rect 675392 113212 675444 113218
rect 675392 113154 675444 113160
rect 675404 112639 675432 113154
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675404 109546 675432 109603
rect 675392 109540 675444 109546
rect 675392 109482 675444 109488
rect 675312 108959 675418 108973
rect 675312 108945 675432 108959
rect 675404 108458 675432 108945
rect 675392 108452 675444 108458
rect 675392 108394 675444 108400
rect 675312 108310 675418 108338
rect 673736 101720 673788 101726
rect 673736 101662 673788 101668
rect 673644 46980 673696 46986
rect 673644 46922 673696 46928
rect 673552 45620 673604 45626
rect 673552 45562 673604 45568
rect 673748 45558 673776 101662
rect 675312 100314 675340 108310
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675404 101726 675432 102151
rect 675392 101720 675444 101726
rect 675392 101662 675444 101668
rect 675407 100927 675887 100983
rect 675312 100286 675418 100314
rect 673736 45552 673788 45558
rect 673736 45494 673788 45500
rect 579896 42764 579948 42770
rect 579896 42706 579948 42712
rect 673460 42764 673512 42770
rect 673460 42706 673512 42712
rect 527916 41948 527968 41954
rect 527916 41890 527968 41896
rect 527928 41834 527956 41890
rect 526720 41812 526838 41818
rect 526772 41806 526838 41812
rect 527928 41806 528678 41834
rect 526720 41754 526772 41760
rect 529295 41713 529351 42193
rect 579908 41886 579936 42706
rect 568856 41880 568908 41886
rect 568856 41822 568908 41828
rect 579896 41880 579948 41886
rect 579896 41822 579948 41828
rect 568868 39681 568896 41822
rect 568854 39672 568910 39681
rect 568854 39607 568910 39616
rect 256238 39536 256294 39545
rect 256238 39471 256294 39480
<< via2 >>
rect 342166 997464 342222 997520
rect 585046 997464 585102 997520
rect 42430 870032 42486 870088
rect 44822 870032 44878 870088
rect 677598 818372 677654 818408
rect 677598 818352 677600 818372
rect 677600 818352 677652 818372
rect 677652 818352 677654 818372
rect 677690 513748 677692 513768
rect 677692 513748 677744 513768
rect 677744 513748 677746 513768
rect 677690 513712 677746 513748
rect 677506 425584 677562 425640
rect 44178 110472 44234 110528
rect 44822 110472 44878 110528
rect 44178 71848 44234 71904
rect 44822 71848 44878 71904
rect 93766 40160 93822 40216
rect 135166 40196 135168 40216
rect 135168 40196 135220 40216
rect 135220 40196 135222 40216
rect 135166 40160 135222 40196
rect 151726 46824 151782 46880
rect 188526 46824 188582 46880
rect 143538 40432 143594 40488
rect 143078 40160 143134 40216
rect 143538 40196 143540 40216
rect 143540 40196 143592 40216
rect 143592 40196 143594 40216
rect 143538 40160 143594 40196
rect 151726 40432 151782 40488
rect 404910 44240 404966 44296
rect 411074 44376 411130 44432
rect 412914 44240 412970 44296
rect 419722 44240 419778 44296
rect 459650 44240 459706 44296
rect 465814 44376 465870 44432
rect 467654 44240 467710 44296
rect 474462 44376 474518 44432
rect 514482 44240 514538 44296
rect 522486 44376 522542 44432
rect 518806 44240 518862 44296
rect 524970 44240 525026 44296
rect 568854 39616 568910 39672
rect 256238 39480 256294 39536
<< metal3 >>
rect 82144 997600 87144 1014070
rect 133544 997600 138544 1014070
rect 184944 997600 189944 1014070
rect 240478 997600 254800 1000736
rect 292078 997600 306400 1000736
rect 342161 997522 342227 997525
rect 343590 997522 343650 997628
rect 393878 997600 408200 1000736
rect 478744 997600 483744 1014070
rect 530144 997600 535144 1014070
rect 342161 997520 343650 997522
rect 342161 997464 342166 997520
rect 342222 997464 343650 997520
rect 342161 997462 343650 997464
rect 585041 997522 585107 997525
rect 585734 997522 585794 997628
rect 631944 997600 636944 1014070
rect 585041 997520 585794 997522
rect 585041 997464 585046 997520
rect 585102 997464 585794 997520
rect 585041 997462 585794 997464
rect 342161 997459 342227 997462
rect 585041 997459 585107 997462
rect 23530 960144 40000 965144
rect 677600 958656 694070 963656
rect 42425 870090 42491 870093
rect 44817 870090 44883 870093
rect 39622 870088 44883 870090
rect 39622 870032 42430 870088
rect 42486 870032 44822 870088
rect 44878 870032 44883 870088
rect 39622 870030 44883 870032
rect 39622 869924 39682 870030
rect 42425 870027 42491 870030
rect 44817 870027 44883 870030
rect 677593 818410 677659 818413
rect 677734 818410 677794 818652
rect 677593 818408 677794 818410
rect 677593 818352 677598 818408
rect 677654 818352 677794 818408
rect 677593 818350 677794 818352
rect 677593 818347 677659 818350
rect 677734 513773 677794 514012
rect 677685 513768 677794 513773
rect 677685 513712 677690 513768
rect 677746 513712 677794 513768
rect 677685 513710 677794 513712
rect 677685 513707 677751 513710
rect 678000 469900 685920 474700
rect 31680 440900 39600 445700
rect 677501 425642 677567 425645
rect 677734 425642 677794 425748
rect 677501 425640 677794 425642
rect 677501 425584 677506 425640
rect 677562 425584 677794 425640
rect 677501 425582 677794 425584
rect 677501 425579 677567 425582
rect 44173 110530 44239 110533
rect 44817 110530 44883 110533
rect 39652 110528 44883 110530
rect 39652 110472 44178 110528
rect 44234 110472 44822 110528
rect 44878 110472 44883 110528
rect 39652 110470 44883 110472
rect 44173 110467 44239 110470
rect 44817 110467 44883 110470
rect 44173 71906 44239 71909
rect 44817 71906 44883 71909
rect 39468 71904 44883 71906
rect 39468 71848 44178 71904
rect 44234 71848 44822 71904
rect 44878 71848 44883 71904
rect 39468 71846 44883 71848
rect 44173 71843 44239 71846
rect 44817 71843 44883 71846
rect 151721 46882 151787 46885
rect 188521 46882 188587 46885
rect 151721 46880 188587 46882
rect 151721 46824 151726 46880
rect 151782 46824 188526 46880
rect 188582 46824 188587 46880
rect 151721 46822 188587 46824
rect 151721 46819 151787 46822
rect 188521 46819 188587 46822
rect 411069 44434 411135 44437
rect 465809 44434 465875 44437
rect 474457 44434 474523 44437
rect 522481 44434 522547 44437
rect 411069 44432 419550 44434
rect 411069 44376 411074 44432
rect 411130 44376 419550 44432
rect 411069 44374 419550 44376
rect 411069 44371 411135 44374
rect 404905 44298 404971 44301
rect 412909 44298 412975 44301
rect 404905 44296 412975 44298
rect 404905 44240 404910 44296
rect 404966 44240 412914 44296
rect 412970 44240 412975 44296
rect 404905 44238 412975 44240
rect 419490 44298 419550 44374
rect 465809 44432 474523 44434
rect 465809 44376 465814 44432
rect 465870 44376 474462 44432
rect 474518 44376 474523 44432
rect 465809 44374 474523 44376
rect 465809 44371 465875 44374
rect 474457 44371 474523 44374
rect 516090 44432 522547 44434
rect 516090 44376 522486 44432
rect 522542 44376 522547 44432
rect 516090 44374 522547 44376
rect 419717 44298 419783 44301
rect 419490 44296 419783 44298
rect 419490 44240 419722 44296
rect 419778 44240 419783 44296
rect 419490 44238 419783 44240
rect 404905 44235 404971 44238
rect 412909 44235 412975 44238
rect 419717 44235 419783 44238
rect 459645 44298 459711 44301
rect 467649 44298 467715 44301
rect 459645 44296 467715 44298
rect 459645 44240 459650 44296
rect 459706 44240 467654 44296
rect 467710 44240 467715 44296
rect 459645 44238 467715 44240
rect 459645 44235 459711 44238
rect 467649 44235 467715 44238
rect 514477 44298 514543 44301
rect 516090 44298 516150 44374
rect 522481 44371 522547 44374
rect 514477 44296 516150 44298
rect 514477 44240 514482 44296
rect 514538 44240 516150 44296
rect 514477 44238 516150 44240
rect 518801 44298 518867 44301
rect 524965 44298 525031 44301
rect 518801 44296 525031 44298
rect 518801 44240 518806 44296
rect 518862 44240 524970 44296
rect 525026 44240 525031 44296
rect 518801 44238 525031 44240
rect 514477 44235 514543 44238
rect 518801 44235 518867 44238
rect 524965 44235 525031 44238
rect 143533 40490 143599 40493
rect 151721 40490 151787 40493
rect 143533 40488 151787 40490
rect 143533 40432 143538 40488
rect 143594 40432 151726 40488
rect 151782 40432 151787 40488
rect 143533 40430 151787 40432
rect 143533 40427 143599 40430
rect 145790 40354 145850 40430
rect 151721 40427 151787 40430
rect 145790 40294 145898 40354
rect 93761 40218 93827 40221
rect 135161 40218 135227 40221
rect 91142 40216 93827 40218
rect 91142 40160 93766 40216
rect 93822 40160 93827 40216
rect 91142 40158 93827 40160
rect 91142 39644 91202 40158
rect 93761 40155 93827 40158
rect 133094 40216 135227 40218
rect 133094 40160 135166 40216
rect 135222 40160 135227 40216
rect 133094 40158 135227 40160
rect 133094 39984 133154 40158
rect 135161 40155 135227 40158
rect 143073 40218 143139 40221
rect 143533 40218 143599 40221
rect 143073 40216 143458 40218
rect 143073 40160 143078 40216
rect 143134 40160 143458 40216
rect 143073 40158 143458 40160
rect 143073 40155 143139 40158
rect 141667 38031 141813 39999
rect 143398 39984 143458 40158
rect 143533 40216 144010 40218
rect 143533 40160 143538 40216
rect 143594 40160 144010 40216
rect 143533 40158 144010 40160
rect 143533 40155 143599 40158
rect 143950 39984 144010 40158
rect 145838 40014 145898 40294
rect 145820 39954 145898 40014
rect 568849 39674 568915 39677
rect 568849 39672 569204 39674
rect 568849 39616 568854 39672
rect 568910 39616 569204 39672
rect 568849 39614 569204 39616
rect 568849 39611 568915 39614
rect 256233 39538 256299 39541
rect 251406 39536 256299 39538
rect 251406 39480 256238 39536
rect 256294 39480 256299 39536
rect 251406 39478 256299 39480
rect 251406 39372 251466 39478
rect 256233 39475 256299 39478
<< metal4 >>
rect 679377 459800 680307 460054
rect 680587 459800 681277 459992
rect 688881 459800 688947 474800
rect 7 455645 4843 456093
rect 28653 440800 28719 455800
rect 32933 455546 33623 455800
rect 36323 455607 37013 455799
rect 37293 455546 38223 455800
rect 38503 455546 39593 455800
rect 132600 36323 132792 37013
rect 132600 30762 132868 31674
rect 132600 28653 147600 28719
<< metal5 >>
rect 78610 1018624 90778 1030788
rect 130010 1018624 142178 1030788
rect 181410 1018624 193578 1030788
rect 231810 1018624 243978 1030788
rect 283410 1018624 295578 1030788
rect 334810 1018624 346978 1030788
rect 385210 1018624 397378 1030788
rect 475210 1018624 487378 1030788
rect 526610 1018624 538778 1030788
rect 577010 1018624 589178 1030788
rect 628410 1018624 640578 1030788
rect 6811 956610 18975 968778
rect 698624 955022 710788 967190
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876180
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786620 19088 799160
rect 698512 774440 711002 786980
rect 6598 743420 19088 755960
rect 698512 729440 711002 741980
rect 6598 700220 19088 712760
rect 698512 684440 711002 696980
rect 6598 657020 19088 669560
rect 698512 639240 711002 651780
rect 6598 613820 19088 626360
rect 698512 594240 711002 606780
rect 6598 570620 19088 583160
rect 698512 549040 711002 561580
rect 6598 527420 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399820 19088 412360
rect 698512 371840 711002 384380
rect 6598 356620 19088 369160
rect 698512 326640 711002 339180
rect 6598 313420 19088 325960
rect 6598 270220 19088 282760
rect 698512 281640 711002 294180
rect 6598 227020 19088 239560
rect 698512 236640 711002 249180
rect 6598 183820 19088 196360
rect 698512 191440 711002 203980
rect 698512 146440 711002 158980
rect 6811 111610 18975 123778
rect 698512 101240 711002 113780
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200180 19088
rect 243266 6167 254146 19619
rect 296240 6598 308780 19088
rect 351040 6598 363580 19088
rect 405840 6598 418380 19088
rect 460640 6598 473180 19088
rect 515440 6598 527980 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use sky130_ef_io__corner_pad  mgmt_corner\[0\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_148 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_352
timestamp 1624635410
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1624635410
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1
timestamp 1624635410
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_152 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_151
timestamp 1624635410
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_150 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_149 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_159
timestamp 1624635410
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1624635410
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1624635410
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1624635410
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_163
timestamp 1624635410
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_162
timestamp 1624635410
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_161
timestamp 1624635410
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_160
timestamp 1624635410
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  mgmt_vssa_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 93800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_165
timestamp 1624635410
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_167
timestamp 1624635410
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_166
timestamp 1624635410
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1624635410
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_169
timestamp 1624635410
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_168
timestamp 1624635410
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1624635410
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1624635410
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1624635410
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1624635410
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1624635410
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_176
timestamp 1624635410
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_180
timestamp 1624635410
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_179
timestamp 1624635410
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_178
timestamp 1624635410
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_177
timestamp 1624635410
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_fd_io__top_xres4v2  resetb_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 147600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1624635410
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_186
timestamp 1624635410
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_185
timestamp 1624635410
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_184
timestamp 1624635410
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_183
timestamp 1624635410
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_182
timestamp 1624635410
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1624635410
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1624635410
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1624635410
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_195
timestamp 1624635410
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_194
timestamp 1624635410
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_193
timestamp 1624635410
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1624635410
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1624635410
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_197
timestamp 1624635410
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_196
timestamp 1624635410
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 202400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1624635410
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_203
timestamp 1624635410
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_202
timestamp 1624635410
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_201
timestamp 1624635410
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_200
timestamp 1624635410
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_199
timestamp 1624635410
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1624635410
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1624635410
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1624635410
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1624635410
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_214
timestamp 1624635410
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_213
timestamp 1624635410
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_212
timestamp 1624635410
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_211
timestamp 1624635410
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_210
timestamp 1624635410
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1624635410
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_clamped_pad  mgmt_vssd_lvclmap_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 256200 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1624635410
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1624635410
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_220
timestamp 1624635410
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_219
timestamp 1624635410
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_218
timestamp 1624635410
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_217
timestamp 1624635410
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_216
timestamp 1624635410
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1624635410
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1624635410
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1624635410
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1624635410
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_231
timestamp 1624635410
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_230
timestamp 1624635410
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_229
timestamp 1624635410
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_228
timestamp 1624635410
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_227
timestamp 1624635410
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1624635410
transform -1 0 311000 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_233
timestamp 1624635410
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_234
timestamp 1624635410
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1624635410
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_237
timestamp 1624635410
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_236
timestamp 1624635410
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_235
timestamp 1624635410
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1624635410
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1624635410
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1624635410
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1624635410
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_248
timestamp 1624635410
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_247
timestamp 1624635410
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_246
timestamp 1624635410
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_245
timestamp 1624635410
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_244
timestamp 1624635410
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1624635410
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1624635410
transform -1 0 365800 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_251
timestamp 1624635410
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_250
timestamp 1624635410
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1624635410
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1624635410
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_254
timestamp 1624635410
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_253
timestamp 1624635410
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_252
timestamp 1624635410
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1624635410
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1624635410
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1624635410
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1624635410
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_265
timestamp 1624635410
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_264
timestamp 1624635410
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_263
timestamp 1624635410
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_262
timestamp 1624635410
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_261
timestamp 1624635410
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1624635410
transform -1 0 420600 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_267
timestamp 1624635410
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1624635410
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1624635410
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1624635410
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_271
timestamp 1624635410
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_270
timestamp 1624635410
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_269
timestamp 1624635410
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_268
timestamp 1624635410
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_278
timestamp 1624635410
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1624635410
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1624635410
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1624635410
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_282
timestamp 1624635410
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_281
timestamp 1624635410
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_280
timestamp 1624635410
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_279
timestamp 1624635410
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1624635410
transform -1 0 475400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_284
timestamp 1624635410
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_285
timestamp 1624635410
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1624635410
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_288
timestamp 1624635410
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_287
timestamp 1624635410
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_286
timestamp 1624635410
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1624635410
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1624635410
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1624635410
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1624635410
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1624635410
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_299
timestamp 1624635410
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_298
timestamp 1624635410
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_297
timestamp 1624635410
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_296
timestamp 1624635410
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_295
timestamp 1624635410
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1624635410
transform -1 0 530200 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1624635410
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_305
timestamp 1624635410
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_304
timestamp 1624635410
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_303
timestamp 1624635410
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_302
timestamp 1624635410
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_301
timestamp 1624635410
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1624635410
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1624635410
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_312
timestamp 1624635410
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1624635410
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1624635410
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1624635410
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_316
timestamp 1624635410
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_315
timestamp 1624635410
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_314
timestamp 1624635410
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_313
timestamp 1624635410
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 584000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_320
timestamp 1624635410
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_319
timestamp 1624635410
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_318
timestamp 1624635410
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1624635410
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1624635410
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1624635410
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1624635410
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_322
timestamp 1624635410
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_321
timestamp 1624635410
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_330
timestamp 1624635410
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_329
timestamp 1624635410
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1624635410
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1624635410
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_333
timestamp 1624635410
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_332
timestamp 1624635410
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_331
timestamp 1624635410
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  mgmt_vdda_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_335
timestamp 1624635410
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_338
timestamp 1624635410
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_337
timestamp 1624635410
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_336
timestamp 1624635410
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1624635410
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_339
timestamp 1624635410
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1624635410
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1624635410
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1624635410
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1624635410
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1624635410
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_346
timestamp 1624635410
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_347
timestamp 1624635410
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1624635410
transform 0 1 676800 -1 0 40000
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_5um  FILLER_348
timestamp 1624635410
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_349
timestamp 1624635410
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_350
timestamp 1624635410
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_351
timestamp 1624635410
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_580
timestamp 1624635410
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_356
timestamp 1624635410
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_355
timestamp 1624635410
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_354
timestamp 1624635410
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_353
timestamp 1624635410
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_360
timestamp 1624635410
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_359
timestamp 1624635410
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_358
timestamp 1624635410
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_357
timestamp 1624635410
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_clamped_pad  mgmt_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 -1 39593 1 0 68000
box 0 -2107 17239 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_362
timestamp 1624635410
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_581
timestamp 1624635410
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_582
timestamp 1624635410
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_583
timestamp 1624635410
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_584
timestamp 1624635410
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1624635410
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1624635410
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_1 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 1 678007 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 1 678007 -1 0 70000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_587
timestamp 1624635410
transform 0 1 678007 -1 0 69000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_590
timestamp 1624635410
transform 0 1 678007 -1 0 75000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_591
timestamp 1624635410
transform 0 1 678007 -1 0 79000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_592
timestamp 1624635410
transform 0 1 678007 -1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_593
timestamp 1624635410
transform 0 1 678007 -1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_366
timestamp 1624635410
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_365
timestamp 1624635410
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_364
timestamp 1624635410
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_363
timestamp 1624635410
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_370
timestamp 1624635410
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_369
timestamp 1624635410
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_368
timestamp 1624635410
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_367
timestamp 1624635410
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_2
timestamp 1624635410
transform 0 -1 39593 1 0 126200
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1624635410
transform 0 -1 39593 1 0 125200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[0\]
timestamp 1624635410
transform 0 1 675407 -1 0 116000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_594
timestamp 1624635410
transform 0 1 678007 -1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1624635410
transform 0 1 678007 -1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1624635410
transform 0 1 678007 -1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_597
timestamp 1624635410
transform 0 1 678007 -1 0 100000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_599
timestamp 1624635410
transform 0 1 678007 -1 0 120000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_600
timestamp 1624635410
transform 0 1 678007 -1 0 124000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_601
timestamp 1624635410
transform 0 1 678007 -1 0 128000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_374
timestamp 1624635410
transform 0 -1 39593 1 0 127200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1624635410
transform 0 -1 39593 1 0 131200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_376
timestamp 1624635410
transform 0 -1 39593 1 0 135200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_377
timestamp 1624635410
transform 0 -1 39593 1 0 139200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_378
timestamp 1624635410
transform 0 -1 39593 1 0 143200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_379
timestamp 1624635410
transform 0 -1 39593 1 0 147200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_380
timestamp 1624635410
transform 0 -1 39593 1 0 151200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_381
timestamp 1624635410
transform 0 -1 39593 1 0 155200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_382
timestamp 1624635410
transform 0 -1 39593 1 0 159200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_383
timestamp 1624635410
transform 0 -1 39593 1 0 163200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1624635410
transform 0 -1 39593 1 0 167200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[1\]
timestamp 1624635410
transform 0 1 675407 -1 0 161200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_602
timestamp 1624635410
transform 0 1 678007 -1 0 132000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_603
timestamp 1624635410
transform 0 1 678007 -1 0 136000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_604
timestamp 1624635410
transform 0 1 678007 -1 0 140000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1624635410
transform 0 1 678007 -1 0 144000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_606
timestamp 1624635410
transform 0 1 678007 -1 0 145000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_607
timestamp 1624635410
transform 0 1 678007 -1 0 145200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_609
timestamp 1624635410
transform 0 1 678007 -1 0 165200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_610
timestamp 1624635410
transform 0 1 678007 -1 0 169200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_389
timestamp 1624635410
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_388
timestamp 1624635410
transform 0 -1 39593 1 0 181200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_387
timestamp 1624635410
transform 0 -1 39593 1 0 179200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_386
timestamp 1624635410
transform 0 -1 39593 1 0 175200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_385
timestamp 1624635410
transform 0 -1 39593 1 0 171200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[12\]
timestamp 1624635410
transform 0 -1 42193 1 0 181600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_391
timestamp 1624635410
transform 0 -1 39593 1 0 197600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1624635410
transform 0 -1 39593 1 0 209600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_393
timestamp 1624635410
transform 0 -1 39593 1 0 205600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_392
timestamp 1624635410
transform 0 -1 39593 1 0 201600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[2\]
timestamp 1624635410
transform 0 1 675407 -1 0 206200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_611
timestamp 1624635410
transform 0 1 678007 -1 0 173200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_612
timestamp 1624635410
transform 0 1 678007 -1 0 177200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_613
timestamp 1624635410
transform 0 1 678007 -1 0 181200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_614
timestamp 1624635410
transform 0 1 678007 -1 0 185200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1624635410
transform 0 1 678007 -1 0 189200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_616
timestamp 1624635410
transform 0 1 678007 -1 0 190200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1624635410
transform 0 1 678007 -1 0 210200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_619
timestamp 1624635410
transform 0 1 678007 -1 0 214200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_399
timestamp 1624635410
transform 0 -1 39593 1 0 224600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_398
timestamp 1624635410
transform 0 -1 39593 1 0 223600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_397
timestamp 1624635410
transform 0 -1 39593 1 0 221600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_396
timestamp 1624635410
transform 0 -1 39593 1 0 217600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_395
timestamp 1624635410
transform 0 -1 39593 1 0 213600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[11\]
timestamp 1624635410
transform 0 -1 42193 1 0 224800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_401
timestamp 1624635410
transform 0 -1 39593 1 0 240800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_404
timestamp 1624635410
transform 0 -1 39593 1 0 252800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_403
timestamp 1624635410
transform 0 -1 39593 1 0 248800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_402
timestamp 1624635410
transform 0 -1 39593 1 0 244800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[3\]
timestamp 1624635410
transform 0 1 675407 -1 0 251400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_620
timestamp 1624635410
transform 0 1 678007 -1 0 218200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_621
timestamp 1624635410
transform 0 1 678007 -1 0 222200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_622
timestamp 1624635410
transform 0 1 678007 -1 0 226200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_623
timestamp 1624635410
transform 0 1 678007 -1 0 230200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1624635410
transform 0 1 678007 -1 0 234200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_625
timestamp 1624635410
transform 0 1 678007 -1 0 235200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_626
timestamp 1624635410
transform 0 1 678007 -1 0 235400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1624635410
transform 0 1 678007 -1 0 255400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[10\]
timestamp 1624635410
transform 0 -1 42193 1 0 268000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1624635410
transform 0 -1 39593 1 0 256800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_406
timestamp 1624635410
transform 0 -1 39593 1 0 260800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_407
timestamp 1624635410
transform 0 -1 39593 1 0 264800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_408
timestamp 1624635410
transform 0 -1 39593 1 0 266800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_409
timestamp 1624635410
transform 0 -1 39593 1 0 267800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_411
timestamp 1624635410
transform 0 -1 39593 1 0 284000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_412
timestamp 1624635410
transform 0 -1 39593 1 0 288000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_413
timestamp 1624635410
transform 0 -1 39593 1 0 292000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[4\]
timestamp 1624635410
transform 0 1 675407 -1 0 296400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_629
timestamp 1624635410
transform 0 1 678007 -1 0 259400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_630
timestamp 1624635410
transform 0 1 678007 -1 0 263400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_631
timestamp 1624635410
transform 0 1 678007 -1 0 267400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_632
timestamp 1624635410
transform 0 1 678007 -1 0 271400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_633
timestamp 1624635410
transform 0 1 678007 -1 0 275400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1624635410
transform 0 1 678007 -1 0 279400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_635
timestamp 1624635410
transform 0 1 678007 -1 0 280400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_419
timestamp 1624635410
transform 0 -1 39593 1 0 311000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_418
timestamp 1624635410
transform 0 -1 39593 1 0 310000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_417
timestamp 1624635410
transform 0 -1 39593 1 0 308000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1624635410
transform 0 -1 39593 1 0 304000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1624635410
transform 0 -1 39593 1 0 300000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_414
timestamp 1624635410
transform 0 -1 39593 1 0 296000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[9\]
timestamp 1624635410
transform 0 -1 42193 1 0 311200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_421
timestamp 1624635410
transform 0 -1 39593 1 0 327200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_423
timestamp 1624635410
transform 0 -1 39593 1 0 335200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_422
timestamp 1624635410
transform 0 -1 39593 1 0 331200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[5\]
timestamp 1624635410
transform 0 1 675407 -1 0 341400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1624635410
transform 0 1 678007 -1 0 300400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_638
timestamp 1624635410
transform 0 1 678007 -1 0 304400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_639
timestamp 1624635410
transform 0 1 678007 -1 0 308400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_640
timestamp 1624635410
transform 0 1 678007 -1 0 312400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_641
timestamp 1624635410
transform 0 1 678007 -1 0 316400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_642
timestamp 1624635410
transform 0 1 678007 -1 0 320400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1624635410
transform 0 1 678007 -1 0 324400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_644
timestamp 1624635410
transform 0 1 678007 -1 0 325400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_428
timestamp 1624635410
transform 0 -1 39593 1 0 353200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_427
timestamp 1624635410
transform 0 -1 39593 1 0 351200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1624635410
transform 0 -1 39593 1 0 347200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1624635410
transform 0 -1 39593 1 0 343200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_424
timestamp 1624635410
transform 0 -1 39593 1 0 339200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_429
timestamp 1624635410
transform 0 -1 39593 1 0 354200
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[8\]
timestamp 1624635410
transform 0 -1 42193 1 0 354400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_433
timestamp 1624635410
transform 0 -1 39593 1 0 378400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_432
timestamp 1624635410
transform 0 -1 39593 1 0 374400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_431
timestamp 1624635410
transform 0 -1 39593 1 0 370400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_649
timestamp 1624635410
transform 0 1 678007 -1 0 357400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_648
timestamp 1624635410
transform 0 1 678007 -1 0 353400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_647
timestamp 1624635410
transform 0 1 678007 -1 0 349400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1624635410
transform 0 1 678007 -1 0 345400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_653
timestamp 1624635410
transform 0 1 678007 -1 0 370400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_652
timestamp 1624635410
transform 0 1 678007 -1 0 369400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_651
timestamp 1624635410
transform 0 1 678007 -1 0 365400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_650
timestamp 1624635410
transform 0 1 678007 -1 0 361400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_654
timestamp 1624635410
transform 0 1 678007 -1 0 370600
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[6\]
timestamp 1624635410
transform 0 1 675407 -1 0 386600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_437
timestamp 1624635410
transform 0 -1 39593 1 0 394400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1624635410
transform 0 -1 39593 1 0 390400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1624635410
transform 0 -1 39593 1 0 386400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_434
timestamp 1624635410
transform 0 -1 39593 1 0 382400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_439
timestamp 1624635410
transform 0 -1 39593 1 0 397400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_438
timestamp 1624635410
transform 0 -1 39593 1 0 396400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[7\]
timestamp 1624635410
transform 0 -1 42193 1 0 397600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_443
timestamp 1624635410
transform 0 -1 39593 1 0 421600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_442
timestamp 1624635410
transform 0 -1 39593 1 0 417600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_441
timestamp 1624635410
transform 0 -1 39593 1 0 413600
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1624635410
transform 0 1 678007 -1 0 430600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1624635410
transform 0 1 678007 -1 0 390600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_657
timestamp 1624635410
transform 0 1 678007 -1 0 394600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_658
timestamp 1624635410
transform 0 1 678007 -1 0 398600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_659
timestamp 1624635410
transform 0 1 678007 -1 0 402600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_660
timestamp 1624635410
transform 0 1 678007 -1 0 406600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_661
timestamp 1624635410
transform 0 1 678007 -1 0 410600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1624635410
transform 0 1 678007 -1 0 414600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_663
timestamp 1624635410
transform 0 1 678007 -1 0 415600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_449
timestamp 1624635410
transform 0 -1 39593 1 0 440600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_448
timestamp 1624635410
transform 0 -1 39593 1 0 439600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_447
timestamp 1624635410
transform 0 -1 39593 1 0 437600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1624635410
transform 0 -1 39593 1 0 433600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1624635410
transform 0 -1 39593 1 0 429600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_444
timestamp 1624635410
transform 0 -1 39593 1 0 425600
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_clamped2_pad  user2_vssd_lvclmap_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 -1 39593 1 0 440800
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_452
timestamp 1624635410
transform 0 -1 39593 1 0 459800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_451
timestamp 1624635410
transform 0 -1 39593 1 0 455800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_453
timestamp 1624635410
transform 0 -1 39593 1 0 463800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_667
timestamp 1624635410
transform 0 1 678007 -1 0 442600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1624635410
transform 0 1 678007 -1 0 438600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1624635410
transform 0 1 678007 -1 0 434600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_673
timestamp 1624635410
transform 0 1 678007 -1 0 459800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_672
timestamp 1624635410
transform 0 1 678007 -1 0 459600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1624635410
transform 0 1 678007 -1 0 458600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_670
timestamp 1624635410
transform 0 1 678007 -1 0 454600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_669
timestamp 1624635410
transform 0 1 678007 -1 0 450600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_668
timestamp 1624635410
transform 0 1 678007 -1 0 446600
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_clamped2_pad  user1_vssd_lvclmap_pad
timestamp 1624635410
transform 0 1 678007 -1 0 474800
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1624635410
transform 0 -1 39593 1 0 475800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1624635410
transform 0 -1 39593 1 0 471800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_454
timestamp 1624635410
transform 0 -1 39593 1 0 467800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_459
timestamp 1624635410
transform 0 -1 39593 1 0 482800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_458
timestamp 1624635410
transform 0 -1 39593 1 0 481800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_457
timestamp 1624635410
transform 0 -1 39593 1 0 479800
box 0 0 2000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user2_vdda_hvclamp_pad
timestamp 1624635410
transform 0 -1 39593 1 0 483000
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_463
timestamp 1624635410
transform 0 -1 39593 1 0 506000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_462
timestamp 1624635410
transform 0 -1 39593 1 0 502000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_461
timestamp 1624635410
transform 0 -1 39593 1 0 498000
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1624635410
transform 0 1 678007 -1 0 518800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1624635410
transform 0 1 678007 -1 0 478800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_676
timestamp 1624635410
transform 0 1 678007 -1 0 482800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_677
timestamp 1624635410
transform 0 1 678007 -1 0 486800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_678
timestamp 1624635410
transform 0 1 678007 -1 0 490800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_679
timestamp 1624635410
transform 0 1 678007 -1 0 494800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_680
timestamp 1624635410
transform 0 1 678007 -1 0 498800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1624635410
transform 0 1 678007 -1 0 502800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_682
timestamp 1624635410
transform 0 1 678007 -1 0 503800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[6\]
timestamp 1624635410
transform 0 -1 42193 1 0 525200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_464
timestamp 1624635410
transform 0 -1 39593 1 0 510000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1624635410
transform 0 -1 39593 1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1624635410
transform 0 -1 39593 1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_467
timestamp 1624635410
transform 0 -1 39593 1 0 522000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_468
timestamp 1624635410
transform 0 -1 39593 1 0 524000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_469
timestamp 1624635410
transform 0 -1 39593 1 0 525000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_471
timestamp 1624635410
transform 0 -1 39593 1 0 541200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_472
timestamp 1624635410
transform 0 -1 39593 1 0 545200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[7\]
timestamp 1624635410
transform 0 1 675407 -1 0 563800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1624635410
transform 0 1 678007 -1 0 522800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_685
timestamp 1624635410
transform 0 1 678007 -1 0 526800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_686
timestamp 1624635410
transform 0 1 678007 -1 0 530800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_687
timestamp 1624635410
transform 0 1 678007 -1 0 534800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_688
timestamp 1624635410
transform 0 1 678007 -1 0 538800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_689
timestamp 1624635410
transform 0 1 678007 -1 0 542800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1624635410
transform 0 1 678007 -1 0 546800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_691
timestamp 1624635410
transform 0 1 678007 -1 0 547800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1624635410
transform 0 -1 39593 1 0 561200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1624635410
transform 0 -1 39593 1 0 557200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_474
timestamp 1624635410
transform 0 -1 39593 1 0 553200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_473
timestamp 1624635410
transform 0 -1 39593 1 0 549200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_479
timestamp 1624635410
transform 0 -1 39593 1 0 568200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_478
timestamp 1624635410
transform 0 -1 39593 1 0 567200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_477
timestamp 1624635410
transform 0 -1 39593 1 0 565200
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[5\]
timestamp 1624635410
transform 0 -1 42193 1 0 568400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_482
timestamp 1624635410
transform 0 -1 39593 1 0 588400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_481
timestamp 1624635410
transform 0 -1 39593 1 0 584400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1624635410
transform 0 1 678007 -1 0 567800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1624635410
transform 0 1 678007 -1 0 571800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_695
timestamp 1624635410
transform 0 1 678007 -1 0 575800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_696
timestamp 1624635410
transform 0 1 678007 -1 0 579800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_697
timestamp 1624635410
transform 0 1 678007 -1 0 583800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_698
timestamp 1624635410
transform 0 1 678007 -1 0 587800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_699
timestamp 1624635410
transform 0 1 678007 -1 0 591800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1624635410
transform 0 -1 39593 1 0 604400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1624635410
transform 0 -1 39593 1 0 600400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_484
timestamp 1624635410
transform 0 -1 39593 1 0 596400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_483
timestamp 1624635410
transform 0 -1 39593 1 0 592400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_489
timestamp 1624635410
transform 0 -1 39593 1 0 611400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_488
timestamp 1624635410
transform 0 -1 39593 1 0 610400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_487
timestamp 1624635410
transform 0 -1 39593 1 0 608400
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[4\]
timestamp 1624635410
transform 0 -1 42193 1 0 611600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_492
timestamp 1624635410
transform 0 -1 39593 1 0 631600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_491
timestamp 1624635410
transform 0 -1 39593 1 0 627600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[8\]
timestamp 1624635410
transform 0 1 675407 -1 0 609000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_700
timestamp 1624635410
transform 0 1 678007 -1 0 592800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_701
timestamp 1624635410
transform 0 1 678007 -1 0 593000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1624635410
transform 0 1 678007 -1 0 613000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_704
timestamp 1624635410
transform 0 1 678007 -1 0 617000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_705
timestamp 1624635410
transform 0 1 678007 -1 0 621000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_706
timestamp 1624635410
transform 0 1 678007 -1 0 625000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_707
timestamp 1624635410
transform 0 1 678007 -1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_708
timestamp 1624635410
transform 0 1 678007 -1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1624635410
transform 0 -1 39593 1 0 647600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1624635410
transform 0 -1 39593 1 0 643600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_494
timestamp 1624635410
transform 0 -1 39593 1 0 639600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_493
timestamp 1624635410
transform 0 -1 39593 1 0 635600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_499
timestamp 1624635410
transform 0 -1 39593 1 0 654600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_498
timestamp 1624635410
transform 0 -1 39593 1 0 653600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_497
timestamp 1624635410
transform 0 -1 39593 1 0 651600
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[3\]
timestamp 1624635410
transform 0 -1 42193 1 0 654800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_502
timestamp 1624635410
transform 0 -1 39593 1 0 674800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_501
timestamp 1624635410
transform 0 -1 39593 1 0 670800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[9\]
timestamp 1624635410
transform 0 1 675407 -1 0 654000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1624635410
transform 0 1 678007 -1 0 637000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_710
timestamp 1624635410
transform 0 1 678007 -1 0 638000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1624635410
transform 0 1 678007 -1 0 658000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1624635410
transform 0 1 678007 -1 0 662000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_714
timestamp 1624635410
transform 0 1 678007 -1 0 666000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_715
timestamp 1624635410
transform 0 1 678007 -1 0 670000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_716
timestamp 1624635410
transform 0 1 678007 -1 0 674000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_717
timestamp 1624635410
transform 0 1 678007 -1 0 678000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[2\]
timestamp 1624635410
transform 0 -1 42193 1 0 698000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_503
timestamp 1624635410
transform 0 -1 39593 1 0 678800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_504
timestamp 1624635410
transform 0 -1 39593 1 0 682800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1624635410
transform 0 -1 39593 1 0 686800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1624635410
transform 0 -1 39593 1 0 690800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_507
timestamp 1624635410
transform 0 -1 39593 1 0 694800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_508
timestamp 1624635410
transform 0 -1 39593 1 0 696800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_509
timestamp 1624635410
transform 0 -1 39593 1 0 697800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_511
timestamp 1624635410
transform 0 -1 39593 1 0 714000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[10\]
timestamp 1624635410
transform 0 1 675407 -1 0 699200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1624635410
transform 0 1 678007 -1 0 682000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_719
timestamp 1624635410
transform 0 1 678007 -1 0 683000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_720
timestamp 1624635410
transform 0 1 678007 -1 0 683200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1624635410
transform 0 1 678007 -1 0 703200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_723
timestamp 1624635410
transform 0 1 678007 -1 0 707200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_724
timestamp 1624635410
transform 0 1 678007 -1 0 711200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_725
timestamp 1624635410
transform 0 1 678007 -1 0 715200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_726
timestamp 1624635410
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1624635410
transform 0 -1 39593 1 0 730000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_514
timestamp 1624635410
transform 0 -1 39593 1 0 726000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_513
timestamp 1624635410
transform 0 -1 39593 1 0 722000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_512
timestamp 1624635410
transform 0 -1 39593 1 0 718000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_519
timestamp 1624635410
transform 0 -1 39593 1 0 741000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_518
timestamp 1624635410
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_517
timestamp 1624635410
transform 0 -1 39593 1 0 738000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1624635410
transform 0 -1 39593 1 0 734000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[1\]
timestamp 1624635410
transform 0 -1 42193 1 0 741200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_521
timestamp 1624635410
transform 0 -1 39593 1 0 757200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[11\]
timestamp 1624635410
transform 0 1 675407 -1 0 744200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_727
timestamp 1624635410
transform 0 1 678007 -1 0 723200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1624635410
transform 0 1 678007 -1 0 727200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_729
timestamp 1624635410
transform 0 1 678007 -1 0 728200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1624635410
transform 0 1 678007 -1 0 748200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_732
timestamp 1624635410
transform 0 1 678007 -1 0 752200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_733
timestamp 1624635410
transform 0 1 678007 -1 0 756200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_734
timestamp 1624635410
transform 0 1 678007 -1 0 760200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1624635410
transform 0 -1 39593 1 0 773200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_524
timestamp 1624635410
transform 0 -1 39593 1 0 769200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_523
timestamp 1624635410
transform 0 -1 39593 1 0 765200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_522
timestamp 1624635410
transform 0 -1 39593 1 0 761200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_529
timestamp 1624635410
transform 0 -1 39593 1 0 784200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_528
timestamp 1624635410
transform 0 -1 39593 1 0 783200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_527
timestamp 1624635410
transform 0 -1 39593 1 0 781200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1624635410
transform 0 -1 39593 1 0 777200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[0\]
timestamp 1624635410
transform 0 -1 42193 1 0 784400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_531
timestamp 1624635410
transform 0 -1 39593 1 0 800400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[12\]
timestamp 1624635410
transform 0 1 675407 -1 0 789200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_735
timestamp 1624635410
transform 0 1 678007 -1 0 764200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_736
timestamp 1624635410
transform 0 1 678007 -1 0 768200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1624635410
transform 0 1 678007 -1 0 772200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_738
timestamp 1624635410
transform 0 1 678007 -1 0 773200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1624635410
transform 0 1 678007 -1 0 793200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1624635410
transform 0 1 678007 -1 0 797200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_742
timestamp 1624635410
transform 0 1 678007 -1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_743
timestamp 1624635410
transform 0 1 678007 -1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1624635410
transform 0 -1 39593 1 0 816400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_534
timestamp 1624635410
transform 0 -1 39593 1 0 812400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_533
timestamp 1624635410
transform 0 -1 39593 1 0 808400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_532
timestamp 1624635410
transform 0 -1 39593 1 0 804400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_539
timestamp 1624635410
transform 0 -1 39593 1 0 827400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_538
timestamp 1624635410
transform 0 -1 39593 1 0 826400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_537
timestamp 1624635410
transform 0 -1 39593 1 0 824400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1624635410
transform 0 -1 39593 1 0 820400
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user2_vssa_hvclamp_pad
timestamp 1624635410
transform 0 -1 39593 1 0 827600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_541
timestamp 1624635410
transform 0 -1 39593 1 0 842600
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1624635410
transform 0 1 678007 -1 0 833400
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_744
timestamp 1624635410
transform 0 1 678007 -1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_745
timestamp 1624635410
transform 0 1 678007 -1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_746
timestamp 1624635410
transform 0 1 678007 -1 0 817200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_747
timestamp 1624635410
transform 0 1 678007 -1 0 818200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_748
timestamp 1624635410
transform 0 1 678007 -1 0 818400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1624635410
transform 0 1 678007 -1 0 837400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_751
timestamp 1624635410
transform 0 1 678007 -1 0 841400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_752
timestamp 1624635410
transform 0 1 678007 -1 0 845400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1624635410
transform 0 -1 39593 1 0 858600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_544
timestamp 1624635410
transform 0 -1 39593 1 0 854600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_543
timestamp 1624635410
transform 0 -1 39593 1 0 850600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_542
timestamp 1624635410
transform 0 -1 39593 1 0 846600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_549
timestamp 1624635410
transform 0 -1 39593 1 0 869600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_548
timestamp 1624635410
transform 0 -1 39593 1 0 868600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_547
timestamp 1624635410
transform 0 -1 39593 1 0 866600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1624635410
transform 0 -1 39593 1 0 862600
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1624635410
transform 0 -1 39593 1 0 869800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_551
timestamp 1624635410
transform 0 -1 39593 1 0 884800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[13\]
timestamp 1624635410
transform 0 1 675407 -1 0 878400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_753
timestamp 1624635410
transform 0 1 678007 -1 0 849400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_754
timestamp 1624635410
transform 0 1 678007 -1 0 853400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_755
timestamp 1624635410
transform 0 1 678007 -1 0 857400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1624635410
transform 0 1 678007 -1 0 861400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_757
timestamp 1624635410
transform 0 1 678007 -1 0 862400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1624635410
transform 0 1 678007 -1 0 882400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1624635410
transform 0 1 678007 -1 0 886400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1624635410
transform 0 -1 39593 1 0 904800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1624635410
transform 0 -1 39593 1 0 900800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_554
timestamp 1624635410
transform 0 -1 39593 1 0 896800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_553
timestamp 1624635410
transform 0 -1 39593 1 0 892800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_552
timestamp 1624635410
transform 0 -1 39593 1 0 888800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_559
timestamp 1624635410
transform 0 -1 39593 1 0 911800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_558
timestamp 1624635410
transform 0 -1 39593 1 0 910800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_557
timestamp 1624635410
transform 0 -1 39593 1 0 908800
box 0 0 2000 39593
use sky130_ef_io__vccd_lvc_clamped2_pad  user2_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 -1 39593 1 0 912000
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_561
timestamp 1624635410
transform 0 -1 39593 1 0 927000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1624635410
transform 0 1 678007 -1 0 906400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_764
timestamp 1624635410
transform 0 1 678007 -1 0 902400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_763
timestamp 1624635410
transform 0 1 678007 -1 0 898400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_762
timestamp 1624635410
transform 0 1 678007 -1 0 894400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_761
timestamp 1624635410
transform 0 1 678007 -1 0 890400
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_clamped2_pad  user1_vccd_lvclamp_pad
timestamp 1624635410
transform 0 1 678007 -1 0 922600
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1624635410
transform 0 1 678007 -1 0 926600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_767
timestamp 1624635410
transform 0 1 678007 -1 0 907600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_766
timestamp 1624635410
transform 0 1 678007 -1 0 907400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_770
timestamp 1624635410
transform 0 1 678007 -1 0 930600
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[3\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 -1 40000 1 0 955200
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_562
timestamp 1624635410
transform 0 -1 39593 1 0 931000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_563
timestamp 1624635410
transform 0 -1 39593 1 0 935000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_564
timestamp 1624635410
transform 0 -1 39593 1 0 939000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1624635410
transform 0 -1 39593 1 0 943000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1624635410
transform 0 -1 39593 1 0 947000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1624635410
transform 0 -1 39593 1 0 951000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_568
timestamp 1624635410
transform 0 -1 39593 1 0 955000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_570
timestamp 1624635410
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[0\]
timestamp 1624635410
transform 0 1 677600 -1 0 968600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_771
timestamp 1624635410
transform 0 1 678007 -1 0 934600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_772
timestamp 1624635410
transform 0 1 678007 -1 0 938600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_773
timestamp 1624635410
transform 0 1 678007 -1 0 942600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_774
timestamp 1624635410
transform 0 1 678007 -1 0 946600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1624635410
transform 0 1 678007 -1 0 950600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_776
timestamp 1624635410
transform 0 1 678007 -1 0 952600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_777
timestamp 1624635410
transform 0 1 678007 -1 0 953600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_779
timestamp 1624635410
transform 0 1 678007 -1 0 972600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1624635410
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_574
timestamp 1624635410
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_573
timestamp 1624635410
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_572
timestamp 1624635410
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_571
timestamp 1624635410
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_579
timestamp 1624635410
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_578
timestamp 1624635410
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_577
timestamp 1624635410
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_576
timestamp 1624635410
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_5
timestamp 1624635410
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1624635410
transform 0 -1 40800 1 0 997600
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1624635410
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1624635410
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1624635410
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1624635410
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1624635410
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1624635410
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1624635410
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15
timestamp 1624635410
transform 1 0 77000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_14
timestamp 1624635410
transform 1 0 76800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_13
timestamp 1624635410
transform 1 0 72800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[2\]
timestamp 1624635410
transform 1 0 77200 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_17
timestamp 1624635410
transform 1 0 92200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1624635410
transform 1 0 96200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1624635410
transform 1 0 100200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1624635410
transform 1 0 104200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1624635410
transform 1 0 108200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1624635410
transform 1 0 112200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1624635410
transform 1 0 116200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1624635410
transform 1 0 120200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1624635410
transform 1 0 124200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_27
timestamp 1624635410
transform 1 0 128400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_26
timestamp 1624635410
transform 1 0 128200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[1\]
timestamp 1624635410
transform 1 0 128600 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1624635410
transform 1 0 155600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1624635410
transform 1 0 151600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_30
timestamp 1624635410
transform 1 0 147600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_29
timestamp 1624635410
transform 1 0 143600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1624635410
transform 1 0 167600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1624635410
transform 1 0 163600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1624635410
transform 1 0 159600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[0\]
timestamp 1624635410
transform 1 0 180000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1624635410
transform 1 0 171600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1624635410
transform 1 0 175600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_38
timestamp 1624635410
transform 1 0 179600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_39
timestamp 1624635410
transform 1 0 179800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_41
timestamp 1624635410
transform 1 0 195000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_42
timestamp 1624635410
transform 1 0 199000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_43
timestamp 1624635410
transform 1 0 203000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1624635410
transform 1 0 207000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__top_power_hvc  user2_analog_pad_with_clamp\[1\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 1 0 221000 0 1 998007
box 0 -407 33800 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1624635410
transform 1 0 211000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1624635410
transform 1 0 215000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_47
timestamp 1624635410
transform 1 0 219000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_57
timestamp 1624635410
transform 1 0 272400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_56
timestamp 1624635410
transform 1 0 272200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1624635410
transform 1 0 272000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1624635410
transform 1 0 271800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_53
timestamp 1624635410
transform 1 0 270800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_52
timestamp 1624635410
transform 1 0 266800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1624635410
transform 1 0 262800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1624635410
transform 1 0 258800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1624635410
transform 1 0 254800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__top_power_hvc  user2_analog_pad_with_clamp\[0\]
timestamp 1624635410
transform 1 0 272600 0 1 998007
box 0 -407 33800 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[1\]
timestamp 1624635410
transform 1 0 333400 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_59
timestamp 1624635410
transform 1 0 306400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1624635410
transform 1 0 310400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1624635410
transform 1 0 314400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1624635410
transform 1 0 318400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1624635410
transform 1 0 322400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1624635410
transform 1 0 326400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_65
timestamp 1624635410
transform 1 0 330400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_66
timestamp 1624635410
transform 1 0 332400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__top_power_hvc  user1_analog_pad_with_clamp
timestamp 1624635410
transform 1 0 374400 0 1 998007
box 0 -407 33800 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_68
timestamp 1624635410
transform 1 0 348400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_69
timestamp 1624635410
transform 1 0 352400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_70
timestamp 1624635410
transform 1 0 356400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1624635410
transform 1 0 360400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1624635410
transform 1 0 364400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1624635410
transform 1 0 368400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0
timestamp 1624635410
transform 1 0 372400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_0
timestamp 1624635410
transform 1 0 373400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_77
timestamp 1624635410
transform 1 0 408200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1624635410
transform 1 0 412200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_79
timestamp 1624635410
transform 1 0 416200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_80
timestamp 1624635410
transform 1 0 420200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_81
timestamp 1624635410
transform 1 0 424200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_82
timestamp 1624635410
transform 1 0 428200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_83
timestamp 1624635410
transform 1 0 432200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_84
timestamp 1624635410
transform 1 0 436200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_85
timestamp 1624635410
transform 1 0 440200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1624635410
transform 1 0 444200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1624635410
transform 1 0 448200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1624635410
transform 1 0 452200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1624635410
transform 1 0 456200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1624635410
transform 1 0 460200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_96
timestamp 1624635410
transform 1 0 473600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1624635410
transform 1 0 473400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_94
timestamp 1624635410
transform 1 0 473200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_93
timestamp 1624635410
transform 1 0 472200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_92
timestamp 1624635410
transform 1 0 468200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1624635410
transform 1 0 464200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[3\]
timestamp 1624635410
transform 1 0 473800 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_99
timestamp 1624635410
transform 1 0 492800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_98
timestamp 1624635410
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1624635410
transform 1 0 504800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1624635410
transform 1 0 500800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1624635410
transform 1 0 496800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_106
timestamp 1624635410
transform 1 0 520800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_105
timestamp 1624635410
transform 1 0 516800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1624635410
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1624635410
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_108
timestamp 1624635410
transform 1 0 525000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_107
timestamp 1624635410
transform 1 0 524800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[2\]
timestamp 1624635410
transform 1 0 525200 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1624635410
transform 1 0 548200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1624635410
transform 1 0 544200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_110
timestamp 1624635410
transform 1 0 540200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1624635410
transform 1 0 560200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1624635410
transform 1 0 556200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1624635410
transform 1 0 552200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_121
timestamp 1624635410
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_120
timestamp 1624635410
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_119
timestamp 1624635410
transform 1 0 574200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_118
timestamp 1624635410
transform 1 0 572200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_117
timestamp 1624635410
transform 1 0 568200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_116
timestamp 1624635410
transform 1 0 564200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1624635410
transform 1 0 575600 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_123
timestamp 1624635410
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_126
timestamp 1624635410
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1624635410
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_124
timestamp 1624635410
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_130
timestamp 1624635410
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_129
timestamp 1624635410
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_128
timestamp 1624635410
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_127
timestamp 1624635410
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_133
timestamp 1624635410
transform 1 0 626800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_132
timestamp 1624635410
transform 1 0 626600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1624635410
transform 1 0 622600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[1\]
timestamp 1624635410
transform 1 0 627000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_135
timestamp 1624635410
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_136
timestamp 1624635410
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_137
timestamp 1624635410
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_138
timestamp 1624635410
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_139
timestamp 1624635410
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_140
timestamp 1624635410
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_141
timestamp 1624635410
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_142
timestamp 1624635410
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_143
timestamp 1624635410
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1624635410
transform 0 1 678007 -1 0 992600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_783
timestamp 1624635410
transform 0 1 678007 -1 0 988600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_782
timestamp 1624635410
transform 0 1 678007 -1 0 984600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_781
timestamp 1624635410
transform 0 1 678007 -1 0 980600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_780
timestamp 1624635410
transform 0 1 678007 -1 0 976600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_786
timestamp 1624635410
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1624635410
transform 0 1 678007 -1 0 996600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_147
timestamp 1624635410
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_146
timestamp 1624635410
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_145
timestamp 1624635410
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_144
timestamp 1624635410
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__corner_pad  user1_corner
timestamp 1624635410
transform 1 0 677600 0 1 996800
box 0 0 40000 40800
<< labels >>
rlabel metal5 s 187640 6598 200180 19088 6 clock
port 0 nsew signal input
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 1 nsew signal tristate
rlabel metal2 s 194043 41713 194099 42193 6 por
port 2 nsew signal input
rlabel metal5 s 351040 6598 363580 19088 6 flash_clk
port 3 nsew signal tristate
rlabel metal2 s 361767 41713 361823 42193 6 flash_clk_core
port 4 nsew signal input
rlabel metal2 s 357443 41713 357499 42193 6 flash_clk_ieb_core
port 5 nsew signal input
rlabel metal2 s 364895 41713 364951 42193 6 flash_clk_oeb_core
port 6 nsew signal input
rlabel metal5 s 296240 6598 308780 19088 6 flash_csb
port 7 nsew signal tristate
rlabel metal2 s 306967 41713 307023 42193 6 flash_csb_core
port 8 nsew signal input
rlabel metal2 s 302643 41713 302699 42193 6 flash_csb_ieb_core
port 9 nsew signal input
rlabel metal2 s 310095 41713 310151 42193 6 flash_csb_oeb_core
port 10 nsew signal input
rlabel metal5 s 405840 6598 418380 19088 6 flash_io0
port 11 nsew signal bidirectional
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 12 nsew signal tristate
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 13 nsew signal input
rlabel metal2 s 412243 41713 412299 42193 6 flash_io0_ieb_core
port 14 nsew signal input
rlabel metal2 s 419695 41713 419751 42193 6 flash_io0_oeb_core
port 15 nsew signal input
rlabel metal5 s 460640 6598 473180 19088 6 flash_io1
port 16 nsew signal bidirectional
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 17 nsew signal tristate
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 18 nsew signal input
rlabel metal2 s 467043 41713 467099 42193 6 flash_io1_ieb_core
port 19 nsew signal input
rlabel metal2 s 474495 41713 474551 42193 6 flash_io1_oeb_core
port 20 nsew signal input
rlabel metal5 s 515440 6598 527980 19088 6 gpio
port 21 nsew signal bidirectional
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 22 nsew signal tristate
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 23 nsew signal input
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 24 nsew signal input
rlabel metal2 s 524971 41713 525027 42193 6 gpio_mode1_core
port 25 nsew signal input
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 26 nsew signal input
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 27 nsew signal input
rlabel metal5 s 6167 70054 19619 80934 6 vccd_pad
port 28 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18975 6 vdda_pad
port 29 nsew signal bidirectional
rlabel metal5 s 6811 111610 18975 123778 6 vddio_pad
port 30 nsew signal bidirectional
rlabel metal5 s 6811 871210 18975 883378 6 vddio_pad2
port 31 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18975 6 vssa_pad
port 32 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19619 6 vssd_pad
port 33 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18975 6 vssio_pad
port 34 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030788 6 vssio_pad2
port 35 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113780 6 mprj_io[0]
port 36 nsew signal bidirectional
rlabel metal2 s 675407 105803 675887 105859 6 mprj_io_analog_en[0]
port 37 nsew signal input
rlabel metal2 s 675407 107091 675887 107147 6 mprj_io_analog_pol[0]
port 38 nsew signal input
rlabel metal2 s 675407 110127 675887 110183 6 mprj_io_analog_sel[0]
port 39 nsew signal input
rlabel metal2 s 675407 106447 675887 106503 6 mprj_io_dm[0]
port 40 nsew signal input
rlabel metal2 s 675407 104607 675887 104663 6 mprj_io_dm[1]
port 41 nsew signal input
rlabel metal2 s 675407 110771 675887 110827 6 mprj_io_dm[2]
port 42 nsew signal input
rlabel metal2 s 675407 111415 675887 111471 6 mprj_io_holdover[0]
port 43 nsew signal input
rlabel metal2 s 675407 114451 675887 114507 6 mprj_io_ib_mode_sel[0]
port 44 nsew signal input
rlabel metal2 s 675407 107643 675887 107699 6 mprj_io_inp_dis[0]
port 45 nsew signal input
rlabel metal2 s 675407 115095 675887 115151 6 mprj_io_oeb[0]
port 46 nsew signal input
rlabel metal2 s 675407 111967 675887 112023 6 mprj_io_out[0]
port 47 nsew signal input
rlabel metal2 s 675407 102767 675887 102823 6 mprj_io_slow_sel[0]
port 48 nsew signal input
rlabel metal2 s 675407 113807 675887 113863 6 mprj_io_vtrip_sel[0]
port 49 nsew signal input
rlabel metal2 s 675407 100927 675887 100983 6 mprj_io_in[0]
port 50 nsew signal tristate
rlabel metal2 s 675407 115647 675887 115703 6 mprj_io_in_3v3[0]
port 51 nsew signal tristate
rlabel metal2 s 675407 686611 675887 686667 6 mprj_gpio_analog[3]
port 52 nsew signal bidirectional
rlabel metal2 s 675407 688451 675887 688507 6 mprj_gpio_noesd[3]
port 53 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696980 6 mprj_io[10]
port 54 nsew signal bidirectional
rlabel metal2 s 675407 689003 675887 689059 6 mprj_io_analog_en[10]
port 55 nsew signal input
rlabel metal2 s 675407 690291 675887 690347 6 mprj_io_analog_pol[10]
port 56 nsew signal input
rlabel metal2 s 675407 693327 675887 693383 6 mprj_io_analog_sel[10]
port 57 nsew signal input
rlabel metal2 s 675407 689647 675887 689703 6 mprj_io_dm[30]
port 58 nsew signal input
rlabel metal2 s 675407 687807 675887 687863 6 mprj_io_dm[31]
port 59 nsew signal input
rlabel metal2 s 675407 693971 675887 694027 6 mprj_io_dm[32]
port 60 nsew signal input
rlabel metal2 s 675407 694615 675887 694671 6 mprj_io_holdover[10]
port 61 nsew signal input
rlabel metal2 s 675407 697651 675887 697707 6 mprj_io_ib_mode_sel[10]
port 62 nsew signal input
rlabel metal2 s 675407 690843 675887 690899 6 mprj_io_inp_dis[10]
port 63 nsew signal input
rlabel metal2 s 675407 698295 675887 698351 6 mprj_io_oeb[10]
port 64 nsew signal input
rlabel metal2 s 675407 695167 675887 695223 6 mprj_io_out[10]
port 65 nsew signal input
rlabel metal2 s 675407 685967 675887 686023 6 mprj_io_slow_sel[10]
port 66 nsew signal input
rlabel metal2 s 675407 697007 675887 697063 6 mprj_io_vtrip_sel[10]
port 67 nsew signal input
rlabel metal2 s 675407 684127 675887 684183 6 mprj_io_in[10]
port 68 nsew signal tristate
rlabel metal2 s 675407 698847 675887 698903 6 mprj_io_in_3v3[10]
port 69 nsew signal tristate
rlabel metal2 s 675407 731611 675887 731667 6 mprj_gpio_analog[4]
port 70 nsew signal bidirectional
rlabel metal2 s 675407 733451 675887 733507 6 mprj_gpio_noesd[4]
port 71 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741980 6 mprj_io[11]
port 72 nsew signal bidirectional
rlabel metal2 s 675407 734003 675887 734059 6 mprj_io_analog_en[11]
port 73 nsew signal input
rlabel metal2 s 675407 735291 675887 735347 6 mprj_io_analog_pol[11]
port 74 nsew signal input
rlabel metal2 s 675407 738327 675887 738383 6 mprj_io_analog_sel[11]
port 75 nsew signal input
rlabel metal2 s 675407 734647 675887 734703 6 mprj_io_dm[33]
port 76 nsew signal input
rlabel metal2 s 675407 732807 675887 732863 6 mprj_io_dm[34]
port 77 nsew signal input
rlabel metal2 s 675407 738971 675887 739027 6 mprj_io_dm[35]
port 78 nsew signal input
rlabel metal2 s 675407 739615 675887 739671 6 mprj_io_holdover[11]
port 79 nsew signal input
rlabel metal2 s 675407 742651 675887 742707 6 mprj_io_ib_mode_sel[11]
port 80 nsew signal input
rlabel metal2 s 675407 735843 675887 735899 6 mprj_io_inp_dis[11]
port 81 nsew signal input
rlabel metal2 s 675407 743295 675887 743351 6 mprj_io_oeb[11]
port 82 nsew signal input
rlabel metal2 s 675407 740167 675887 740223 6 mprj_io_out[11]
port 83 nsew signal input
rlabel metal2 s 675407 730967 675887 731023 6 mprj_io_slow_sel[11]
port 84 nsew signal input
rlabel metal2 s 675407 742007 675887 742063 6 mprj_io_vtrip_sel[11]
port 85 nsew signal input
rlabel metal2 s 675407 729127 675887 729183 6 mprj_io_in[11]
port 86 nsew signal tristate
rlabel metal2 s 675407 743847 675887 743903 6 mprj_io_in_3v3[11]
port 87 nsew signal tristate
rlabel metal2 s 675407 776611 675887 776667 6 mprj_gpio_analog[5]
port 88 nsew signal bidirectional
rlabel metal2 s 675407 778451 675887 778507 6 mprj_gpio_noesd[5]
port 89 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786980 6 mprj_io[12]
port 90 nsew signal bidirectional
rlabel metal2 s 675407 779003 675887 779059 6 mprj_io_analog_en[12]
port 91 nsew signal input
rlabel metal2 s 675407 780291 675887 780347 6 mprj_io_analog_pol[12]
port 92 nsew signal input
rlabel metal2 s 675407 783327 675887 783383 6 mprj_io_analog_sel[12]
port 93 nsew signal input
rlabel metal2 s 675407 779647 675887 779703 6 mprj_io_dm[36]
port 94 nsew signal input
rlabel metal2 s 675407 777807 675887 777863 6 mprj_io_dm[37]
port 95 nsew signal input
rlabel metal2 s 675407 783971 675887 784027 6 mprj_io_dm[38]
port 96 nsew signal input
rlabel metal2 s 675407 784615 675887 784671 6 mprj_io_holdover[12]
port 97 nsew signal input
rlabel metal2 s 675407 787651 675887 787707 6 mprj_io_ib_mode_sel[12]
port 98 nsew signal input
rlabel metal2 s 675407 780843 675887 780899 6 mprj_io_inp_dis[12]
port 99 nsew signal input
rlabel metal2 s 675407 788295 675887 788351 6 mprj_io_oeb[12]
port 100 nsew signal input
rlabel metal2 s 675407 785167 675887 785223 6 mprj_io_out[12]
port 101 nsew signal input
rlabel metal2 s 675407 775967 675887 776023 6 mprj_io_slow_sel[12]
port 102 nsew signal input
rlabel metal2 s 675407 787007 675887 787063 6 mprj_io_vtrip_sel[12]
port 103 nsew signal input
rlabel metal2 s 675407 774127 675887 774183 6 mprj_io_in[12]
port 104 nsew signal tristate
rlabel metal2 s 675407 788847 675887 788903 6 mprj_io_in_3v3[12]
port 105 nsew signal tristate
rlabel metal2 s 675407 865811 675887 865867 6 mprj_gpio_analog[6]
port 106 nsew signal bidirectional
rlabel metal2 s 675407 867651 675887 867707 6 mprj_gpio_noesd[6]
port 107 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876180 6 mprj_io[13]
port 108 nsew signal bidirectional
rlabel metal2 s 675407 868203 675887 868259 6 mprj_io_analog_en[13]
port 109 nsew signal input
rlabel metal2 s 675407 869491 675887 869547 6 mprj_io_analog_pol[13]
port 110 nsew signal input
rlabel metal2 s 675407 872527 675887 872583 6 mprj_io_analog_sel[13]
port 111 nsew signal input
rlabel metal2 s 675407 868847 675887 868903 6 mprj_io_dm[39]
port 112 nsew signal input
rlabel metal2 s 675407 867007 675887 867063 6 mprj_io_dm[40]
port 113 nsew signal input
rlabel metal2 s 675407 873171 675887 873227 6 mprj_io_dm[41]
port 114 nsew signal input
rlabel metal2 s 675407 873815 675887 873871 6 mprj_io_holdover[13]
port 115 nsew signal input
rlabel metal2 s 675407 876851 675887 876907 6 mprj_io_ib_mode_sel[13]
port 116 nsew signal input
rlabel metal2 s 675407 870043 675887 870099 6 mprj_io_inp_dis[13]
port 117 nsew signal input
rlabel metal2 s 675407 877495 675887 877551 6 mprj_io_oeb[13]
port 118 nsew signal input
rlabel metal2 s 675407 874367 675887 874423 6 mprj_io_out[13]
port 119 nsew signal input
rlabel metal2 s 675407 865167 675887 865223 6 mprj_io_slow_sel[13]
port 120 nsew signal input
rlabel metal2 s 675407 876207 675887 876263 6 mprj_io_vtrip_sel[13]
port 121 nsew signal input
rlabel metal2 s 675407 863327 675887 863383 6 mprj_io_in[13]
port 122 nsew signal tristate
rlabel metal2 s 675407 878047 675887 878103 6 mprj_io_in_3v3[13]
port 123 nsew signal tristate
rlabel metal5 s 698512 146440 711002 158980 6 mprj_io[1]
port 124 nsew signal bidirectional
rlabel metal2 s 675407 151003 675887 151059 6 mprj_io_analog_en[1]
port 125 nsew signal input
rlabel metal2 s 675407 152291 675887 152347 6 mprj_io_analog_pol[1]
port 126 nsew signal input
rlabel metal2 s 675407 155327 675887 155383 6 mprj_io_analog_sel[1]
port 127 nsew signal input
rlabel metal2 s 675407 151647 675887 151703 6 mprj_io_dm[3]
port 128 nsew signal input
rlabel metal2 s 675407 149807 675887 149863 6 mprj_io_dm[4]
port 129 nsew signal input
rlabel metal2 s 675407 155971 675887 156027 6 mprj_io_dm[5]
port 130 nsew signal input
rlabel metal2 s 675407 156615 675887 156671 6 mprj_io_holdover[1]
port 131 nsew signal input
rlabel metal2 s 675407 159651 675887 159707 6 mprj_io_ib_mode_sel[1]
port 132 nsew signal input
rlabel metal2 s 675407 152843 675887 152899 6 mprj_io_inp_dis[1]
port 133 nsew signal input
rlabel metal2 s 675407 160295 675887 160351 6 mprj_io_oeb[1]
port 134 nsew signal input
rlabel metal2 s 675407 157167 675887 157223 6 mprj_io_out[1]
port 135 nsew signal input
rlabel metal2 s 675407 147967 675887 148023 6 mprj_io_slow_sel[1]
port 136 nsew signal input
rlabel metal2 s 675407 159007 675887 159063 6 mprj_io_vtrip_sel[1]
port 137 nsew signal input
rlabel metal2 s 675407 146127 675887 146183 6 mprj_io_in[1]
port 138 nsew signal tristate
rlabel metal2 s 675407 160847 675887 160903 6 mprj_io_in_3v3[1]
port 139 nsew signal tristate
rlabel metal5 s 698512 191440 711002 203980 6 mprj_io[2]
port 140 nsew signal bidirectional
rlabel metal2 s 675407 196003 675887 196059 6 mprj_io_analog_en[2]
port 141 nsew signal input
rlabel metal2 s 675407 197291 675887 197347 6 mprj_io_analog_pol[2]
port 142 nsew signal input
rlabel metal2 s 675407 200327 675887 200383 6 mprj_io_analog_sel[2]
port 143 nsew signal input
rlabel metal2 s 675407 196647 675887 196703 6 mprj_io_dm[6]
port 144 nsew signal input
rlabel metal2 s 675407 194807 675887 194863 6 mprj_io_dm[7]
port 145 nsew signal input
rlabel metal2 s 675407 200971 675887 201027 6 mprj_io_dm[8]
port 146 nsew signal input
rlabel metal2 s 675407 201615 675887 201671 6 mprj_io_holdover[2]
port 147 nsew signal input
rlabel metal2 s 675407 204651 675887 204707 6 mprj_io_ib_mode_sel[2]
port 148 nsew signal input
rlabel metal2 s 675407 197843 675887 197899 6 mprj_io_inp_dis[2]
port 149 nsew signal input
rlabel metal2 s 675407 205295 675887 205351 6 mprj_io_oeb[2]
port 150 nsew signal input
rlabel metal2 s 675407 202167 675887 202223 6 mprj_io_out[2]
port 151 nsew signal input
rlabel metal2 s 675407 192967 675887 193023 6 mprj_io_slow_sel[2]
port 152 nsew signal input
rlabel metal2 s 675407 204007 675887 204063 6 mprj_io_vtrip_sel[2]
port 153 nsew signal input
rlabel metal2 s 675407 191127 675887 191183 6 mprj_io_in[2]
port 154 nsew signal tristate
rlabel metal2 s 675407 205847 675887 205903 6 mprj_io_in_3v3[2]
port 155 nsew signal tristate
rlabel metal5 s 698512 236640 711002 249180 6 mprj_io[3]
port 156 nsew signal bidirectional
rlabel metal2 s 675407 241203 675887 241259 6 mprj_io_analog_en[3]
port 157 nsew signal input
rlabel metal2 s 675407 242491 675887 242547 6 mprj_io_analog_pol[3]
port 158 nsew signal input
rlabel metal2 s 675407 245527 675887 245583 6 mprj_io_analog_sel[3]
port 159 nsew signal input
rlabel metal2 s 675407 240007 675887 240063 6 mprj_io_dm[10]
port 160 nsew signal input
rlabel metal2 s 675407 246171 675887 246227 6 mprj_io_dm[11]
port 161 nsew signal input
rlabel metal2 s 675407 241847 675887 241903 6 mprj_io_dm[9]
port 162 nsew signal input
rlabel metal2 s 675407 246815 675887 246871 6 mprj_io_holdover[3]
port 163 nsew signal input
rlabel metal2 s 675407 249851 675887 249907 6 mprj_io_ib_mode_sel[3]
port 164 nsew signal input
rlabel metal2 s 675407 243043 675887 243099 6 mprj_io_inp_dis[3]
port 165 nsew signal input
rlabel metal2 s 675407 250495 675887 250551 6 mprj_io_oeb[3]
port 166 nsew signal input
rlabel metal2 s 675407 247367 675887 247423 6 mprj_io_out[3]
port 167 nsew signal input
rlabel metal2 s 675407 238167 675887 238223 6 mprj_io_slow_sel[3]
port 168 nsew signal input
rlabel metal2 s 675407 249207 675887 249263 6 mprj_io_vtrip_sel[3]
port 169 nsew signal input
rlabel metal2 s 675407 236327 675887 236383 6 mprj_io_in[3]
port 170 nsew signal tristate
rlabel metal2 s 675407 251047 675887 251103 6 mprj_io_in_3v3[3]
port 171 nsew signal tristate
rlabel metal5 s 698512 281640 711002 294180 6 mprj_io[4]
port 172 nsew signal bidirectional
rlabel metal2 s 675407 286203 675887 286259 6 mprj_io_analog_en[4]
port 173 nsew signal input
rlabel metal2 s 675407 287491 675887 287547 6 mprj_io_analog_pol[4]
port 174 nsew signal input
rlabel metal2 s 675407 290527 675887 290583 6 mprj_io_analog_sel[4]
port 175 nsew signal input
rlabel metal2 s 675407 286847 675887 286903 6 mprj_io_dm[12]
port 176 nsew signal input
rlabel metal2 s 675407 285007 675887 285063 6 mprj_io_dm[13]
port 177 nsew signal input
rlabel metal2 s 675407 291171 675887 291227 6 mprj_io_dm[14]
port 178 nsew signal input
rlabel metal2 s 675407 291815 675887 291871 6 mprj_io_holdover[4]
port 179 nsew signal input
rlabel metal2 s 675407 294851 675887 294907 6 mprj_io_ib_mode_sel[4]
port 180 nsew signal input
rlabel metal2 s 675407 288043 675887 288099 6 mprj_io_inp_dis[4]
port 181 nsew signal input
rlabel metal2 s 675407 295495 675887 295551 6 mprj_io_oeb[4]
port 182 nsew signal input
rlabel metal2 s 675407 292367 675887 292423 6 mprj_io_out[4]
port 183 nsew signal input
rlabel metal2 s 675407 283167 675887 283223 6 mprj_io_slow_sel[4]
port 184 nsew signal input
rlabel metal2 s 675407 294207 675887 294263 6 mprj_io_vtrip_sel[4]
port 185 nsew signal input
rlabel metal2 s 675407 281327 675887 281383 6 mprj_io_in[4]
port 186 nsew signal tristate
rlabel metal2 s 675407 296047 675887 296103 6 mprj_io_in_3v3[4]
port 187 nsew signal tristate
rlabel metal5 s 698512 326640 711002 339180 6 mprj_io[5]
port 188 nsew signal bidirectional
rlabel metal2 s 675407 331203 675887 331259 6 mprj_io_analog_en[5]
port 189 nsew signal input
rlabel metal2 s 675407 332491 675887 332547 6 mprj_io_analog_pol[5]
port 190 nsew signal input
rlabel metal2 s 675407 335527 675887 335583 6 mprj_io_analog_sel[5]
port 191 nsew signal input
rlabel metal2 s 675407 331847 675887 331903 6 mprj_io_dm[15]
port 192 nsew signal input
rlabel metal2 s 675407 330007 675887 330063 6 mprj_io_dm[16]
port 193 nsew signal input
rlabel metal2 s 675407 336171 675887 336227 6 mprj_io_dm[17]
port 194 nsew signal input
rlabel metal2 s 675407 336815 675887 336871 6 mprj_io_holdover[5]
port 195 nsew signal input
rlabel metal2 s 675407 339851 675887 339907 6 mprj_io_ib_mode_sel[5]
port 196 nsew signal input
rlabel metal2 s 675407 333043 675887 333099 6 mprj_io_inp_dis[5]
port 197 nsew signal input
rlabel metal2 s 675407 340495 675887 340551 6 mprj_io_oeb[5]
port 198 nsew signal input
rlabel metal2 s 675407 337367 675887 337423 6 mprj_io_out[5]
port 199 nsew signal input
rlabel metal2 s 675407 328167 675887 328223 6 mprj_io_slow_sel[5]
port 200 nsew signal input
rlabel metal2 s 675407 339207 675887 339263 6 mprj_io_vtrip_sel[5]
port 201 nsew signal input
rlabel metal2 s 675407 326327 675887 326383 6 mprj_io_in[5]
port 202 nsew signal tristate
rlabel metal2 s 675407 341047 675887 341103 6 mprj_io_in_3v3[5]
port 203 nsew signal tristate
rlabel metal5 s 698512 371840 711002 384380 6 mprj_io[6]
port 204 nsew signal bidirectional
rlabel metal2 s 675407 376403 675887 376459 6 mprj_io_analog_en[6]
port 205 nsew signal input
rlabel metal2 s 675407 377691 675887 377747 6 mprj_io_analog_pol[6]
port 206 nsew signal input
rlabel metal2 s 675407 380727 675887 380783 6 mprj_io_analog_sel[6]
port 207 nsew signal input
rlabel metal2 s 675407 377047 675887 377103 6 mprj_io_dm[18]
port 208 nsew signal input
rlabel metal2 s 675407 375207 675887 375263 6 mprj_io_dm[19]
port 209 nsew signal input
rlabel metal2 s 675407 381371 675887 381427 6 mprj_io_dm[20]
port 210 nsew signal input
rlabel metal2 s 675407 382015 675887 382071 6 mprj_io_holdover[6]
port 211 nsew signal input
rlabel metal2 s 675407 385051 675887 385107 6 mprj_io_ib_mode_sel[6]
port 212 nsew signal input
rlabel metal2 s 675407 378243 675887 378299 6 mprj_io_inp_dis[6]
port 213 nsew signal input
rlabel metal2 s 675407 385695 675887 385751 6 mprj_io_oeb[6]
port 214 nsew signal input
rlabel metal2 s 675407 382567 675887 382623 6 mprj_io_out[6]
port 215 nsew signal input
rlabel metal2 s 675407 373367 675887 373423 6 mprj_io_slow_sel[6]
port 216 nsew signal input
rlabel metal2 s 675407 384407 675887 384463 6 mprj_io_vtrip_sel[6]
port 217 nsew signal input
rlabel metal2 s 675407 371527 675887 371583 6 mprj_io_in[6]
port 218 nsew signal tristate
rlabel metal2 s 675407 386247 675887 386303 6 mprj_io_in_3v3[6]
port 219 nsew signal tristate
rlabel metal2 s 675407 551211 675887 551267 6 mprj_gpio_analog[0]
port 220 nsew signal bidirectional
rlabel metal2 s 675407 553051 675887 553107 6 mprj_gpio_noesd[0]
port 221 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561580 6 mprj_io[7]
port 222 nsew signal bidirectional
rlabel metal2 s 675407 553603 675887 553659 6 mprj_io_analog_en[7]
port 223 nsew signal input
rlabel metal2 s 675407 554891 675887 554947 6 mprj_io_analog_pol[7]
port 224 nsew signal input
rlabel metal2 s 675407 557927 675887 557983 6 mprj_io_analog_sel[7]
port 225 nsew signal input
rlabel metal2 s 675407 554247 675887 554303 6 mprj_io_dm[21]
port 226 nsew signal input
rlabel metal2 s 675407 552407 675887 552463 6 mprj_io_dm[22]
port 227 nsew signal input
rlabel metal2 s 675407 558571 675887 558627 6 mprj_io_dm[23]
port 228 nsew signal input
rlabel metal2 s 675407 559215 675887 559271 6 mprj_io_holdover[7]
port 229 nsew signal input
rlabel metal2 s 675407 562251 675887 562307 6 mprj_io_ib_mode_sel[7]
port 230 nsew signal input
rlabel metal2 s 675407 555443 675887 555499 6 mprj_io_inp_dis[7]
port 231 nsew signal input
rlabel metal2 s 675407 562895 675887 562951 6 mprj_io_oeb[7]
port 232 nsew signal input
rlabel metal2 s 675407 559767 675887 559823 6 mprj_io_out[7]
port 233 nsew signal input
rlabel metal2 s 675407 550567 675887 550623 6 mprj_io_slow_sel[7]
port 234 nsew signal input
rlabel metal2 s 675407 561607 675887 561663 6 mprj_io_vtrip_sel[7]
port 235 nsew signal input
rlabel metal2 s 675407 548727 675887 548783 6 mprj_io_in[7]
port 236 nsew signal tristate
rlabel metal2 s 675407 563447 675887 563503 6 mprj_io_in_3v3[7]
port 237 nsew signal tristate
rlabel metal2 s 675407 596411 675887 596467 6 mprj_gpio_analog[1]
port 238 nsew signal bidirectional
rlabel metal2 s 675407 598251 675887 598307 6 mprj_gpio_noesd[1]
port 239 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606780 6 mprj_io[8]
port 240 nsew signal bidirectional
rlabel metal2 s 675407 598803 675887 598859 6 mprj_io_analog_en[8]
port 241 nsew signal input
rlabel metal2 s 675407 600091 675887 600147 6 mprj_io_analog_pol[8]
port 242 nsew signal input
rlabel metal2 s 675407 603127 675887 603183 6 mprj_io_analog_sel[8]
port 243 nsew signal input
rlabel metal2 s 675407 599447 675887 599503 6 mprj_io_dm[24]
port 244 nsew signal input
rlabel metal2 s 675407 597607 675887 597663 6 mprj_io_dm[25]
port 245 nsew signal input
rlabel metal2 s 675407 603771 675887 603827 6 mprj_io_dm[26]
port 246 nsew signal input
rlabel metal2 s 675407 604415 675887 604471 6 mprj_io_holdover[8]
port 247 nsew signal input
rlabel metal2 s 675407 607451 675887 607507 6 mprj_io_ib_mode_sel[8]
port 248 nsew signal input
rlabel metal2 s 675407 600643 675887 600699 6 mprj_io_inp_dis[8]
port 249 nsew signal input
rlabel metal2 s 675407 608095 675887 608151 6 mprj_io_oeb[8]
port 250 nsew signal input
rlabel metal2 s 675407 604967 675887 605023 6 mprj_io_out[8]
port 251 nsew signal input
rlabel metal2 s 675407 595767 675887 595823 6 mprj_io_slow_sel[8]
port 252 nsew signal input
rlabel metal2 s 675407 606807 675887 606863 6 mprj_io_vtrip_sel[8]
port 253 nsew signal input
rlabel metal2 s 675407 593927 675887 593983 6 mprj_io_in[8]
port 254 nsew signal tristate
rlabel metal2 s 675407 608647 675887 608703 6 mprj_io_in_3v3[8]
port 255 nsew signal tristate
rlabel metal2 s 675407 641411 675887 641467 6 mprj_gpio_analog[2]
port 256 nsew signal bidirectional
rlabel metal2 s 675407 643251 675887 643307 6 mprj_gpio_noesd[2]
port 257 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651780 6 mprj_io[9]
port 258 nsew signal bidirectional
rlabel metal2 s 675407 643803 675887 643859 6 mprj_io_analog_en[9]
port 259 nsew signal input
rlabel metal2 s 675407 645091 675887 645147 6 mprj_io_analog_pol[9]
port 260 nsew signal input
rlabel metal2 s 675407 648127 675887 648183 6 mprj_io_analog_sel[9]
port 261 nsew signal input
rlabel metal2 s 675407 644447 675887 644503 6 mprj_io_dm[27]
port 262 nsew signal input
rlabel metal2 s 675407 642607 675887 642663 6 mprj_io_dm[28]
port 263 nsew signal input
rlabel metal2 s 675407 648771 675887 648827 6 mprj_io_dm[29]
port 264 nsew signal input
rlabel metal2 s 675407 649415 675887 649471 6 mprj_io_holdover[9]
port 265 nsew signal input
rlabel metal2 s 675407 652451 675887 652507 6 mprj_io_ib_mode_sel[9]
port 266 nsew signal input
rlabel metal2 s 675407 645643 675887 645699 6 mprj_io_inp_dis[9]
port 267 nsew signal input
rlabel metal2 s 675407 653095 675887 653151 6 mprj_io_oeb[9]
port 268 nsew signal input
rlabel metal2 s 675407 649967 675887 650023 6 mprj_io_out[9]
port 269 nsew signal input
rlabel metal2 s 675407 640767 675887 640823 6 mprj_io_slow_sel[9]
port 270 nsew signal input
rlabel metal2 s 675407 651807 675887 651863 6 mprj_io_vtrip_sel[9]
port 271 nsew signal input
rlabel metal2 s 675407 638927 675887 638983 6 mprj_io_in[9]
port 272 nsew signal tristate
rlabel metal2 s 675407 653647 675887 653703 6 mprj_io_in_3v3[9]
port 273 nsew signal tristate
rlabel metal2 s 41713 796933 42193 796989 6 mprj_gpio_analog[7]
port 274 nsew signal bidirectional
rlabel metal2 s 41713 795093 42193 795149 6 mprj_gpio_noesd[7]
port 275 nsew signal bidirectional
rlabel metal5 s 6598 786620 19088 799160 6 mprj_io[25]
port 276 nsew signal bidirectional
rlabel metal2 s 41713 794541 42193 794597 6 mprj_io_analog_en[14]
port 277 nsew signal input
rlabel metal2 s 41713 793253 42193 793309 6 mprj_io_analog_pol[14]
port 278 nsew signal input
rlabel metal2 s 41713 790217 42193 790273 6 mprj_io_analog_sel[14]
port 279 nsew signal input
rlabel metal2 s 41713 793897 42193 793953 6 mprj_io_dm[42]
port 280 nsew signal input
rlabel metal2 s 41713 795737 42193 795793 6 mprj_io_dm[43]
port 281 nsew signal input
rlabel metal2 s 41713 789573 42193 789629 6 mprj_io_dm[44]
port 282 nsew signal input
rlabel metal2 s 41713 788929 42193 788985 6 mprj_io_holdover[14]
port 283 nsew signal input
rlabel metal2 s 41713 785893 42193 785949 6 mprj_io_ib_mode_sel[14]
port 284 nsew signal input
rlabel metal2 s 41713 792701 42193 792757 6 mprj_io_inp_dis[14]
port 285 nsew signal input
rlabel metal2 s 41713 785249 42193 785305 6 mprj_io_oeb[14]
port 286 nsew signal input
rlabel metal2 s 41713 788377 42193 788433 6 mprj_io_out[14]
port 287 nsew signal input
rlabel metal2 s 41713 797577 42193 797633 6 mprj_io_slow_sel[14]
port 288 nsew signal input
rlabel metal2 s 41713 786537 42193 786593 6 mprj_io_vtrip_sel[14]
port 289 nsew signal input
rlabel metal2 s 41713 799417 42193 799473 6 mprj_io_in[14]
port 290 nsew signal tristate
rlabel metal2 s 41713 784697 42193 784753 6 mprj_io_in_3v3[14]
port 291 nsew signal tristate
rlabel metal2 s 41713 280533 42193 280589 6 mprj_gpio_analog[17]
port 292 nsew signal bidirectional
rlabel metal2 s 41713 278693 42193 278749 6 mprj_gpio_noesd[17]
port 293 nsew signal bidirectional
rlabel metal5 s 6598 270220 19088 282760 6 mprj_io[35]
port 294 nsew signal bidirectional
rlabel metal2 s 41713 278141 42193 278197 6 mprj_io_analog_en[24]
port 295 nsew signal input
rlabel metal2 s 41713 276853 42193 276909 6 mprj_io_analog_pol[24]
port 296 nsew signal input
rlabel metal2 s 41713 273817 42193 273873 6 mprj_io_analog_sel[24]
port 297 nsew signal input
rlabel metal2 s 41713 277497 42193 277553 6 mprj_io_dm[72]
port 298 nsew signal input
rlabel metal2 s 41713 279337 42193 279393 6 mprj_io_dm[73]
port 299 nsew signal input
rlabel metal2 s 41713 273173 42193 273229 6 mprj_io_dm[74]
port 300 nsew signal input
rlabel metal2 s 41713 272529 42193 272585 6 mprj_io_holdover[24]
port 301 nsew signal input
rlabel metal2 s 41713 269493 42193 269549 6 mprj_io_ib_mode_sel[24]
port 302 nsew signal input
rlabel metal2 s 41713 276301 42193 276357 6 mprj_io_inp_dis[24]
port 303 nsew signal input
rlabel metal2 s 41713 268849 42193 268905 6 mprj_io_oeb[24]
port 304 nsew signal input
rlabel metal2 s 41713 271977 42193 272033 6 mprj_io_out[24]
port 305 nsew signal input
rlabel metal2 s 41713 281177 42193 281233 6 mprj_io_slow_sel[24]
port 306 nsew signal input
rlabel metal2 s 41713 270137 42193 270193 6 mprj_io_vtrip_sel[24]
port 307 nsew signal input
rlabel metal2 s 41713 283017 42193 283073 6 mprj_io_in[24]
port 308 nsew signal tristate
rlabel metal2 s 41713 268297 42193 268353 6 mprj_io_in_3v3[24]
port 309 nsew signal tristate
rlabel metal5 s 6598 227020 19088 239560 6 mprj_io[36]
port 310 nsew signal bidirectional
rlabel metal2 s 41713 234941 42193 234997 6 mprj_io_analog_en[25]
port 311 nsew signal input
rlabel metal2 s 41713 233653 42193 233709 6 mprj_io_analog_pol[25]
port 312 nsew signal input
rlabel metal2 s 41713 230617 42193 230673 6 mprj_io_analog_sel[25]
port 313 nsew signal input
rlabel metal2 s 41713 234297 42193 234353 6 mprj_io_dm[75]
port 314 nsew signal input
rlabel metal2 s 41713 236137 42193 236193 6 mprj_io_dm[76]
port 315 nsew signal input
rlabel metal2 s 41713 229973 42193 230029 6 mprj_io_dm[77]
port 316 nsew signal input
rlabel metal2 s 41713 229329 42193 229385 6 mprj_io_holdover[25]
port 317 nsew signal input
rlabel metal2 s 41713 226293 42193 226349 6 mprj_io_ib_mode_sel[25]
port 318 nsew signal input
rlabel metal2 s 41713 233101 42193 233157 6 mprj_io_inp_dis[25]
port 319 nsew signal input
rlabel metal2 s 41713 225649 42193 225705 6 mprj_io_oeb[25]
port 320 nsew signal input
rlabel metal2 s 41713 228777 42193 228833 6 mprj_io_out[25]
port 321 nsew signal input
rlabel metal2 s 41713 237977 42193 238033 6 mprj_io_slow_sel[25]
port 322 nsew signal input
rlabel metal2 s 41713 226937 42193 226993 6 mprj_io_vtrip_sel[25]
port 323 nsew signal input
rlabel metal2 s 41713 239817 42193 239873 6 mprj_io_in[25]
port 324 nsew signal tristate
rlabel metal2 s 41713 225097 42193 225153 6 mprj_io_in_3v3[25]
port 325 nsew signal tristate
rlabel metal5 s 6598 183820 19088 196360 6 mprj_io[37]
port 326 nsew signal bidirectional
rlabel metal2 s 41713 191741 42193 191797 6 mprj_io_analog_en[26]
port 327 nsew signal input
rlabel metal2 s 41713 190453 42193 190509 6 mprj_io_analog_pol[26]
port 328 nsew signal input
rlabel metal2 s 41713 187417 42193 187473 6 mprj_io_analog_sel[26]
port 329 nsew signal input
rlabel metal2 s 41713 191097 42193 191153 6 mprj_io_dm[78]
port 330 nsew signal input
rlabel metal2 s 41713 192937 42193 192993 6 mprj_io_dm[79]
port 331 nsew signal input
rlabel metal2 s 41713 186773 42193 186829 6 mprj_io_dm[80]
port 332 nsew signal input
rlabel metal2 s 41713 186129 42193 186185 6 mprj_io_holdover[26]
port 333 nsew signal input
rlabel metal2 s 41713 183093 42193 183149 6 mprj_io_ib_mode_sel[26]
port 334 nsew signal input
rlabel metal2 s 41713 189901 42193 189957 6 mprj_io_inp_dis[26]
port 335 nsew signal input
rlabel metal2 s 41713 182449 42193 182505 6 mprj_io_oeb[26]
port 336 nsew signal input
rlabel metal2 s 41713 185577 42193 185633 6 mprj_io_out[26]
port 337 nsew signal input
rlabel metal2 s 41713 194777 42193 194833 6 mprj_io_slow_sel[26]
port 338 nsew signal input
rlabel metal2 s 41713 183737 42193 183793 6 mprj_io_vtrip_sel[26]
port 339 nsew signal input
rlabel metal2 s 41713 196617 42193 196673 6 mprj_io_in[26]
port 340 nsew signal tristate
rlabel metal2 s 41713 181897 42193 181953 6 mprj_io_in_3v3[26]
port 341 nsew signal tristate
rlabel metal2 s 41713 753733 42193 753789 6 mprj_gpio_analog[8]
port 342 nsew signal bidirectional
rlabel metal2 s 41713 751893 42193 751949 6 mprj_gpio_noesd[8]
port 343 nsew signal bidirectional
rlabel metal5 s 6598 743420 19088 755960 6 mprj_io[26]
port 344 nsew signal bidirectional
rlabel metal2 s 41713 751341 42193 751397 6 mprj_io_analog_en[15]
port 345 nsew signal input
rlabel metal2 s 41713 750053 42193 750109 6 mprj_io_analog_pol[15]
port 346 nsew signal input
rlabel metal2 s 41713 747017 42193 747073 6 mprj_io_analog_sel[15]
port 347 nsew signal input
rlabel metal2 s 41713 750697 42193 750753 6 mprj_io_dm[45]
port 348 nsew signal input
rlabel metal2 s 41713 752537 42193 752593 6 mprj_io_dm[46]
port 349 nsew signal input
rlabel metal2 s 41713 746373 42193 746429 6 mprj_io_dm[47]
port 350 nsew signal input
rlabel metal2 s 41713 745729 42193 745785 6 mprj_io_holdover[15]
port 351 nsew signal input
rlabel metal2 s 41713 742693 42193 742749 6 mprj_io_ib_mode_sel[15]
port 352 nsew signal input
rlabel metal2 s 41713 749501 42193 749557 6 mprj_io_inp_dis[15]
port 353 nsew signal input
rlabel metal2 s 41713 742049 42193 742105 6 mprj_io_oeb[15]
port 354 nsew signal input
rlabel metal2 s 41713 745177 42193 745233 6 mprj_io_out[15]
port 355 nsew signal input
rlabel metal2 s 41713 754377 42193 754433 6 mprj_io_slow_sel[15]
port 356 nsew signal input
rlabel metal2 s 41713 743337 42193 743393 6 mprj_io_vtrip_sel[15]
port 357 nsew signal input
rlabel metal2 s 41713 756217 42193 756273 6 mprj_io_in[15]
port 358 nsew signal tristate
rlabel metal2 s 41713 741497 42193 741553 6 mprj_io_in_3v3[15]
port 359 nsew signal tristate
rlabel metal2 s 41713 710533 42193 710589 6 mprj_gpio_analog[9]
port 360 nsew signal bidirectional
rlabel metal2 s 41713 708693 42193 708749 6 mprj_gpio_noesd[9]
port 361 nsew signal bidirectional
rlabel metal5 s 6598 700220 19088 712760 6 mprj_io[27]
port 362 nsew signal bidirectional
rlabel metal2 s 41713 708141 42193 708197 6 mprj_io_analog_en[16]
port 363 nsew signal input
rlabel metal2 s 41713 706853 42193 706909 6 mprj_io_analog_pol[16]
port 364 nsew signal input
rlabel metal2 s 41713 703817 42193 703873 6 mprj_io_analog_sel[16]
port 365 nsew signal input
rlabel metal2 s 41713 707497 42193 707553 6 mprj_io_dm[48]
port 366 nsew signal input
rlabel metal2 s 41713 709337 42193 709393 6 mprj_io_dm[49]
port 367 nsew signal input
rlabel metal2 s 41713 703173 42193 703229 6 mprj_io_dm[50]
port 368 nsew signal input
rlabel metal2 s 41713 702529 42193 702585 6 mprj_io_holdover[16]
port 369 nsew signal input
rlabel metal2 s 41713 699493 42193 699549 6 mprj_io_ib_mode_sel[16]
port 370 nsew signal input
rlabel metal2 s 41713 706301 42193 706357 6 mprj_io_inp_dis[16]
port 371 nsew signal input
rlabel metal2 s 41713 698849 42193 698905 6 mprj_io_oeb[16]
port 372 nsew signal input
rlabel metal2 s 41713 701977 42193 702033 6 mprj_io_out[16]
port 373 nsew signal input
rlabel metal2 s 41713 711177 42193 711233 6 mprj_io_slow_sel[16]
port 374 nsew signal input
rlabel metal2 s 41713 700137 42193 700193 6 mprj_io_vtrip_sel[16]
port 375 nsew signal input
rlabel metal2 s 41713 713017 42193 713073 6 mprj_io_in[16]
port 376 nsew signal tristate
rlabel metal2 s 41713 698297 42193 698353 6 mprj_io_in_3v3[16]
port 377 nsew signal tristate
rlabel metal2 s 41713 667333 42193 667389 6 mprj_gpio_analog[10]
port 378 nsew signal bidirectional
rlabel metal2 s 41713 665493 42193 665549 6 mprj_gpio_noesd[10]
port 379 nsew signal bidirectional
rlabel metal5 s 6598 657020 19088 669560 6 mprj_io[28]
port 380 nsew signal bidirectional
rlabel metal2 s 41713 664941 42193 664997 6 mprj_io_analog_en[17]
port 381 nsew signal input
rlabel metal2 s 41713 663653 42193 663709 6 mprj_io_analog_pol[17]
port 382 nsew signal input
rlabel metal2 s 41713 660617 42193 660673 6 mprj_io_analog_sel[17]
port 383 nsew signal input
rlabel metal2 s 41713 664297 42193 664353 6 mprj_io_dm[51]
port 384 nsew signal input
rlabel metal2 s 41713 666137 42193 666193 6 mprj_io_dm[52]
port 385 nsew signal input
rlabel metal2 s 41713 659973 42193 660029 6 mprj_io_dm[53]
port 386 nsew signal input
rlabel metal2 s 41713 659329 42193 659385 6 mprj_io_holdover[17]
port 387 nsew signal input
rlabel metal2 s 41713 656293 42193 656349 6 mprj_io_ib_mode_sel[17]
port 388 nsew signal input
rlabel metal2 s 41713 663101 42193 663157 6 mprj_io_inp_dis[17]
port 389 nsew signal input
rlabel metal2 s 41713 655649 42193 655705 6 mprj_io_oeb[17]
port 390 nsew signal input
rlabel metal2 s 41713 658777 42193 658833 6 mprj_io_out[17]
port 391 nsew signal input
rlabel metal2 s 41713 667977 42193 668033 6 mprj_io_slow_sel[17]
port 392 nsew signal input
rlabel metal2 s 41713 656937 42193 656993 6 mprj_io_vtrip_sel[17]
port 393 nsew signal input
rlabel metal2 s 41713 669817 42193 669873 6 mprj_io_in[17]
port 394 nsew signal tristate
rlabel metal2 s 41713 655097 42193 655153 6 mprj_io_in_3v3[17]
port 395 nsew signal tristate
rlabel metal2 s 41713 624133 42193 624189 6 mprj_gpio_analog[11]
port 396 nsew signal bidirectional
rlabel metal2 s 41713 622293 42193 622349 6 mprj_gpio_noesd[11]
port 397 nsew signal bidirectional
rlabel metal5 s 6598 613820 19088 626360 6 mprj_io[29]
port 398 nsew signal bidirectional
rlabel metal2 s 41713 621741 42193 621797 6 mprj_io_analog_en[18]
port 399 nsew signal input
rlabel metal2 s 41713 620453 42193 620509 6 mprj_io_analog_pol[18]
port 400 nsew signal input
rlabel metal2 s 41713 617417 42193 617473 6 mprj_io_analog_sel[18]
port 401 nsew signal input
rlabel metal2 s 41713 621097 42193 621153 6 mprj_io_dm[54]
port 402 nsew signal input
rlabel metal2 s 41713 622937 42193 622993 6 mprj_io_dm[55]
port 403 nsew signal input
rlabel metal2 s 41713 616773 42193 616829 6 mprj_io_dm[56]
port 404 nsew signal input
rlabel metal2 s 41713 616129 42193 616185 6 mprj_io_holdover[18]
port 405 nsew signal input
rlabel metal2 s 41713 613093 42193 613149 6 mprj_io_ib_mode_sel[18]
port 406 nsew signal input
rlabel metal2 s 41713 619901 42193 619957 6 mprj_io_inp_dis[18]
port 407 nsew signal input
rlabel metal2 s 41713 612449 42193 612505 6 mprj_io_oeb[18]
port 408 nsew signal input
rlabel metal2 s 41713 615577 42193 615633 6 mprj_io_out[18]
port 409 nsew signal input
rlabel metal2 s 41713 624777 42193 624833 6 mprj_io_slow_sel[18]
port 410 nsew signal input
rlabel metal2 s 41713 613737 42193 613793 6 mprj_io_vtrip_sel[18]
port 411 nsew signal input
rlabel metal2 s 41713 626617 42193 626673 6 mprj_io_in[18]
port 412 nsew signal tristate
rlabel metal2 s 41713 611897 42193 611953 6 mprj_io_in_3v3[18]
port 413 nsew signal tristate
rlabel metal2 s 41713 580933 42193 580989 6 mprj_gpio_analog[12]
port 414 nsew signal bidirectional
rlabel metal2 s 41713 579093 42193 579149 6 mprj_gpio_noesd[12]
port 415 nsew signal bidirectional
rlabel metal5 s 6598 570620 19088 583160 6 mprj_io[30]
port 416 nsew signal bidirectional
rlabel metal2 s 41713 578541 42193 578597 6 mprj_io_analog_en[19]
port 417 nsew signal input
rlabel metal2 s 41713 577253 42193 577309 6 mprj_io_analog_pol[19]
port 418 nsew signal input
rlabel metal2 s 41713 574217 42193 574273 6 mprj_io_analog_sel[19]
port 419 nsew signal input
rlabel metal2 s 41713 577897 42193 577953 6 mprj_io_dm[57]
port 420 nsew signal input
rlabel metal2 s 41713 579737 42193 579793 6 mprj_io_dm[58]
port 421 nsew signal input
rlabel metal2 s 41713 573573 42193 573629 6 mprj_io_dm[59]
port 422 nsew signal input
rlabel metal2 s 41713 572929 42193 572985 6 mprj_io_holdover[19]
port 423 nsew signal input
rlabel metal2 s 41713 569893 42193 569949 6 mprj_io_ib_mode_sel[19]
port 424 nsew signal input
rlabel metal2 s 41713 576701 42193 576757 6 mprj_io_inp_dis[19]
port 425 nsew signal input
rlabel metal2 s 41713 569249 42193 569305 6 mprj_io_oeb[19]
port 426 nsew signal input
rlabel metal2 s 41713 572377 42193 572433 6 mprj_io_out[19]
port 427 nsew signal input
rlabel metal2 s 41713 581577 42193 581633 6 mprj_io_slow_sel[19]
port 428 nsew signal input
rlabel metal2 s 41713 570537 42193 570593 6 mprj_io_vtrip_sel[19]
port 429 nsew signal input
rlabel metal2 s 41713 583417 42193 583473 6 mprj_io_in[19]
port 430 nsew signal tristate
rlabel metal2 s 41713 568697 42193 568753 6 mprj_io_in_3v3[19]
port 431 nsew signal tristate
rlabel metal2 s 41713 537733 42193 537789 6 mprj_gpio_analog[13]
port 432 nsew signal bidirectional
rlabel metal2 s 41713 535893 42193 535949 6 mprj_gpio_noesd[13]
port 433 nsew signal bidirectional
rlabel metal5 s 6598 527420 19088 539960 6 mprj_io[31]
port 434 nsew signal bidirectional
rlabel metal2 s 41713 535341 42193 535397 6 mprj_io_analog_en[20]
port 435 nsew signal input
rlabel metal2 s 41713 534053 42193 534109 6 mprj_io_analog_pol[20]
port 436 nsew signal input
rlabel metal2 s 41713 531017 42193 531073 6 mprj_io_analog_sel[20]
port 437 nsew signal input
rlabel metal2 s 41713 534697 42193 534753 6 mprj_io_dm[60]
port 438 nsew signal input
rlabel metal2 s 41713 536537 42193 536593 6 mprj_io_dm[61]
port 439 nsew signal input
rlabel metal2 s 41713 530373 42193 530429 6 mprj_io_dm[62]
port 440 nsew signal input
rlabel metal2 s 41713 529729 42193 529785 6 mprj_io_holdover[20]
port 441 nsew signal input
rlabel metal2 s 41713 526693 42193 526749 6 mprj_io_ib_mode_sel[20]
port 442 nsew signal input
rlabel metal2 s 41713 533501 42193 533557 6 mprj_io_inp_dis[20]
port 443 nsew signal input
rlabel metal2 s 41713 526049 42193 526105 6 mprj_io_oeb[20]
port 444 nsew signal input
rlabel metal2 s 41713 529177 42193 529233 6 mprj_io_out[20]
port 445 nsew signal input
rlabel metal2 s 41713 538377 42193 538433 6 mprj_io_slow_sel[20]
port 446 nsew signal input
rlabel metal2 s 41713 527337 42193 527393 6 mprj_io_vtrip_sel[20]
port 447 nsew signal input
rlabel metal2 s 41713 540217 42193 540273 6 mprj_io_in[20]
port 448 nsew signal tristate
rlabel metal2 s 41713 525497 42193 525553 6 mprj_io_in_3v3[20]
port 449 nsew signal tristate
rlabel metal2 s 41713 410133 42193 410189 6 mprj_gpio_analog[14]
port 450 nsew signal bidirectional
rlabel metal2 s 41713 408293 42193 408349 6 mprj_gpio_noesd[14]
port 451 nsew signal bidirectional
rlabel metal5 s 6598 399820 19088 412360 6 mprj_io[32]
port 452 nsew signal bidirectional
rlabel metal2 s 41713 407741 42193 407797 6 mprj_io_analog_en[21]
port 453 nsew signal input
rlabel metal2 s 41713 406453 42193 406509 6 mprj_io_analog_pol[21]
port 454 nsew signal input
rlabel metal2 s 41713 403417 42193 403473 6 mprj_io_analog_sel[21]
port 455 nsew signal input
rlabel metal2 s 41713 407097 42193 407153 6 mprj_io_dm[63]
port 456 nsew signal input
rlabel metal2 s 41713 408937 42193 408993 6 mprj_io_dm[64]
port 457 nsew signal input
rlabel metal2 s 41713 402773 42193 402829 6 mprj_io_dm[65]
port 458 nsew signal input
rlabel metal2 s 41713 402129 42193 402185 6 mprj_io_holdover[21]
port 459 nsew signal input
rlabel metal2 s 41713 399093 42193 399149 6 mprj_io_ib_mode_sel[21]
port 460 nsew signal input
rlabel metal2 s 41713 405901 42193 405957 6 mprj_io_inp_dis[21]
port 461 nsew signal input
rlabel metal2 s 41713 398449 42193 398505 6 mprj_io_oeb[21]
port 462 nsew signal input
rlabel metal2 s 41713 401577 42193 401633 6 mprj_io_out[21]
port 463 nsew signal input
rlabel metal2 s 41713 410777 42193 410833 6 mprj_io_slow_sel[21]
port 464 nsew signal input
rlabel metal2 s 41713 399737 42193 399793 6 mprj_io_vtrip_sel[21]
port 465 nsew signal input
rlabel metal2 s 41713 412617 42193 412673 6 mprj_io_in[21]
port 466 nsew signal tristate
rlabel metal2 s 41713 397897 42193 397953 6 mprj_io_in_3v3[21]
port 467 nsew signal tristate
rlabel metal2 s 41713 366933 42193 366989 6 mprj_gpio_analog[15]
port 468 nsew signal bidirectional
rlabel metal2 s 41713 365093 42193 365149 6 mprj_gpio_noesd[15]
port 469 nsew signal bidirectional
rlabel metal5 s 6598 356620 19088 369160 6 mprj_io[33]
port 470 nsew signal bidirectional
rlabel metal2 s 41713 364541 42193 364597 6 mprj_io_analog_en[22]
port 471 nsew signal input
rlabel metal2 s 41713 363253 42193 363309 6 mprj_io_analog_pol[22]
port 472 nsew signal input
rlabel metal2 s 41713 360217 42193 360273 6 mprj_io_analog_sel[22]
port 473 nsew signal input
rlabel metal2 s 41713 363897 42193 363953 6 mprj_io_dm[66]
port 474 nsew signal input
rlabel metal2 s 41713 365737 42193 365793 6 mprj_io_dm[67]
port 475 nsew signal input
rlabel metal2 s 41713 359573 42193 359629 6 mprj_io_dm[68]
port 476 nsew signal input
rlabel metal2 s 41713 358929 42193 358985 6 mprj_io_holdover[22]
port 477 nsew signal input
rlabel metal2 s 41713 355893 42193 355949 6 mprj_io_ib_mode_sel[22]
port 478 nsew signal input
rlabel metal2 s 41713 362701 42193 362757 6 mprj_io_inp_dis[22]
port 479 nsew signal input
rlabel metal2 s 41713 355249 42193 355305 6 mprj_io_oeb[22]
port 480 nsew signal input
rlabel metal2 s 41713 358377 42193 358433 6 mprj_io_out[22]
port 481 nsew signal input
rlabel metal2 s 41713 367577 42193 367633 6 mprj_io_slow_sel[22]
port 482 nsew signal input
rlabel metal2 s 41713 356537 42193 356593 6 mprj_io_vtrip_sel[22]
port 483 nsew signal input
rlabel metal2 s 41713 369417 42193 369473 6 mprj_io_in[22]
port 484 nsew signal tristate
rlabel metal2 s 41713 354697 42193 354753 6 mprj_io_in_3v3[22]
port 485 nsew signal tristate
rlabel metal2 s 41713 323733 42193 323789 6 mprj_gpio_analog[16]
port 486 nsew signal bidirectional
rlabel metal2 s 41713 321893 42193 321949 6 mprj_gpio_noesd[16]
port 487 nsew signal bidirectional
rlabel metal5 s 6598 313420 19088 325960 6 mprj_io[34]
port 488 nsew signal bidirectional
rlabel metal2 s 41713 321341 42193 321397 6 mprj_io_analog_en[23]
port 489 nsew signal input
rlabel metal2 s 41713 320053 42193 320109 6 mprj_io_analog_pol[23]
port 490 nsew signal input
rlabel metal2 s 41713 317017 42193 317073 6 mprj_io_analog_sel[23]
port 491 nsew signal input
rlabel metal2 s 41713 320697 42193 320753 6 mprj_io_dm[69]
port 492 nsew signal input
rlabel metal2 s 41713 322537 42193 322593 6 mprj_io_dm[70]
port 493 nsew signal input
rlabel metal2 s 41713 316373 42193 316429 6 mprj_io_dm[71]
port 494 nsew signal input
rlabel metal2 s 41713 315729 42193 315785 6 mprj_io_holdover[23]
port 495 nsew signal input
rlabel metal2 s 41713 312693 42193 312749 6 mprj_io_ib_mode_sel[23]
port 496 nsew signal input
rlabel metal2 s 41713 319501 42193 319557 6 mprj_io_inp_dis[23]
port 497 nsew signal input
rlabel metal2 s 41713 312049 42193 312105 6 mprj_io_oeb[23]
port 498 nsew signal input
rlabel metal2 s 41713 315177 42193 315233 6 mprj_io_out[23]
port 499 nsew signal input
rlabel metal2 s 41713 324377 42193 324433 6 mprj_io_slow_sel[23]
port 500 nsew signal input
rlabel metal2 s 41713 313337 42193 313393 6 mprj_io_vtrip_sel[23]
port 501 nsew signal input
rlabel metal2 s 41713 326217 42193 326273 6 mprj_io_in[23]
port 502 nsew signal tristate
rlabel metal2 s 41713 311497 42193 311553 6 mprj_io_in_3v3[23]
port 503 nsew signal tristate
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 504 nsew signal input
rlabel metal5 s 136713 7143 144149 18309 6 resetb
port 505 nsew signal input
rlabel metal3 s 141667 38031 141813 39999 6 resetb_core_h
port 506 nsew signal tristate
rlabel metal4 s 132600 36323 132792 37013 6 vdda
port 507 nsew signal bidirectional
rlabel metal4 s 132600 28653 147600 28719 6 vssa
port 508 nsew signal bidirectional
rlabel metal4 s 132600 30762 132868 31674 6 vssd
port 509 nsew signal bidirectional
rlabel metal3 s 677600 958656 694070 963656 6 mprj_analog[0]
port 510 nsew signal bidirectional
rlabel metal5 s 698624 955022 710788 967190 6 mprj_io[15]
port 511 nsew signal bidirectional
rlabel metal3 s 631944 997600 636944 1014070 6 mprj_analog[1]
port 512 nsew signal bidirectional
rlabel metal5 s 628410 1018624 640578 1030788 6 mprj_io[16]
port 513 nsew signal bidirectional
rlabel metal3 s 530144 997600 535144 1014070 6 mprj_analog[2]
port 514 nsew signal bidirectional
rlabel metal5 s 526610 1018624 538778 1030788 6 mprj_io[17]
port 515 nsew signal bidirectional
rlabel metal3 s 478744 997600 483744 1014070 6 mprj_analog[3]
port 516 nsew signal bidirectional
rlabel metal5 s 475210 1018624 487378 1030788 6 mprj_io[18]
port 517 nsew signal bidirectional
rlabel metal3 s 393878 997600 408200 1000736 6 mprj_analog[4]
port 518 nsew signal bidirectional
rlabel metal2 s 393878 997600 398658 1002732 6 mprj_clamp_high[0]
port 519 nsew signal input
rlabel metal2 s 383899 997600 388679 998010 6 mprj_clamp_low[0]
port 520 nsew signal input
rlabel metal5 s 385210 1018624 397378 1030788 6 mprj_io[14]
port 521 nsew signal bidirectional
rlabel metal5 s 697980 909666 711432 920546 6 vccd1_pad
port 522 nsew signal bidirectional
rlabel metal5 s 698624 819822 710788 831990 6 vdda1_pad
port 523 nsew signal bidirectional
rlabel metal5 s 698624 505222 710788 517390 6 vdda1_pad2
port 524 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030788 6 vssa1_pad
port 525 nsew signal bidirectional
rlabel metal5 s 698624 417022 710788 429190 6 vssa1_pad2
port 526 nsew signal bidirectional
rlabel metal4 s 679377 459800 680307 460054 6 vccd1
port 527 nsew signal bidirectional
rlabel metal4 s 680587 459800 681277 459992 6 vdda1
port 528 nsew signal bidirectional
rlabel metal4 s 688881 459800 688947 474800 6 vssa1
port 529 nsew signal bidirectional
rlabel metal3 s 678000 469900 685920 474700 6 vssd1
port 530 nsew signal bidirectional
rlabel metal5 s 697980 461866 711432 472746 6 vssd1_pad
port 531 nsew signal bidirectional
rlabel metal3 s 184944 997600 189944 1014070 6 mprj_analog[7]
port 532 nsew signal bidirectional
rlabel metal5 s 181410 1018624 193578 1030788 6 mprj_io[21]
port 533 nsew signal bidirectional
rlabel metal3 s 133544 997600 138544 1014070 6 mprj_analog[8]
port 534 nsew signal bidirectional
rlabel metal5 s 130010 1018624 142178 1030788 6 mprj_io[22]
port 535 nsew signal bidirectional
rlabel metal3 s 82144 997600 87144 1014070 6 mprj_analog[9]
port 536 nsew signal bidirectional
rlabel metal5 s 78610 1018624 90778 1030788 6 mprj_io[23]
port 537 nsew signal bidirectional
rlabel metal3 s 23530 960144 40000 965144 6 mprj_analog[10]
port 538 nsew signal bidirectional
rlabel metal5 s 6811 956610 18975 968778 6 mprj_io[24]
port 539 nsew signal bidirectional
rlabel metal3 s 292078 997600 306400 1000736 6 mprj_analog[5]
port 540 nsew signal bidirectional
rlabel metal2 s 292078 997600 296858 1002732 6 mprj_clamp_high[1]
port 541 nsew signal input
rlabel metal2 s 282099 997600 286879 998010 6 mprj_clamp_low[1]
port 542 nsew signal input
rlabel metal5 s 283410 1018624 295578 1030788 6 mprj_io[19]
port 543 nsew signal bidirectional
rlabel metal3 s 240478 997600 254800 1000736 6 mprj_analog[6]
port 544 nsew signal bidirectional
rlabel metal2 s 240478 997600 245258 1002732 6 mprj_clamp_high[2]
port 545 nsew signal input
rlabel metal2 s 230499 997600 235279 998010 6 mprj_clamp_low[2]
port 546 nsew signal input
rlabel metal5 s 231810 1018624 243978 1030788 6 mprj_io[20]
port 547 nsew signal bidirectional
rlabel metal5 s 6167 914054 19619 924934 6 vccd2_pad
port 548 nsew signal bidirectional
rlabel metal5 s 6811 484410 18975 496578 6 vdda2_pad
port 549 nsew signal bidirectional
rlabel metal5 s 6811 829010 18975 841178 6 vssa2_pad
port 550 nsew signal bidirectional
rlabel metal4 s 38503 455546 39593 455800 6 vccd
port 551 nsew signal bidirectional
rlabel metal4 s 37293 455546 38223 455800 6 vccd2
port 552 nsew signal bidirectional
rlabel metal4 s 36323 455607 37013 455799 6 vdda2
port 553 nsew signal bidirectional
rlabel metal4 s 32933 455546 33623 455800 6 vddio
port 554 nsew signal bidirectional
rlabel metal4 s 28653 440800 28719 455800 6 vssa2
port 555 nsew signal bidirectional
rlabel metal3 s 31680 440900 39600 445700 6 vssd2
port 556 nsew signal bidirectional
rlabel metal5 s 6167 442854 19619 453734 6 vssd2_pad
port 557 nsew signal bidirectional
rlabel metal4 s 7 455645 4843 456093 6 vssio
port 558 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
