VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_protect
  CLASS BLOCK ;
  FOREIGN mgmt_protect ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 90.000 ;
  PIN caravel_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 15.000 0.300 15.600 ;
    END
  END caravel_clk
  PIN caravel_clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 44.920 0.300 45.520 ;
    END
  END caravel_clk2
  PIN caravel_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 74.840 0.300 75.440 ;
    END
  END caravel_rstn
  PIN la_data_in_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 89.700 9.570 92.000 ;
    END
  END la_data_in_core[0]
  PIN la_data_in_core[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 89.700 227.610 92.000 ;
    END
  END la_data_in_core[100]
  PIN la_data_in_core[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 89.700 229.910 92.000 ;
    END
  END la_data_in_core[101]
  PIN la_data_in_core[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 89.700 232.210 92.000 ;
    END
  END la_data_in_core[102]
  PIN la_data_in_core[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 89.700 234.050 92.000 ;
    END
  END la_data_in_core[103]
  PIN la_data_in_core[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 89.700 236.350 92.000 ;
    END
  END la_data_in_core[104]
  PIN la_data_in_core[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 89.700 238.650 92.000 ;
    END
  END la_data_in_core[105]
  PIN la_data_in_core[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 89.700 240.950 92.000 ;
    END
  END la_data_in_core[106]
  PIN la_data_in_core[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 89.700 242.790 92.000 ;
    END
  END la_data_in_core[107]
  PIN la_data_in_core[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 89.700 245.090 92.000 ;
    END
  END la_data_in_core[108]
  PIN la_data_in_core[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 89.700 247.390 92.000 ;
    END
  END la_data_in_core[109]
  PIN la_data_in_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 89.700 31.650 92.000 ;
    END
  END la_data_in_core[10]
  PIN la_data_in_core[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 89.700 249.230 92.000 ;
    END
  END la_data_in_core[110]
  PIN la_data_in_core[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 89.700 251.530 92.000 ;
    END
  END la_data_in_core[111]
  PIN la_data_in_core[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 89.700 253.830 92.000 ;
    END
  END la_data_in_core[112]
  PIN la_data_in_core[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 89.700 256.130 92.000 ;
    END
  END la_data_in_core[113]
  PIN la_data_in_core[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 89.700 257.970 92.000 ;
    END
  END la_data_in_core[114]
  PIN la_data_in_core[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 89.700 260.270 92.000 ;
    END
  END la_data_in_core[115]
  PIN la_data_in_core[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 89.700 262.570 92.000 ;
    END
  END la_data_in_core[116]
  PIN la_data_in_core[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 89.700 264.870 92.000 ;
    END
  END la_data_in_core[117]
  PIN la_data_in_core[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 89.700 266.710 92.000 ;
    END
  END la_data_in_core[118]
  PIN la_data_in_core[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 89.700 269.010 92.000 ;
    END
  END la_data_in_core[119]
  PIN la_data_in_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 89.700 33.950 92.000 ;
    END
  END la_data_in_core[11]
  PIN la_data_in_core[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 89.700 271.310 92.000 ;
    END
  END la_data_in_core[120]
  PIN la_data_in_core[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 89.700 273.610 92.000 ;
    END
  END la_data_in_core[121]
  PIN la_data_in_core[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 89.700 275.450 92.000 ;
    END
  END la_data_in_core[122]
  PIN la_data_in_core[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 89.700 277.750 92.000 ;
    END
  END la_data_in_core[123]
  PIN la_data_in_core[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 89.700 280.050 92.000 ;
    END
  END la_data_in_core[124]
  PIN la_data_in_core[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 89.700 281.890 92.000 ;
    END
  END la_data_in_core[125]
  PIN la_data_in_core[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 89.700 284.190 92.000 ;
    END
  END la_data_in_core[126]
  PIN la_data_in_core[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 89.700 286.490 92.000 ;
    END
  END la_data_in_core[127]
  PIN la_data_in_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 89.700 35.790 92.000 ;
    END
  END la_data_in_core[12]
  PIN la_data_in_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 89.700 38.090 92.000 ;
    END
  END la_data_in_core[13]
  PIN la_data_in_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 89.700 40.390 92.000 ;
    END
  END la_data_in_core[14]
  PIN la_data_in_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 89.700 42.230 92.000 ;
    END
  END la_data_in_core[15]
  PIN la_data_in_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 89.700 44.530 92.000 ;
    END
  END la_data_in_core[16]
  PIN la_data_in_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 89.700 46.830 92.000 ;
    END
  END la_data_in_core[17]
  PIN la_data_in_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 89.700 49.130 92.000 ;
    END
  END la_data_in_core[18]
  PIN la_data_in_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 89.700 50.970 92.000 ;
    END
  END la_data_in_core[19]
  PIN la_data_in_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 89.700 11.870 92.000 ;
    END
  END la_data_in_core[1]
  PIN la_data_in_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 89.700 53.270 92.000 ;
    END
  END la_data_in_core[20]
  PIN la_data_in_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 89.700 55.570 92.000 ;
    END
  END la_data_in_core[21]
  PIN la_data_in_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 89.700 57.870 92.000 ;
    END
  END la_data_in_core[22]
  PIN la_data_in_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 89.700 59.710 92.000 ;
    END
  END la_data_in_core[23]
  PIN la_data_in_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 89.700 62.010 92.000 ;
    END
  END la_data_in_core[24]
  PIN la_data_in_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 89.700 64.310 92.000 ;
    END
  END la_data_in_core[25]
  PIN la_data_in_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 89.700 66.610 92.000 ;
    END
  END la_data_in_core[26]
  PIN la_data_in_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 89.700 68.450 92.000 ;
    END
  END la_data_in_core[27]
  PIN la_data_in_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 89.700 70.750 92.000 ;
    END
  END la_data_in_core[28]
  PIN la_data_in_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 89.700 73.050 92.000 ;
    END
  END la_data_in_core[29]
  PIN la_data_in_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 89.700 14.170 92.000 ;
    END
  END la_data_in_core[2]
  PIN la_data_in_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 89.700 75.350 92.000 ;
    END
  END la_data_in_core[30]
  PIN la_data_in_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 89.700 77.190 92.000 ;
    END
  END la_data_in_core[31]
  PIN la_data_in_core[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 89.700 79.490 92.000 ;
    END
  END la_data_in_core[32]
  PIN la_data_in_core[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 89.700 81.790 92.000 ;
    END
  END la_data_in_core[33]
  PIN la_data_in_core[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 89.700 83.630 92.000 ;
    END
  END la_data_in_core[34]
  PIN la_data_in_core[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 89.700 85.930 92.000 ;
    END
  END la_data_in_core[35]
  PIN la_data_in_core[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 89.700 88.230 92.000 ;
    END
  END la_data_in_core[36]
  PIN la_data_in_core[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 89.700 90.530 92.000 ;
    END
  END la_data_in_core[37]
  PIN la_data_in_core[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 89.700 92.370 92.000 ;
    END
  END la_data_in_core[38]
  PIN la_data_in_core[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 89.700 94.670 92.000 ;
    END
  END la_data_in_core[39]
  PIN la_data_in_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 89.700 16.470 92.000 ;
    END
  END la_data_in_core[3]
  PIN la_data_in_core[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 89.700 96.970 92.000 ;
    END
  END la_data_in_core[40]
  PIN la_data_in_core[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 89.700 99.270 92.000 ;
    END
  END la_data_in_core[41]
  PIN la_data_in_core[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 89.700 101.110 92.000 ;
    END
  END la_data_in_core[42]
  PIN la_data_in_core[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 89.700 103.410 92.000 ;
    END
  END la_data_in_core[43]
  PIN la_data_in_core[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 89.700 105.710 92.000 ;
    END
  END la_data_in_core[44]
  PIN la_data_in_core[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 89.700 108.010 92.000 ;
    END
  END la_data_in_core[45]
  PIN la_data_in_core[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 89.700 109.850 92.000 ;
    END
  END la_data_in_core[46]
  PIN la_data_in_core[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 89.700 112.150 92.000 ;
    END
  END la_data_in_core[47]
  PIN la_data_in_core[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 89.700 114.450 92.000 ;
    END
  END la_data_in_core[48]
  PIN la_data_in_core[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 89.700 116.750 92.000 ;
    END
  END la_data_in_core[49]
  PIN la_data_in_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 89.700 18.310 92.000 ;
    END
  END la_data_in_core[4]
  PIN la_data_in_core[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 89.700 118.590 92.000 ;
    END
  END la_data_in_core[50]
  PIN la_data_in_core[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 89.700 120.890 92.000 ;
    END
  END la_data_in_core[51]
  PIN la_data_in_core[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 89.700 123.190 92.000 ;
    END
  END la_data_in_core[52]
  PIN la_data_in_core[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 89.700 125.030 92.000 ;
    END
  END la_data_in_core[53]
  PIN la_data_in_core[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 89.700 127.330 92.000 ;
    END
  END la_data_in_core[54]
  PIN la_data_in_core[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 89.700 129.630 92.000 ;
    END
  END la_data_in_core[55]
  PIN la_data_in_core[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 89.700 131.930 92.000 ;
    END
  END la_data_in_core[56]
  PIN la_data_in_core[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 89.700 133.770 92.000 ;
    END
  END la_data_in_core[57]
  PIN la_data_in_core[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 89.700 136.070 92.000 ;
    END
  END la_data_in_core[58]
  PIN la_data_in_core[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 89.700 138.370 92.000 ;
    END
  END la_data_in_core[59]
  PIN la_data_in_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 89.700 20.610 92.000 ;
    END
  END la_data_in_core[5]
  PIN la_data_in_core[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 89.700 140.670 92.000 ;
    END
  END la_data_in_core[60]
  PIN la_data_in_core[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 89.700 142.510 92.000 ;
    END
  END la_data_in_core[61]
  PIN la_data_in_core[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 89.700 144.810 92.000 ;
    END
  END la_data_in_core[62]
  PIN la_data_in_core[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 89.700 147.110 92.000 ;
    END
  END la_data_in_core[63]
  PIN la_data_in_core[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 89.700 149.410 92.000 ;
    END
  END la_data_in_core[64]
  PIN la_data_in_core[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 89.700 151.250 92.000 ;
    END
  END la_data_in_core[65]
  PIN la_data_in_core[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 89.700 153.550 92.000 ;
    END
  END la_data_in_core[66]
  PIN la_data_in_core[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 89.700 155.850 92.000 ;
    END
  END la_data_in_core[67]
  PIN la_data_in_core[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 89.700 158.150 92.000 ;
    END
  END la_data_in_core[68]
  PIN la_data_in_core[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 89.700 159.990 92.000 ;
    END
  END la_data_in_core[69]
  PIN la_data_in_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 89.700 22.910 92.000 ;
    END
  END la_data_in_core[6]
  PIN la_data_in_core[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 89.700 162.290 92.000 ;
    END
  END la_data_in_core[70]
  PIN la_data_in_core[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 89.700 164.590 92.000 ;
    END
  END la_data_in_core[71]
  PIN la_data_in_core[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 89.700 166.430 92.000 ;
    END
  END la_data_in_core[72]
  PIN la_data_in_core[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 89.700 168.730 92.000 ;
    END
  END la_data_in_core[73]
  PIN la_data_in_core[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 89.700 171.030 92.000 ;
    END
  END la_data_in_core[74]
  PIN la_data_in_core[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 89.700 173.330 92.000 ;
    END
  END la_data_in_core[75]
  PIN la_data_in_core[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 89.700 175.170 92.000 ;
    END
  END la_data_in_core[76]
  PIN la_data_in_core[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 89.700 177.470 92.000 ;
    END
  END la_data_in_core[77]
  PIN la_data_in_core[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 89.700 179.770 92.000 ;
    END
  END la_data_in_core[78]
  PIN la_data_in_core[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 89.700 182.070 92.000 ;
    END
  END la_data_in_core[79]
  PIN la_data_in_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 89.700 25.210 92.000 ;
    END
  END la_data_in_core[7]
  PIN la_data_in_core[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 89.700 183.910 92.000 ;
    END
  END la_data_in_core[80]
  PIN la_data_in_core[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 89.700 186.210 92.000 ;
    END
  END la_data_in_core[81]
  PIN la_data_in_core[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 89.700 188.510 92.000 ;
    END
  END la_data_in_core[82]
  PIN la_data_in_core[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 89.700 190.810 92.000 ;
    END
  END la_data_in_core[83]
  PIN la_data_in_core[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 89.700 192.650 92.000 ;
    END
  END la_data_in_core[84]
  PIN la_data_in_core[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 89.700 194.950 92.000 ;
    END
  END la_data_in_core[85]
  PIN la_data_in_core[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 89.700 197.250 92.000 ;
    END
  END la_data_in_core[86]
  PIN la_data_in_core[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 89.700 199.550 92.000 ;
    END
  END la_data_in_core[87]
  PIN la_data_in_core[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 89.700 201.390 92.000 ;
    END
  END la_data_in_core[88]
  PIN la_data_in_core[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 89.700 203.690 92.000 ;
    END
  END la_data_in_core[89]
  PIN la_data_in_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 89.700 27.050 92.000 ;
    END
  END la_data_in_core[8]
  PIN la_data_in_core[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 89.700 205.990 92.000 ;
    END
  END la_data_in_core[90]
  PIN la_data_in_core[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 89.700 207.830 92.000 ;
    END
  END la_data_in_core[91]
  PIN la_data_in_core[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 89.700 210.130 92.000 ;
    END
  END la_data_in_core[92]
  PIN la_data_in_core[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 89.700 212.430 92.000 ;
    END
  END la_data_in_core[93]
  PIN la_data_in_core[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 89.700 214.730 92.000 ;
    END
  END la_data_in_core[94]
  PIN la_data_in_core[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 89.700 216.570 92.000 ;
    END
  END la_data_in_core[95]
  PIN la_data_in_core[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 89.700 218.870 92.000 ;
    END
  END la_data_in_core[96]
  PIN la_data_in_core[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 89.700 221.170 92.000 ;
    END
  END la_data_in_core[97]
  PIN la_data_in_core[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 89.700 223.470 92.000 ;
    END
  END la_data_in_core[98]
  PIN la_data_in_core[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 89.700 225.310 92.000 ;
    END
  END la_data_in_core[99]
  PIN la_data_in_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 89.700 29.350 92.000 ;
    END
  END la_data_in_core[9]
  PIN la_data_in_mprj[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 -2.000 280.050 0.300 ;
    END
  END la_data_in_mprj[0]
  PIN la_data_in_mprj[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 -2.000 497.630 0.300 ;
    END
  END la_data_in_mprj[100]
  PIN la_data_in_mprj[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 -2.000 499.930 0.300 ;
    END
  END la_data_in_mprj[101]
  PIN la_data_in_mprj[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 -2.000 502.230 0.300 ;
    END
  END la_data_in_mprj[102]
  PIN la_data_in_mprj[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 -2.000 504.530 0.300 ;
    END
  END la_data_in_mprj[103]
  PIN la_data_in_mprj[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 -2.000 506.370 0.300 ;
    END
  END la_data_in_mprj[104]
  PIN la_data_in_mprj[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 -2.000 508.670 0.300 ;
    END
  END la_data_in_mprj[105]
  PIN la_data_in_mprj[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 -2.000 510.970 0.300 ;
    END
  END la_data_in_mprj[106]
  PIN la_data_in_mprj[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 -2.000 513.270 0.300 ;
    END
  END la_data_in_mprj[107]
  PIN la_data_in_mprj[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 -2.000 515.110 0.300 ;
    END
  END la_data_in_mprj[108]
  PIN la_data_in_mprj[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 -2.000 517.410 0.300 ;
    END
  END la_data_in_mprj[109]
  PIN la_data_in_mprj[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 -2.000 301.670 0.300 ;
    END
  END la_data_in_mprj[10]
  PIN la_data_in_mprj[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 -2.000 519.710 0.300 ;
    END
  END la_data_in_mprj[110]
  PIN la_data_in_mprj[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 -2.000 521.550 0.300 ;
    END
  END la_data_in_mprj[111]
  PIN la_data_in_mprj[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 -2.000 523.850 0.300 ;
    END
  END la_data_in_mprj[112]
  PIN la_data_in_mprj[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 -2.000 526.150 0.300 ;
    END
  END la_data_in_mprj[113]
  PIN la_data_in_mprj[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 -2.000 528.450 0.300 ;
    END
  END la_data_in_mprj[114]
  PIN la_data_in_mprj[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 -2.000 530.290 0.300 ;
    END
  END la_data_in_mprj[115]
  PIN la_data_in_mprj[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 -2.000 532.590 0.300 ;
    END
  END la_data_in_mprj[116]
  PIN la_data_in_mprj[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 -2.000 534.890 0.300 ;
    END
  END la_data_in_mprj[117]
  PIN la_data_in_mprj[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 -2.000 537.190 0.300 ;
    END
  END la_data_in_mprj[118]
  PIN la_data_in_mprj[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 -2.000 539.030 0.300 ;
    END
  END la_data_in_mprj[119]
  PIN la_data_in_mprj[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 -2.000 303.970 0.300 ;
    END
  END la_data_in_mprj[11]
  PIN la_data_in_mprj[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 -2.000 541.330 0.300 ;
    END
  END la_data_in_mprj[120]
  PIN la_data_in_mprj[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 -2.000 543.630 0.300 ;
    END
  END la_data_in_mprj[121]
  PIN la_data_in_mprj[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 -2.000 545.930 0.300 ;
    END
  END la_data_in_mprj[122]
  PIN la_data_in_mprj[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 -2.000 547.770 0.300 ;
    END
  END la_data_in_mprj[123]
  PIN la_data_in_mprj[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 -2.000 550.070 0.300 ;
    END
  END la_data_in_mprj[124]
  PIN la_data_in_mprj[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 -2.000 552.370 0.300 ;
    END
  END la_data_in_mprj[125]
  PIN la_data_in_mprj[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 -2.000 554.670 0.300 ;
    END
  END la_data_in_mprj[126]
  PIN la_data_in_mprj[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 -2.000 556.510 0.300 ;
    END
  END la_data_in_mprj[127]
  PIN la_data_in_mprj[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 -2.000 306.270 0.300 ;
    END
  END la_data_in_mprj[12]
  PIN la_data_in_mprj[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 -2.000 308.110 0.300 ;
    END
  END la_data_in_mprj[13]
  PIN la_data_in_mprj[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 -2.000 310.410 0.300 ;
    END
  END la_data_in_mprj[14]
  PIN la_data_in_mprj[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 -2.000 312.710 0.300 ;
    END
  END la_data_in_mprj[15]
  PIN la_data_in_mprj[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 -2.000 315.010 0.300 ;
    END
  END la_data_in_mprj[16]
  PIN la_data_in_mprj[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 -2.000 316.850 0.300 ;
    END
  END la_data_in_mprj[17]
  PIN la_data_in_mprj[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 -2.000 319.150 0.300 ;
    END
  END la_data_in_mprj[18]
  PIN la_data_in_mprj[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 -2.000 321.450 0.300 ;
    END
  END la_data_in_mprj[19]
  PIN la_data_in_mprj[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 -2.000 281.890 0.300 ;
    END
  END la_data_in_mprj[1]
  PIN la_data_in_mprj[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 -2.000 323.290 0.300 ;
    END
  END la_data_in_mprj[20]
  PIN la_data_in_mprj[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 -2.000 325.590 0.300 ;
    END
  END la_data_in_mprj[21]
  PIN la_data_in_mprj[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 -2.000 327.890 0.300 ;
    END
  END la_data_in_mprj[22]
  PIN la_data_in_mprj[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 -2.000 330.190 0.300 ;
    END
  END la_data_in_mprj[23]
  PIN la_data_in_mprj[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 -2.000 332.030 0.300 ;
    END
  END la_data_in_mprj[24]
  PIN la_data_in_mprj[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 -2.000 334.330 0.300 ;
    END
  END la_data_in_mprj[25]
  PIN la_data_in_mprj[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 -2.000 336.630 0.300 ;
    END
  END la_data_in_mprj[26]
  PIN la_data_in_mprj[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 -2.000 338.930 0.300 ;
    END
  END la_data_in_mprj[27]
  PIN la_data_in_mprj[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 -2.000 340.770 0.300 ;
    END
  END la_data_in_mprj[28]
  PIN la_data_in_mprj[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 -2.000 343.070 0.300 ;
    END
  END la_data_in_mprj[29]
  PIN la_data_in_mprj[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 -2.000 284.190 0.300 ;
    END
  END la_data_in_mprj[2]
  PIN la_data_in_mprj[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 -2.000 345.370 0.300 ;
    END
  END la_data_in_mprj[30]
  PIN la_data_in_mprj[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 -2.000 347.670 0.300 ;
    END
  END la_data_in_mprj[31]
  PIN la_data_in_mprj[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 -2.000 349.510 0.300 ;
    END
  END la_data_in_mprj[32]
  PIN la_data_in_mprj[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 -2.000 351.810 0.300 ;
    END
  END la_data_in_mprj[33]
  PIN la_data_in_mprj[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 -2.000 354.110 0.300 ;
    END
  END la_data_in_mprj[34]
  PIN la_data_in_mprj[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 -2.000 356.410 0.300 ;
    END
  END la_data_in_mprj[35]
  PIN la_data_in_mprj[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 -2.000 358.250 0.300 ;
    END
  END la_data_in_mprj[36]
  PIN la_data_in_mprj[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 -2.000 360.550 0.300 ;
    END
  END la_data_in_mprj[37]
  PIN la_data_in_mprj[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 -2.000 362.850 0.300 ;
    END
  END la_data_in_mprj[38]
  PIN la_data_in_mprj[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 -2.000 364.690 0.300 ;
    END
  END la_data_in_mprj[39]
  PIN la_data_in_mprj[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 -2.000 286.490 0.300 ;
    END
  END la_data_in_mprj[3]
  PIN la_data_in_mprj[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 -2.000 366.990 0.300 ;
    END
  END la_data_in_mprj[40]
  PIN la_data_in_mprj[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 -2.000 369.290 0.300 ;
    END
  END la_data_in_mprj[41]
  PIN la_data_in_mprj[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 -2.000 371.590 0.300 ;
    END
  END la_data_in_mprj[42]
  PIN la_data_in_mprj[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 -2.000 373.430 0.300 ;
    END
  END la_data_in_mprj[43]
  PIN la_data_in_mprj[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 -2.000 375.730 0.300 ;
    END
  END la_data_in_mprj[44]
  PIN la_data_in_mprj[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 -2.000 378.030 0.300 ;
    END
  END la_data_in_mprj[45]
  PIN la_data_in_mprj[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 -2.000 380.330 0.300 ;
    END
  END la_data_in_mprj[46]
  PIN la_data_in_mprj[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 -2.000 382.170 0.300 ;
    END
  END la_data_in_mprj[47]
  PIN la_data_in_mprj[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 -2.000 384.470 0.300 ;
    END
  END la_data_in_mprj[48]
  PIN la_data_in_mprj[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 -2.000 386.770 0.300 ;
    END
  END la_data_in_mprj[49]
  PIN la_data_in_mprj[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 -2.000 288.790 0.300 ;
    END
  END la_data_in_mprj[4]
  PIN la_data_in_mprj[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 -2.000 389.070 0.300 ;
    END
  END la_data_in_mprj[50]
  PIN la_data_in_mprj[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 -2.000 390.910 0.300 ;
    END
  END la_data_in_mprj[51]
  PIN la_data_in_mprj[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 -2.000 393.210 0.300 ;
    END
  END la_data_in_mprj[52]
  PIN la_data_in_mprj[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 -2.000 395.510 0.300 ;
    END
  END la_data_in_mprj[53]
  PIN la_data_in_mprj[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 -2.000 397.810 0.300 ;
    END
  END la_data_in_mprj[54]
  PIN la_data_in_mprj[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 -2.000 399.650 0.300 ;
    END
  END la_data_in_mprj[55]
  PIN la_data_in_mprj[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 -2.000 401.950 0.300 ;
    END
  END la_data_in_mprj[56]
  PIN la_data_in_mprj[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 -2.000 404.250 0.300 ;
    END
  END la_data_in_mprj[57]
  PIN la_data_in_mprj[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 -2.000 406.090 0.300 ;
    END
  END la_data_in_mprj[58]
  PIN la_data_in_mprj[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 -2.000 408.390 0.300 ;
    END
  END la_data_in_mprj[59]
  PIN la_data_in_mprj[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 -2.000 290.630 0.300 ;
    END
  END la_data_in_mprj[5]
  PIN la_data_in_mprj[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 -2.000 410.690 0.300 ;
    END
  END la_data_in_mprj[60]
  PIN la_data_in_mprj[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 -2.000 412.990 0.300 ;
    END
  END la_data_in_mprj[61]
  PIN la_data_in_mprj[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 -2.000 414.830 0.300 ;
    END
  END la_data_in_mprj[62]
  PIN la_data_in_mprj[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 -2.000 417.130 0.300 ;
    END
  END la_data_in_mprj[63]
  PIN la_data_in_mprj[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 -2.000 419.430 0.300 ;
    END
  END la_data_in_mprj[64]
  PIN la_data_in_mprj[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 -2.000 421.730 0.300 ;
    END
  END la_data_in_mprj[65]
  PIN la_data_in_mprj[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 -2.000 423.570 0.300 ;
    END
  END la_data_in_mprj[66]
  PIN la_data_in_mprj[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 -2.000 425.870 0.300 ;
    END
  END la_data_in_mprj[67]
  PIN la_data_in_mprj[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 -2.000 428.170 0.300 ;
    END
  END la_data_in_mprj[68]
  PIN la_data_in_mprj[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 -2.000 430.470 0.300 ;
    END
  END la_data_in_mprj[69]
  PIN la_data_in_mprj[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 -2.000 292.930 0.300 ;
    END
  END la_data_in_mprj[6]
  PIN la_data_in_mprj[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 -2.000 432.310 0.300 ;
    END
  END la_data_in_mprj[70]
  PIN la_data_in_mprj[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 -2.000 434.610 0.300 ;
    END
  END la_data_in_mprj[71]
  PIN la_data_in_mprj[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 -2.000 436.910 0.300 ;
    END
  END la_data_in_mprj[72]
  PIN la_data_in_mprj[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 -2.000 439.210 0.300 ;
    END
  END la_data_in_mprj[73]
  PIN la_data_in_mprj[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 -2.000 441.050 0.300 ;
    END
  END la_data_in_mprj[74]
  PIN la_data_in_mprj[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 -2.000 443.350 0.300 ;
    END
  END la_data_in_mprj[75]
  PIN la_data_in_mprj[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 -2.000 445.650 0.300 ;
    END
  END la_data_in_mprj[76]
  PIN la_data_in_mprj[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 -2.000 447.490 0.300 ;
    END
  END la_data_in_mprj[77]
  PIN la_data_in_mprj[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 -2.000 449.790 0.300 ;
    END
  END la_data_in_mprj[78]
  PIN la_data_in_mprj[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 -2.000 452.090 0.300 ;
    END
  END la_data_in_mprj[79]
  PIN la_data_in_mprj[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 -2.000 295.230 0.300 ;
    END
  END la_data_in_mprj[7]
  PIN la_data_in_mprj[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 -2.000 454.390 0.300 ;
    END
  END la_data_in_mprj[80]
  PIN la_data_in_mprj[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 -2.000 456.230 0.300 ;
    END
  END la_data_in_mprj[81]
  PIN la_data_in_mprj[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 -2.000 458.530 0.300 ;
    END
  END la_data_in_mprj[82]
  PIN la_data_in_mprj[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 -2.000 460.830 0.300 ;
    END
  END la_data_in_mprj[83]
  PIN la_data_in_mprj[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 -2.000 463.130 0.300 ;
    END
  END la_data_in_mprj[84]
  PIN la_data_in_mprj[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 -2.000 464.970 0.300 ;
    END
  END la_data_in_mprj[85]
  PIN la_data_in_mprj[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 -2.000 467.270 0.300 ;
    END
  END la_data_in_mprj[86]
  PIN la_data_in_mprj[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 -2.000 469.570 0.300 ;
    END
  END la_data_in_mprj[87]
  PIN la_data_in_mprj[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 -2.000 471.870 0.300 ;
    END
  END la_data_in_mprj[88]
  PIN la_data_in_mprj[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 -2.000 473.710 0.300 ;
    END
  END la_data_in_mprj[89]
  PIN la_data_in_mprj[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 -2.000 297.530 0.300 ;
    END
  END la_data_in_mprj[8]
  PIN la_data_in_mprj[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 -2.000 476.010 0.300 ;
    END
  END la_data_in_mprj[90]
  PIN la_data_in_mprj[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 -2.000 478.310 0.300 ;
    END
  END la_data_in_mprj[91]
  PIN la_data_in_mprj[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 -2.000 480.610 0.300 ;
    END
  END la_data_in_mprj[92]
  PIN la_data_in_mprj[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 -2.000 482.450 0.300 ;
    END
  END la_data_in_mprj[93]
  PIN la_data_in_mprj[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 -2.000 484.750 0.300 ;
    END
  END la_data_in_mprj[94]
  PIN la_data_in_mprj[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 -2.000 487.050 0.300 ;
    END
  END la_data_in_mprj[95]
  PIN la_data_in_mprj[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 -2.000 488.890 0.300 ;
    END
  END la_data_in_mprj[96]
  PIN la_data_in_mprj[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 -2.000 491.190 0.300 ;
    END
  END la_data_in_mprj[97]
  PIN la_data_in_mprj[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 -2.000 493.490 0.300 ;
    END
  END la_data_in_mprj[98]
  PIN la_data_in_mprj[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 -2.000 495.790 0.300 ;
    END
  END la_data_in_mprj[99]
  PIN la_data_in_mprj[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 -2.000 299.370 0.300 ;
    END
  END la_data_in_mprj[9]
  PIN la_data_out_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 89.700 288.790 92.000 ;
    END
  END la_data_out_core[0]
  PIN la_data_out_core[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 89.700 506.370 92.000 ;
    END
  END la_data_out_core[100]
  PIN la_data_out_core[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 89.700 508.670 92.000 ;
    END
  END la_data_out_core[101]
  PIN la_data_out_core[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 89.700 510.970 92.000 ;
    END
  END la_data_out_core[102]
  PIN la_data_out_core[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 89.700 513.270 92.000 ;
    END
  END la_data_out_core[103]
  PIN la_data_out_core[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 89.700 515.110 92.000 ;
    END
  END la_data_out_core[104]
  PIN la_data_out_core[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 89.700 517.410 92.000 ;
    END
  END la_data_out_core[105]
  PIN la_data_out_core[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 89.700 519.710 92.000 ;
    END
  END la_data_out_core[106]
  PIN la_data_out_core[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 89.700 521.550 92.000 ;
    END
  END la_data_out_core[107]
  PIN la_data_out_core[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 89.700 523.850 92.000 ;
    END
  END la_data_out_core[108]
  PIN la_data_out_core[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 89.700 526.150 92.000 ;
    END
  END la_data_out_core[109]
  PIN la_data_out_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 89.700 310.410 92.000 ;
    END
  END la_data_out_core[10]
  PIN la_data_out_core[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 89.700 528.450 92.000 ;
    END
  END la_data_out_core[110]
  PIN la_data_out_core[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 89.700 530.290 92.000 ;
    END
  END la_data_out_core[111]
  PIN la_data_out_core[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 89.700 532.590 92.000 ;
    END
  END la_data_out_core[112]
  PIN la_data_out_core[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 89.700 534.890 92.000 ;
    END
  END la_data_out_core[113]
  PIN la_data_out_core[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 89.700 537.190 92.000 ;
    END
  END la_data_out_core[114]
  PIN la_data_out_core[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 89.700 539.030 92.000 ;
    END
  END la_data_out_core[115]
  PIN la_data_out_core[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 89.700 541.330 92.000 ;
    END
  END la_data_out_core[116]
  PIN la_data_out_core[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 89.700 543.630 92.000 ;
    END
  END la_data_out_core[117]
  PIN la_data_out_core[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 89.700 545.930 92.000 ;
    END
  END la_data_out_core[118]
  PIN la_data_out_core[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 89.700 547.770 92.000 ;
    END
  END la_data_out_core[119]
  PIN la_data_out_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 89.700 312.710 92.000 ;
    END
  END la_data_out_core[11]
  PIN la_data_out_core[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 89.700 550.070 92.000 ;
    END
  END la_data_out_core[120]
  PIN la_data_out_core[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 89.700 552.370 92.000 ;
    END
  END la_data_out_core[121]
  PIN la_data_out_core[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 89.700 554.670 92.000 ;
    END
  END la_data_out_core[122]
  PIN la_data_out_core[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 89.700 556.510 92.000 ;
    END
  END la_data_out_core[123]
  PIN la_data_out_core[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 89.700 558.810 92.000 ;
    END
  END la_data_out_core[124]
  PIN la_data_out_core[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 89.700 561.110 92.000 ;
    END
  END la_data_out_core[125]
  PIN la_data_out_core[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 89.700 562.950 92.000 ;
    END
  END la_data_out_core[126]
  PIN la_data_out_core[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 89.700 565.250 92.000 ;
    END
  END la_data_out_core[127]
  PIN la_data_out_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 89.700 315.010 92.000 ;
    END
  END la_data_out_core[12]
  PIN la_data_out_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 89.700 316.850 92.000 ;
    END
  END la_data_out_core[13]
  PIN la_data_out_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 89.700 319.150 92.000 ;
    END
  END la_data_out_core[14]
  PIN la_data_out_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 89.700 321.450 92.000 ;
    END
  END la_data_out_core[15]
  PIN la_data_out_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 89.700 323.290 92.000 ;
    END
  END la_data_out_core[16]
  PIN la_data_out_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 89.700 325.590 92.000 ;
    END
  END la_data_out_core[17]
  PIN la_data_out_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 89.700 327.890 92.000 ;
    END
  END la_data_out_core[18]
  PIN la_data_out_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 89.700 330.190 92.000 ;
    END
  END la_data_out_core[19]
  PIN la_data_out_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 89.700 290.630 92.000 ;
    END
  END la_data_out_core[1]
  PIN la_data_out_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 89.700 332.030 92.000 ;
    END
  END la_data_out_core[20]
  PIN la_data_out_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 89.700 334.330 92.000 ;
    END
  END la_data_out_core[21]
  PIN la_data_out_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 89.700 336.630 92.000 ;
    END
  END la_data_out_core[22]
  PIN la_data_out_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 89.700 338.930 92.000 ;
    END
  END la_data_out_core[23]
  PIN la_data_out_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 89.700 340.770 92.000 ;
    END
  END la_data_out_core[24]
  PIN la_data_out_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 89.700 343.070 92.000 ;
    END
  END la_data_out_core[25]
  PIN la_data_out_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 89.700 345.370 92.000 ;
    END
  END la_data_out_core[26]
  PIN la_data_out_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 89.700 347.670 92.000 ;
    END
  END la_data_out_core[27]
  PIN la_data_out_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 89.700 349.510 92.000 ;
    END
  END la_data_out_core[28]
  PIN la_data_out_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 89.700 351.810 92.000 ;
    END
  END la_data_out_core[29]
  PIN la_data_out_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 89.700 292.930 92.000 ;
    END
  END la_data_out_core[2]
  PIN la_data_out_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 89.700 354.110 92.000 ;
    END
  END la_data_out_core[30]
  PIN la_data_out_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 89.700 356.410 92.000 ;
    END
  END la_data_out_core[31]
  PIN la_data_out_core[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 89.700 358.250 92.000 ;
    END
  END la_data_out_core[32]
  PIN la_data_out_core[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 89.700 360.550 92.000 ;
    END
  END la_data_out_core[33]
  PIN la_data_out_core[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 89.700 362.850 92.000 ;
    END
  END la_data_out_core[34]
  PIN la_data_out_core[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 89.700 364.690 92.000 ;
    END
  END la_data_out_core[35]
  PIN la_data_out_core[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 89.700 366.990 92.000 ;
    END
  END la_data_out_core[36]
  PIN la_data_out_core[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 89.700 369.290 92.000 ;
    END
  END la_data_out_core[37]
  PIN la_data_out_core[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 89.700 371.590 92.000 ;
    END
  END la_data_out_core[38]
  PIN la_data_out_core[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 89.700 373.430 92.000 ;
    END
  END la_data_out_core[39]
  PIN la_data_out_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 89.700 295.230 92.000 ;
    END
  END la_data_out_core[3]
  PIN la_data_out_core[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 89.700 375.730 92.000 ;
    END
  END la_data_out_core[40]
  PIN la_data_out_core[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 89.700 378.030 92.000 ;
    END
  END la_data_out_core[41]
  PIN la_data_out_core[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 89.700 380.330 92.000 ;
    END
  END la_data_out_core[42]
  PIN la_data_out_core[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 89.700 382.170 92.000 ;
    END
  END la_data_out_core[43]
  PIN la_data_out_core[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 89.700 384.470 92.000 ;
    END
  END la_data_out_core[44]
  PIN la_data_out_core[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 89.700 386.770 92.000 ;
    END
  END la_data_out_core[45]
  PIN la_data_out_core[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 89.700 389.070 92.000 ;
    END
  END la_data_out_core[46]
  PIN la_data_out_core[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 89.700 390.910 92.000 ;
    END
  END la_data_out_core[47]
  PIN la_data_out_core[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 89.700 393.210 92.000 ;
    END
  END la_data_out_core[48]
  PIN la_data_out_core[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 89.700 395.510 92.000 ;
    END
  END la_data_out_core[49]
  PIN la_data_out_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 89.700 297.530 92.000 ;
    END
  END la_data_out_core[4]
  PIN la_data_out_core[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 89.700 397.810 92.000 ;
    END
  END la_data_out_core[50]
  PIN la_data_out_core[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 89.700 399.650 92.000 ;
    END
  END la_data_out_core[51]
  PIN la_data_out_core[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 89.700 401.950 92.000 ;
    END
  END la_data_out_core[52]
  PIN la_data_out_core[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 89.700 404.250 92.000 ;
    END
  END la_data_out_core[53]
  PIN la_data_out_core[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 89.700 406.090 92.000 ;
    END
  END la_data_out_core[54]
  PIN la_data_out_core[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 89.700 408.390 92.000 ;
    END
  END la_data_out_core[55]
  PIN la_data_out_core[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 89.700 410.690 92.000 ;
    END
  END la_data_out_core[56]
  PIN la_data_out_core[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 89.700 412.990 92.000 ;
    END
  END la_data_out_core[57]
  PIN la_data_out_core[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 89.700 414.830 92.000 ;
    END
  END la_data_out_core[58]
  PIN la_data_out_core[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 89.700 417.130 92.000 ;
    END
  END la_data_out_core[59]
  PIN la_data_out_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 89.700 299.370 92.000 ;
    END
  END la_data_out_core[5]
  PIN la_data_out_core[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 89.700 419.430 92.000 ;
    END
  END la_data_out_core[60]
  PIN la_data_out_core[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 89.700 421.730 92.000 ;
    END
  END la_data_out_core[61]
  PIN la_data_out_core[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 89.700 423.570 92.000 ;
    END
  END la_data_out_core[62]
  PIN la_data_out_core[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 89.700 425.870 92.000 ;
    END
  END la_data_out_core[63]
  PIN la_data_out_core[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 89.700 428.170 92.000 ;
    END
  END la_data_out_core[64]
  PIN la_data_out_core[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 89.700 430.470 92.000 ;
    END
  END la_data_out_core[65]
  PIN la_data_out_core[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 89.700 432.310 92.000 ;
    END
  END la_data_out_core[66]
  PIN la_data_out_core[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 89.700 434.610 92.000 ;
    END
  END la_data_out_core[67]
  PIN la_data_out_core[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 89.700 436.910 92.000 ;
    END
  END la_data_out_core[68]
  PIN la_data_out_core[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 89.700 439.210 92.000 ;
    END
  END la_data_out_core[69]
  PIN la_data_out_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 89.700 301.670 92.000 ;
    END
  END la_data_out_core[6]
  PIN la_data_out_core[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 89.700 441.050 92.000 ;
    END
  END la_data_out_core[70]
  PIN la_data_out_core[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 89.700 443.350 92.000 ;
    END
  END la_data_out_core[71]
  PIN la_data_out_core[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 89.700 445.650 92.000 ;
    END
  END la_data_out_core[72]
  PIN la_data_out_core[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 89.700 447.490 92.000 ;
    END
  END la_data_out_core[73]
  PIN la_data_out_core[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 89.700 449.790 92.000 ;
    END
  END la_data_out_core[74]
  PIN la_data_out_core[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 89.700 452.090 92.000 ;
    END
  END la_data_out_core[75]
  PIN la_data_out_core[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 89.700 454.390 92.000 ;
    END
  END la_data_out_core[76]
  PIN la_data_out_core[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 89.700 456.230 92.000 ;
    END
  END la_data_out_core[77]
  PIN la_data_out_core[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 89.700 458.530 92.000 ;
    END
  END la_data_out_core[78]
  PIN la_data_out_core[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 89.700 460.830 92.000 ;
    END
  END la_data_out_core[79]
  PIN la_data_out_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 89.700 303.970 92.000 ;
    END
  END la_data_out_core[7]
  PIN la_data_out_core[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 89.700 463.130 92.000 ;
    END
  END la_data_out_core[80]
  PIN la_data_out_core[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 89.700 464.970 92.000 ;
    END
  END la_data_out_core[81]
  PIN la_data_out_core[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 89.700 467.270 92.000 ;
    END
  END la_data_out_core[82]
  PIN la_data_out_core[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 89.700 469.570 92.000 ;
    END
  END la_data_out_core[83]
  PIN la_data_out_core[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 89.700 471.870 92.000 ;
    END
  END la_data_out_core[84]
  PIN la_data_out_core[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 89.700 473.710 92.000 ;
    END
  END la_data_out_core[85]
  PIN la_data_out_core[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 89.700 476.010 92.000 ;
    END
  END la_data_out_core[86]
  PIN la_data_out_core[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 89.700 478.310 92.000 ;
    END
  END la_data_out_core[87]
  PIN la_data_out_core[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 89.700 480.610 92.000 ;
    END
  END la_data_out_core[88]
  PIN la_data_out_core[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 89.700 482.450 92.000 ;
    END
  END la_data_out_core[89]
  PIN la_data_out_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 89.700 306.270 92.000 ;
    END
  END la_data_out_core[8]
  PIN la_data_out_core[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 89.700 484.750 92.000 ;
    END
  END la_data_out_core[90]
  PIN la_data_out_core[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 89.700 487.050 92.000 ;
    END
  END la_data_out_core[91]
  PIN la_data_out_core[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 89.700 488.890 92.000 ;
    END
  END la_data_out_core[92]
  PIN la_data_out_core[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 89.700 491.190 92.000 ;
    END
  END la_data_out_core[93]
  PIN la_data_out_core[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 89.700 493.490 92.000 ;
    END
  END la_data_out_core[94]
  PIN la_data_out_core[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 89.700 495.790 92.000 ;
    END
  END la_data_out_core[95]
  PIN la_data_out_core[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 89.700 497.630 92.000 ;
    END
  END la_data_out_core[96]
  PIN la_data_out_core[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 89.700 499.930 92.000 ;
    END
  END la_data_out_core[97]
  PIN la_data_out_core[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 89.700 502.230 92.000 ;
    END
  END la_data_out_core[98]
  PIN la_data_out_core[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 89.700 504.530 92.000 ;
    END
  END la_data_out_core[99]
  PIN la_data_out_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 89.700 308.110 92.000 ;
    END
  END la_data_out_core[9]
  PIN la_data_out_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 -2.000 1.290 0.300 ;
    END
  END la_data_out_mprj[0]
  PIN la_data_out_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 -2.000 218.870 0.300 ;
    END
  END la_data_out_mprj[100]
  PIN la_data_out_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 -2.000 221.170 0.300 ;
    END
  END la_data_out_mprj[101]
  PIN la_data_out_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 -2.000 223.470 0.300 ;
    END
  END la_data_out_mprj[102]
  PIN la_data_out_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 -2.000 225.310 0.300 ;
    END
  END la_data_out_mprj[103]
  PIN la_data_out_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 -2.000 227.610 0.300 ;
    END
  END la_data_out_mprj[104]
  PIN la_data_out_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 -2.000 229.910 0.300 ;
    END
  END la_data_out_mprj[105]
  PIN la_data_out_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 -2.000 232.210 0.300 ;
    END
  END la_data_out_mprj[106]
  PIN la_data_out_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 -2.000 234.050 0.300 ;
    END
  END la_data_out_mprj[107]
  PIN la_data_out_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 -2.000 236.350 0.300 ;
    END
  END la_data_out_mprj[108]
  PIN la_data_out_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 -2.000 238.650 0.300 ;
    END
  END la_data_out_mprj[109]
  PIN la_data_out_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 -2.000 22.910 0.300 ;
    END
  END la_data_out_mprj[10]
  PIN la_data_out_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 -2.000 240.950 0.300 ;
    END
  END la_data_out_mprj[110]
  PIN la_data_out_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 -2.000 242.790 0.300 ;
    END
  END la_data_out_mprj[111]
  PIN la_data_out_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 -2.000 245.090 0.300 ;
    END
  END la_data_out_mprj[112]
  PIN la_data_out_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 -2.000 247.390 0.300 ;
    END
  END la_data_out_mprj[113]
  PIN la_data_out_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 -2.000 249.230 0.300 ;
    END
  END la_data_out_mprj[114]
  PIN la_data_out_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 -2.000 251.530 0.300 ;
    END
  END la_data_out_mprj[115]
  PIN la_data_out_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 -2.000 253.830 0.300 ;
    END
  END la_data_out_mprj[116]
  PIN la_data_out_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 -2.000 256.130 0.300 ;
    END
  END la_data_out_mprj[117]
  PIN la_data_out_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 -2.000 257.970 0.300 ;
    END
  END la_data_out_mprj[118]
  PIN la_data_out_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 -2.000 260.270 0.300 ;
    END
  END la_data_out_mprj[119]
  PIN la_data_out_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 -2.000 25.210 0.300 ;
    END
  END la_data_out_mprj[11]
  PIN la_data_out_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 -2.000 262.570 0.300 ;
    END
  END la_data_out_mprj[120]
  PIN la_data_out_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 -2.000 264.870 0.300 ;
    END
  END la_data_out_mprj[121]
  PIN la_data_out_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 -2.000 266.710 0.300 ;
    END
  END la_data_out_mprj[122]
  PIN la_data_out_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 -2.000 269.010 0.300 ;
    END
  END la_data_out_mprj[123]
  PIN la_data_out_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 -2.000 271.310 0.300 ;
    END
  END la_data_out_mprj[124]
  PIN la_data_out_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 -2.000 273.610 0.300 ;
    END
  END la_data_out_mprj[125]
  PIN la_data_out_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 -2.000 275.450 0.300 ;
    END
  END la_data_out_mprj[126]
  PIN la_data_out_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 -2.000 277.750 0.300 ;
    END
  END la_data_out_mprj[127]
  PIN la_data_out_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 -2.000 27.050 0.300 ;
    END
  END la_data_out_mprj[12]
  PIN la_data_out_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 -2.000 29.350 0.300 ;
    END
  END la_data_out_mprj[13]
  PIN la_data_out_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 -2.000 31.650 0.300 ;
    END
  END la_data_out_mprj[14]
  PIN la_data_out_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 -2.000 33.950 0.300 ;
    END
  END la_data_out_mprj[15]
  PIN la_data_out_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 -2.000 35.790 0.300 ;
    END
  END la_data_out_mprj[16]
  PIN la_data_out_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 -2.000 38.090 0.300 ;
    END
  END la_data_out_mprj[17]
  PIN la_data_out_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 -2.000 40.390 0.300 ;
    END
  END la_data_out_mprj[18]
  PIN la_data_out_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 -2.000 42.230 0.300 ;
    END
  END la_data_out_mprj[19]
  PIN la_data_out_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 -2.000 3.130 0.300 ;
    END
  END la_data_out_mprj[1]
  PIN la_data_out_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 -2.000 44.530 0.300 ;
    END
  END la_data_out_mprj[20]
  PIN la_data_out_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 -2.000 46.830 0.300 ;
    END
  END la_data_out_mprj[21]
  PIN la_data_out_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 -2.000 49.130 0.300 ;
    END
  END la_data_out_mprj[22]
  PIN la_data_out_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 -2.000 50.970 0.300 ;
    END
  END la_data_out_mprj[23]
  PIN la_data_out_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 -2.000 53.270 0.300 ;
    END
  END la_data_out_mprj[24]
  PIN la_data_out_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 -2.000 55.570 0.300 ;
    END
  END la_data_out_mprj[25]
  PIN la_data_out_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 -2.000 57.870 0.300 ;
    END
  END la_data_out_mprj[26]
  PIN la_data_out_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 -2.000 59.710 0.300 ;
    END
  END la_data_out_mprj[27]
  PIN la_data_out_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 -2.000 62.010 0.300 ;
    END
  END la_data_out_mprj[28]
  PIN la_data_out_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 -2.000 64.310 0.300 ;
    END
  END la_data_out_mprj[29]
  PIN la_data_out_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 -2.000 5.430 0.300 ;
    END
  END la_data_out_mprj[2]
  PIN la_data_out_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 -2.000 66.610 0.300 ;
    END
  END la_data_out_mprj[30]
  PIN la_data_out_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 -2.000 68.450 0.300 ;
    END
  END la_data_out_mprj[31]
  PIN la_data_out_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 -2.000 70.750 0.300 ;
    END
  END la_data_out_mprj[32]
  PIN la_data_out_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 -2.000 73.050 0.300 ;
    END
  END la_data_out_mprj[33]
  PIN la_data_out_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 -2.000 75.350 0.300 ;
    END
  END la_data_out_mprj[34]
  PIN la_data_out_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 -2.000 77.190 0.300 ;
    END
  END la_data_out_mprj[35]
  PIN la_data_out_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 -2.000 79.490 0.300 ;
    END
  END la_data_out_mprj[36]
  PIN la_data_out_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 -2.000 81.790 0.300 ;
    END
  END la_data_out_mprj[37]
  PIN la_data_out_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 -2.000 83.630 0.300 ;
    END
  END la_data_out_mprj[38]
  PIN la_data_out_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 -2.000 85.930 0.300 ;
    END
  END la_data_out_mprj[39]
  PIN la_data_out_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 -2.000 7.730 0.300 ;
    END
  END la_data_out_mprj[3]
  PIN la_data_out_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 -2.000 88.230 0.300 ;
    END
  END la_data_out_mprj[40]
  PIN la_data_out_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 -2.000 90.530 0.300 ;
    END
  END la_data_out_mprj[41]
  PIN la_data_out_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 -2.000 92.370 0.300 ;
    END
  END la_data_out_mprj[42]
  PIN la_data_out_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 -2.000 94.670 0.300 ;
    END
  END la_data_out_mprj[43]
  PIN la_data_out_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 -2.000 96.970 0.300 ;
    END
  END la_data_out_mprj[44]
  PIN la_data_out_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 -2.000 99.270 0.300 ;
    END
  END la_data_out_mprj[45]
  PIN la_data_out_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 -2.000 101.110 0.300 ;
    END
  END la_data_out_mprj[46]
  PIN la_data_out_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 -2.000 103.410 0.300 ;
    END
  END la_data_out_mprj[47]
  PIN la_data_out_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 -2.000 105.710 0.300 ;
    END
  END la_data_out_mprj[48]
  PIN la_data_out_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 -2.000 108.010 0.300 ;
    END
  END la_data_out_mprj[49]
  PIN la_data_out_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 -2.000 9.570 0.300 ;
    END
  END la_data_out_mprj[4]
  PIN la_data_out_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 -2.000 109.850 0.300 ;
    END
  END la_data_out_mprj[50]
  PIN la_data_out_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 -2.000 112.150 0.300 ;
    END
  END la_data_out_mprj[51]
  PIN la_data_out_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 -2.000 114.450 0.300 ;
    END
  END la_data_out_mprj[52]
  PIN la_data_out_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 -2.000 116.750 0.300 ;
    END
  END la_data_out_mprj[53]
  PIN la_data_out_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 -2.000 118.590 0.300 ;
    END
  END la_data_out_mprj[54]
  PIN la_data_out_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 -2.000 120.890 0.300 ;
    END
  END la_data_out_mprj[55]
  PIN la_data_out_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 -2.000 123.190 0.300 ;
    END
  END la_data_out_mprj[56]
  PIN la_data_out_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 -2.000 125.030 0.300 ;
    END
  END la_data_out_mprj[57]
  PIN la_data_out_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 -2.000 127.330 0.300 ;
    END
  END la_data_out_mprj[58]
  PIN la_data_out_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 -2.000 129.630 0.300 ;
    END
  END la_data_out_mprj[59]
  PIN la_data_out_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 -2.000 11.870 0.300 ;
    END
  END la_data_out_mprj[5]
  PIN la_data_out_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 -2.000 131.930 0.300 ;
    END
  END la_data_out_mprj[60]
  PIN la_data_out_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 -2.000 133.770 0.300 ;
    END
  END la_data_out_mprj[61]
  PIN la_data_out_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 -2.000 136.070 0.300 ;
    END
  END la_data_out_mprj[62]
  PIN la_data_out_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 -2.000 138.370 0.300 ;
    END
  END la_data_out_mprj[63]
  PIN la_data_out_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 -2.000 140.670 0.300 ;
    END
  END la_data_out_mprj[64]
  PIN la_data_out_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 -2.000 142.510 0.300 ;
    END
  END la_data_out_mprj[65]
  PIN la_data_out_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 -2.000 144.810 0.300 ;
    END
  END la_data_out_mprj[66]
  PIN la_data_out_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 -2.000 147.110 0.300 ;
    END
  END la_data_out_mprj[67]
  PIN la_data_out_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 -2.000 149.410 0.300 ;
    END
  END la_data_out_mprj[68]
  PIN la_data_out_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 -2.000 151.250 0.300 ;
    END
  END la_data_out_mprj[69]
  PIN la_data_out_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 -2.000 14.170 0.300 ;
    END
  END la_data_out_mprj[6]
  PIN la_data_out_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 -2.000 153.550 0.300 ;
    END
  END la_data_out_mprj[70]
  PIN la_data_out_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 -2.000 155.850 0.300 ;
    END
  END la_data_out_mprj[71]
  PIN la_data_out_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 -2.000 158.150 0.300 ;
    END
  END la_data_out_mprj[72]
  PIN la_data_out_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 -2.000 159.990 0.300 ;
    END
  END la_data_out_mprj[73]
  PIN la_data_out_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 -2.000 162.290 0.300 ;
    END
  END la_data_out_mprj[74]
  PIN la_data_out_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 -2.000 164.590 0.300 ;
    END
  END la_data_out_mprj[75]
  PIN la_data_out_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 -2.000 166.430 0.300 ;
    END
  END la_data_out_mprj[76]
  PIN la_data_out_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 -2.000 168.730 0.300 ;
    END
  END la_data_out_mprj[77]
  PIN la_data_out_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 -2.000 171.030 0.300 ;
    END
  END la_data_out_mprj[78]
  PIN la_data_out_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 -2.000 173.330 0.300 ;
    END
  END la_data_out_mprj[79]
  PIN la_data_out_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 -2.000 16.470 0.300 ;
    END
  END la_data_out_mprj[7]
  PIN la_data_out_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 -2.000 175.170 0.300 ;
    END
  END la_data_out_mprj[80]
  PIN la_data_out_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 -2.000 177.470 0.300 ;
    END
  END la_data_out_mprj[81]
  PIN la_data_out_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 -2.000 179.770 0.300 ;
    END
  END la_data_out_mprj[82]
  PIN la_data_out_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 -2.000 182.070 0.300 ;
    END
  END la_data_out_mprj[83]
  PIN la_data_out_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 -2.000 183.910 0.300 ;
    END
  END la_data_out_mprj[84]
  PIN la_data_out_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 -2.000 186.210 0.300 ;
    END
  END la_data_out_mprj[85]
  PIN la_data_out_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 -2.000 188.510 0.300 ;
    END
  END la_data_out_mprj[86]
  PIN la_data_out_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 -2.000 190.810 0.300 ;
    END
  END la_data_out_mprj[87]
  PIN la_data_out_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 -2.000 192.650 0.300 ;
    END
  END la_data_out_mprj[88]
  PIN la_data_out_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 -2.000 194.950 0.300 ;
    END
  END la_data_out_mprj[89]
  PIN la_data_out_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 -2.000 18.310 0.300 ;
    END
  END la_data_out_mprj[8]
  PIN la_data_out_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 -2.000 197.250 0.300 ;
    END
  END la_data_out_mprj[90]
  PIN la_data_out_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 -2.000 199.550 0.300 ;
    END
  END la_data_out_mprj[91]
  PIN la_data_out_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 -2.000 201.390 0.300 ;
    END
  END la_data_out_mprj[92]
  PIN la_data_out_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 -2.000 203.690 0.300 ;
    END
  END la_data_out_mprj[93]
  PIN la_data_out_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 -2.000 205.990 0.300 ;
    END
  END la_data_out_mprj[94]
  PIN la_data_out_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 -2.000 207.830 0.300 ;
    END
  END la_data_out_mprj[95]
  PIN la_data_out_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 -2.000 210.130 0.300 ;
    END
  END la_data_out_mprj[96]
  PIN la_data_out_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 -2.000 212.430 0.300 ;
    END
  END la_data_out_mprj[97]
  PIN la_data_out_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 -2.000 214.730 0.300 ;
    END
  END la_data_out_mprj[98]
  PIN la_data_out_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 -2.000 216.570 0.300 ;
    END
  END la_data_out_mprj[99]
  PIN la_data_out_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 -2.000 20.610 0.300 ;
    END
  END la_data_out_mprj[9]
  PIN la_oen_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 89.700 567.550 92.000 ;
    END
  END la_oen_core[0]
  PIN la_oen_core[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 89.700 785.590 92.000 ;
    END
  END la_oen_core[100]
  PIN la_oen_core[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 89.700 787.430 92.000 ;
    END
  END la_oen_core[101]
  PIN la_oen_core[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 89.700 789.730 92.000 ;
    END
  END la_oen_core[102]
  PIN la_oen_core[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.750 89.700 792.030 92.000 ;
    END
  END la_oen_core[103]
  PIN la_oen_core[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 89.700 794.330 92.000 ;
    END
  END la_oen_core[104]
  PIN la_oen_core[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 89.700 796.170 92.000 ;
    END
  END la_oen_core[105]
  PIN la_oen_core[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 89.700 798.470 92.000 ;
    END
  END la_oen_core[106]
  PIN la_oen_core[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 89.700 800.770 92.000 ;
    END
  END la_oen_core[107]
  PIN la_oen_core[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 89.700 802.610 92.000 ;
    END
  END la_oen_core[108]
  PIN la_oen_core[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 89.700 804.910 92.000 ;
    END
  END la_oen_core[109]
  PIN la_oen_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 89.700 589.170 92.000 ;
    END
  END la_oen_core[10]
  PIN la_oen_core[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.930 89.700 807.210 92.000 ;
    END
  END la_oen_core[110]
  PIN la_oen_core[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 89.700 809.510 92.000 ;
    END
  END la_oen_core[111]
  PIN la_oen_core[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 89.700 811.350 92.000 ;
    END
  END la_oen_core[112]
  PIN la_oen_core[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 89.700 813.650 92.000 ;
    END
  END la_oen_core[113]
  PIN la_oen_core[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 89.700 815.950 92.000 ;
    END
  END la_oen_core[114]
  PIN la_oen_core[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 89.700 818.250 92.000 ;
    END
  END la_oen_core[115]
  PIN la_oen_core[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 89.700 820.090 92.000 ;
    END
  END la_oen_core[116]
  PIN la_oen_core[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 89.700 822.390 92.000 ;
    END
  END la_oen_core[117]
  PIN la_oen_core[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 89.700 824.690 92.000 ;
    END
  END la_oen_core[118]
  PIN la_oen_core[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 89.700 826.990 92.000 ;
    END
  END la_oen_core[119]
  PIN la_oen_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 89.700 591.470 92.000 ;
    END
  END la_oen_core[11]
  PIN la_oen_core[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 89.700 828.830 92.000 ;
    END
  END la_oen_core[120]
  PIN la_oen_core[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 89.700 831.130 92.000 ;
    END
  END la_oen_core[121]
  PIN la_oen_core[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 89.700 833.430 92.000 ;
    END
  END la_oen_core[122]
  PIN la_oen_core[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 89.700 835.730 92.000 ;
    END
  END la_oen_core[123]
  PIN la_oen_core[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 89.700 837.570 92.000 ;
    END
  END la_oen_core[124]
  PIN la_oen_core[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 89.700 839.870 92.000 ;
    END
  END la_oen_core[125]
  PIN la_oen_core[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 89.700 842.170 92.000 ;
    END
  END la_oen_core[126]
  PIN la_oen_core[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 89.700 844.010 92.000 ;
    END
  END la_oen_core[127]
  PIN la_oen_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 89.700 593.770 92.000 ;
    END
  END la_oen_core[12]
  PIN la_oen_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 89.700 596.070 92.000 ;
    END
  END la_oen_core[13]
  PIN la_oen_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 89.700 597.910 92.000 ;
    END
  END la_oen_core[14]
  PIN la_oen_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 89.700 600.210 92.000 ;
    END
  END la_oen_core[15]
  PIN la_oen_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 89.700 602.510 92.000 ;
    END
  END la_oen_core[16]
  PIN la_oen_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 89.700 604.350 92.000 ;
    END
  END la_oen_core[17]
  PIN la_oen_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 89.700 606.650 92.000 ;
    END
  END la_oen_core[18]
  PIN la_oen_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 89.700 608.950 92.000 ;
    END
  END la_oen_core[19]
  PIN la_oen_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 89.700 569.850 92.000 ;
    END
  END la_oen_core[1]
  PIN la_oen_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 89.700 611.250 92.000 ;
    END
  END la_oen_core[20]
  PIN la_oen_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 89.700 613.090 92.000 ;
    END
  END la_oen_core[21]
  PIN la_oen_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 89.700 615.390 92.000 ;
    END
  END la_oen_core[22]
  PIN la_oen_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 89.700 617.690 92.000 ;
    END
  END la_oen_core[23]
  PIN la_oen_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 89.700 619.990 92.000 ;
    END
  END la_oen_core[24]
  PIN la_oen_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 89.700 621.830 92.000 ;
    END
  END la_oen_core[25]
  PIN la_oen_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 89.700 624.130 92.000 ;
    END
  END la_oen_core[26]
  PIN la_oen_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 89.700 626.430 92.000 ;
    END
  END la_oen_core[27]
  PIN la_oen_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 89.700 628.730 92.000 ;
    END
  END la_oen_core[28]
  PIN la_oen_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 89.700 630.570 92.000 ;
    END
  END la_oen_core[29]
  PIN la_oen_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 89.700 571.690 92.000 ;
    END
  END la_oen_core[2]
  PIN la_oen_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 89.700 632.870 92.000 ;
    END
  END la_oen_core[30]
  PIN la_oen_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 89.700 635.170 92.000 ;
    END
  END la_oen_core[31]
  PIN la_oen_core[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 89.700 637.470 92.000 ;
    END
  END la_oen_core[32]
  PIN la_oen_core[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 89.700 639.310 92.000 ;
    END
  END la_oen_core[33]
  PIN la_oen_core[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 89.700 641.610 92.000 ;
    END
  END la_oen_core[34]
  PIN la_oen_core[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 89.700 643.910 92.000 ;
    END
  END la_oen_core[35]
  PIN la_oen_core[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 89.700 645.750 92.000 ;
    END
  END la_oen_core[36]
  PIN la_oen_core[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 89.700 648.050 92.000 ;
    END
  END la_oen_core[37]
  PIN la_oen_core[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 89.700 650.350 92.000 ;
    END
  END la_oen_core[38]
  PIN la_oen_core[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 89.700 652.650 92.000 ;
    END
  END la_oen_core[39]
  PIN la_oen_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 89.700 573.990 92.000 ;
    END
  END la_oen_core[3]
  PIN la_oen_core[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 89.700 654.490 92.000 ;
    END
  END la_oen_core[40]
  PIN la_oen_core[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 89.700 656.790 92.000 ;
    END
  END la_oen_core[41]
  PIN la_oen_core[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 89.700 659.090 92.000 ;
    END
  END la_oen_core[42]
  PIN la_oen_core[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 89.700 661.390 92.000 ;
    END
  END la_oen_core[43]
  PIN la_oen_core[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.950 89.700 663.230 92.000 ;
    END
  END la_oen_core[44]
  PIN la_oen_core[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 89.700 665.530 92.000 ;
    END
  END la_oen_core[45]
  PIN la_oen_core[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 89.700 667.830 92.000 ;
    END
  END la_oen_core[46]
  PIN la_oen_core[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 89.700 670.130 92.000 ;
    END
  END la_oen_core[47]
  PIN la_oen_core[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 89.700 671.970 92.000 ;
    END
  END la_oen_core[48]
  PIN la_oen_core[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 89.700 674.270 92.000 ;
    END
  END la_oen_core[49]
  PIN la_oen_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 89.700 576.290 92.000 ;
    END
  END la_oen_core[4]
  PIN la_oen_core[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 89.700 676.570 92.000 ;
    END
  END la_oen_core[50]
  PIN la_oen_core[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 89.700 678.870 92.000 ;
    END
  END la_oen_core[51]
  PIN la_oen_core[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 89.700 680.710 92.000 ;
    END
  END la_oen_core[52]
  PIN la_oen_core[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 89.700 683.010 92.000 ;
    END
  END la_oen_core[53]
  PIN la_oen_core[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 89.700 685.310 92.000 ;
    END
  END la_oen_core[54]
  PIN la_oen_core[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 89.700 687.150 92.000 ;
    END
  END la_oen_core[55]
  PIN la_oen_core[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 89.700 689.450 92.000 ;
    END
  END la_oen_core[56]
  PIN la_oen_core[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 89.700 691.750 92.000 ;
    END
  END la_oen_core[57]
  PIN la_oen_core[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 89.700 694.050 92.000 ;
    END
  END la_oen_core[58]
  PIN la_oen_core[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 89.700 695.890 92.000 ;
    END
  END la_oen_core[59]
  PIN la_oen_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 89.700 578.590 92.000 ;
    END
  END la_oen_core[5]
  PIN la_oen_core[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 89.700 698.190 92.000 ;
    END
  END la_oen_core[60]
  PIN la_oen_core[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 89.700 700.490 92.000 ;
    END
  END la_oen_core[61]
  PIN la_oen_core[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 89.700 702.790 92.000 ;
    END
  END la_oen_core[62]
  PIN la_oen_core[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 89.700 704.630 92.000 ;
    END
  END la_oen_core[63]
  PIN la_oen_core[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 89.700 706.930 92.000 ;
    END
  END la_oen_core[64]
  PIN la_oen_core[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 89.700 709.230 92.000 ;
    END
  END la_oen_core[65]
  PIN la_oen_core[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 89.700 711.530 92.000 ;
    END
  END la_oen_core[66]
  PIN la_oen_core[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 89.700 713.370 92.000 ;
    END
  END la_oen_core[67]
  PIN la_oen_core[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 89.700 715.670 92.000 ;
    END
  END la_oen_core[68]
  PIN la_oen_core[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 89.700 717.970 92.000 ;
    END
  END la_oen_core[69]
  PIN la_oen_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 89.700 580.430 92.000 ;
    END
  END la_oen_core[6]
  PIN la_oen_core[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 89.700 720.270 92.000 ;
    END
  END la_oen_core[70]
  PIN la_oen_core[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 89.700 722.110 92.000 ;
    END
  END la_oen_core[71]
  PIN la_oen_core[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 89.700 724.410 92.000 ;
    END
  END la_oen_core[72]
  PIN la_oen_core[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 89.700 726.710 92.000 ;
    END
  END la_oen_core[73]
  PIN la_oen_core[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 89.700 728.550 92.000 ;
    END
  END la_oen_core[74]
  PIN la_oen_core[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 89.700 730.850 92.000 ;
    END
  END la_oen_core[75]
  PIN la_oen_core[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 89.700 733.150 92.000 ;
    END
  END la_oen_core[76]
  PIN la_oen_core[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 89.700 735.450 92.000 ;
    END
  END la_oen_core[77]
  PIN la_oen_core[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 89.700 737.290 92.000 ;
    END
  END la_oen_core[78]
  PIN la_oen_core[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 89.700 739.590 92.000 ;
    END
  END la_oen_core[79]
  PIN la_oen_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 89.700 582.730 92.000 ;
    END
  END la_oen_core[7]
  PIN la_oen_core[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 89.700 741.890 92.000 ;
    END
  END la_oen_core[80]
  PIN la_oen_core[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 89.700 744.190 92.000 ;
    END
  END la_oen_core[81]
  PIN la_oen_core[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 89.700 746.030 92.000 ;
    END
  END la_oen_core[82]
  PIN la_oen_core[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 89.700 748.330 92.000 ;
    END
  END la_oen_core[83]
  PIN la_oen_core[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 89.700 750.630 92.000 ;
    END
  END la_oen_core[84]
  PIN la_oen_core[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 89.700 752.930 92.000 ;
    END
  END la_oen_core[85]
  PIN la_oen_core[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 89.700 754.770 92.000 ;
    END
  END la_oen_core[86]
  PIN la_oen_core[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 89.700 757.070 92.000 ;
    END
  END la_oen_core[87]
  PIN la_oen_core[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 89.700 759.370 92.000 ;
    END
  END la_oen_core[88]
  PIN la_oen_core[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 89.700 761.210 92.000 ;
    END
  END la_oen_core[89]
  PIN la_oen_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 89.700 585.030 92.000 ;
    END
  END la_oen_core[8]
  PIN la_oen_core[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 89.700 763.510 92.000 ;
    END
  END la_oen_core[90]
  PIN la_oen_core[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 89.700 765.810 92.000 ;
    END
  END la_oen_core[91]
  PIN la_oen_core[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 89.700 768.110 92.000 ;
    END
  END la_oen_core[92]
  PIN la_oen_core[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 89.700 769.950 92.000 ;
    END
  END la_oen_core[93]
  PIN la_oen_core[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 89.700 772.250 92.000 ;
    END
  END la_oen_core[94]
  PIN la_oen_core[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 89.700 774.550 92.000 ;
    END
  END la_oen_core[95]
  PIN la_oen_core[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 89.700 776.850 92.000 ;
    END
  END la_oen_core[96]
  PIN la_oen_core[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 89.700 778.690 92.000 ;
    END
  END la_oen_core[97]
  PIN la_oen_core[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 89.700 780.990 92.000 ;
    END
  END la_oen_core[98]
  PIN la_oen_core[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 89.700 783.290 92.000 ;
    END
  END la_oen_core[99]
  PIN la_oen_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 89.700 587.330 92.000 ;
    END
  END la_oen_core[9]
  PIN la_oen_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 -2.000 558.810 0.300 ;
    END
  END la_oen_mprj[0]
  PIN la_oen_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 -2.000 776.850 0.300 ;
    END
  END la_oen_mprj[100]
  PIN la_oen_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 -2.000 778.690 0.300 ;
    END
  END la_oen_mprj[101]
  PIN la_oen_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 -2.000 780.990 0.300 ;
    END
  END la_oen_mprj[102]
  PIN la_oen_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 -2.000 783.290 0.300 ;
    END
  END la_oen_mprj[103]
  PIN la_oen_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 -2.000 785.590 0.300 ;
    END
  END la_oen_mprj[104]
  PIN la_oen_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 -2.000 787.430 0.300 ;
    END
  END la_oen_mprj[105]
  PIN la_oen_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 -2.000 789.730 0.300 ;
    END
  END la_oen_mprj[106]
  PIN la_oen_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.750 -2.000 792.030 0.300 ;
    END
  END la_oen_mprj[107]
  PIN la_oen_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 -2.000 794.330 0.300 ;
    END
  END la_oen_mprj[108]
  PIN la_oen_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 -2.000 796.170 0.300 ;
    END
  END la_oen_mprj[109]
  PIN la_oen_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 -2.000 580.430 0.300 ;
    END
  END la_oen_mprj[10]
  PIN la_oen_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 -2.000 798.470 0.300 ;
    END
  END la_oen_mprj[110]
  PIN la_oen_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 -2.000 800.770 0.300 ;
    END
  END la_oen_mprj[111]
  PIN la_oen_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 -2.000 802.610 0.300 ;
    END
  END la_oen_mprj[112]
  PIN la_oen_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 -2.000 804.910 0.300 ;
    END
  END la_oen_mprj[113]
  PIN la_oen_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.930 -2.000 807.210 0.300 ;
    END
  END la_oen_mprj[114]
  PIN la_oen_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 -2.000 809.510 0.300 ;
    END
  END la_oen_mprj[115]
  PIN la_oen_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 -2.000 811.350 0.300 ;
    END
  END la_oen_mprj[116]
  PIN la_oen_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 -2.000 813.650 0.300 ;
    END
  END la_oen_mprj[117]
  PIN la_oen_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 -2.000 815.950 0.300 ;
    END
  END la_oen_mprj[118]
  PIN la_oen_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 -2.000 818.250 0.300 ;
    END
  END la_oen_mprj[119]
  PIN la_oen_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 -2.000 582.730 0.300 ;
    END
  END la_oen_mprj[11]
  PIN la_oen_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 -2.000 820.090 0.300 ;
    END
  END la_oen_mprj[120]
  PIN la_oen_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 -2.000 822.390 0.300 ;
    END
  END la_oen_mprj[121]
  PIN la_oen_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 -2.000 824.690 0.300 ;
    END
  END la_oen_mprj[122]
  PIN la_oen_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 -2.000 826.990 0.300 ;
    END
  END la_oen_mprj[123]
  PIN la_oen_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 -2.000 828.830 0.300 ;
    END
  END la_oen_mprj[124]
  PIN la_oen_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 -2.000 831.130 0.300 ;
    END
  END la_oen_mprj[125]
  PIN la_oen_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 -2.000 833.430 0.300 ;
    END
  END la_oen_mprj[126]
  PIN la_oen_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 -2.000 835.730 0.300 ;
    END
  END la_oen_mprj[127]
  PIN la_oen_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 -2.000 585.030 0.300 ;
    END
  END la_oen_mprj[12]
  PIN la_oen_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 -2.000 587.330 0.300 ;
    END
  END la_oen_mprj[13]
  PIN la_oen_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 -2.000 589.170 0.300 ;
    END
  END la_oen_mprj[14]
  PIN la_oen_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 -2.000 591.470 0.300 ;
    END
  END la_oen_mprj[15]
  PIN la_oen_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 -2.000 593.770 0.300 ;
    END
  END la_oen_mprj[16]
  PIN la_oen_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 -2.000 596.070 0.300 ;
    END
  END la_oen_mprj[17]
  PIN la_oen_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 -2.000 597.910 0.300 ;
    END
  END la_oen_mprj[18]
  PIN la_oen_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 -2.000 600.210 0.300 ;
    END
  END la_oen_mprj[19]
  PIN la_oen_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 -2.000 561.110 0.300 ;
    END
  END la_oen_mprj[1]
  PIN la_oen_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 -2.000 602.510 0.300 ;
    END
  END la_oen_mprj[20]
  PIN la_oen_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 -2.000 604.350 0.300 ;
    END
  END la_oen_mprj[21]
  PIN la_oen_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 -2.000 606.650 0.300 ;
    END
  END la_oen_mprj[22]
  PIN la_oen_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 -2.000 608.950 0.300 ;
    END
  END la_oen_mprj[23]
  PIN la_oen_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 -2.000 611.250 0.300 ;
    END
  END la_oen_mprj[24]
  PIN la_oen_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 -2.000 613.090 0.300 ;
    END
  END la_oen_mprj[25]
  PIN la_oen_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 -2.000 615.390 0.300 ;
    END
  END la_oen_mprj[26]
  PIN la_oen_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 -2.000 617.690 0.300 ;
    END
  END la_oen_mprj[27]
  PIN la_oen_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 -2.000 619.990 0.300 ;
    END
  END la_oen_mprj[28]
  PIN la_oen_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 -2.000 621.830 0.300 ;
    END
  END la_oen_mprj[29]
  PIN la_oen_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 -2.000 562.950 0.300 ;
    END
  END la_oen_mprj[2]
  PIN la_oen_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 -2.000 624.130 0.300 ;
    END
  END la_oen_mprj[30]
  PIN la_oen_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 -2.000 626.430 0.300 ;
    END
  END la_oen_mprj[31]
  PIN la_oen_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 -2.000 628.730 0.300 ;
    END
  END la_oen_mprj[32]
  PIN la_oen_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 -2.000 630.570 0.300 ;
    END
  END la_oen_mprj[33]
  PIN la_oen_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 -2.000 632.870 0.300 ;
    END
  END la_oen_mprj[34]
  PIN la_oen_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 -2.000 635.170 0.300 ;
    END
  END la_oen_mprj[35]
  PIN la_oen_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 -2.000 637.470 0.300 ;
    END
  END la_oen_mprj[36]
  PIN la_oen_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 -2.000 639.310 0.300 ;
    END
  END la_oen_mprj[37]
  PIN la_oen_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 -2.000 641.610 0.300 ;
    END
  END la_oen_mprj[38]
  PIN la_oen_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 -2.000 643.910 0.300 ;
    END
  END la_oen_mprj[39]
  PIN la_oen_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 -2.000 565.250 0.300 ;
    END
  END la_oen_mprj[3]
  PIN la_oen_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 -2.000 645.750 0.300 ;
    END
  END la_oen_mprj[40]
  PIN la_oen_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 -2.000 648.050 0.300 ;
    END
  END la_oen_mprj[41]
  PIN la_oen_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 -2.000 650.350 0.300 ;
    END
  END la_oen_mprj[42]
  PIN la_oen_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 -2.000 652.650 0.300 ;
    END
  END la_oen_mprj[43]
  PIN la_oen_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 -2.000 654.490 0.300 ;
    END
  END la_oen_mprj[44]
  PIN la_oen_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 -2.000 656.790 0.300 ;
    END
  END la_oen_mprj[45]
  PIN la_oen_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 -2.000 659.090 0.300 ;
    END
  END la_oen_mprj[46]
  PIN la_oen_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 -2.000 661.390 0.300 ;
    END
  END la_oen_mprj[47]
  PIN la_oen_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.950 -2.000 663.230 0.300 ;
    END
  END la_oen_mprj[48]
  PIN la_oen_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 -2.000 665.530 0.300 ;
    END
  END la_oen_mprj[49]
  PIN la_oen_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 -2.000 567.550 0.300 ;
    END
  END la_oen_mprj[4]
  PIN la_oen_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 -2.000 667.830 0.300 ;
    END
  END la_oen_mprj[50]
  PIN la_oen_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 -2.000 670.130 0.300 ;
    END
  END la_oen_mprj[51]
  PIN la_oen_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 -2.000 671.970 0.300 ;
    END
  END la_oen_mprj[52]
  PIN la_oen_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 -2.000 674.270 0.300 ;
    END
  END la_oen_mprj[53]
  PIN la_oen_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 -2.000 676.570 0.300 ;
    END
  END la_oen_mprj[54]
  PIN la_oen_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 -2.000 678.870 0.300 ;
    END
  END la_oen_mprj[55]
  PIN la_oen_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 -2.000 680.710 0.300 ;
    END
  END la_oen_mprj[56]
  PIN la_oen_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 -2.000 683.010 0.300 ;
    END
  END la_oen_mprj[57]
  PIN la_oen_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 -2.000 685.310 0.300 ;
    END
  END la_oen_mprj[58]
  PIN la_oen_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 -2.000 687.150 0.300 ;
    END
  END la_oen_mprj[59]
  PIN la_oen_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 -2.000 569.850 0.300 ;
    END
  END la_oen_mprj[5]
  PIN la_oen_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 -2.000 689.450 0.300 ;
    END
  END la_oen_mprj[60]
  PIN la_oen_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 -2.000 691.750 0.300 ;
    END
  END la_oen_mprj[61]
  PIN la_oen_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 -2.000 694.050 0.300 ;
    END
  END la_oen_mprj[62]
  PIN la_oen_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 -2.000 695.890 0.300 ;
    END
  END la_oen_mprj[63]
  PIN la_oen_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 -2.000 698.190 0.300 ;
    END
  END la_oen_mprj[64]
  PIN la_oen_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 -2.000 700.490 0.300 ;
    END
  END la_oen_mprj[65]
  PIN la_oen_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 -2.000 702.790 0.300 ;
    END
  END la_oen_mprj[66]
  PIN la_oen_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 -2.000 704.630 0.300 ;
    END
  END la_oen_mprj[67]
  PIN la_oen_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 -2.000 706.930 0.300 ;
    END
  END la_oen_mprj[68]
  PIN la_oen_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 -2.000 709.230 0.300 ;
    END
  END la_oen_mprj[69]
  PIN la_oen_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 -2.000 571.690 0.300 ;
    END
  END la_oen_mprj[6]
  PIN la_oen_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 -2.000 711.530 0.300 ;
    END
  END la_oen_mprj[70]
  PIN la_oen_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 -2.000 713.370 0.300 ;
    END
  END la_oen_mprj[71]
  PIN la_oen_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 -2.000 715.670 0.300 ;
    END
  END la_oen_mprj[72]
  PIN la_oen_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 -2.000 717.970 0.300 ;
    END
  END la_oen_mprj[73]
  PIN la_oen_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 -2.000 720.270 0.300 ;
    END
  END la_oen_mprj[74]
  PIN la_oen_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 -2.000 722.110 0.300 ;
    END
  END la_oen_mprj[75]
  PIN la_oen_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 -2.000 724.410 0.300 ;
    END
  END la_oen_mprj[76]
  PIN la_oen_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 -2.000 726.710 0.300 ;
    END
  END la_oen_mprj[77]
  PIN la_oen_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 -2.000 728.550 0.300 ;
    END
  END la_oen_mprj[78]
  PIN la_oen_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 -2.000 730.850 0.300 ;
    END
  END la_oen_mprj[79]
  PIN la_oen_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 -2.000 573.990 0.300 ;
    END
  END la_oen_mprj[7]
  PIN la_oen_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 -2.000 733.150 0.300 ;
    END
  END la_oen_mprj[80]
  PIN la_oen_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 -2.000 735.450 0.300 ;
    END
  END la_oen_mprj[81]
  PIN la_oen_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 -2.000 737.290 0.300 ;
    END
  END la_oen_mprj[82]
  PIN la_oen_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 -2.000 739.590 0.300 ;
    END
  END la_oen_mprj[83]
  PIN la_oen_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 -2.000 741.890 0.300 ;
    END
  END la_oen_mprj[84]
  PIN la_oen_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 -2.000 744.190 0.300 ;
    END
  END la_oen_mprj[85]
  PIN la_oen_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 -2.000 746.030 0.300 ;
    END
  END la_oen_mprj[86]
  PIN la_oen_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 -2.000 748.330 0.300 ;
    END
  END la_oen_mprj[87]
  PIN la_oen_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 -2.000 750.630 0.300 ;
    END
  END la_oen_mprj[88]
  PIN la_oen_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 -2.000 752.930 0.300 ;
    END
  END la_oen_mprj[89]
  PIN la_oen_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 -2.000 576.290 0.300 ;
    END
  END la_oen_mprj[8]
  PIN la_oen_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 -2.000 754.770 0.300 ;
    END
  END la_oen_mprj[90]
  PIN la_oen_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 -2.000 757.070 0.300 ;
    END
  END la_oen_mprj[91]
  PIN la_oen_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 -2.000 759.370 0.300 ;
    END
  END la_oen_mprj[92]
  PIN la_oen_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 -2.000 761.210 0.300 ;
    END
  END la_oen_mprj[93]
  PIN la_oen_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 -2.000 763.510 0.300 ;
    END
  END la_oen_mprj[94]
  PIN la_oen_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 -2.000 765.810 0.300 ;
    END
  END la_oen_mprj[95]
  PIN la_oen_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 -2.000 768.110 0.300 ;
    END
  END la_oen_mprj[96]
  PIN la_oen_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 -2.000 769.950 0.300 ;
    END
  END la_oen_mprj[97]
  PIN la_oen_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 -2.000 772.250 0.300 ;
    END
  END la_oen_mprj[98]
  PIN la_oen_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 -2.000 774.550 0.300 ;
    END
  END la_oen_mprj[99]
  PIN la_oen_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 -2.000 578.590 0.300 ;
    END
  END la_oen_mprj[9]
  PIN mprj_adr_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 -2.000 844.010 0.300 ;
    END
  END mprj_adr_o_core[0]
  PIN mprj_adr_o_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 -2.000 896.450 0.300 ;
    END
  END mprj_adr_o_core[10]
  PIN mprj_adr_o_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 -2.000 901.050 0.300 ;
    END
  END mprj_adr_o_core[11]
  PIN mprj_adr_o_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 -2.000 905.190 0.300 ;
    END
  END mprj_adr_o_core[12]
  PIN mprj_adr_o_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 -2.000 909.790 0.300 ;
    END
  END mprj_adr_o_core[13]
  PIN mprj_adr_o_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 -2.000 913.930 0.300 ;
    END
  END mprj_adr_o_core[14]
  PIN mprj_adr_o_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 -2.000 918.530 0.300 ;
    END
  END mprj_adr_o_core[15]
  PIN mprj_adr_o_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 -2.000 922.670 0.300 ;
    END
  END mprj_adr_o_core[16]
  PIN mprj_adr_o_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.530 -2.000 926.810 0.300 ;
    END
  END mprj_adr_o_core[17]
  PIN mprj_adr_o_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 -2.000 931.410 0.300 ;
    END
  END mprj_adr_o_core[18]
  PIN mprj_adr_o_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.270 -2.000 935.550 0.300 ;
    END
  END mprj_adr_o_core[19]
  PIN mprj_adr_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 -2.000 850.910 0.300 ;
    END
  END mprj_adr_o_core[1]
  PIN mprj_adr_o_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 -2.000 940.150 0.300 ;
    END
  END mprj_adr_o_core[20]
  PIN mprj_adr_o_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 -2.000 944.290 0.300 ;
    END
  END mprj_adr_o_core[21]
  PIN mprj_adr_o_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 -2.000 948.890 0.300 ;
    END
  END mprj_adr_o_core[22]
  PIN mprj_adr_o_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 -2.000 953.030 0.300 ;
    END
  END mprj_adr_o_core[23]
  PIN mprj_adr_o_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 -2.000 957.630 0.300 ;
    END
  END mprj_adr_o_core[24]
  PIN mprj_adr_o_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 -2.000 961.770 0.300 ;
    END
  END mprj_adr_o_core[25]
  PIN mprj_adr_o_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 -2.000 966.370 0.300 ;
    END
  END mprj_adr_o_core[26]
  PIN mprj_adr_o_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 -2.000 970.510 0.300 ;
    END
  END mprj_adr_o_core[27]
  PIN mprj_adr_o_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.830 -2.000 975.110 0.300 ;
    END
  END mprj_adr_o_core[28]
  PIN mprj_adr_o_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 -2.000 979.250 0.300 ;
    END
  END mprj_adr_o_core[29]
  PIN mprj_adr_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070 -2.000 857.350 0.300 ;
    END
  END mprj_adr_o_core[2]
  PIN mprj_adr_o_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.570 -2.000 983.850 0.300 ;
    END
  END mprj_adr_o_core[30]
  PIN mprj_adr_o_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.710 -2.000 987.990 0.300 ;
    END
  END mprj_adr_o_core[31]
  PIN mprj_adr_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 -2.000 863.790 0.300 ;
    END
  END mprj_adr_o_core[3]
  PIN mprj_adr_o_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 -2.000 870.230 0.300 ;
    END
  END mprj_adr_o_core[4]
  PIN mprj_adr_o_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 -2.000 874.830 0.300 ;
    END
  END mprj_adr_o_core[5]
  PIN mprj_adr_o_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 -2.000 878.970 0.300 ;
    END
  END mprj_adr_o_core[6]
  PIN mprj_adr_o_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 -2.000 883.570 0.300 ;
    END
  END mprj_adr_o_core[7]
  PIN mprj_adr_o_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 -2.000 887.710 0.300 ;
    END
  END mprj_adr_o_core[8]
  PIN mprj_adr_o_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 -2.000 892.310 0.300 ;
    END
  END mprj_adr_o_core[9]
  PIN mprj_adr_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 89.700 852.750 92.000 ;
    END
  END mprj_adr_o_user[0]
  PIN mprj_adr_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 89.700 905.190 92.000 ;
    END
  END mprj_adr_o_user[10]
  PIN mprj_adr_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 89.700 909.790 92.000 ;
    END
  END mprj_adr_o_user[11]
  PIN mprj_adr_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 89.700 913.930 92.000 ;
    END
  END mprj_adr_o_user[12]
  PIN mprj_adr_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 89.700 918.530 92.000 ;
    END
  END mprj_adr_o_user[13]
  PIN mprj_adr_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 89.700 922.670 92.000 ;
    END
  END mprj_adr_o_user[14]
  PIN mprj_adr_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.530 89.700 926.810 92.000 ;
    END
  END mprj_adr_o_user[15]
  PIN mprj_adr_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 89.700 931.410 92.000 ;
    END
  END mprj_adr_o_user[16]
  PIN mprj_adr_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.270 89.700 935.550 92.000 ;
    END
  END mprj_adr_o_user[17]
  PIN mprj_adr_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 89.700 940.150 92.000 ;
    END
  END mprj_adr_o_user[18]
  PIN mprj_adr_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 89.700 944.290 92.000 ;
    END
  END mprj_adr_o_user[19]
  PIN mprj_adr_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 89.700 859.650 92.000 ;
    END
  END mprj_adr_o_user[1]
  PIN mprj_adr_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 89.700 948.890 92.000 ;
    END
  END mprj_adr_o_user[20]
  PIN mprj_adr_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 89.700 953.030 92.000 ;
    END
  END mprj_adr_o_user[21]
  PIN mprj_adr_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 89.700 957.630 92.000 ;
    END
  END mprj_adr_o_user[22]
  PIN mprj_adr_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 89.700 961.770 92.000 ;
    END
  END mprj_adr_o_user[23]
  PIN mprj_adr_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 89.700 966.370 92.000 ;
    END
  END mprj_adr_o_user[24]
  PIN mprj_adr_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 89.700 970.510 92.000 ;
    END
  END mprj_adr_o_user[25]
  PIN mprj_adr_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.830 89.700 975.110 92.000 ;
    END
  END mprj_adr_o_user[26]
  PIN mprj_adr_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 89.700 979.250 92.000 ;
    END
  END mprj_adr_o_user[27]
  PIN mprj_adr_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.570 89.700 983.850 92.000 ;
    END
  END mprj_adr_o_user[28]
  PIN mprj_adr_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.710 89.700 987.990 92.000 ;
    END
  END mprj_adr_o_user[29]
  PIN mprj_adr_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 89.700 866.090 92.000 ;
    END
  END mprj_adr_o_user[2]
  PIN mprj_adr_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 89.700 992.590 92.000 ;
    END
  END mprj_adr_o_user[30]
  PIN mprj_adr_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 89.700 996.730 92.000 ;
    END
  END mprj_adr_o_user[31]
  PIN mprj_adr_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 89.700 872.530 92.000 ;
    END
  END mprj_adr_o_user[3]
  PIN mprj_adr_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 89.700 878.970 92.000 ;
    END
  END mprj_adr_o_user[4]
  PIN mprj_adr_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 89.700 883.570 92.000 ;
    END
  END mprj_adr_o_user[5]
  PIN mprj_adr_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 89.700 887.710 92.000 ;
    END
  END mprj_adr_o_user[6]
  PIN mprj_adr_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 89.700 892.310 92.000 ;
    END
  END mprj_adr_o_user[7]
  PIN mprj_adr_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 89.700 896.450 92.000 ;
    END
  END mprj_adr_o_user[8]
  PIN mprj_adr_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 89.700 901.050 92.000 ;
    END
  END mprj_adr_o_user[9]
  PIN mprj_cyc_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 -2.000 837.570 0.300 ;
    END
  END mprj_cyc_o_core
  PIN mprj_cyc_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 89.700 846.310 92.000 ;
    END
  END mprj_cyc_o_user
  PIN mprj_dat_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 -2.000 846.310 0.300 ;
    END
  END mprj_dat_o_core[0]
  PIN mprj_dat_o_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 -2.000 898.750 0.300 ;
    END
  END mprj_dat_o_core[10]
  PIN mprj_dat_o_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 -2.000 902.890 0.300 ;
    END
  END mprj_dat_o_core[11]
  PIN mprj_dat_o_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 -2.000 907.490 0.300 ;
    END
  END mprj_dat_o_core[12]
  PIN mprj_dat_o_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 -2.000 911.630 0.300 ;
    END
  END mprj_dat_o_core[13]
  PIN mprj_dat_o_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 -2.000 916.230 0.300 ;
    END
  END mprj_dat_o_core[14]
  PIN mprj_dat_o_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 -2.000 920.370 0.300 ;
    END
  END mprj_dat_o_core[15]
  PIN mprj_dat_o_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 -2.000 924.970 0.300 ;
    END
  END mprj_dat_o_core[16]
  PIN mprj_dat_o_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 -2.000 929.110 0.300 ;
    END
  END mprj_dat_o_core[17]
  PIN mprj_dat_o_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 -2.000 933.710 0.300 ;
    END
  END mprj_dat_o_core[18]
  PIN mprj_dat_o_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 -2.000 937.850 0.300 ;
    END
  END mprj_dat_o_core[19]
  PIN mprj_dat_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 -2.000 852.750 0.300 ;
    END
  END mprj_dat_o_core[1]
  PIN mprj_dat_o_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 -2.000 942.450 0.300 ;
    END
  END mprj_dat_o_core[20]
  PIN mprj_dat_o_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 -2.000 946.590 0.300 ;
    END
  END mprj_dat_o_core[21]
  PIN mprj_dat_o_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 -2.000 951.190 0.300 ;
    END
  END mprj_dat_o_core[22]
  PIN mprj_dat_o_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 -2.000 955.330 0.300 ;
    END
  END mprj_dat_o_core[23]
  PIN mprj_dat_o_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 -2.000 959.930 0.300 ;
    END
  END mprj_dat_o_core[24]
  PIN mprj_dat_o_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 -2.000 964.070 0.300 ;
    END
  END mprj_dat_o_core[25]
  PIN mprj_dat_o_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 -2.000 968.210 0.300 ;
    END
  END mprj_dat_o_core[26]
  PIN mprj_dat_o_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 -2.000 972.810 0.300 ;
    END
  END mprj_dat_o_core[27]
  PIN mprj_dat_o_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 -2.000 976.950 0.300 ;
    END
  END mprj_dat_o_core[28]
  PIN mprj_dat_o_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 -2.000 981.550 0.300 ;
    END
  END mprj_dat_o_core[29]
  PIN mprj_dat_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 -2.000 859.650 0.300 ;
    END
  END mprj_dat_o_core[2]
  PIN mprj_dat_o_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 -2.000 985.690 0.300 ;
    END
  END mprj_dat_o_core[30]
  PIN mprj_dat_o_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 -2.000 990.290 0.300 ;
    END
  END mprj_dat_o_core[31]
  PIN mprj_dat_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 -2.000 866.090 0.300 ;
    END
  END mprj_dat_o_core[3]
  PIN mprj_dat_o_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 -2.000 872.530 0.300 ;
    END
  END mprj_dat_o_core[4]
  PIN mprj_dat_o_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.850 -2.000 877.130 0.300 ;
    END
  END mprj_dat_o_core[5]
  PIN mprj_dat_o_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 -2.000 881.270 0.300 ;
    END
  END mprj_dat_o_core[6]
  PIN mprj_dat_o_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 -2.000 885.410 0.300 ;
    END
  END mprj_dat_o_core[7]
  PIN mprj_dat_o_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 -2.000 890.010 0.300 ;
    END
  END mprj_dat_o_core[8]
  PIN mprj_dat_o_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 -2.000 894.150 0.300 ;
    END
  END mprj_dat_o_core[9]
  PIN mprj_dat_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 89.700 855.050 92.000 ;
    END
  END mprj_dat_o_user[0]
  PIN mprj_dat_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 89.700 907.490 92.000 ;
    END
  END mprj_dat_o_user[10]
  PIN mprj_dat_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 89.700 911.630 92.000 ;
    END
  END mprj_dat_o_user[11]
  PIN mprj_dat_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 89.700 916.230 92.000 ;
    END
  END mprj_dat_o_user[12]
  PIN mprj_dat_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 89.700 920.370 92.000 ;
    END
  END mprj_dat_o_user[13]
  PIN mprj_dat_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 89.700 924.970 92.000 ;
    END
  END mprj_dat_o_user[14]
  PIN mprj_dat_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 89.700 929.110 92.000 ;
    END
  END mprj_dat_o_user[15]
  PIN mprj_dat_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 89.700 933.710 92.000 ;
    END
  END mprj_dat_o_user[16]
  PIN mprj_dat_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 89.700 937.850 92.000 ;
    END
  END mprj_dat_o_user[17]
  PIN mprj_dat_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 89.700 942.450 92.000 ;
    END
  END mprj_dat_o_user[18]
  PIN mprj_dat_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 89.700 946.590 92.000 ;
    END
  END mprj_dat_o_user[19]
  PIN mprj_dat_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 89.700 861.490 92.000 ;
    END
  END mprj_dat_o_user[1]
  PIN mprj_dat_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 89.700 951.190 92.000 ;
    END
  END mprj_dat_o_user[20]
  PIN mprj_dat_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 89.700 955.330 92.000 ;
    END
  END mprj_dat_o_user[21]
  PIN mprj_dat_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 89.700 959.930 92.000 ;
    END
  END mprj_dat_o_user[22]
  PIN mprj_dat_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 89.700 964.070 92.000 ;
    END
  END mprj_dat_o_user[23]
  PIN mprj_dat_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 89.700 968.210 92.000 ;
    END
  END mprj_dat_o_user[24]
  PIN mprj_dat_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 89.700 972.810 92.000 ;
    END
  END mprj_dat_o_user[25]
  PIN mprj_dat_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 89.700 976.950 92.000 ;
    END
  END mprj_dat_o_user[26]
  PIN mprj_dat_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 89.700 981.550 92.000 ;
    END
  END mprj_dat_o_user[27]
  PIN mprj_dat_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 89.700 985.690 92.000 ;
    END
  END mprj_dat_o_user[28]
  PIN mprj_dat_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 89.700 990.290 92.000 ;
    END
  END mprj_dat_o_user[29]
  PIN mprj_dat_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 89.700 868.390 92.000 ;
    END
  END mprj_dat_o_user[2]
  PIN mprj_dat_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 89.700 994.430 92.000 ;
    END
  END mprj_dat_o_user[30]
  PIN mprj_dat_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 89.700 999.030 92.000 ;
    END
  END mprj_dat_o_user[31]
  PIN mprj_dat_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 89.700 874.830 92.000 ;
    END
  END mprj_dat_o_user[3]
  PIN mprj_dat_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 89.700 881.270 92.000 ;
    END
  END mprj_dat_o_user[4]
  PIN mprj_dat_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 89.700 885.410 92.000 ;
    END
  END mprj_dat_o_user[5]
  PIN mprj_dat_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 89.700 890.010 92.000 ;
    END
  END mprj_dat_o_user[6]
  PIN mprj_dat_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 89.700 894.150 92.000 ;
    END
  END mprj_dat_o_user[7]
  PIN mprj_dat_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 89.700 898.750 92.000 ;
    END
  END mprj_dat_o_user[8]
  PIN mprj_dat_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 89.700 902.890 92.000 ;
    END
  END mprj_dat_o_user[9]
  PIN mprj_sel_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 -2.000 848.610 0.300 ;
    END
  END mprj_sel_o_core[0]
  PIN mprj_sel_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 -2.000 855.050 0.300 ;
    END
  END mprj_sel_o_core[1]
  PIN mprj_sel_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 -2.000 861.490 0.300 ;
    END
  END mprj_sel_o_core[2]
  PIN mprj_sel_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 -2.000 868.390 0.300 ;
    END
  END mprj_sel_o_core[3]
  PIN mprj_sel_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070 89.700 857.350 92.000 ;
    END
  END mprj_sel_o_user[0]
  PIN mprj_sel_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 89.700 863.790 92.000 ;
    END
  END mprj_sel_o_user[1]
  PIN mprj_sel_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 89.700 870.230 92.000 ;
    END
  END mprj_sel_o_user[2]
  PIN mprj_sel_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.850 89.700 877.130 92.000 ;
    END
  END mprj_sel_o_user[3]
  PIN mprj_stb_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 -2.000 839.870 0.300 ;
    END
  END mprj_stb_o_core
  PIN mprj_stb_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 89.700 848.610 92.000 ;
    END
  END mprj_stb_o_user
  PIN mprj_we_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 -2.000 842.170 0.300 ;
    END
  END mprj_we_o_core
  PIN mprj_we_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 89.700 850.910 92.000 ;
    END
  END mprj_we_o_user
  PIN user1_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 -2.000 992.590 0.300 ;
    END
  END user1_vcc_powergood
  PIN user1_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 -2.000 994.430 0.300 ;
    END
  END user1_vdd_powergood
  PIN user2_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 -2.000 996.730 0.300 ;
    END
  END user2_vcc_powergood
  PIN user2_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 -2.000 999.030 0.300 ;
    END
  END user2_vdd_powergood
  PIN user_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 89.700 1.290 92.000 ;
    END
  END user_clock
  PIN user_clock2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 89.700 3.130 92.000 ;
    END
  END user_clock2
  PIN user_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 89.700 5.430 92.000 ;
    END
  END user_reset
  PIN user_resetn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 89.700 7.730 92.000 ;
    END
  END user_resetn
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -1.930 90.870 1001.510 91.770 ;
        RECT -1.930 -2.010 1001.510 -1.110 ;
      LAYER via3 ;
        RECT -1.840 91.360 -1.520 91.680 ;
        RECT -1.440 91.360 -1.120 91.680 ;
        RECT 20.160 91.360 20.480 91.680 ;
        RECT 20.560 91.360 20.880 91.680 ;
        RECT 170.160 91.360 170.480 91.680 ;
        RECT 170.560 91.360 170.880 91.680 ;
        RECT 320.160 91.360 320.480 91.680 ;
        RECT 320.560 91.360 320.880 91.680 ;
        RECT 470.160 91.360 470.480 91.680 ;
        RECT 470.560 91.360 470.880 91.680 ;
        RECT 620.160 91.360 620.480 91.680 ;
        RECT 620.560 91.360 620.880 91.680 ;
        RECT 770.160 91.360 770.480 91.680 ;
        RECT 770.560 91.360 770.880 91.680 ;
        RECT 920.160 91.360 920.480 91.680 ;
        RECT 920.560 91.360 920.880 91.680 ;
        RECT 1000.700 91.360 1001.020 91.680 ;
        RECT 1001.100 91.360 1001.420 91.680 ;
        RECT -1.840 90.960 -1.520 91.280 ;
        RECT -1.440 90.960 -1.120 91.280 ;
        RECT 20.160 90.960 20.480 91.280 ;
        RECT 20.560 90.960 20.880 91.280 ;
        RECT 170.160 90.960 170.480 91.280 ;
        RECT 170.560 90.960 170.880 91.280 ;
        RECT 320.160 90.960 320.480 91.280 ;
        RECT 320.560 90.960 320.880 91.280 ;
        RECT 470.160 90.960 470.480 91.280 ;
        RECT 470.560 90.960 470.880 91.280 ;
        RECT 620.160 90.960 620.480 91.280 ;
        RECT 620.560 90.960 620.880 91.280 ;
        RECT 770.160 90.960 770.480 91.280 ;
        RECT 770.560 90.960 770.880 91.280 ;
        RECT 920.160 90.960 920.480 91.280 ;
        RECT 920.560 90.960 920.880 91.280 ;
        RECT 1000.700 90.960 1001.020 91.280 ;
        RECT 1001.100 90.960 1001.420 91.280 ;
        RECT -1.840 -1.520 -1.520 -1.200 ;
        RECT -1.440 -1.520 -1.120 -1.200 ;
        RECT 20.160 -1.520 20.480 -1.200 ;
        RECT 20.560 -1.520 20.880 -1.200 ;
        RECT 170.160 -1.520 170.480 -1.200 ;
        RECT 170.560 -1.520 170.880 -1.200 ;
        RECT 320.160 -1.520 320.480 -1.200 ;
        RECT 320.560 -1.520 320.880 -1.200 ;
        RECT 470.160 -1.520 470.480 -1.200 ;
        RECT 470.560 -1.520 470.880 -1.200 ;
        RECT 620.160 -1.520 620.480 -1.200 ;
        RECT 620.560 -1.520 620.880 -1.200 ;
        RECT 770.160 -1.520 770.480 -1.200 ;
        RECT 770.560 -1.520 770.880 -1.200 ;
        RECT 920.160 -1.520 920.480 -1.200 ;
        RECT 920.560 -1.520 920.880 -1.200 ;
        RECT 1000.700 -1.520 1001.020 -1.200 ;
        RECT 1001.100 -1.520 1001.420 -1.200 ;
        RECT -1.840 -1.920 -1.520 -1.600 ;
        RECT -1.440 -1.920 -1.120 -1.600 ;
        RECT 20.160 -1.920 20.480 -1.600 ;
        RECT 20.560 -1.920 20.880 -1.600 ;
        RECT 170.160 -1.920 170.480 -1.600 ;
        RECT 170.560 -1.920 170.880 -1.600 ;
        RECT 320.160 -1.920 320.480 -1.600 ;
        RECT 320.560 -1.920 320.880 -1.600 ;
        RECT 470.160 -1.920 470.480 -1.600 ;
        RECT 470.560 -1.920 470.880 -1.600 ;
        RECT 620.160 -1.920 620.480 -1.600 ;
        RECT 620.560 -1.920 620.880 -1.600 ;
        RECT 770.160 -1.920 770.480 -1.600 ;
        RECT 770.560 -1.920 770.880 -1.600 ;
        RECT 920.160 -1.920 920.480 -1.600 ;
        RECT 920.560 -1.920 920.880 -1.600 ;
        RECT 1000.700 -1.920 1001.020 -1.600 ;
        RECT 1001.100 -1.920 1001.420 -1.600 ;
      LAYER met4 ;
        RECT -1.930 -2.010 -1.030 91.770 ;
        RECT 20.070 89.700 20.970 93.090 ;
        RECT 170.070 89.700 170.970 93.090 ;
        RECT 320.070 89.700 320.970 93.090 ;
        RECT 470.070 89.700 470.970 93.090 ;
        RECT 620.070 89.700 620.970 93.090 ;
        RECT 770.070 89.700 770.970 93.090 ;
        RECT 920.070 89.700 920.970 93.090 ;
        RECT 20.070 -3.330 20.970 0.300 ;
        RECT 170.070 -3.330 170.970 0.300 ;
        RECT 320.070 -3.330 320.970 0.300 ;
        RECT 470.070 -3.330 470.970 0.300 ;
        RECT 620.070 -3.330 620.970 0.300 ;
        RECT 770.070 -3.330 770.970 0.300 ;
        RECT 920.070 -3.330 920.970 0.300 ;
        RECT 1000.610 -2.010 1001.510 91.770 ;
    END
  END vccd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -3.250 92.190 1002.830 93.090 ;
        RECT -3.250 -3.330 1002.830 -2.430 ;
      LAYER via3 ;
        RECT -3.160 92.680 -2.840 93.000 ;
        RECT -2.760 92.680 -2.440 93.000 ;
        RECT 95.160 92.680 95.480 93.000 ;
        RECT 95.560 92.680 95.880 93.000 ;
        RECT 245.160 92.680 245.480 93.000 ;
        RECT 245.560 92.680 245.880 93.000 ;
        RECT 395.160 92.680 395.480 93.000 ;
        RECT 395.560 92.680 395.880 93.000 ;
        RECT 545.160 92.680 545.480 93.000 ;
        RECT 545.560 92.680 545.880 93.000 ;
        RECT 695.160 92.680 695.480 93.000 ;
        RECT 695.560 92.680 695.880 93.000 ;
        RECT 845.160 92.680 845.480 93.000 ;
        RECT 845.560 92.680 845.880 93.000 ;
        RECT 1002.020 92.680 1002.340 93.000 ;
        RECT 1002.420 92.680 1002.740 93.000 ;
        RECT -3.160 92.280 -2.840 92.600 ;
        RECT -2.760 92.280 -2.440 92.600 ;
        RECT 95.160 92.280 95.480 92.600 ;
        RECT 95.560 92.280 95.880 92.600 ;
        RECT 245.160 92.280 245.480 92.600 ;
        RECT 245.560 92.280 245.880 92.600 ;
        RECT 395.160 92.280 395.480 92.600 ;
        RECT 395.560 92.280 395.880 92.600 ;
        RECT 545.160 92.280 545.480 92.600 ;
        RECT 545.560 92.280 545.880 92.600 ;
        RECT 695.160 92.280 695.480 92.600 ;
        RECT 695.560 92.280 695.880 92.600 ;
        RECT 845.160 92.280 845.480 92.600 ;
        RECT 845.560 92.280 845.880 92.600 ;
        RECT 1002.020 92.280 1002.340 92.600 ;
        RECT 1002.420 92.280 1002.740 92.600 ;
        RECT -3.160 -2.840 -2.840 -2.520 ;
        RECT -2.760 -2.840 -2.440 -2.520 ;
        RECT 95.160 -2.840 95.480 -2.520 ;
        RECT 95.560 -2.840 95.880 -2.520 ;
        RECT 245.160 -2.840 245.480 -2.520 ;
        RECT 245.560 -2.840 245.880 -2.520 ;
        RECT 395.160 -2.840 395.480 -2.520 ;
        RECT 395.560 -2.840 395.880 -2.520 ;
        RECT 545.160 -2.840 545.480 -2.520 ;
        RECT 545.560 -2.840 545.880 -2.520 ;
        RECT 695.160 -2.840 695.480 -2.520 ;
        RECT 695.560 -2.840 695.880 -2.520 ;
        RECT 845.160 -2.840 845.480 -2.520 ;
        RECT 845.560 -2.840 845.880 -2.520 ;
        RECT 1002.020 -2.840 1002.340 -2.520 ;
        RECT 1002.420 -2.840 1002.740 -2.520 ;
        RECT -3.160 -3.240 -2.840 -2.920 ;
        RECT -2.760 -3.240 -2.440 -2.920 ;
        RECT 95.160 -3.240 95.480 -2.920 ;
        RECT 95.560 -3.240 95.880 -2.920 ;
        RECT 245.160 -3.240 245.480 -2.920 ;
        RECT 245.560 -3.240 245.880 -2.920 ;
        RECT 395.160 -3.240 395.480 -2.920 ;
        RECT 395.560 -3.240 395.880 -2.920 ;
        RECT 545.160 -3.240 545.480 -2.920 ;
        RECT 545.560 -3.240 545.880 -2.920 ;
        RECT 695.160 -3.240 695.480 -2.920 ;
        RECT 695.560 -3.240 695.880 -2.920 ;
        RECT 845.160 -3.240 845.480 -2.920 ;
        RECT 845.560 -3.240 845.880 -2.920 ;
        RECT 1002.020 -3.240 1002.340 -2.920 ;
        RECT 1002.420 -3.240 1002.740 -2.920 ;
      LAYER met4 ;
        RECT -3.250 -3.330 -2.350 93.090 ;
        RECT 95.070 89.700 95.970 93.090 ;
        RECT 245.070 89.700 245.970 93.090 ;
        RECT 395.070 89.700 395.970 93.090 ;
        RECT 545.070 89.700 545.970 93.090 ;
        RECT 695.070 89.700 695.970 93.090 ;
        RECT 845.070 89.700 845.970 93.090 ;
        RECT 95.070 -3.330 95.970 0.300 ;
        RECT 245.070 -3.330 245.970 0.300 ;
        RECT 395.070 -3.330 395.970 0.300 ;
        RECT 545.070 -3.330 545.970 0.300 ;
        RECT 695.070 -3.330 695.970 0.300 ;
        RECT 845.070 -3.330 845.970 0.300 ;
        RECT 1001.930 -3.330 1002.830 93.090 ;
    END
  END vssd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -4.570 93.510 1004.150 94.410 ;
        RECT -4.570 -4.650 1004.150 -3.750 ;
      LAYER via3 ;
        RECT -4.480 94.000 -4.160 94.320 ;
        RECT -4.080 94.000 -3.760 94.320 ;
        RECT 24.260 94.000 24.580 94.320 ;
        RECT 24.660 94.000 24.980 94.320 ;
        RECT 174.260 94.000 174.580 94.320 ;
        RECT 174.660 94.000 174.980 94.320 ;
        RECT 324.260 94.000 324.580 94.320 ;
        RECT 324.660 94.000 324.980 94.320 ;
        RECT 474.260 94.000 474.580 94.320 ;
        RECT 474.660 94.000 474.980 94.320 ;
        RECT 624.260 94.000 624.580 94.320 ;
        RECT 624.660 94.000 624.980 94.320 ;
        RECT 774.260 94.000 774.580 94.320 ;
        RECT 774.660 94.000 774.980 94.320 ;
        RECT 924.260 94.000 924.580 94.320 ;
        RECT 924.660 94.000 924.980 94.320 ;
        RECT 1003.340 94.000 1003.660 94.320 ;
        RECT 1003.740 94.000 1004.060 94.320 ;
        RECT -4.480 93.600 -4.160 93.920 ;
        RECT -4.080 93.600 -3.760 93.920 ;
        RECT 24.260 93.600 24.580 93.920 ;
        RECT 24.660 93.600 24.980 93.920 ;
        RECT 174.260 93.600 174.580 93.920 ;
        RECT 174.660 93.600 174.980 93.920 ;
        RECT 324.260 93.600 324.580 93.920 ;
        RECT 324.660 93.600 324.980 93.920 ;
        RECT 474.260 93.600 474.580 93.920 ;
        RECT 474.660 93.600 474.980 93.920 ;
        RECT 624.260 93.600 624.580 93.920 ;
        RECT 624.660 93.600 624.980 93.920 ;
        RECT 774.260 93.600 774.580 93.920 ;
        RECT 774.660 93.600 774.980 93.920 ;
        RECT 924.260 93.600 924.580 93.920 ;
        RECT 924.660 93.600 924.980 93.920 ;
        RECT 1003.340 93.600 1003.660 93.920 ;
        RECT 1003.740 93.600 1004.060 93.920 ;
        RECT -4.480 -4.160 -4.160 -3.840 ;
        RECT -4.080 -4.160 -3.760 -3.840 ;
        RECT 24.260 -4.160 24.580 -3.840 ;
        RECT 24.660 -4.160 24.980 -3.840 ;
        RECT 174.260 -4.160 174.580 -3.840 ;
        RECT 174.660 -4.160 174.980 -3.840 ;
        RECT 324.260 -4.160 324.580 -3.840 ;
        RECT 324.660 -4.160 324.980 -3.840 ;
        RECT 474.260 -4.160 474.580 -3.840 ;
        RECT 474.660 -4.160 474.980 -3.840 ;
        RECT 624.260 -4.160 624.580 -3.840 ;
        RECT 624.660 -4.160 624.980 -3.840 ;
        RECT 774.260 -4.160 774.580 -3.840 ;
        RECT 774.660 -4.160 774.980 -3.840 ;
        RECT 924.260 -4.160 924.580 -3.840 ;
        RECT 924.660 -4.160 924.980 -3.840 ;
        RECT 1003.340 -4.160 1003.660 -3.840 ;
        RECT 1003.740 -4.160 1004.060 -3.840 ;
        RECT -4.480 -4.560 -4.160 -4.240 ;
        RECT -4.080 -4.560 -3.760 -4.240 ;
        RECT 24.260 -4.560 24.580 -4.240 ;
        RECT 24.660 -4.560 24.980 -4.240 ;
        RECT 174.260 -4.560 174.580 -4.240 ;
        RECT 174.660 -4.560 174.980 -4.240 ;
        RECT 324.260 -4.560 324.580 -4.240 ;
        RECT 324.660 -4.560 324.980 -4.240 ;
        RECT 474.260 -4.560 474.580 -4.240 ;
        RECT 474.660 -4.560 474.980 -4.240 ;
        RECT 624.260 -4.560 624.580 -4.240 ;
        RECT 624.660 -4.560 624.980 -4.240 ;
        RECT 774.260 -4.560 774.580 -4.240 ;
        RECT 774.660 -4.560 774.980 -4.240 ;
        RECT 924.260 -4.560 924.580 -4.240 ;
        RECT 924.660 -4.560 924.980 -4.240 ;
        RECT 1003.340 -4.560 1003.660 -4.240 ;
        RECT 1003.740 -4.560 1004.060 -4.240 ;
      LAYER met4 ;
        RECT -4.570 -4.650 -3.670 94.410 ;
        RECT 24.170 89.700 25.070 95.730 ;
        RECT 174.170 89.700 175.070 95.730 ;
        RECT 324.170 89.700 325.070 95.730 ;
        RECT 474.170 89.700 475.070 95.730 ;
        RECT 624.170 89.700 625.070 95.730 ;
        RECT 774.170 89.700 775.070 95.730 ;
        RECT 924.170 89.700 925.070 95.730 ;
        RECT 24.170 -5.970 25.070 0.300 ;
        RECT 174.170 -5.970 175.070 0.300 ;
        RECT 324.170 -5.970 325.070 0.300 ;
        RECT 474.170 -5.970 475.070 0.300 ;
        RECT 624.170 -5.970 625.070 0.300 ;
        RECT 774.170 -5.970 775.070 0.300 ;
        RECT 924.170 -5.970 925.070 0.300 ;
        RECT 1003.250 -4.650 1004.150 94.410 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -5.890 94.830 1005.470 95.730 ;
        RECT -5.890 -5.970 1005.470 -5.070 ;
      LAYER via3 ;
        RECT -5.800 95.320 -5.480 95.640 ;
        RECT -5.400 95.320 -5.080 95.640 ;
        RECT 99.260 95.320 99.580 95.640 ;
        RECT 99.660 95.320 99.980 95.640 ;
        RECT 249.260 95.320 249.580 95.640 ;
        RECT 249.660 95.320 249.980 95.640 ;
        RECT 399.260 95.320 399.580 95.640 ;
        RECT 399.660 95.320 399.980 95.640 ;
        RECT 549.260 95.320 549.580 95.640 ;
        RECT 549.660 95.320 549.980 95.640 ;
        RECT 699.260 95.320 699.580 95.640 ;
        RECT 699.660 95.320 699.980 95.640 ;
        RECT 849.260 95.320 849.580 95.640 ;
        RECT 849.660 95.320 849.980 95.640 ;
        RECT 1004.660 95.320 1004.980 95.640 ;
        RECT 1005.060 95.320 1005.380 95.640 ;
        RECT -5.800 94.920 -5.480 95.240 ;
        RECT -5.400 94.920 -5.080 95.240 ;
        RECT 99.260 94.920 99.580 95.240 ;
        RECT 99.660 94.920 99.980 95.240 ;
        RECT 249.260 94.920 249.580 95.240 ;
        RECT 249.660 94.920 249.980 95.240 ;
        RECT 399.260 94.920 399.580 95.240 ;
        RECT 399.660 94.920 399.980 95.240 ;
        RECT 549.260 94.920 549.580 95.240 ;
        RECT 549.660 94.920 549.980 95.240 ;
        RECT 699.260 94.920 699.580 95.240 ;
        RECT 699.660 94.920 699.980 95.240 ;
        RECT 849.260 94.920 849.580 95.240 ;
        RECT 849.660 94.920 849.980 95.240 ;
        RECT 1004.660 94.920 1004.980 95.240 ;
        RECT 1005.060 94.920 1005.380 95.240 ;
        RECT -5.800 -5.480 -5.480 -5.160 ;
        RECT -5.400 -5.480 -5.080 -5.160 ;
        RECT 99.260 -5.480 99.580 -5.160 ;
        RECT 99.660 -5.480 99.980 -5.160 ;
        RECT 249.260 -5.480 249.580 -5.160 ;
        RECT 249.660 -5.480 249.980 -5.160 ;
        RECT 399.260 -5.480 399.580 -5.160 ;
        RECT 399.660 -5.480 399.980 -5.160 ;
        RECT 549.260 -5.480 549.580 -5.160 ;
        RECT 549.660 -5.480 549.980 -5.160 ;
        RECT 699.260 -5.480 699.580 -5.160 ;
        RECT 699.660 -5.480 699.980 -5.160 ;
        RECT 849.260 -5.480 849.580 -5.160 ;
        RECT 849.660 -5.480 849.980 -5.160 ;
        RECT 1004.660 -5.480 1004.980 -5.160 ;
        RECT 1005.060 -5.480 1005.380 -5.160 ;
        RECT -5.800 -5.880 -5.480 -5.560 ;
        RECT -5.400 -5.880 -5.080 -5.560 ;
        RECT 99.260 -5.880 99.580 -5.560 ;
        RECT 99.660 -5.880 99.980 -5.560 ;
        RECT 249.260 -5.880 249.580 -5.560 ;
        RECT 249.660 -5.880 249.980 -5.560 ;
        RECT 399.260 -5.880 399.580 -5.560 ;
        RECT 399.660 -5.880 399.980 -5.560 ;
        RECT 549.260 -5.880 549.580 -5.560 ;
        RECT 549.660 -5.880 549.980 -5.560 ;
        RECT 699.260 -5.880 699.580 -5.560 ;
        RECT 699.660 -5.880 699.980 -5.560 ;
        RECT 849.260 -5.880 849.580 -5.560 ;
        RECT 849.660 -5.880 849.980 -5.560 ;
        RECT 1004.660 -5.880 1004.980 -5.560 ;
        RECT 1005.060 -5.880 1005.380 -5.560 ;
      LAYER met4 ;
        RECT -5.890 -5.970 -4.990 95.730 ;
        RECT 99.170 89.700 100.070 95.730 ;
        RECT 249.170 89.700 250.070 95.730 ;
        RECT 399.170 89.700 400.070 95.730 ;
        RECT 549.170 89.700 550.070 95.730 ;
        RECT 699.170 89.700 700.070 95.730 ;
        RECT 849.170 89.700 850.070 95.730 ;
        RECT 99.170 -5.970 100.070 0.300 ;
        RECT 249.170 -5.970 250.070 0.300 ;
        RECT 399.170 -5.970 400.070 0.300 ;
        RECT 549.170 -5.970 550.070 0.300 ;
        RECT 699.170 -5.970 700.070 0.300 ;
        RECT 849.170 -5.970 850.070 0.300 ;
        RECT 1004.570 -5.970 1005.470 95.730 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -7.210 96.150 1006.790 97.050 ;
        RECT -7.210 -7.290 1006.790 -6.390 ;
      LAYER via3 ;
        RECT -7.120 96.640 -6.800 96.960 ;
        RECT -6.720 96.640 -6.400 96.960 ;
        RECT 28.360 96.640 28.680 96.960 ;
        RECT 28.760 96.640 29.080 96.960 ;
        RECT 178.360 96.640 178.680 96.960 ;
        RECT 178.760 96.640 179.080 96.960 ;
        RECT 328.360 96.640 328.680 96.960 ;
        RECT 328.760 96.640 329.080 96.960 ;
        RECT 478.360 96.640 478.680 96.960 ;
        RECT 478.760 96.640 479.080 96.960 ;
        RECT 628.360 96.640 628.680 96.960 ;
        RECT 628.760 96.640 629.080 96.960 ;
        RECT 778.360 96.640 778.680 96.960 ;
        RECT 778.760 96.640 779.080 96.960 ;
        RECT 928.360 96.640 928.680 96.960 ;
        RECT 928.760 96.640 929.080 96.960 ;
        RECT 1005.980 96.640 1006.300 96.960 ;
        RECT 1006.380 96.640 1006.700 96.960 ;
        RECT -7.120 96.240 -6.800 96.560 ;
        RECT -6.720 96.240 -6.400 96.560 ;
        RECT 28.360 96.240 28.680 96.560 ;
        RECT 28.760 96.240 29.080 96.560 ;
        RECT 178.360 96.240 178.680 96.560 ;
        RECT 178.760 96.240 179.080 96.560 ;
        RECT 328.360 96.240 328.680 96.560 ;
        RECT 328.760 96.240 329.080 96.560 ;
        RECT 478.360 96.240 478.680 96.560 ;
        RECT 478.760 96.240 479.080 96.560 ;
        RECT 628.360 96.240 628.680 96.560 ;
        RECT 628.760 96.240 629.080 96.560 ;
        RECT 778.360 96.240 778.680 96.560 ;
        RECT 778.760 96.240 779.080 96.560 ;
        RECT 928.360 96.240 928.680 96.560 ;
        RECT 928.760 96.240 929.080 96.560 ;
        RECT 1005.980 96.240 1006.300 96.560 ;
        RECT 1006.380 96.240 1006.700 96.560 ;
        RECT -7.120 -6.800 -6.800 -6.480 ;
        RECT -6.720 -6.800 -6.400 -6.480 ;
        RECT 28.360 -6.800 28.680 -6.480 ;
        RECT 28.760 -6.800 29.080 -6.480 ;
        RECT 178.360 -6.800 178.680 -6.480 ;
        RECT 178.760 -6.800 179.080 -6.480 ;
        RECT 328.360 -6.800 328.680 -6.480 ;
        RECT 328.760 -6.800 329.080 -6.480 ;
        RECT 478.360 -6.800 478.680 -6.480 ;
        RECT 478.760 -6.800 479.080 -6.480 ;
        RECT 628.360 -6.800 628.680 -6.480 ;
        RECT 628.760 -6.800 629.080 -6.480 ;
        RECT 778.360 -6.800 778.680 -6.480 ;
        RECT 778.760 -6.800 779.080 -6.480 ;
        RECT 928.360 -6.800 928.680 -6.480 ;
        RECT 928.760 -6.800 929.080 -6.480 ;
        RECT 1005.980 -6.800 1006.300 -6.480 ;
        RECT 1006.380 -6.800 1006.700 -6.480 ;
        RECT -7.120 -7.200 -6.800 -6.880 ;
        RECT -6.720 -7.200 -6.400 -6.880 ;
        RECT 28.360 -7.200 28.680 -6.880 ;
        RECT 28.760 -7.200 29.080 -6.880 ;
        RECT 178.360 -7.200 178.680 -6.880 ;
        RECT 178.760 -7.200 179.080 -6.880 ;
        RECT 328.360 -7.200 328.680 -6.880 ;
        RECT 328.760 -7.200 329.080 -6.880 ;
        RECT 478.360 -7.200 478.680 -6.880 ;
        RECT 478.760 -7.200 479.080 -6.880 ;
        RECT 628.360 -7.200 628.680 -6.880 ;
        RECT 628.760 -7.200 629.080 -6.880 ;
        RECT 778.360 -7.200 778.680 -6.880 ;
        RECT 778.760 -7.200 779.080 -6.880 ;
        RECT 928.360 -7.200 928.680 -6.880 ;
        RECT 928.760 -7.200 929.080 -6.880 ;
        RECT 1005.980 -7.200 1006.300 -6.880 ;
        RECT 1006.380 -7.200 1006.700 -6.880 ;
      LAYER met4 ;
        RECT -7.210 -7.290 -6.310 97.050 ;
        RECT 28.270 89.700 29.170 98.370 ;
        RECT 178.270 89.700 179.170 98.370 ;
        RECT 328.270 89.700 329.170 98.370 ;
        RECT 478.270 89.700 479.170 98.370 ;
        RECT 628.270 89.700 629.170 98.370 ;
        RECT 778.270 89.700 779.170 98.370 ;
        RECT 928.270 89.700 929.170 98.370 ;
        RECT 28.270 -8.610 29.170 0.300 ;
        RECT 178.270 -8.610 179.170 0.300 ;
        RECT 328.270 -8.610 329.170 0.300 ;
        RECT 478.270 -8.610 479.170 0.300 ;
        RECT 628.270 -8.610 629.170 0.300 ;
        RECT 778.270 -8.610 779.170 0.300 ;
        RECT 928.270 -8.610 929.170 0.300 ;
        RECT 1005.890 -7.290 1006.790 97.050 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -8.530 97.470 1008.110 98.370 ;
        RECT -8.530 -8.610 1008.110 -7.710 ;
      LAYER via3 ;
        RECT -8.440 97.960 -8.120 98.280 ;
        RECT -8.040 97.960 -7.720 98.280 ;
        RECT 103.360 97.960 103.680 98.280 ;
        RECT 103.760 97.960 104.080 98.280 ;
        RECT 253.360 97.960 253.680 98.280 ;
        RECT 253.760 97.960 254.080 98.280 ;
        RECT 403.360 97.960 403.680 98.280 ;
        RECT 403.760 97.960 404.080 98.280 ;
        RECT 553.360 97.960 553.680 98.280 ;
        RECT 553.760 97.960 554.080 98.280 ;
        RECT 703.360 97.960 703.680 98.280 ;
        RECT 703.760 97.960 704.080 98.280 ;
        RECT 853.360 97.960 853.680 98.280 ;
        RECT 853.760 97.960 854.080 98.280 ;
        RECT 1007.300 97.960 1007.620 98.280 ;
        RECT 1007.700 97.960 1008.020 98.280 ;
        RECT -8.440 97.560 -8.120 97.880 ;
        RECT -8.040 97.560 -7.720 97.880 ;
        RECT 103.360 97.560 103.680 97.880 ;
        RECT 103.760 97.560 104.080 97.880 ;
        RECT 253.360 97.560 253.680 97.880 ;
        RECT 253.760 97.560 254.080 97.880 ;
        RECT 403.360 97.560 403.680 97.880 ;
        RECT 403.760 97.560 404.080 97.880 ;
        RECT 553.360 97.560 553.680 97.880 ;
        RECT 553.760 97.560 554.080 97.880 ;
        RECT 703.360 97.560 703.680 97.880 ;
        RECT 703.760 97.560 704.080 97.880 ;
        RECT 853.360 97.560 853.680 97.880 ;
        RECT 853.760 97.560 854.080 97.880 ;
        RECT 1007.300 97.560 1007.620 97.880 ;
        RECT 1007.700 97.560 1008.020 97.880 ;
        RECT -8.440 -8.120 -8.120 -7.800 ;
        RECT -8.040 -8.120 -7.720 -7.800 ;
        RECT 103.360 -8.120 103.680 -7.800 ;
        RECT 103.760 -8.120 104.080 -7.800 ;
        RECT 253.360 -8.120 253.680 -7.800 ;
        RECT 253.760 -8.120 254.080 -7.800 ;
        RECT 403.360 -8.120 403.680 -7.800 ;
        RECT 403.760 -8.120 404.080 -7.800 ;
        RECT 553.360 -8.120 553.680 -7.800 ;
        RECT 553.760 -8.120 554.080 -7.800 ;
        RECT 703.360 -8.120 703.680 -7.800 ;
        RECT 703.760 -8.120 704.080 -7.800 ;
        RECT 853.360 -8.120 853.680 -7.800 ;
        RECT 853.760 -8.120 854.080 -7.800 ;
        RECT 1007.300 -8.120 1007.620 -7.800 ;
        RECT 1007.700 -8.120 1008.020 -7.800 ;
        RECT -8.440 -8.520 -8.120 -8.200 ;
        RECT -8.040 -8.520 -7.720 -8.200 ;
        RECT 103.360 -8.520 103.680 -8.200 ;
        RECT 103.760 -8.520 104.080 -8.200 ;
        RECT 253.360 -8.520 253.680 -8.200 ;
        RECT 253.760 -8.520 254.080 -8.200 ;
        RECT 403.360 -8.520 403.680 -8.200 ;
        RECT 403.760 -8.520 404.080 -8.200 ;
        RECT 553.360 -8.520 553.680 -8.200 ;
        RECT 553.760 -8.520 554.080 -8.200 ;
        RECT 703.360 -8.520 703.680 -8.200 ;
        RECT 703.760 -8.520 704.080 -8.200 ;
        RECT 853.360 -8.520 853.680 -8.200 ;
        RECT 853.760 -8.520 854.080 -8.200 ;
        RECT 1007.300 -8.520 1007.620 -8.200 ;
        RECT 1007.700 -8.520 1008.020 -8.200 ;
      LAYER met4 ;
        RECT -8.530 -8.610 -7.630 98.370 ;
        RECT 103.270 89.700 104.170 98.370 ;
        RECT 253.270 89.700 254.170 98.370 ;
        RECT 403.270 89.700 404.170 98.370 ;
        RECT 553.270 89.700 554.170 98.370 ;
        RECT 703.270 89.700 704.170 98.370 ;
        RECT 853.270 89.700 854.170 98.370 ;
        RECT 103.270 -8.610 104.170 0.300 ;
        RECT 253.270 -8.610 254.170 0.300 ;
        RECT 403.270 -8.610 404.170 0.300 ;
        RECT 553.270 -8.610 554.170 0.300 ;
        RECT 703.270 -8.610 704.170 0.300 ;
        RECT 853.270 -8.610 854.170 0.300 ;
        RECT 1007.210 -8.610 1008.110 98.370 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -9.850 98.790 1009.430 99.690 ;
        RECT -9.850 -9.930 1009.430 -9.030 ;
      LAYER via3 ;
        RECT -9.760 99.280 -9.440 99.600 ;
        RECT -9.360 99.280 -9.040 99.600 ;
        RECT 32.460 99.280 32.780 99.600 ;
        RECT 32.860 99.280 33.180 99.600 ;
        RECT 182.460 99.280 182.780 99.600 ;
        RECT 182.860 99.280 183.180 99.600 ;
        RECT 332.460 99.280 332.780 99.600 ;
        RECT 332.860 99.280 333.180 99.600 ;
        RECT 482.460 99.280 482.780 99.600 ;
        RECT 482.860 99.280 483.180 99.600 ;
        RECT 632.460 99.280 632.780 99.600 ;
        RECT 632.860 99.280 633.180 99.600 ;
        RECT 782.460 99.280 782.780 99.600 ;
        RECT 782.860 99.280 783.180 99.600 ;
        RECT 932.460 99.280 932.780 99.600 ;
        RECT 932.860 99.280 933.180 99.600 ;
        RECT 1008.620 99.280 1008.940 99.600 ;
        RECT 1009.020 99.280 1009.340 99.600 ;
        RECT -9.760 98.880 -9.440 99.200 ;
        RECT -9.360 98.880 -9.040 99.200 ;
        RECT 32.460 98.880 32.780 99.200 ;
        RECT 32.860 98.880 33.180 99.200 ;
        RECT 182.460 98.880 182.780 99.200 ;
        RECT 182.860 98.880 183.180 99.200 ;
        RECT 332.460 98.880 332.780 99.200 ;
        RECT 332.860 98.880 333.180 99.200 ;
        RECT 482.460 98.880 482.780 99.200 ;
        RECT 482.860 98.880 483.180 99.200 ;
        RECT 632.460 98.880 632.780 99.200 ;
        RECT 632.860 98.880 633.180 99.200 ;
        RECT 782.460 98.880 782.780 99.200 ;
        RECT 782.860 98.880 783.180 99.200 ;
        RECT 932.460 98.880 932.780 99.200 ;
        RECT 932.860 98.880 933.180 99.200 ;
        RECT 1008.620 98.880 1008.940 99.200 ;
        RECT 1009.020 98.880 1009.340 99.200 ;
        RECT -9.760 -9.440 -9.440 -9.120 ;
        RECT -9.360 -9.440 -9.040 -9.120 ;
        RECT 32.460 -9.440 32.780 -9.120 ;
        RECT 32.860 -9.440 33.180 -9.120 ;
        RECT 182.460 -9.440 182.780 -9.120 ;
        RECT 182.860 -9.440 183.180 -9.120 ;
        RECT 332.460 -9.440 332.780 -9.120 ;
        RECT 332.860 -9.440 333.180 -9.120 ;
        RECT 482.460 -9.440 482.780 -9.120 ;
        RECT 482.860 -9.440 483.180 -9.120 ;
        RECT 632.460 -9.440 632.780 -9.120 ;
        RECT 632.860 -9.440 633.180 -9.120 ;
        RECT 782.460 -9.440 782.780 -9.120 ;
        RECT 782.860 -9.440 783.180 -9.120 ;
        RECT 932.460 -9.440 932.780 -9.120 ;
        RECT 932.860 -9.440 933.180 -9.120 ;
        RECT 1008.620 -9.440 1008.940 -9.120 ;
        RECT 1009.020 -9.440 1009.340 -9.120 ;
        RECT -9.760 -9.840 -9.440 -9.520 ;
        RECT -9.360 -9.840 -9.040 -9.520 ;
        RECT 32.460 -9.840 32.780 -9.520 ;
        RECT 32.860 -9.840 33.180 -9.520 ;
        RECT 182.460 -9.840 182.780 -9.520 ;
        RECT 182.860 -9.840 183.180 -9.520 ;
        RECT 332.460 -9.840 332.780 -9.520 ;
        RECT 332.860 -9.840 333.180 -9.520 ;
        RECT 482.460 -9.840 482.780 -9.520 ;
        RECT 482.860 -9.840 483.180 -9.520 ;
        RECT 632.460 -9.840 632.780 -9.520 ;
        RECT 632.860 -9.840 633.180 -9.520 ;
        RECT 782.460 -9.840 782.780 -9.520 ;
        RECT 782.860 -9.840 783.180 -9.520 ;
        RECT 932.460 -9.840 932.780 -9.520 ;
        RECT 932.860 -9.840 933.180 -9.520 ;
        RECT 1008.620 -9.840 1008.940 -9.520 ;
        RECT 1009.020 -9.840 1009.340 -9.520 ;
      LAYER met4 ;
        RECT -9.850 -9.930 -8.950 99.690 ;
        RECT 32.370 89.700 33.270 101.010 ;
        RECT 182.370 89.700 183.270 101.010 ;
        RECT 332.370 89.700 333.270 101.010 ;
        RECT 482.370 89.700 483.270 101.010 ;
        RECT 632.370 89.700 633.270 101.010 ;
        RECT 782.370 89.700 783.270 101.010 ;
        RECT 932.370 89.700 933.270 101.010 ;
        RECT 32.370 -11.250 33.270 0.300 ;
        RECT 182.370 -11.250 183.270 0.300 ;
        RECT 332.370 -11.250 333.270 0.300 ;
        RECT 482.370 -11.250 483.270 0.300 ;
        RECT 632.370 -11.250 633.270 0.300 ;
        RECT 782.370 -11.250 783.270 0.300 ;
        RECT 932.370 -11.250 933.270 0.300 ;
        RECT 1008.530 -9.930 1009.430 99.690 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -11.170 100.110 1010.750 101.010 ;
        RECT -11.170 -11.250 1010.750 -10.350 ;
      LAYER via3 ;
        RECT -11.080 100.600 -10.760 100.920 ;
        RECT -10.680 100.600 -10.360 100.920 ;
        RECT 107.460 100.600 107.780 100.920 ;
        RECT 107.860 100.600 108.180 100.920 ;
        RECT 257.460 100.600 257.780 100.920 ;
        RECT 257.860 100.600 258.180 100.920 ;
        RECT 407.460 100.600 407.780 100.920 ;
        RECT 407.860 100.600 408.180 100.920 ;
        RECT 557.460 100.600 557.780 100.920 ;
        RECT 557.860 100.600 558.180 100.920 ;
        RECT 707.460 100.600 707.780 100.920 ;
        RECT 707.860 100.600 708.180 100.920 ;
        RECT 857.460 100.600 857.780 100.920 ;
        RECT 857.860 100.600 858.180 100.920 ;
        RECT 1009.940 100.600 1010.260 100.920 ;
        RECT 1010.340 100.600 1010.660 100.920 ;
        RECT -11.080 100.200 -10.760 100.520 ;
        RECT -10.680 100.200 -10.360 100.520 ;
        RECT 107.460 100.200 107.780 100.520 ;
        RECT 107.860 100.200 108.180 100.520 ;
        RECT 257.460 100.200 257.780 100.520 ;
        RECT 257.860 100.200 258.180 100.520 ;
        RECT 407.460 100.200 407.780 100.520 ;
        RECT 407.860 100.200 408.180 100.520 ;
        RECT 557.460 100.200 557.780 100.520 ;
        RECT 557.860 100.200 558.180 100.520 ;
        RECT 707.460 100.200 707.780 100.520 ;
        RECT 707.860 100.200 708.180 100.520 ;
        RECT 857.460 100.200 857.780 100.520 ;
        RECT 857.860 100.200 858.180 100.520 ;
        RECT 1009.940 100.200 1010.260 100.520 ;
        RECT 1010.340 100.200 1010.660 100.520 ;
        RECT -11.080 -10.760 -10.760 -10.440 ;
        RECT -10.680 -10.760 -10.360 -10.440 ;
        RECT 107.460 -10.760 107.780 -10.440 ;
        RECT 107.860 -10.760 108.180 -10.440 ;
        RECT 257.460 -10.760 257.780 -10.440 ;
        RECT 257.860 -10.760 258.180 -10.440 ;
        RECT 407.460 -10.760 407.780 -10.440 ;
        RECT 407.860 -10.760 408.180 -10.440 ;
        RECT 557.460 -10.760 557.780 -10.440 ;
        RECT 557.860 -10.760 558.180 -10.440 ;
        RECT 707.460 -10.760 707.780 -10.440 ;
        RECT 707.860 -10.760 708.180 -10.440 ;
        RECT 857.460 -10.760 857.780 -10.440 ;
        RECT 857.860 -10.760 858.180 -10.440 ;
        RECT 1009.940 -10.760 1010.260 -10.440 ;
        RECT 1010.340 -10.760 1010.660 -10.440 ;
        RECT -11.080 -11.160 -10.760 -10.840 ;
        RECT -10.680 -11.160 -10.360 -10.840 ;
        RECT 107.460 -11.160 107.780 -10.840 ;
        RECT 107.860 -11.160 108.180 -10.840 ;
        RECT 257.460 -11.160 257.780 -10.840 ;
        RECT 257.860 -11.160 258.180 -10.840 ;
        RECT 407.460 -11.160 407.780 -10.840 ;
        RECT 407.860 -11.160 408.180 -10.840 ;
        RECT 557.460 -11.160 557.780 -10.840 ;
        RECT 557.860 -11.160 558.180 -10.840 ;
        RECT 707.460 -11.160 707.780 -10.840 ;
        RECT 707.860 -11.160 708.180 -10.840 ;
        RECT 857.460 -11.160 857.780 -10.840 ;
        RECT 857.860 -11.160 858.180 -10.840 ;
        RECT 1009.940 -11.160 1010.260 -10.840 ;
        RECT 1010.340 -11.160 1010.660 -10.840 ;
      LAYER met4 ;
        RECT -11.170 -11.250 -10.270 101.010 ;
        RECT 107.370 89.700 108.270 101.010 ;
        RECT 257.370 89.700 258.270 101.010 ;
        RECT 407.370 89.700 408.270 101.010 ;
        RECT 557.370 89.700 558.270 101.010 ;
        RECT 707.370 89.700 708.270 101.010 ;
        RECT 857.370 89.700 858.270 101.010 ;
        RECT 107.370 -11.250 108.270 0.300 ;
        RECT 257.370 -11.250 258.270 0.300 ;
        RECT 407.370 -11.250 408.270 0.300 ;
        RECT 557.370 -11.250 558.270 0.300 ;
        RECT 707.370 -11.250 708.270 0.300 ;
        RECT 857.370 -11.250 858.270 0.300 ;
        RECT 1009.850 -11.250 1010.750 101.010 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -12.490 101.430 1012.070 102.330 ;
        RECT -12.490 -12.570 1012.070 -11.670 ;
      LAYER via3 ;
        RECT -12.400 101.920 -12.080 102.240 ;
        RECT -12.000 101.920 -11.680 102.240 ;
        RECT 36.560 101.920 36.880 102.240 ;
        RECT 36.960 101.920 37.280 102.240 ;
        RECT 186.560 101.920 186.880 102.240 ;
        RECT 186.960 101.920 187.280 102.240 ;
        RECT 336.560 101.920 336.880 102.240 ;
        RECT 336.960 101.920 337.280 102.240 ;
        RECT 486.560 101.920 486.880 102.240 ;
        RECT 486.960 101.920 487.280 102.240 ;
        RECT 636.560 101.920 636.880 102.240 ;
        RECT 636.960 101.920 637.280 102.240 ;
        RECT 786.560 101.920 786.880 102.240 ;
        RECT 786.960 101.920 787.280 102.240 ;
        RECT 936.560 101.920 936.880 102.240 ;
        RECT 936.960 101.920 937.280 102.240 ;
        RECT 1011.260 101.920 1011.580 102.240 ;
        RECT 1011.660 101.920 1011.980 102.240 ;
        RECT -12.400 101.520 -12.080 101.840 ;
        RECT -12.000 101.520 -11.680 101.840 ;
        RECT 36.560 101.520 36.880 101.840 ;
        RECT 36.960 101.520 37.280 101.840 ;
        RECT 186.560 101.520 186.880 101.840 ;
        RECT 186.960 101.520 187.280 101.840 ;
        RECT 336.560 101.520 336.880 101.840 ;
        RECT 336.960 101.520 337.280 101.840 ;
        RECT 486.560 101.520 486.880 101.840 ;
        RECT 486.960 101.520 487.280 101.840 ;
        RECT 636.560 101.520 636.880 101.840 ;
        RECT 636.960 101.520 637.280 101.840 ;
        RECT 786.560 101.520 786.880 101.840 ;
        RECT 786.960 101.520 787.280 101.840 ;
        RECT 936.560 101.520 936.880 101.840 ;
        RECT 936.960 101.520 937.280 101.840 ;
        RECT 1011.260 101.520 1011.580 101.840 ;
        RECT 1011.660 101.520 1011.980 101.840 ;
        RECT -12.400 -12.080 -12.080 -11.760 ;
        RECT -12.000 -12.080 -11.680 -11.760 ;
        RECT 36.560 -12.080 36.880 -11.760 ;
        RECT 36.960 -12.080 37.280 -11.760 ;
        RECT 186.560 -12.080 186.880 -11.760 ;
        RECT 186.960 -12.080 187.280 -11.760 ;
        RECT 336.560 -12.080 336.880 -11.760 ;
        RECT 336.960 -12.080 337.280 -11.760 ;
        RECT 486.560 -12.080 486.880 -11.760 ;
        RECT 486.960 -12.080 487.280 -11.760 ;
        RECT 636.560 -12.080 636.880 -11.760 ;
        RECT 636.960 -12.080 637.280 -11.760 ;
        RECT 786.560 -12.080 786.880 -11.760 ;
        RECT 786.960 -12.080 787.280 -11.760 ;
        RECT 936.560 -12.080 936.880 -11.760 ;
        RECT 936.960 -12.080 937.280 -11.760 ;
        RECT 1011.260 -12.080 1011.580 -11.760 ;
        RECT 1011.660 -12.080 1011.980 -11.760 ;
        RECT -12.400 -12.480 -12.080 -12.160 ;
        RECT -12.000 -12.480 -11.680 -12.160 ;
        RECT 36.560 -12.480 36.880 -12.160 ;
        RECT 36.960 -12.480 37.280 -12.160 ;
        RECT 186.560 -12.480 186.880 -12.160 ;
        RECT 186.960 -12.480 187.280 -12.160 ;
        RECT 336.560 -12.480 336.880 -12.160 ;
        RECT 336.960 -12.480 337.280 -12.160 ;
        RECT 486.560 -12.480 486.880 -12.160 ;
        RECT 486.960 -12.480 487.280 -12.160 ;
        RECT 636.560 -12.480 636.880 -12.160 ;
        RECT 636.960 -12.480 637.280 -12.160 ;
        RECT 786.560 -12.480 786.880 -12.160 ;
        RECT 786.960 -12.480 787.280 -12.160 ;
        RECT 936.560 -12.480 936.880 -12.160 ;
        RECT 936.960 -12.480 937.280 -12.160 ;
        RECT 1011.260 -12.480 1011.580 -12.160 ;
        RECT 1011.660 -12.480 1011.980 -12.160 ;
      LAYER met4 ;
        RECT -12.490 -12.570 -11.590 102.330 ;
        RECT 36.470 89.700 37.370 103.650 ;
        RECT 186.470 89.700 187.370 103.650 ;
        RECT 336.470 89.700 337.370 103.650 ;
        RECT 486.470 89.700 487.370 103.650 ;
        RECT 636.470 89.700 637.370 103.650 ;
        RECT 786.470 89.700 787.370 103.650 ;
        RECT 936.470 89.700 937.370 103.650 ;
        RECT 36.470 -13.890 37.370 0.300 ;
        RECT 186.470 -13.890 187.370 0.300 ;
        RECT 336.470 -13.890 337.370 0.300 ;
        RECT 486.470 -13.890 487.370 0.300 ;
        RECT 636.470 -13.890 637.370 0.300 ;
        RECT 786.470 -13.890 787.370 0.300 ;
        RECT 936.470 -13.890 937.370 0.300 ;
        RECT 1011.170 -12.570 1012.070 102.330 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -13.810 102.750 1013.390 103.650 ;
        RECT -13.810 -13.890 1013.390 -12.990 ;
      LAYER via3 ;
        RECT -13.720 103.240 -13.400 103.560 ;
        RECT -13.320 103.240 -13.000 103.560 ;
        RECT 111.560 103.240 111.880 103.560 ;
        RECT 111.960 103.240 112.280 103.560 ;
        RECT 261.560 103.240 261.880 103.560 ;
        RECT 261.960 103.240 262.280 103.560 ;
        RECT 411.560 103.240 411.880 103.560 ;
        RECT 411.960 103.240 412.280 103.560 ;
        RECT 561.560 103.240 561.880 103.560 ;
        RECT 561.960 103.240 562.280 103.560 ;
        RECT 711.560 103.240 711.880 103.560 ;
        RECT 711.960 103.240 712.280 103.560 ;
        RECT 861.560 103.240 861.880 103.560 ;
        RECT 861.960 103.240 862.280 103.560 ;
        RECT 1012.580 103.240 1012.900 103.560 ;
        RECT 1012.980 103.240 1013.300 103.560 ;
        RECT -13.720 102.840 -13.400 103.160 ;
        RECT -13.320 102.840 -13.000 103.160 ;
        RECT 111.560 102.840 111.880 103.160 ;
        RECT 111.960 102.840 112.280 103.160 ;
        RECT 261.560 102.840 261.880 103.160 ;
        RECT 261.960 102.840 262.280 103.160 ;
        RECT 411.560 102.840 411.880 103.160 ;
        RECT 411.960 102.840 412.280 103.160 ;
        RECT 561.560 102.840 561.880 103.160 ;
        RECT 561.960 102.840 562.280 103.160 ;
        RECT 711.560 102.840 711.880 103.160 ;
        RECT 711.960 102.840 712.280 103.160 ;
        RECT 861.560 102.840 861.880 103.160 ;
        RECT 861.960 102.840 862.280 103.160 ;
        RECT 1012.580 102.840 1012.900 103.160 ;
        RECT 1012.980 102.840 1013.300 103.160 ;
        RECT -13.720 -13.400 -13.400 -13.080 ;
        RECT -13.320 -13.400 -13.000 -13.080 ;
        RECT 111.560 -13.400 111.880 -13.080 ;
        RECT 111.960 -13.400 112.280 -13.080 ;
        RECT 261.560 -13.400 261.880 -13.080 ;
        RECT 261.960 -13.400 262.280 -13.080 ;
        RECT 411.560 -13.400 411.880 -13.080 ;
        RECT 411.960 -13.400 412.280 -13.080 ;
        RECT 561.560 -13.400 561.880 -13.080 ;
        RECT 561.960 -13.400 562.280 -13.080 ;
        RECT 711.560 -13.400 711.880 -13.080 ;
        RECT 711.960 -13.400 712.280 -13.080 ;
        RECT 861.560 -13.400 861.880 -13.080 ;
        RECT 861.960 -13.400 862.280 -13.080 ;
        RECT 1012.580 -13.400 1012.900 -13.080 ;
        RECT 1012.980 -13.400 1013.300 -13.080 ;
        RECT -13.720 -13.800 -13.400 -13.480 ;
        RECT -13.320 -13.800 -13.000 -13.480 ;
        RECT 111.560 -13.800 111.880 -13.480 ;
        RECT 111.960 -13.800 112.280 -13.480 ;
        RECT 261.560 -13.800 261.880 -13.480 ;
        RECT 261.960 -13.800 262.280 -13.480 ;
        RECT 411.560 -13.800 411.880 -13.480 ;
        RECT 411.960 -13.800 412.280 -13.480 ;
        RECT 561.560 -13.800 561.880 -13.480 ;
        RECT 561.960 -13.800 562.280 -13.480 ;
        RECT 711.560 -13.800 711.880 -13.480 ;
        RECT 711.960 -13.800 712.280 -13.480 ;
        RECT 861.560 -13.800 861.880 -13.480 ;
        RECT 861.960 -13.800 862.280 -13.480 ;
        RECT 1012.580 -13.800 1012.900 -13.480 ;
        RECT 1012.980 -13.800 1013.300 -13.480 ;
      LAYER met4 ;
        RECT -13.810 -13.890 -12.910 103.650 ;
        RECT 111.470 89.700 112.370 103.650 ;
        RECT 261.470 89.700 262.370 103.650 ;
        RECT 411.470 89.700 412.370 103.650 ;
        RECT 561.470 89.700 562.370 103.650 ;
        RECT 711.470 89.700 712.370 103.650 ;
        RECT 861.470 89.700 862.370 103.650 ;
        RECT 111.470 -13.890 112.370 0.300 ;
        RECT 261.470 -13.890 262.370 0.300 ;
        RECT 411.470 -13.890 412.370 0.300 ;
        RECT 561.470 -13.890 562.370 0.300 ;
        RECT 711.470 -13.890 712.370 0.300 ;
        RECT 861.470 -13.890 862.370 0.300 ;
        RECT 1012.490 -13.890 1013.390 103.650 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 279.365 89.700 279.535 90.015 ;
        RECT 322.145 89.845 328.295 90.015 ;
        RECT 350.665 89.845 351.755 90.015 ;
        RECT 322.145 89.700 322.315 89.845 ;
        RECT 351.585 89.700 351.755 89.845 ;
        RECT 399.425 89.845 400.975 90.015 ;
        RECT 399.425 89.700 399.595 89.845 ;
        RECT 400.805 89.700 400.975 89.845 ;
        RECT 462.905 89.845 465.375 90.015 ;
        RECT 565.485 89.845 569.795 90.015 ;
        RECT 462.905 89.700 463.075 89.845 ;
        RECT 465.205 89.700 465.375 89.845 ;
        RECT 569.625 89.700 569.795 89.845 ;
        RECT 593.085 89.700 593.255 90.015 ;
        RECT 5.520 3.145 994.060 89.700 ;
      LAYER mcon ;
        RECT 279.365 89.845 279.535 90.015 ;
        RECT 328.125 89.845 328.295 90.015 ;
        RECT 593.085 89.845 593.255 90.015 ;
      LAYER met1 ;
        RECT 279.305 90.000 279.595 90.045 ;
        RECT 328.065 90.000 328.355 90.045 ;
        RECT 344.150 90.000 344.470 90.060 ;
        RECT 279.305 89.860 327.360 90.000 ;
        RECT 279.305 89.815 279.595 89.860 ;
        RECT 203.850 89.700 204.170 89.720 ;
        RECT 326.685 89.700 326.975 89.705 ;
        RECT 327.220 89.700 327.360 89.860 ;
        RECT 328.065 89.860 344.470 90.000 ;
        RECT 328.065 89.815 328.355 89.860 ;
        RECT 344.150 89.800 344.470 89.860 ;
        RECT 345.530 90.000 345.850 90.060 ;
        RECT 350.605 90.000 350.895 90.045 ;
        RECT 345.530 89.860 350.895 90.000 ;
        RECT 345.530 89.800 345.850 89.860 ;
        RECT 350.605 89.815 350.895 89.860 ;
        RECT 351.050 90.000 351.370 90.060 ;
        RECT 565.425 90.000 565.715 90.045 ;
        RECT 351.050 89.860 565.715 90.000 ;
        RECT 351.050 89.800 351.370 89.860 ;
        RECT 565.425 89.815 565.715 89.860 ;
        RECT 565.870 90.000 566.190 90.060 ;
        RECT 593.025 90.000 593.315 90.045 ;
        RECT 565.870 89.860 593.315 90.000 ;
        RECT 565.870 89.800 566.190 89.860 ;
        RECT 593.025 89.815 593.315 89.860 ;
        RECT 327.605 89.700 327.895 89.705 ;
        RECT 373.590 89.700 373.910 89.720 ;
        RECT 374.050 89.700 374.370 89.720 ;
        RECT 399.365 89.700 399.655 89.705 ;
        RECT 400.745 89.700 401.035 89.705 ;
        RECT 448.585 89.700 448.875 89.705 ;
        RECT 449.030 89.700 449.350 89.720 ;
        RECT 459.610 89.700 459.930 89.720 ;
        RECT 460.085 89.700 460.375 89.705 ;
        RECT 463.765 89.700 464.055 89.705 ;
        RECT 506.990 89.700 507.310 89.720 ;
        RECT 509.290 89.700 509.610 89.720 ;
        RECT 518.490 89.700 518.810 89.720 ;
        RECT 631.650 89.700 631.970 89.720 ;
        RECT 0.990 3.100 999.050 89.700 ;
      LAYER via ;
        RECT 203.880 89.460 204.140 89.720 ;
        RECT 344.180 89.800 344.440 90.060 ;
        RECT 345.560 89.800 345.820 90.060 ;
        RECT 351.080 89.800 351.340 90.060 ;
        RECT 565.900 89.800 566.160 90.060 ;
        RECT 373.620 89.460 373.880 89.720 ;
        RECT 374.080 89.460 374.340 89.720 ;
        RECT 449.060 89.460 449.320 89.720 ;
        RECT 459.640 89.460 459.900 89.720 ;
        RECT 507.020 89.460 507.280 89.720 ;
        RECT 509.320 89.460 509.580 89.720 ;
        RECT 518.520 89.460 518.780 89.720 ;
        RECT 631.680 89.460 631.940 89.720 ;
      LAYER met2 ;
        RECT 344.180 89.770 344.440 90.090 ;
        RECT 345.560 89.770 345.820 90.090 ;
        RECT 351.080 89.770 351.340 90.090 ;
        RECT 565.900 89.770 566.160 90.090 ;
        RECT 203.880 89.700 204.140 89.750 ;
        RECT 344.240 89.700 344.380 89.770 ;
        RECT 345.620 89.700 345.760 89.770 ;
        RECT 351.140 89.700 351.280 89.770 ;
        RECT 373.620 89.700 373.880 89.750 ;
        RECT 374.080 89.700 374.340 89.750 ;
        RECT 449.060 89.700 449.320 89.750 ;
        RECT 459.640 89.700 459.900 89.750 ;
        RECT 507.020 89.700 507.280 89.750 ;
        RECT 509.320 89.700 509.580 89.750 ;
        RECT 518.520 89.700 518.780 89.750 ;
        RECT 565.960 89.700 566.100 89.770 ;
        RECT 631.680 89.700 631.940 89.750 ;
        RECT 1.010 0.300 999.030 89.700 ;
      LAYER met3 ;
        RECT 0.300 4.255 973.295 89.585 ;
      LAYER met4 ;
        RECT 20.070 0.300 965.705 89.700 ;
  END
END mgmt_protect
END LIBRARY

