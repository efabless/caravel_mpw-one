magic
tech sky130A
magscale 1 2
timestamp 1607746021
<< obsli1 >>
rect 1380 1071 58604 3281
<< obsm1 >>
rect 566 1040 59326 3664
<< metal2 >>
rect 570 3800 626 4600
rect 754 3800 810 4600
rect 1122 3800 1178 4600
rect 1306 3800 1362 4600
rect 1674 3800 1730 4600
rect 1858 3800 1914 4600
rect 2226 3800 2282 4600
rect 2410 3800 2466 4600
rect 2778 3800 2834 4600
rect 2962 3800 3018 4600
rect 3146 3800 3202 4600
rect 3514 3800 3570 4600
rect 3698 3800 3754 4600
rect 4066 3800 4122 4600
rect 4250 3800 4306 4600
rect 4618 3800 4674 4600
rect 4802 3800 4858 4600
rect 5170 3800 5226 4600
rect 5354 3800 5410 4600
rect 5538 3800 5594 4600
rect 5906 3800 5962 4600
rect 6090 3800 6146 4600
rect 6458 3800 6514 4600
rect 6642 3800 6698 4600
rect 7010 3800 7066 4600
rect 7194 3800 7250 4600
rect 7562 3800 7618 4600
rect 7746 3800 7802 4600
rect 7930 3800 7986 4600
rect 8298 3800 8354 4600
rect 8482 3800 8538 4600
rect 8850 3800 8906 4600
rect 9034 3800 9090 4600
rect 9402 3800 9458 4600
rect 9586 3800 9642 4600
rect 9954 3800 10010 4600
rect 10138 3800 10194 4600
rect 10322 3800 10378 4600
rect 10690 3800 10746 4600
rect 10874 3800 10930 4600
rect 11242 3800 11298 4600
rect 11426 3800 11482 4600
rect 11794 3800 11850 4600
rect 11978 3800 12034 4600
rect 12162 3800 12218 4600
rect 12530 3800 12586 4600
rect 12714 3800 12770 4600
rect 13082 3800 13138 4600
rect 13266 3800 13322 4600
rect 13634 3800 13690 4600
rect 13818 3800 13874 4600
rect 14186 3800 14242 4600
rect 14370 3800 14426 4600
rect 14554 3800 14610 4600
rect 14922 3800 14978 4600
rect 15106 3800 15162 4600
rect 15474 3800 15530 4600
rect 15658 3800 15714 4600
rect 16026 3800 16082 4600
rect 16210 3800 16266 4600
rect 16578 3800 16634 4600
rect 16762 3800 16818 4600
rect 16946 3800 17002 4600
rect 17314 3800 17370 4600
rect 17498 3800 17554 4600
rect 17866 3800 17922 4600
rect 18050 3800 18106 4600
rect 18418 3800 18474 4600
rect 18602 3800 18658 4600
rect 18970 3800 19026 4600
rect 19154 3800 19210 4600
rect 19338 3800 19394 4600
rect 19706 3800 19762 4600
rect 19890 3800 19946 4600
rect 20258 3800 20314 4600
rect 20442 3800 20498 4600
rect 20810 3800 20866 4600
rect 20994 3800 21050 4600
rect 21362 3800 21418 4600
rect 21546 3800 21602 4600
rect 21730 3800 21786 4600
rect 22098 3800 22154 4600
rect 22282 3800 22338 4600
rect 22650 3800 22706 4600
rect 22834 3800 22890 4600
rect 23202 3800 23258 4600
rect 23386 3800 23442 4600
rect 23754 3800 23810 4600
rect 23938 3800 23994 4600
rect 24122 3800 24178 4600
rect 24490 3800 24546 4600
rect 24674 3800 24730 4600
rect 25042 3800 25098 4600
rect 25226 3800 25282 4600
rect 25594 3800 25650 4600
rect 25778 3800 25834 4600
rect 25962 3800 26018 4600
rect 26330 3800 26386 4600
rect 26514 3800 26570 4600
rect 26882 3800 26938 4600
rect 27066 3800 27122 4600
rect 27434 3800 27490 4600
rect 27618 3800 27674 4600
rect 27986 3800 28042 4600
rect 28170 3800 28226 4600
rect 28354 3800 28410 4600
rect 28722 3800 28778 4600
rect 28906 3800 28962 4600
rect 29274 3800 29330 4600
rect 29458 3800 29514 4600
rect 29826 3800 29882 4600
rect 30010 3800 30066 4600
rect 30378 3800 30434 4600
rect 30562 3800 30618 4600
rect 30746 3800 30802 4600
rect 31114 3800 31170 4600
rect 31298 3800 31354 4600
rect 31666 3800 31722 4600
rect 31850 3800 31906 4600
rect 32218 3800 32274 4600
rect 32402 3800 32458 4600
rect 32770 3800 32826 4600
rect 32954 3800 33010 4600
rect 33138 3800 33194 4600
rect 33506 3800 33562 4600
rect 33690 3800 33746 4600
rect 34058 3800 34114 4600
rect 34242 3800 34298 4600
rect 34610 3800 34666 4600
rect 34794 3800 34850 4600
rect 35162 3800 35218 4600
rect 35346 3800 35402 4600
rect 35530 3800 35586 4600
rect 35898 3800 35954 4600
rect 36082 3800 36138 4600
rect 36450 3800 36506 4600
rect 36634 3800 36690 4600
rect 37002 3800 37058 4600
rect 37186 3800 37242 4600
rect 37554 3800 37610 4600
rect 37738 3800 37794 4600
rect 37922 3800 37978 4600
rect 38290 3800 38346 4600
rect 38474 3800 38530 4600
rect 38842 3800 38898 4600
rect 39026 3800 39082 4600
rect 39394 3800 39450 4600
rect 39578 3800 39634 4600
rect 39762 3800 39818 4600
rect 40130 3800 40186 4600
rect 40314 3800 40370 4600
rect 40682 3800 40738 4600
rect 40866 3800 40922 4600
rect 41234 3800 41290 4600
rect 41418 3800 41474 4600
rect 41786 3800 41842 4600
rect 41970 3800 42026 4600
rect 42154 3800 42210 4600
rect 42522 3800 42578 4600
rect 42706 3800 42762 4600
rect 43074 3800 43130 4600
rect 43258 3800 43314 4600
rect 43626 3800 43682 4600
rect 43810 3800 43866 4600
rect 44178 3800 44234 4600
rect 44362 3800 44418 4600
rect 44546 3800 44602 4600
rect 44914 3800 44970 4600
rect 45098 3800 45154 4600
rect 45466 3800 45522 4600
rect 45650 3800 45706 4600
rect 46018 3800 46074 4600
rect 46202 3800 46258 4600
rect 46570 3800 46626 4600
rect 46754 3800 46810 4600
rect 46938 3800 46994 4600
rect 47306 3800 47362 4600
rect 47490 3800 47546 4600
rect 47858 3800 47914 4600
rect 48042 3800 48098 4600
rect 48410 3800 48466 4600
rect 48594 3800 48650 4600
rect 48962 3800 49018 4600
rect 49146 3800 49202 4600
rect 49330 3800 49386 4600
rect 49698 3800 49754 4600
rect 49882 3800 49938 4600
rect 50250 3800 50306 4600
rect 50434 3800 50490 4600
rect 50802 3800 50858 4600
rect 50986 3800 51042 4600
rect 51354 3800 51410 4600
rect 51538 3800 51594 4600
rect 51722 3800 51778 4600
rect 52090 3800 52146 4600
rect 52274 3800 52330 4600
rect 52642 3800 52698 4600
rect 52826 3800 52882 4600
rect 53194 3800 53250 4600
rect 53378 3800 53434 4600
rect 53562 3800 53618 4600
rect 53930 3800 53986 4600
rect 54114 3800 54170 4600
rect 54482 3800 54538 4600
rect 54666 3800 54722 4600
rect 55034 3800 55090 4600
rect 55218 3800 55274 4600
rect 55586 3800 55642 4600
rect 55770 3800 55826 4600
rect 55954 3800 56010 4600
rect 56322 3800 56378 4600
rect 56506 3800 56562 4600
rect 56874 3800 56930 4600
rect 57058 3800 57114 4600
rect 57426 3800 57482 4600
rect 57610 3800 57666 4600
rect 57978 3800 58034 4600
rect 58162 3800 58218 4600
rect 58346 3800 58402 4600
rect 58714 3800 58770 4600
rect 58898 3800 58954 4600
rect 59266 3800 59322 4600
rect 3350 1040 3410 3312
rect 11350 1040 11410 3312
rect 19350 1040 19410 3312
rect 27350 1040 27410 3312
rect 35350 1040 35410 3312
rect 43350 1040 43410 3312
rect 51350 1040 51410 3312
rect 570 0 626 800
rect 754 0 810 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2594 0 2650 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 25962 0 26018 800
rect 26146 0 26202 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27618 0 27674 800
rect 27802 0 27858 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31298 0 31354 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38474 0 38530 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43442 0 43498 800
rect 43810 0 43866 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44546 0 44602 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45650 0 45706 800
rect 45834 0 45890 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48594 0 48650 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49514 0 49570 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50618 0 50674 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53378 0 53434 800
rect 53562 0 53618 800
rect 53746 0 53802 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55586 0 55642 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59082 0 59138 800
<< obsm2 >>
rect 682 3744 698 3800
rect 866 3744 1066 3800
rect 1234 3744 1250 3800
rect 1418 3744 1618 3800
rect 1786 3744 1802 3800
rect 1970 3744 2170 3800
rect 2338 3744 2354 3800
rect 2522 3744 2722 3800
rect 2890 3744 2906 3800
rect 3074 3744 3090 3800
rect 3258 3744 3458 3800
rect 3626 3744 3642 3800
rect 3810 3744 4010 3800
rect 4178 3744 4194 3800
rect 4362 3744 4562 3800
rect 4730 3744 4746 3800
rect 4914 3744 5114 3800
rect 5282 3744 5298 3800
rect 5466 3744 5482 3800
rect 5650 3744 5850 3800
rect 6018 3744 6034 3800
rect 6202 3744 6402 3800
rect 6570 3744 6586 3800
rect 6754 3744 6954 3800
rect 7122 3744 7138 3800
rect 7306 3744 7506 3800
rect 7674 3744 7690 3800
rect 7858 3744 7874 3800
rect 8042 3744 8242 3800
rect 8410 3744 8426 3800
rect 8594 3744 8794 3800
rect 8962 3744 8978 3800
rect 9146 3744 9346 3800
rect 9514 3744 9530 3800
rect 9698 3744 9898 3800
rect 10066 3744 10082 3800
rect 10250 3744 10266 3800
rect 10434 3744 10634 3800
rect 10802 3744 10818 3800
rect 10986 3744 11186 3800
rect 11354 3744 11370 3800
rect 11538 3744 11738 3800
rect 11906 3744 11922 3800
rect 12090 3744 12106 3800
rect 12274 3744 12474 3800
rect 12642 3744 12658 3800
rect 12826 3744 13026 3800
rect 13194 3744 13210 3800
rect 13378 3744 13578 3800
rect 13746 3744 13762 3800
rect 13930 3744 14130 3800
rect 14298 3744 14314 3800
rect 14482 3744 14498 3800
rect 14666 3744 14866 3800
rect 15034 3744 15050 3800
rect 15218 3744 15418 3800
rect 15586 3744 15602 3800
rect 15770 3744 15970 3800
rect 16138 3744 16154 3800
rect 16322 3744 16522 3800
rect 16690 3744 16706 3800
rect 16874 3744 16890 3800
rect 17058 3744 17258 3800
rect 17426 3744 17442 3800
rect 17610 3744 17810 3800
rect 17978 3744 17994 3800
rect 18162 3744 18362 3800
rect 18530 3744 18546 3800
rect 18714 3744 18914 3800
rect 19082 3744 19098 3800
rect 19266 3744 19282 3800
rect 19450 3744 19650 3800
rect 19818 3744 19834 3800
rect 20002 3744 20202 3800
rect 20370 3744 20386 3800
rect 20554 3744 20754 3800
rect 20922 3744 20938 3800
rect 21106 3744 21306 3800
rect 21474 3744 21490 3800
rect 21658 3744 21674 3800
rect 21842 3744 22042 3800
rect 22210 3744 22226 3800
rect 22394 3744 22594 3800
rect 22762 3744 22778 3800
rect 22946 3744 23146 3800
rect 23314 3744 23330 3800
rect 23498 3744 23698 3800
rect 23866 3744 23882 3800
rect 24050 3744 24066 3800
rect 24234 3744 24434 3800
rect 24602 3744 24618 3800
rect 24786 3744 24986 3800
rect 25154 3744 25170 3800
rect 25338 3744 25538 3800
rect 25706 3744 25722 3800
rect 25890 3744 25906 3800
rect 26074 3744 26274 3800
rect 26442 3744 26458 3800
rect 26626 3744 26826 3800
rect 26994 3744 27010 3800
rect 27178 3744 27378 3800
rect 27546 3744 27562 3800
rect 27730 3744 27930 3800
rect 28098 3744 28114 3800
rect 28282 3744 28298 3800
rect 28466 3744 28666 3800
rect 28834 3744 28850 3800
rect 29018 3744 29218 3800
rect 29386 3744 29402 3800
rect 29570 3744 29770 3800
rect 29938 3744 29954 3800
rect 30122 3744 30322 3800
rect 30490 3744 30506 3800
rect 30674 3744 30690 3800
rect 30858 3744 31058 3800
rect 31226 3744 31242 3800
rect 31410 3744 31610 3800
rect 31778 3744 31794 3800
rect 31962 3744 32162 3800
rect 32330 3744 32346 3800
rect 32514 3744 32714 3800
rect 32882 3744 32898 3800
rect 33066 3744 33082 3800
rect 33250 3744 33450 3800
rect 33618 3744 33634 3800
rect 33802 3744 34002 3800
rect 34170 3744 34186 3800
rect 34354 3744 34554 3800
rect 34722 3744 34738 3800
rect 34906 3744 35106 3800
rect 35274 3744 35290 3800
rect 35458 3744 35474 3800
rect 35642 3744 35842 3800
rect 36010 3744 36026 3800
rect 36194 3744 36394 3800
rect 36562 3744 36578 3800
rect 36746 3744 36946 3800
rect 37114 3744 37130 3800
rect 37298 3744 37498 3800
rect 37666 3744 37682 3800
rect 37850 3744 37866 3800
rect 38034 3744 38234 3800
rect 38402 3744 38418 3800
rect 38586 3744 38786 3800
rect 38954 3744 38970 3800
rect 39138 3744 39338 3800
rect 39506 3744 39522 3800
rect 39690 3744 39706 3800
rect 39874 3744 40074 3800
rect 40242 3744 40258 3800
rect 40426 3744 40626 3800
rect 40794 3744 40810 3800
rect 40978 3744 41178 3800
rect 41346 3744 41362 3800
rect 41530 3744 41730 3800
rect 41898 3744 41914 3800
rect 42082 3744 42098 3800
rect 42266 3744 42466 3800
rect 42634 3744 42650 3800
rect 42818 3744 43018 3800
rect 43186 3744 43202 3800
rect 43370 3744 43570 3800
rect 43738 3744 43754 3800
rect 43922 3744 44122 3800
rect 44290 3744 44306 3800
rect 44474 3744 44490 3800
rect 44658 3744 44858 3800
rect 45026 3744 45042 3800
rect 45210 3744 45410 3800
rect 45578 3744 45594 3800
rect 45762 3744 45962 3800
rect 46130 3744 46146 3800
rect 46314 3744 46514 3800
rect 46682 3744 46698 3800
rect 46866 3744 46882 3800
rect 47050 3744 47250 3800
rect 47418 3744 47434 3800
rect 47602 3744 47802 3800
rect 47970 3744 47986 3800
rect 48154 3744 48354 3800
rect 48522 3744 48538 3800
rect 48706 3744 48906 3800
rect 49074 3744 49090 3800
rect 49258 3744 49274 3800
rect 49442 3744 49642 3800
rect 49810 3744 49826 3800
rect 49994 3744 50194 3800
rect 50362 3744 50378 3800
rect 50546 3744 50746 3800
rect 50914 3744 50930 3800
rect 51098 3744 51298 3800
rect 51466 3744 51482 3800
rect 51650 3744 51666 3800
rect 51834 3744 52034 3800
rect 52202 3744 52218 3800
rect 52386 3744 52586 3800
rect 52754 3744 52770 3800
rect 52938 3744 53138 3800
rect 53306 3744 53322 3800
rect 53490 3744 53506 3800
rect 53674 3744 53874 3800
rect 54042 3744 54058 3800
rect 54226 3744 54426 3800
rect 54594 3744 54610 3800
rect 54778 3744 54978 3800
rect 55146 3744 55162 3800
rect 55330 3744 55530 3800
rect 55698 3744 55714 3800
rect 55882 3744 55898 3800
rect 56066 3744 56266 3800
rect 56434 3744 56450 3800
rect 56618 3744 56818 3800
rect 56986 3744 57002 3800
rect 57170 3744 57370 3800
rect 57538 3744 57554 3800
rect 57722 3744 57922 3800
rect 58090 3744 58106 3800
rect 58274 3744 58290 3800
rect 58458 3744 58658 3800
rect 58826 3744 58842 3800
rect 59010 3744 59210 3800
rect 572 3368 59320 3744
rect 572 984 3294 3368
rect 3466 984 11294 3368
rect 11466 984 19294 3368
rect 19466 984 27294 3368
rect 27466 984 35294 3368
rect 35466 984 43294 3368
rect 43466 984 51294 3368
rect 51466 984 59320 3368
rect 572 856 59320 984
rect 682 800 698 856
rect 866 800 882 856
rect 1050 800 1250 856
rect 1418 800 1434 856
rect 1602 800 1802 856
rect 1970 800 1986 856
rect 2154 800 2354 856
rect 2522 800 2538 856
rect 2706 800 2722 856
rect 2890 800 3090 856
rect 3258 800 3274 856
rect 3442 800 3642 856
rect 3810 800 3826 856
rect 3994 800 4194 856
rect 4362 800 4378 856
rect 4546 800 4746 856
rect 4914 800 4930 856
rect 5098 800 5114 856
rect 5282 800 5482 856
rect 5650 800 5666 856
rect 5834 800 6034 856
rect 6202 800 6218 856
rect 6386 800 6586 856
rect 6754 800 6770 856
rect 6938 800 7138 856
rect 7306 800 7322 856
rect 7490 800 7506 856
rect 7674 800 7874 856
rect 8042 800 8058 856
rect 8226 800 8426 856
rect 8594 800 8610 856
rect 8778 800 8978 856
rect 9146 800 9162 856
rect 9330 800 9530 856
rect 9698 800 9714 856
rect 9882 800 9898 856
rect 10066 800 10266 856
rect 10434 800 10450 856
rect 10618 800 10818 856
rect 10986 800 11002 856
rect 11170 800 11370 856
rect 11538 800 11554 856
rect 11722 800 11922 856
rect 12090 800 12106 856
rect 12274 800 12290 856
rect 12458 800 12658 856
rect 12826 800 12842 856
rect 13010 800 13210 856
rect 13378 800 13394 856
rect 13562 800 13762 856
rect 13930 800 13946 856
rect 14114 800 14130 856
rect 14298 800 14498 856
rect 14666 800 14682 856
rect 14850 800 15050 856
rect 15218 800 15234 856
rect 15402 800 15602 856
rect 15770 800 15786 856
rect 15954 800 16154 856
rect 16322 800 16338 856
rect 16506 800 16522 856
rect 16690 800 16890 856
rect 17058 800 17074 856
rect 17242 800 17442 856
rect 17610 800 17626 856
rect 17794 800 17994 856
rect 18162 800 18178 856
rect 18346 800 18546 856
rect 18714 800 18730 856
rect 18898 800 18914 856
rect 19082 800 19282 856
rect 19450 800 19466 856
rect 19634 800 19834 856
rect 20002 800 20018 856
rect 20186 800 20386 856
rect 20554 800 20570 856
rect 20738 800 20938 856
rect 21106 800 21122 856
rect 21290 800 21306 856
rect 21474 800 21674 856
rect 21842 800 21858 856
rect 22026 800 22226 856
rect 22394 800 22410 856
rect 22578 800 22778 856
rect 22946 800 22962 856
rect 23130 800 23330 856
rect 23498 800 23514 856
rect 23682 800 23698 856
rect 23866 800 24066 856
rect 24234 800 24250 856
rect 24418 800 24618 856
rect 24786 800 24802 856
rect 24970 800 25170 856
rect 25338 800 25354 856
rect 25522 800 25722 856
rect 25890 800 25906 856
rect 26074 800 26090 856
rect 26258 800 26458 856
rect 26626 800 26642 856
rect 26810 800 27010 856
rect 27178 800 27194 856
rect 27362 800 27562 856
rect 27730 800 27746 856
rect 27914 800 27930 856
rect 28098 800 28298 856
rect 28466 800 28482 856
rect 28650 800 28850 856
rect 29018 800 29034 856
rect 29202 800 29402 856
rect 29570 800 29586 856
rect 29754 800 29954 856
rect 30122 800 30138 856
rect 30306 800 30322 856
rect 30490 800 30690 856
rect 30858 800 30874 856
rect 31042 800 31242 856
rect 31410 800 31426 856
rect 31594 800 31794 856
rect 31962 800 31978 856
rect 32146 800 32346 856
rect 32514 800 32530 856
rect 32698 800 32714 856
rect 32882 800 33082 856
rect 33250 800 33266 856
rect 33434 800 33634 856
rect 33802 800 33818 856
rect 33986 800 34186 856
rect 34354 800 34370 856
rect 34538 800 34738 856
rect 34906 800 34922 856
rect 35090 800 35106 856
rect 35274 800 35474 856
rect 35642 800 35658 856
rect 35826 800 36026 856
rect 36194 800 36210 856
rect 36378 800 36578 856
rect 36746 800 36762 856
rect 36930 800 37130 856
rect 37298 800 37314 856
rect 37482 800 37498 856
rect 37666 800 37866 856
rect 38034 800 38050 856
rect 38218 800 38418 856
rect 38586 800 38602 856
rect 38770 800 38970 856
rect 39138 800 39154 856
rect 39322 800 39522 856
rect 39690 800 39706 856
rect 39874 800 39890 856
rect 40058 800 40258 856
rect 40426 800 40442 856
rect 40610 800 40810 856
rect 40978 800 40994 856
rect 41162 800 41362 856
rect 41530 800 41546 856
rect 41714 800 41730 856
rect 41898 800 42098 856
rect 42266 800 42282 856
rect 42450 800 42650 856
rect 42818 800 42834 856
rect 43002 800 43202 856
rect 43370 800 43386 856
rect 43554 800 43754 856
rect 43922 800 43938 856
rect 44106 800 44122 856
rect 44290 800 44490 856
rect 44658 800 44674 856
rect 44842 800 45042 856
rect 45210 800 45226 856
rect 45394 800 45594 856
rect 45762 800 45778 856
rect 45946 800 46146 856
rect 46314 800 46330 856
rect 46498 800 46514 856
rect 46682 800 46882 856
rect 47050 800 47066 856
rect 47234 800 47434 856
rect 47602 800 47618 856
rect 47786 800 47986 856
rect 48154 800 48170 856
rect 48338 800 48538 856
rect 48706 800 48722 856
rect 48890 800 48906 856
rect 49074 800 49274 856
rect 49442 800 49458 856
rect 49626 800 49826 856
rect 49994 800 50010 856
rect 50178 800 50378 856
rect 50546 800 50562 856
rect 50730 800 50930 856
rect 51098 800 51114 856
rect 51282 800 51298 856
rect 51466 800 51666 856
rect 51834 800 51850 856
rect 52018 800 52218 856
rect 52386 800 52402 856
rect 52570 800 52770 856
rect 52938 800 52954 856
rect 53122 800 53322 856
rect 53490 800 53506 856
rect 53674 800 53690 856
rect 53858 800 54058 856
rect 54226 800 54242 856
rect 54410 800 54610 856
rect 54778 800 54794 856
rect 54962 800 55162 856
rect 55330 800 55346 856
rect 55514 800 55530 856
rect 55698 800 55898 856
rect 56066 800 56082 856
rect 56250 800 56450 856
rect 56618 800 56634 856
rect 56802 800 57002 856
rect 57170 800 57186 856
rect 57354 800 57554 856
rect 57722 800 57738 856
rect 57906 800 57922 856
rect 58090 800 58290 856
rect 58458 800 58474 856
rect 58642 800 58842 856
rect 59010 800 59026 856
rect 59194 800 59320 856
<< metal3 >>
rect 0 3544 800 3664
rect 59200 3544 60000 3664
rect 0 3000 800 3120
rect 0 2728 800 2848
rect 59200 3000 60000 3120
rect 59200 2728 60000 2848
rect 0 2184 800 2304
rect 1380 2290 58604 2350
rect 0 1912 800 2032
rect 59200 2184 60000 2304
rect 59200 1912 60000 2032
rect 59200 1640 60000 1760
rect 0 1368 800 1488
rect 0 1096 800 1216
rect 1380 1210 58604 1270
rect 59200 1096 60000 1216
rect 59200 824 60000 944
<< obsm3 >>
rect 880 3464 59120 3637
rect 800 3200 59200 3464
rect 880 2648 59120 3200
rect 800 2430 59200 2648
rect 800 2384 1300 2430
rect 880 2210 1300 2384
rect 58684 2384 59200 2430
rect 58684 2210 59120 2384
rect 880 1832 59120 2210
rect 800 1568 59120 1832
rect 880 1560 59120 1568
rect 880 1350 59200 1560
rect 880 1130 1300 1350
rect 58684 1296 59200 1350
rect 58684 1130 59120 1296
rect 880 1016 59120 1130
rect 800 851 59120 1016
<< labels >>
rlabel metal2 s 32954 3800 33010 4600 6 HI[0]
port 1 nsew signal output
rlabel metal3 s 59200 1912 60000 2032 6 HI[100]
port 2 nsew signal output
rlabel metal2 s 28906 3800 28962 4600 6 HI[101]
port 3 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 HI[102]
port 4 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 HI[103]
port 5 nsew signal output
rlabel metal2 s 9402 3800 9458 4600 6 HI[104]
port 6 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 HI[105]
port 7 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 HI[106]
port 8 nsew signal output
rlabel metal2 s 20442 3800 20498 4600 6 HI[107]
port 9 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 HI[108]
port 10 nsew signal output
rlabel metal2 s 13082 3800 13138 4600 6 HI[109]
port 11 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 HI[10]
port 12 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 HI[110]
port 13 nsew signal output
rlabel metal2 s 51722 3800 51778 4600 6 HI[111]
port 14 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 HI[112]
port 15 nsew signal output
rlabel metal2 s 28170 3800 28226 4600 6 HI[113]
port 16 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 HI[114]
port 17 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 HI[115]
port 18 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 HI[116]
port 19 nsew signal output
rlabel metal2 s 18970 3800 19026 4600 6 HI[117]
port 20 nsew signal output
rlabel metal2 s 46938 3800 46994 4600 6 HI[118]
port 21 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 HI[119]
port 22 nsew signal output
rlabel metal2 s 38290 3800 38346 4600 6 HI[11]
port 23 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 HI[120]
port 24 nsew signal output
rlabel metal2 s 12714 3800 12770 4600 6 HI[121]
port 25 nsew signal output
rlabel metal2 s 10322 3800 10378 4600 6 HI[122]
port 26 nsew signal output
rlabel metal2 s 14922 3800 14978 4600 6 HI[123]
port 27 nsew signal output
rlabel metal2 s 11794 3800 11850 4600 6 HI[124]
port 28 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 HI[125]
port 29 nsew signal output
rlabel metal2 s 46202 3800 46258 4600 6 HI[126]
port 30 nsew signal output
rlabel metal2 s 37738 3800 37794 4600 6 HI[127]
port 31 nsew signal output
rlabel metal2 s 54482 3800 54538 4600 6 HI[128]
port 32 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 HI[129]
port 33 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 HI[12]
port 34 nsew signal output
rlabel metal2 s 40130 3800 40186 4600 6 HI[130]
port 35 nsew signal output
rlabel metal2 s 19706 3800 19762 4600 6 HI[131]
port 36 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 HI[132]
port 37 nsew signal output
rlabel metal2 s 3698 3800 3754 4600 6 HI[133]
port 38 nsew signal output
rlabel metal2 s 54666 3800 54722 4600 6 HI[134]
port 39 nsew signal output
rlabel metal2 s 43258 3800 43314 4600 6 HI[135]
port 40 nsew signal output
rlabel metal2 s 58346 3800 58402 4600 6 HI[136]
port 41 nsew signal output
rlabel metal2 s 13266 3800 13322 4600 6 HI[137]
port 42 nsew signal output
rlabel metal2 s 4250 3800 4306 4600 6 HI[138]
port 43 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 HI[139]
port 44 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 HI[13]
port 45 nsew signal output
rlabel metal2 s 38842 3800 38898 4600 6 HI[140]
port 46 nsew signal output
rlabel metal2 s 58898 3800 58954 4600 6 HI[141]
port 47 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 HI[142]
port 48 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 HI[143]
port 49 nsew signal output
rlabel metal2 s 6090 3800 6146 4600 6 HI[144]
port 50 nsew signal output
rlabel metal2 s 43810 3800 43866 4600 6 HI[145]
port 51 nsew signal output
rlabel metal2 s 26330 3800 26386 4600 6 HI[146]
port 52 nsew signal output
rlabel metal2 s 59266 3800 59322 4600 6 HI[147]
port 53 nsew signal output
rlabel metal2 s 19154 3800 19210 4600 6 HI[148]
port 54 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 HI[149]
port 55 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 HI[14]
port 56 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 HI[150]
port 57 nsew signal output
rlabel metal2 s 39578 3800 39634 4600 6 HI[151]
port 58 nsew signal output
rlabel metal2 s 34794 3800 34850 4600 6 HI[152]
port 59 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 HI[153]
port 60 nsew signal output
rlabel metal2 s 18602 3800 18658 4600 6 HI[154]
port 61 nsew signal output
rlabel metal2 s 52274 3800 52330 4600 6 HI[155]
port 62 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 HI[156]
port 63 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 HI[157]
port 64 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 HI[158]
port 65 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 HI[159]
port 66 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 HI[15]
port 67 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 HI[160]
port 68 nsew signal output
rlabel metal2 s 53378 3800 53434 4600 6 HI[161]
port 69 nsew signal output
rlabel metal2 s 44178 3800 44234 4600 6 HI[162]
port 70 nsew signal output
rlabel metal2 s 37002 3800 37058 4600 6 HI[163]
port 71 nsew signal output
rlabel metal2 s 7746 3800 7802 4600 6 HI[164]
port 72 nsew signal output
rlabel metal2 s 39026 3800 39082 4600 6 HI[165]
port 73 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 HI[166]
port 74 nsew signal output
rlabel metal2 s 30562 3800 30618 4600 6 HI[167]
port 75 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 HI[168]
port 76 nsew signal output
rlabel metal2 s 5170 3800 5226 4600 6 HI[169]
port 77 nsew signal output
rlabel metal2 s 2962 3800 3018 4600 6 HI[16]
port 78 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 HI[170]
port 79 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 HI[171]
port 80 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 HI[172]
port 81 nsew signal output
rlabel metal2 s 55586 3800 55642 4600 6 HI[173]
port 82 nsew signal output
rlabel metal2 s 42522 3800 42578 4600 6 HI[174]
port 83 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 HI[175]
port 84 nsew signal output
rlabel metal2 s 938 0 994 800 6 HI[176]
port 85 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 HI[177]
port 86 nsew signal output
rlabel metal2 s 21546 3800 21602 4600 6 HI[178]
port 87 nsew signal output
rlabel metal2 s 33138 3800 33194 4600 6 HI[179]
port 88 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 HI[17]
port 89 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 HI[180]
port 90 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 HI[181]
port 91 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 HI[182]
port 92 nsew signal output
rlabel metal2 s 52642 3800 52698 4600 6 HI[183]
port 93 nsew signal output
rlabel metal2 s 24674 3800 24730 4600 6 HI[184]
port 94 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 HI[185]
port 95 nsew signal output
rlabel metal2 s 5354 3800 5410 4600 6 HI[186]
port 96 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 HI[187]
port 97 nsew signal output
rlabel metal2 s 35530 3800 35586 4600 6 HI[188]
port 98 nsew signal output
rlabel metal2 s 41234 3800 41290 4600 6 HI[189]
port 99 nsew signal output
rlabel metal2 s 14370 3800 14426 4600 6 HI[18]
port 100 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 HI[190]
port 101 nsew signal output
rlabel metal2 s 22650 3800 22706 4600 6 HI[191]
port 102 nsew signal output
rlabel metal2 s 12530 3800 12586 4600 6 HI[192]
port 103 nsew signal output
rlabel metal2 s 1674 3800 1730 4600 6 HI[193]
port 104 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 HI[194]
port 105 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 HI[195]
port 106 nsew signal output
rlabel metal2 s 41786 3800 41842 4600 6 HI[196]
port 107 nsew signal output
rlabel metal2 s 23386 3800 23442 4600 6 HI[197]
port 108 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 HI[198]
port 109 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 HI[199]
port 110 nsew signal output
rlabel metal2 s 31666 3800 31722 4600 6 HI[19]
port 111 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 HI[1]
port 112 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 HI[200]
port 113 nsew signal output
rlabel metal3 s 0 1912 800 2032 6 HI[201]
port 114 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 HI[202]
port 115 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 HI[203]
port 116 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 HI[204]
port 117 nsew signal output
rlabel metal2 s 7930 3800 7986 4600 6 HI[205]
port 118 nsew signal output
rlabel metal2 s 34058 3800 34114 4600 6 HI[206]
port 119 nsew signal output
rlabel metal2 s 24122 3800 24178 4600 6 HI[207]
port 120 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 HI[208]
port 121 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 HI[209]
port 122 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 HI[20]
port 123 nsew signal output
rlabel metal2 s 36634 3800 36690 4600 6 HI[210]
port 124 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 HI[211]
port 125 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 HI[212]
port 126 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 HI[213]
port 127 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 HI[214]
port 128 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 HI[215]
port 129 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 HI[216]
port 130 nsew signal output
rlabel metal2 s 8482 3800 8538 4600 6 HI[217]
port 131 nsew signal output
rlabel metal2 s 55218 3800 55274 4600 6 HI[218]
port 132 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 HI[219]
port 133 nsew signal output
rlabel metal2 s 27618 3800 27674 4600 6 HI[21]
port 134 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 HI[220]
port 135 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 HI[221]
port 136 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 HI[222]
port 137 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 HI[223]
port 138 nsew signal output
rlabel metal2 s 44362 3800 44418 4600 6 HI[224]
port 139 nsew signal output
rlabel metal2 s 754 3800 810 4600 6 HI[225]
port 140 nsew signal output
rlabel metal3 s 59200 3000 60000 3120 6 HI[226]
port 141 nsew signal output
rlabel metal2 s 50802 3800 50858 4600 6 HI[227]
port 142 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 HI[228]
port 143 nsew signal output
rlabel metal2 s 47306 3800 47362 4600 6 HI[229]
port 144 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 HI[22]
port 145 nsew signal output
rlabel metal2 s 39394 3800 39450 4600 6 HI[230]
port 146 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 HI[231]
port 147 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 HI[232]
port 148 nsew signal output
rlabel metal2 s 11426 3800 11482 4600 6 HI[233]
port 149 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 HI[234]
port 150 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 HI[235]
port 151 nsew signal output
rlabel metal2 s 4618 3800 4674 4600 6 HI[236]
port 152 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 HI[237]
port 153 nsew signal output
rlabel metal2 s 31298 3800 31354 4600 6 HI[238]
port 154 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 HI[239]
port 155 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 HI[23]
port 156 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 HI[240]
port 157 nsew signal output
rlabel metal2 s 42154 3800 42210 4600 6 HI[241]
port 158 nsew signal output
rlabel metal2 s 56322 3800 56378 4600 6 HI[242]
port 159 nsew signal output
rlabel metal2 s 50986 3800 51042 4600 6 HI[243]
port 160 nsew signal output
rlabel metal2 s 9034 3800 9090 4600 6 HI[244]
port 161 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 HI[245]
port 162 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 HI[246]
port 163 nsew signal output
rlabel metal2 s 7194 3800 7250 4600 6 HI[247]
port 164 nsew signal output
rlabel metal2 s 16946 3800 17002 4600 6 HI[248]
port 165 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 HI[249]
port 166 nsew signal output
rlabel metal2 s 41418 3800 41474 4600 6 HI[24]
port 167 nsew signal output
rlabel metal3 s 59200 3544 60000 3664 6 HI[250]
port 168 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 HI[251]
port 169 nsew signal output
rlabel metal2 s 47858 3800 47914 4600 6 HI[252]
port 170 nsew signal output
rlabel metal2 s 25594 3800 25650 4600 6 HI[253]
port 171 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 HI[254]
port 172 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 HI[255]
port 173 nsew signal output
rlabel metal2 s 45466 3800 45522 4600 6 HI[256]
port 174 nsew signal output
rlabel metal2 s 49330 3800 49386 4600 6 HI[257]
port 175 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 HI[258]
port 176 nsew signal output
rlabel metal2 s 12162 3800 12218 4600 6 HI[259]
port 177 nsew signal output
rlabel metal2 s 21730 3800 21786 4600 6 HI[25]
port 178 nsew signal output
rlabel metal2 s 29826 3800 29882 4600 6 HI[260]
port 179 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 HI[261]
port 180 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 HI[262]
port 181 nsew signal output
rlabel metal2 s 22282 3800 22338 4600 6 HI[263]
port 182 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 HI[264]
port 183 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 HI[265]
port 184 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 HI[266]
port 185 nsew signal output
rlabel metal2 s 25962 3800 26018 4600 6 HI[267]
port 186 nsew signal output
rlabel metal2 s 570 0 626 800 6 HI[268]
port 187 nsew signal output
rlabel metal2 s 48594 3800 48650 4600 6 HI[269]
port 188 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 HI[26]
port 189 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 HI[270]
port 190 nsew signal output
rlabel metal2 s 56874 3800 56930 4600 6 HI[271]
port 191 nsew signal output
rlabel metal2 s 27434 3800 27490 4600 6 HI[272]
port 192 nsew signal output
rlabel metal2 s 37186 3800 37242 4600 6 HI[273]
port 193 nsew signal output
rlabel metal2 s 43074 3800 43130 4600 6 HI[274]
port 194 nsew signal output
rlabel metal2 s 41970 3800 42026 4600 6 HI[275]
port 195 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 HI[276]
port 196 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 HI[277]
port 197 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 HI[278]
port 198 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 HI[279]
port 199 nsew signal output
rlabel metal2 s 28354 3800 28410 4600 6 HI[27]
port 200 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 HI[280]
port 201 nsew signal output
rlabel metal2 s 1306 3800 1362 4600 6 HI[281]
port 202 nsew signal output
rlabel metal2 s 27066 3800 27122 4600 6 HI[282]
port 203 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 HI[283]
port 204 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 HI[284]
port 205 nsew signal output
rlabel metal3 s 59200 2184 60000 2304 6 HI[285]
port 206 nsew signal output
rlabel metal2 s 16026 3800 16082 4600 6 HI[286]
port 207 nsew signal output
rlabel metal2 s 25226 3800 25282 4600 6 HI[287]
port 208 nsew signal output
rlabel metal2 s 40682 3800 40738 4600 6 HI[288]
port 209 nsew signal output
rlabel metal2 s 22098 3800 22154 4600 6 HI[289]
port 210 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 HI[28]
port 211 nsew signal output
rlabel metal2 s 39762 3800 39818 4600 6 HI[290]
port 212 nsew signal output
rlabel metal2 s 7010 3800 7066 4600 6 HI[291]
port 213 nsew signal output
rlabel metal2 s 2410 3800 2466 4600 6 HI[292]
port 214 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 HI[293]
port 215 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 HI[294]
port 216 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 HI[295]
port 217 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 HI[296]
port 218 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 HI[297]
port 219 nsew signal output
rlabel metal2 s 53562 3800 53618 4600 6 HI[298]
port 220 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 HI[299]
port 221 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 HI[29]
port 222 nsew signal output
rlabel metal2 s 42706 3800 42762 4600 6 HI[2]
port 223 nsew signal output
rlabel metal2 s 14554 3800 14610 4600 6 HI[300]
port 224 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 HI[301]
port 225 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 HI[302]
port 226 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 HI[303]
port 227 nsew signal output
rlabel metal2 s 10874 3800 10930 4600 6 HI[304]
port 228 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 HI[305]
port 229 nsew signal output
rlabel metal2 s 4802 3800 4858 4600 6 HI[306]
port 230 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 HI[307]
port 231 nsew signal output
rlabel metal2 s 10690 3800 10746 4600 6 HI[308]
port 232 nsew signal output
rlabel metal2 s 32770 3800 32826 4600 6 HI[309]
port 233 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 HI[30]
port 234 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 HI[310]
port 235 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 HI[311]
port 236 nsew signal output
rlabel metal2 s 2226 3800 2282 4600 6 HI[312]
port 237 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 HI[313]
port 238 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 HI[314]
port 239 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 HI[315]
port 240 nsew signal output
rlabel metal2 s 52826 3800 52882 4600 6 HI[316]
port 241 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 HI[317]
port 242 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 HI[318]
port 243 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 HI[319]
port 244 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 HI[31]
port 245 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 HI[320]
port 246 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 HI[321]
port 247 nsew signal output
rlabel metal2 s 57610 3800 57666 4600 6 HI[322]
port 248 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 HI[323]
port 249 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 HI[324]
port 250 nsew signal output
rlabel metal2 s 23754 3800 23810 4600 6 HI[325]
port 251 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 HI[326]
port 252 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 HI[327]
port 253 nsew signal output
rlabel metal2 s 35898 3800 35954 4600 6 HI[328]
port 254 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 HI[329]
port 255 nsew signal output
rlabel metal2 s 51538 3800 51594 4600 6 HI[32]
port 256 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 HI[330]
port 257 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 HI[331]
port 258 nsew signal output
rlabel metal2 s 33690 3800 33746 4600 6 HI[332]
port 259 nsew signal output
rlabel metal2 s 40866 3800 40922 4600 6 HI[333]
port 260 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 HI[334]
port 261 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 HI[335]
port 262 nsew signal output
rlabel metal2 s 57978 3800 58034 4600 6 HI[336]
port 263 nsew signal output
rlabel metal2 s 45098 3800 45154 4600 6 HI[337]
port 264 nsew signal output
rlabel metal2 s 36450 3800 36506 4600 6 HI[338]
port 265 nsew signal output
rlabel metal2 s 11242 3800 11298 4600 6 HI[339]
port 266 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 HI[33]
port 267 nsew signal output
rlabel metal2 s 32402 3800 32458 4600 6 HI[340]
port 268 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 HI[341]
port 269 nsew signal output
rlabel metal2 s 25042 3800 25098 4600 6 HI[342]
port 270 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 HI[343]
port 271 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 HI[344]
port 272 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 HI[345]
port 273 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 HI[346]
port 274 nsew signal output
rlabel metal2 s 19890 3800 19946 4600 6 HI[347]
port 275 nsew signal output
rlabel metal2 s 23938 3800 23994 4600 6 HI[348]
port 276 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 HI[349]
port 277 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 HI[34]
port 278 nsew signal output
rlabel metal2 s 5906 3800 5962 4600 6 HI[350]
port 279 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 HI[351]
port 280 nsew signal output
rlabel metal2 s 48042 3800 48098 4600 6 HI[352]
port 281 nsew signal output
rlabel metal2 s 16578 3800 16634 4600 6 HI[353]
port 282 nsew signal output
rlabel metal2 s 44914 3800 44970 4600 6 HI[354]
port 283 nsew signal output
rlabel metal2 s 6458 3800 6514 4600 6 HI[355]
port 284 nsew signal output
rlabel metal2 s 50434 3800 50490 4600 6 HI[356]
port 285 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 HI[357]
port 286 nsew signal output
rlabel metal2 s 35346 3800 35402 4600 6 HI[358]
port 287 nsew signal output
rlabel metal2 s 43626 3800 43682 4600 6 HI[359]
port 288 nsew signal output
rlabel metal2 s 54114 3800 54170 4600 6 HI[35]
port 289 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 HI[360]
port 290 nsew signal output
rlabel metal3 s 59200 1640 60000 1760 6 HI[361]
port 291 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 HI[362]
port 292 nsew signal output
rlabel metal3 s 59200 1096 60000 1216 6 HI[363]
port 293 nsew signal output
rlabel metal2 s 29274 3800 29330 4600 6 HI[364]
port 294 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 HI[365]
port 295 nsew signal output
rlabel metal2 s 27986 3800 28042 4600 6 HI[366]
port 296 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 HI[367]
port 297 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 HI[368]
port 298 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 HI[369]
port 299 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 HI[36]
port 300 nsew signal output
rlabel metal2 s 49882 3800 49938 4600 6 HI[370]
port 301 nsew signal output
rlabel metal3 s 0 1096 800 1216 6 HI[371]
port 302 nsew signal output
rlabel metal2 s 21362 3800 21418 4600 6 HI[372]
port 303 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 HI[373]
port 304 nsew signal output
rlabel metal2 s 29458 3800 29514 4600 6 HI[374]
port 305 nsew signal output
rlabel metal2 s 26514 3800 26570 4600 6 HI[375]
port 306 nsew signal output
rlabel metal2 s 53930 3800 53986 4600 6 HI[376]
port 307 nsew signal output
rlabel metal2 s 9586 3800 9642 4600 6 HI[377]
port 308 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 HI[378]
port 309 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 HI[379]
port 310 nsew signal output
rlabel metal2 s 16762 3800 16818 4600 6 HI[37]
port 311 nsew signal output
rlabel metal2 s 38474 3800 38530 4600 6 HI[380]
port 312 nsew signal output
rlabel metal2 s 570 3800 626 4600 6 HI[381]
port 313 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 HI[382]
port 314 nsew signal output
rlabel metal2 s 6642 3800 6698 4600 6 HI[383]
port 315 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 HI[384]
port 316 nsew signal output
rlabel metal2 s 30010 3800 30066 4600 6 HI[385]
port 317 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 HI[386]
port 318 nsew signal output
rlabel metal2 s 45650 3800 45706 4600 6 HI[387]
port 319 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 HI[388]
port 320 nsew signal output
rlabel metal2 s 31850 3800 31906 4600 6 HI[389]
port 321 nsew signal output
rlabel metal2 s 23202 3800 23258 4600 6 HI[38]
port 322 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 HI[390]
port 323 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 HI[391]
port 324 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 HI[392]
port 325 nsew signal output
rlabel metal2 s 47490 3800 47546 4600 6 HI[393]
port 326 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 HI[394]
port 327 nsew signal output
rlabel metal2 s 20994 3800 21050 4600 6 HI[395]
port 328 nsew signal output
rlabel metal2 s 57058 3800 57114 4600 6 HI[396]
port 329 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 HI[397]
port 330 nsew signal output
rlabel metal2 s 28722 3800 28778 4600 6 HI[398]
port 331 nsew signal output
rlabel metal2 s 22834 3800 22890 4600 6 HI[399]
port 332 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 HI[39]
port 333 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 HI[3]
port 334 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 HI[400]
port 335 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 HI[401]
port 336 nsew signal output
rlabel metal2 s 15658 3800 15714 4600 6 HI[402]
port 337 nsew signal output
rlabel metal2 s 7562 3800 7618 4600 6 HI[403]
port 338 nsew signal output
rlabel metal2 s 56506 3800 56562 4600 6 HI[404]
port 339 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 HI[405]
port 340 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 HI[406]
port 341 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 HI[407]
port 342 nsew signal output
rlabel metal2 s 8850 3800 8906 4600 6 HI[408]
port 343 nsew signal output
rlabel metal2 s 37554 3800 37610 4600 6 HI[409]
port 344 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 HI[40]
port 345 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 HI[410]
port 346 nsew signal output
rlabel metal2 s 2410 0 2466 800 6 HI[411]
port 347 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 HI[412]
port 348 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 HI[413]
port 349 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 HI[414]
port 350 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 HI[415]
port 351 nsew signal output
rlabel metal2 s 30378 3800 30434 4600 6 HI[416]
port 352 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 HI[417]
port 353 nsew signal output
rlabel metal2 s 55770 3800 55826 4600 6 HI[418]
port 354 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 HI[419]
port 355 nsew signal output
rlabel metal2 s 34242 3800 34298 4600 6 HI[41]
port 356 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 HI[420]
port 357 nsew signal output
rlabel metal2 s 15106 3800 15162 4600 6 HI[421]
port 358 nsew signal output
rlabel metal2 s 11978 3800 12034 4600 6 HI[422]
port 359 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 HI[423]
port 360 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 HI[424]
port 361 nsew signal output
rlabel metal2 s 58162 3800 58218 4600 6 HI[425]
port 362 nsew signal output
rlabel metal2 s 9954 3800 10010 4600 6 HI[426]
port 363 nsew signal output
rlabel metal2 s 58714 3800 58770 4600 6 HI[427]
port 364 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 HI[428]
port 365 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 HI[429]
port 366 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 HI[42]
port 367 nsew signal output
rlabel metal2 s 36082 3800 36138 4600 6 HI[430]
port 368 nsew signal output
rlabel metal2 s 34610 3800 34666 4600 6 HI[431]
port 369 nsew signal output
rlabel metal2 s 17314 3800 17370 4600 6 HI[432]
port 370 nsew signal output
rlabel metal2 s 18050 3800 18106 4600 6 HI[433]
port 371 nsew signal output
rlabel metal2 s 48410 3800 48466 4600 6 HI[434]
port 372 nsew signal output
rlabel metal2 s 16210 3800 16266 4600 6 HI[435]
port 373 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 HI[436]
port 374 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 HI[437]
port 375 nsew signal output
rlabel metal2 s 55034 3800 55090 4600 6 HI[438]
port 376 nsew signal output
rlabel metal3 s 59200 2728 60000 2848 6 HI[439]
port 377 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 HI[43]
port 378 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 HI[440]
port 379 nsew signal output
rlabel metal2 s 46754 3800 46810 4600 6 HI[441]
port 380 nsew signal output
rlabel metal2 s 13818 3800 13874 4600 6 HI[442]
port 381 nsew signal output
rlabel metal2 s 52090 3800 52146 4600 6 HI[443]
port 382 nsew signal output
rlabel metal2 s 14186 3800 14242 4600 6 HI[444]
port 383 nsew signal output
rlabel metal2 s 25778 3800 25834 4600 6 HI[445]
port 384 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 HI[446]
port 385 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 HI[447]
port 386 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 HI[448]
port 387 nsew signal output
rlabel metal2 s 1490 0 1546 800 6 HI[449]
port 388 nsew signal output
rlabel metal2 s 8298 3800 8354 4600 6 HI[44]
port 389 nsew signal output
rlabel metal2 s 18418 3800 18474 4600 6 HI[450]
port 390 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 HI[451]
port 391 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 HI[452]
port 392 nsew signal output
rlabel metal2 s 5538 3800 5594 4600 6 HI[453]
port 393 nsew signal output
rlabel metal2 s 24490 3800 24546 4600 6 HI[454]
port 394 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 HI[455]
port 395 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 HI[456]
port 396 nsew signal output
rlabel metal2 s 17866 3800 17922 4600 6 HI[457]
port 397 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 HI[458]
port 398 nsew signal output
rlabel metal2 s 40314 3800 40370 4600 6 HI[45]
port 399 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 HI[46]
port 400 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 HI[47]
port 401 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 HI[48]
port 402 nsew signal output
rlabel metal2 s 30746 3800 30802 4600 6 HI[49]
port 403 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 HI[4]
port 404 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 HI[50]
port 405 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 HI[51]
port 406 nsew signal output
rlabel metal2 s 48962 3800 49018 4600 6 HI[52]
port 407 nsew signal output
rlabel metal2 s 20258 3800 20314 4600 6 HI[53]
port 408 nsew signal output
rlabel metal2 s 57426 3800 57482 4600 6 HI[54]
port 409 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 HI[55]
port 410 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 HI[56]
port 411 nsew signal output
rlabel metal2 s 55954 3800 56010 4600 6 HI[57]
port 412 nsew signal output
rlabel metal2 s 19338 3800 19394 4600 6 HI[58]
port 413 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 HI[59]
port 414 nsew signal output
rlabel metal2 s 35162 3800 35218 4600 6 HI[5]
port 415 nsew signal output
rlabel metal2 s 50250 3800 50306 4600 6 HI[60]
port 416 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 HI[61]
port 417 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 HI[62]
port 418 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 HI[63]
port 419 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 HI[64]
port 420 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 HI[65]
port 421 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 HI[66]
port 422 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 HI[67]
port 423 nsew signal output
rlabel metal2 s 754 0 810 800 6 HI[68]
port 424 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 HI[69]
port 425 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 HI[6]
port 426 nsew signal output
rlabel metal2 s 3514 3800 3570 4600 6 HI[70]
port 427 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 HI[71]
port 428 nsew signal output
rlabel metal2 s 4066 3800 4122 4600 6 HI[72]
port 429 nsew signal output
rlabel metal2 s 13634 3800 13690 4600 6 HI[73]
port 430 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 HI[74]
port 431 nsew signal output
rlabel metal2 s 49698 3800 49754 4600 6 HI[75]
port 432 nsew signal output
rlabel metal2 s 44546 3800 44602 4600 6 HI[76]
port 433 nsew signal output
rlabel metal2 s 33506 3800 33562 4600 6 HI[77]
port 434 nsew signal output
rlabel metal2 s 49146 3800 49202 4600 6 HI[78]
port 435 nsew signal output
rlabel metal2 s 46570 3800 46626 4600 6 HI[79]
port 436 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 HI[7]
port 437 nsew signal output
rlabel metal2 s 32218 3800 32274 4600 6 HI[80]
port 438 nsew signal output
rlabel metal2 s 51354 3800 51410 4600 6 HI[81]
port 439 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 HI[82]
port 440 nsew signal output
rlabel metal2 s 17498 3800 17554 4600 6 HI[83]
port 441 nsew signal output
rlabel metal2 s 20810 3800 20866 4600 6 HI[84]
port 442 nsew signal output
rlabel metal2 s 10138 3800 10194 4600 6 HI[85]
port 443 nsew signal output
rlabel metal2 s 31114 3800 31170 4600 6 HI[86]
port 444 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 HI[87]
port 445 nsew signal output
rlabel metal2 s 53194 3800 53250 4600 6 HI[88]
port 446 nsew signal output
rlabel metal2 s 1858 3800 1914 4600 6 HI[89]
port 447 nsew signal output
rlabel metal2 s 37922 3800 37978 4600 6 HI[8]
port 448 nsew signal output
rlabel metal2 s 1122 3800 1178 4600 6 HI[90]
port 449 nsew signal output
rlabel metal2 s 26882 3800 26938 4600 6 HI[91]
port 450 nsew signal output
rlabel metal2 s 3146 3800 3202 4600 6 HI[92]
port 451 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 HI[93]
port 452 nsew signal output
rlabel metal2 s 46018 3800 46074 4600 6 HI[94]
port 453 nsew signal output
rlabel metal2 s 2778 3800 2834 4600 6 HI[95]
port 454 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 HI[96]
port 455 nsew signal output
rlabel metal2 s 15474 3800 15530 4600 6 HI[97]
port 456 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 HI[98]
port 457 nsew signal output
rlabel metal3 s 59200 824 60000 944 6 HI[99]
port 458 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 HI[9]
port 459 nsew signal output
rlabel metal2 s 51350 1040 51410 3312 6 vccd1
port 460 nsew power bidirectional
rlabel metal2 s 35350 1040 35410 3312 6 vccd1
port 461 nsew power bidirectional
rlabel metal2 s 19350 1040 19410 3312 6 vccd1
port 462 nsew power bidirectional
rlabel metal2 s 3350 1040 3410 3312 6 vccd1
port 463 nsew power bidirectional
rlabel metal3 s 1380 1210 58604 1270 6 vccd1
port 464 nsew power bidirectional
rlabel metal2 s 43350 1040 43410 3312 6 vssd1
port 465 nsew ground bidirectional
rlabel metal2 s 27350 1040 27410 3312 6 vssd1
port 466 nsew ground bidirectional
rlabel metal2 s 11350 1040 11410 3312 6 vssd1
port 467 nsew ground bidirectional
rlabel metal3 s 1380 2290 58604 2350 6 vssd1
port 468 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60000 4600
string LEFview TRUE
<< end >>
