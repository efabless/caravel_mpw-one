magic
tech sky130A
magscale 1 2
timestamp 1605708945
<< pdiff >>
rect 80158 1034729 80192 1034755
rect 81392 1034729 81426 1034755
rect 134758 1034729 134792 1034755
rect 135992 1034729 136026 1034755
rect 189358 1034729 189392 1034755
rect 190592 1034729 190626 1034755
rect 243958 1034729 243992 1034755
rect 245192 1034729 245226 1034755
rect 298558 1034729 298592 1034755
rect 299792 1034729 299826 1034755
rect 406558 1034729 406592 1034755
rect 407792 1034729 407826 1034755
rect 461158 1034729 461192 1034755
rect 462392 1034729 462426 1034755
rect 515758 1034729 515792 1034755
rect 516992 1034729 517026 1034755
rect 623958 1034729 623992 1034755
rect 625192 1034729 625226 1034755
rect 85440 1032412 92551 1032434
rect 94386 1031622 94400 1032466
rect 140040 1032412 147151 1032434
rect 148986 1031622 149000 1032466
rect 194640 1032412 201751 1032434
rect 203586 1031622 203600 1032466
rect 249240 1032412 256351 1032434
rect 258186 1031622 258200 1032466
rect 303840 1032412 310951 1032434
rect 312786 1031622 312800 1032466
rect 411840 1032412 418951 1032434
rect 420786 1031622 420800 1032466
rect 466440 1032412 473551 1032434
rect 475386 1031622 475400 1032466
rect 521040 1032412 528151 1032434
rect 529986 1031622 530000 1032466
rect 629240 1032412 636351 1032434
rect 638186 1031622 638200 1032466
rect 94376 1031608 94400 1031622
rect 148976 1031608 149000 1031622
rect 203576 1031608 203600 1031622
rect 258176 1031608 258200 1031622
rect 312776 1031608 312800 1031622
rect 420776 1031608 420800 1031622
rect 475376 1031608 475400 1031622
rect 529976 1031608 530000 1031622
rect 638176 1031608 638200 1031622
rect 80370 1031582 92551 1031598
rect 92594 1031582 94400 1031608
rect 134970 1031582 147151 1031598
rect 147194 1031582 149000 1031608
rect 189570 1031582 201751 1031598
rect 201794 1031582 203600 1031608
rect 244170 1031582 256351 1031598
rect 256394 1031582 258200 1031608
rect 298770 1031582 310951 1031598
rect 310994 1031582 312800 1031608
rect 406770 1031582 418951 1031598
rect 418994 1031582 420800 1031608
rect 461370 1031582 473551 1031598
rect 473594 1031582 475400 1031608
rect 515970 1031582 528151 1031598
rect 528194 1031582 530000 1031608
rect 624170 1031582 636351 1031598
rect 636394 1031582 638200 1031608
rect 81005 1029214 81167 1030214
rect 93291 1029214 93332 1030214
rect 93853 1029214 94063 1030214
rect 135605 1029214 135767 1030214
rect 147891 1029214 147932 1030214
rect 148453 1029214 148663 1030214
rect 190205 1029214 190367 1030214
rect 202491 1029214 202532 1030214
rect 203053 1029214 203263 1030214
rect 244805 1029214 244967 1030214
rect 257091 1029214 257132 1030214
rect 257653 1029214 257863 1030214
rect 299405 1029214 299567 1030214
rect 311691 1029214 311732 1030214
rect 312253 1029214 312463 1030214
rect 407405 1029214 407567 1030214
rect 419691 1029214 419732 1030214
rect 420253 1029214 420463 1030214
rect 462005 1029214 462167 1030214
rect 474291 1029214 474332 1030214
rect 474853 1029214 475063 1030214
rect 516605 1029214 516767 1030214
rect 528891 1029214 528932 1030214
rect 529453 1029214 529663 1030214
rect 624805 1029214 624967 1030214
rect 637091 1029214 637132 1030214
rect 637653 1029214 637863 1030214
rect 81028 1027613 81168 1028613
rect 93291 1027613 93332 1028613
rect 93853 1027613 94063 1028613
rect 135628 1027613 135768 1028613
rect 147891 1027613 147932 1028613
rect 148453 1027613 148663 1028613
rect 190228 1027613 190368 1028613
rect 202491 1027613 202532 1028613
rect 203053 1027613 203263 1028613
rect 244828 1027613 244968 1028613
rect 257091 1027613 257132 1028613
rect 257653 1027613 257863 1028613
rect 299428 1027613 299568 1028613
rect 311691 1027613 311732 1028613
rect 312253 1027613 312463 1028613
rect 407428 1027613 407568 1028613
rect 419691 1027613 419732 1028613
rect 420253 1027613 420463 1028613
rect 462028 1027613 462168 1028613
rect 474291 1027613 474332 1028613
rect 474853 1027613 475063 1028613
rect 516628 1027613 516768 1028613
rect 528891 1027613 528932 1028613
rect 529453 1027613 529663 1028613
rect 624828 1027613 624968 1028613
rect 637091 1027613 637132 1028613
rect 637653 1027613 637863 1028613
rect 79904 1018113 80052 1022859
rect 80569 1020925 80595 1021925
rect 80640 1020925 80742 1021925
rect 93808 1020925 93963 1021925
rect 94133 1020925 94288 1021925
rect 80569 1019325 80595 1020325
rect 80640 1019325 80742 1020325
rect 93808 1019325 93963 1020325
rect 94133 1019325 94288 1020325
rect 134504 1018113 134652 1022859
rect 135169 1020925 135195 1021925
rect 135240 1020925 135342 1021925
rect 148408 1020925 148563 1021925
rect 148733 1020925 148888 1021925
rect 135169 1019325 135195 1020325
rect 135240 1019325 135342 1020325
rect 148408 1019325 148563 1020325
rect 148733 1019325 148888 1020325
rect 189104 1018113 189252 1022859
rect 189769 1020925 189795 1021925
rect 189840 1020925 189942 1021925
rect 203008 1020925 203163 1021925
rect 203333 1020925 203488 1021925
rect 189769 1019325 189795 1020325
rect 189840 1019325 189942 1020325
rect 203008 1019325 203163 1020325
rect 203333 1019325 203488 1020325
rect 243704 1018113 243852 1022859
rect 244369 1020925 244395 1021925
rect 244440 1020925 244542 1021925
rect 257608 1020925 257763 1021925
rect 257933 1020925 258088 1021925
rect 244369 1019325 244395 1020325
rect 244440 1019325 244542 1020325
rect 257608 1019325 257763 1020325
rect 257933 1019325 258088 1020325
rect 298304 1018113 298452 1022859
rect 298969 1020925 298995 1021925
rect 299040 1020925 299142 1021925
rect 312208 1020925 312363 1021925
rect 312533 1020925 312688 1021925
rect 298969 1019325 298995 1020325
rect 299040 1019325 299142 1020325
rect 312208 1019325 312363 1020325
rect 312533 1019325 312688 1020325
rect 406304 1018113 406452 1022859
rect 406969 1020925 406995 1021925
rect 407040 1020925 407142 1021925
rect 420208 1020925 420363 1021925
rect 420533 1020925 420688 1021925
rect 406969 1019325 406995 1020325
rect 407040 1019325 407142 1020325
rect 420208 1019325 420363 1020325
rect 420533 1019325 420688 1020325
rect 460904 1018113 461052 1022859
rect 461569 1020925 461595 1021925
rect 461640 1020925 461742 1021925
rect 474808 1020925 474963 1021925
rect 475133 1020925 475288 1021925
rect 461569 1019325 461595 1020325
rect 461640 1019325 461742 1020325
rect 474808 1019325 474963 1020325
rect 475133 1019325 475288 1020325
rect 515504 1018113 515652 1022859
rect 516169 1020925 516195 1021925
rect 516240 1020925 516342 1021925
rect 529408 1020925 529563 1021925
rect 529733 1020925 529888 1021925
rect 516169 1019325 516195 1020325
rect 516240 1019325 516342 1020325
rect 529408 1019325 529563 1020325
rect 529733 1019325 529888 1020325
rect 623704 1018113 623852 1022859
rect 624369 1020925 624395 1021925
rect 624440 1020925 624542 1021925
rect 637608 1020925 637763 1021925
rect 637933 1020925 638088 1021925
rect 624369 1019325 624395 1020325
rect 624440 1019325 624542 1020325
rect 637608 1019325 637763 1020325
rect 637933 1019325 638088 1020325
rect 80078 1018056 87002 1018087
rect 134678 1018056 141602 1018087
rect 189278 1018056 196202 1018087
rect 243878 1018056 250802 1018087
rect 298478 1018056 305402 1018087
rect 406478 1018056 413402 1018087
rect 461078 1018056 468002 1018087
rect 515678 1018056 522602 1018087
rect 623878 1018056 630802 1018087
rect 87006 1016820 88211 1016824
rect 141606 1016820 142811 1016824
rect 196206 1016820 197411 1016824
rect 250806 1016820 252011 1016824
rect 305406 1016820 306611 1016824
rect 413406 1016820 414611 1016824
rect 468006 1016820 469211 1016824
rect 522606 1016820 523811 1016824
rect 630806 1016820 632011 1016824
rect 80787 1016782 80843 1016794
rect 135387 1016782 135443 1016794
rect 189987 1016782 190043 1016794
rect 244587 1016782 244643 1016794
rect 299187 1016782 299243 1016794
rect 407187 1016782 407243 1016794
rect 461787 1016782 461843 1016794
rect 516387 1016782 516443 1016794
rect 624587 1016782 624643 1016794
rect 87632 1007761 88080 1007767
rect 90678 1007761 91152 1007767
rect 142232 1007761 142680 1007767
rect 145278 1007761 145752 1007767
rect 196832 1007761 197280 1007767
rect 199878 1007761 200352 1007767
rect 251432 1007761 251880 1007767
rect 254478 1007761 254952 1007767
rect 306032 1007761 306480 1007767
rect 309078 1007761 309552 1007767
rect 414032 1007761 414480 1007767
rect 417078 1007761 417552 1007767
rect 468632 1007761 469080 1007767
rect 471678 1007761 472152 1007767
rect 523232 1007761 523680 1007767
rect 526278 1007761 526752 1007767
rect 631432 1007761 631880 1007767
rect 634478 1007761 634952 1007767
rect 85804 1007648 91357 1007651
rect 140404 1007648 145957 1007651
rect 195004 1007648 200557 1007651
rect 249604 1007648 255157 1007651
rect 304204 1007648 309757 1007651
rect 412204 1007648 417757 1007651
rect 466804 1007648 472357 1007651
rect 521404 1007648 526957 1007651
rect 629604 1007648 635157 1007651
rect 86597 1007576 92346 1007588
rect 141197 1007576 146946 1007588
rect 195797 1007576 201546 1007588
rect 250397 1007576 256146 1007588
rect 304997 1007576 310746 1007588
rect 412997 1007576 418746 1007588
rect 467597 1007576 473346 1007588
rect 522197 1007576 527946 1007588
rect 630397 1007576 636146 1007588
rect 86597 1006885 86623 1007576
rect 141197 1006885 141223 1007576
rect 195797 1006885 195823 1007576
rect 250397 1006885 250423 1007576
rect 304997 1006885 305023 1007576
rect 412997 1006885 413023 1007576
rect 467597 1006885 467623 1007576
rect 522197 1006885 522223 1007576
rect 630397 1006885 630423 1007576
rect 86613 1006882 86623 1006885
rect 141213 1006882 141223 1006885
rect 195813 1006882 195823 1006885
rect 250413 1006882 250423 1006885
rect 305013 1006882 305023 1006885
rect 413013 1006882 413023 1006885
rect 467613 1006882 467623 1006885
rect 522213 1006882 522223 1006885
rect 630413 1006882 630423 1006885
rect 82785 1005806 82801 1006122
rect 83989 1005806 84007 1006122
rect 137385 1005806 137401 1006122
rect 138589 1005806 138607 1006122
rect 191985 1005806 192001 1006122
rect 193189 1005806 193207 1006122
rect 246585 1005806 246601 1006122
rect 247789 1005806 247807 1006122
rect 301185 1005806 301201 1006122
rect 302389 1005806 302407 1006122
rect 409185 1005806 409201 1006122
rect 410389 1005806 410407 1006122
rect 463785 1005806 463801 1006122
rect 464989 1005806 465007 1006122
rect 518385 1005806 518401 1006122
rect 519589 1005806 519607 1006122
rect 626585 1005806 626601 1006122
rect 627789 1005806 627807 1006122
rect 82785 1005780 82789 1005806
rect 137385 1005780 137389 1005806
rect 191985 1005780 191989 1005806
rect 246585 1005780 246589 1005806
rect 301185 1005780 301189 1005806
rect 409185 1005780 409189 1005806
rect 463785 1005780 463789 1005806
rect 518385 1005780 518389 1005806
rect 626585 1005780 626589 1005806
rect 82751 1005542 82789 1005780
rect 84009 1005542 84041 1005780
rect 137351 1005542 137389 1005780
rect 138609 1005542 138641 1005780
rect 191951 1005542 191989 1005780
rect 193209 1005542 193241 1005780
rect 246551 1005542 246589 1005780
rect 247809 1005542 247841 1005780
rect 301151 1005542 301189 1005780
rect 302409 1005542 302441 1005780
rect 409151 1005542 409189 1005780
rect 410409 1005542 410441 1005780
rect 463751 1005542 463789 1005780
rect 465009 1005542 465041 1005780
rect 518351 1005542 518389 1005780
rect 519609 1005542 519641 1005780
rect 626551 1005542 626589 1005780
rect 627809 1005542 627841 1005780
rect 83574 1001505 84064 1001532
rect 138174 1001505 138664 1001532
rect 192774 1001505 193264 1001532
rect 247374 1001505 247864 1001532
rect 301974 1001505 302464 1001532
rect 409974 1001505 410464 1001532
rect 464574 1001505 465064 1001532
rect 519174 1001505 519664 1001532
rect 627374 1001505 627864 1001532
rect 88082 998649 88108 998657
rect 91292 998649 91317 998657
rect 142682 998649 142708 998657
rect 145892 998649 145917 998657
rect 197282 998649 197308 998657
rect 200492 998649 200517 998657
rect 251882 998649 251908 998657
rect 255092 998649 255117 998657
rect 306482 998649 306508 998657
rect 309692 998649 309717 998657
rect 414482 998649 414508 998657
rect 417692 998649 417717 998657
rect 469082 998649 469108 998657
rect 472292 998649 472317 998657
rect 523682 998649 523708 998657
rect 526892 998649 526917 998657
rect 631882 998649 631908 998657
rect 635092 998649 635117 998657
rect 5000 968324 5884 968338
rect 5844 968314 5884 968324
rect 5858 966532 5884 968314
rect 15541 968071 16541 968226
rect 17141 968071 18141 968226
rect 7252 967791 8252 968001
rect 8853 967791 9853 968001
rect 15541 967746 16541 967901
rect 17141 967746 18141 967901
rect 7252 967229 8252 967270
rect 8853 967229 9853 967270
rect 5032 959378 5054 966489
rect 2711 955330 2737 955364
rect 5868 954308 5884 966489
rect 29699 964616 29705 965090
rect 20642 960944 20646 962149
rect 29699 961570 29705 962018
rect 7252 954943 8252 955105
rect 8853 954966 9853 955106
rect 15541 954578 16541 954680
rect 17141 954578 18141 954680
rect 15541 954507 16541 954533
rect 17141 954507 18141 954533
rect 2711 954096 2737 954130
rect 19379 954016 19410 960940
rect 29815 959742 29818 965295
rect 29878 960561 29890 966284
rect 38809 965230 38817 965255
rect 697975 965214 702721 965362
rect 696644 964423 696656 964479
rect 685404 962481 685642 962515
rect 685404 962477 685984 962481
rect 685668 962465 685984 962477
rect 38809 962020 38817 962046
rect 681367 961202 681394 961692
rect 685668 961259 685984 961277
rect 685404 961225 685642 961257
rect 29878 960551 30584 960561
rect 29878 960535 30581 960551
rect 686747 958653 687450 958669
rect 686744 958643 687450 958653
rect 31686 957947 31924 957979
rect 31344 957927 31660 957945
rect 35934 957512 35961 958002
rect 678511 957158 678519 957184
rect 31344 956727 31660 956739
rect 31344 956723 31924 956727
rect 31686 956689 31924 956723
rect 20672 954725 20684 954781
rect 14607 953842 19353 953990
rect 678511 953949 678519 953974
rect 687438 952920 687450 958643
rect 687510 953909 687513 959462
rect 697918 958264 697949 965188
rect 714591 965074 714617 965108
rect 699187 964671 700187 964697
rect 700787 964671 701787 964697
rect 699187 964524 700187 964626
rect 700787 964524 701787 964626
rect 707475 964098 708475 964238
rect 709076 964099 710076 964261
rect 687623 957186 687629 957634
rect 696682 957055 696686 958260
rect 687623 954114 687629 954588
rect 711444 952715 711460 964896
rect 714591 963840 714617 963874
rect 712274 952715 712296 959826
rect 707475 951934 708475 951975
rect 709076 951934 710076 951975
rect 699187 951303 700187 951458
rect 700787 951303 701787 951458
rect 707475 951203 708475 951413
rect 709076 951203 710076 951413
rect 699187 950978 700187 951133
rect 700787 950978 701787 951133
rect 711444 950890 711470 952672
rect 711444 950880 711484 950890
rect 711444 950866 712328 950880
rect 35794 916717 39182 916731
rect 678146 916189 681534 916247
rect 35794 912757 39182 912815
rect 678146 912273 681534 912287
rect 697975 873014 702721 873162
rect 696644 872223 696656 872279
rect 685404 870281 685642 870315
rect 685404 870277 685984 870281
rect 685668 870265 685984 870277
rect 681367 869002 681394 869492
rect 685668 869059 685984 869077
rect 685404 869025 685642 869057
rect 686747 866453 687450 866469
rect 686744 866443 687450 866453
rect 678511 864958 678519 864984
rect 678511 861749 678519 861774
rect 687438 860720 687450 866443
rect 687510 861709 687513 867262
rect 697918 866064 697949 872988
rect 714591 872874 714617 872908
rect 699187 872471 700187 872497
rect 700787 872471 701787 872497
rect 699187 872324 700187 872426
rect 700787 872324 701787 872426
rect 707475 871898 708475 872038
rect 709076 871899 710076 872061
rect 687623 864986 687629 865434
rect 696682 864855 696686 866060
rect 687623 861914 687629 862388
rect 711444 860515 711460 872696
rect 714591 871640 714617 871674
rect 712274 860515 712296 867626
rect 707475 859734 708475 859775
rect 709076 859734 710076 859775
rect 699187 859103 700187 859258
rect 700787 859103 701787 859258
rect 707475 859003 708475 859213
rect 709076 859003 710076 859213
rect 699187 858778 700187 858933
rect 700787 858778 701787 858933
rect 711444 858690 711470 860472
rect 711444 858680 711484 858690
rect 711444 858666 712328 858680
rect 5000 793124 5884 793138
rect 5844 793114 5884 793124
rect 5858 791332 5884 793114
rect 15541 792871 16541 793026
rect 17141 792871 18141 793026
rect 7252 792591 8252 792801
rect 8853 792591 9853 792801
rect 15541 792546 16541 792701
rect 17141 792546 18141 792701
rect 7252 792029 8252 792070
rect 8853 792029 9853 792070
rect 5032 784178 5054 791289
rect 2711 780130 2737 780164
rect 5868 779108 5884 791289
rect 29699 789416 29705 789890
rect 20642 785744 20646 786949
rect 29699 786370 29705 786818
rect 7252 779743 8252 779905
rect 8853 779766 9853 779906
rect 15541 779378 16541 779480
rect 17141 779378 18141 779480
rect 15541 779307 16541 779333
rect 17141 779307 18141 779333
rect 2711 778896 2737 778930
rect 19379 778816 19410 785740
rect 29815 784542 29818 790095
rect 29878 785361 29890 791084
rect 38809 790030 38817 790055
rect 38809 786820 38817 786846
rect 29878 785351 30584 785361
rect 29878 785335 30581 785351
rect 31686 782747 31924 782779
rect 31344 782727 31660 782745
rect 35934 782312 35961 782802
rect 31344 781527 31660 781539
rect 31344 781523 31924 781527
rect 31686 781489 31924 781523
rect 697975 780814 702721 780962
rect 696644 780023 696656 780079
rect 20672 779525 20684 779581
rect 14607 778642 19353 778790
rect 685404 778081 685642 778115
rect 685404 778077 685984 778081
rect 685668 778065 685984 778077
rect 681367 776802 681394 777292
rect 685668 776859 685984 776877
rect 685404 776825 685642 776857
rect 686747 774253 687450 774269
rect 686744 774243 687450 774253
rect 678511 772758 678519 772784
rect 678511 769549 678519 769574
rect 687438 768520 687450 774243
rect 687510 769509 687513 775062
rect 697918 773864 697949 780788
rect 714591 780674 714617 780708
rect 699187 780271 700187 780297
rect 700787 780271 701787 780297
rect 699187 780124 700187 780226
rect 700787 780124 701787 780226
rect 707475 779698 708475 779838
rect 709076 779699 710076 779861
rect 687623 772786 687629 773234
rect 696682 772655 696686 773860
rect 687623 769714 687629 770188
rect 711444 768315 711460 780496
rect 714591 779440 714617 779474
rect 712274 768315 712296 775426
rect 707475 767534 708475 767575
rect 709076 767534 710076 767575
rect 699187 766903 700187 767058
rect 700787 766903 701787 767058
rect 707475 766803 708475 767013
rect 709076 766803 710076 767013
rect 699187 766578 700187 766733
rect 700787 766578 701787 766733
rect 711444 766490 711470 768272
rect 711444 766480 711484 766490
rect 711444 766466 712328 766480
rect 5000 748524 5884 748538
rect 5844 748514 5884 748524
rect 5858 746732 5884 748514
rect 15541 748271 16541 748426
rect 17141 748271 18141 748426
rect 7252 747991 8252 748201
rect 8853 747991 9853 748201
rect 15541 747946 16541 748101
rect 17141 747946 18141 748101
rect 7252 747429 8252 747470
rect 8853 747429 9853 747470
rect 5032 739578 5054 746689
rect 2711 735530 2737 735564
rect 5868 734508 5884 746689
rect 29699 744816 29705 745290
rect 20642 741144 20646 742349
rect 29699 741770 29705 742218
rect 7252 735143 8252 735305
rect 8853 735166 9853 735306
rect 15541 734778 16541 734880
rect 17141 734778 18141 734880
rect 15541 734707 16541 734733
rect 17141 734707 18141 734733
rect 2711 734296 2737 734330
rect 19379 734216 19410 741140
rect 29815 739942 29818 745495
rect 29878 740761 29890 746484
rect 38809 745430 38817 745455
rect 38809 742220 38817 742246
rect 29878 740751 30584 740761
rect 29878 740735 30581 740751
rect 31686 738147 31924 738179
rect 31344 738127 31660 738145
rect 35934 737712 35961 738202
rect 31344 736927 31660 736939
rect 31344 736923 31924 736927
rect 31686 736889 31924 736923
rect 20672 734925 20684 734981
rect 697975 734414 702721 734562
rect 14607 734042 19353 734190
rect 696644 733623 696656 733679
rect 685404 731681 685642 731715
rect 685404 731677 685984 731681
rect 685668 731665 685984 731677
rect 681367 730402 681394 730892
rect 685668 730459 685984 730477
rect 685404 730425 685642 730457
rect 686747 727853 687450 727869
rect 686744 727843 687450 727853
rect 678511 726358 678519 726384
rect 678511 723149 678519 723174
rect 687438 722120 687450 727843
rect 687510 723109 687513 728662
rect 697918 727464 697949 734388
rect 714591 734274 714617 734308
rect 699187 733871 700187 733897
rect 700787 733871 701787 733897
rect 699187 733724 700187 733826
rect 700787 733724 701787 733826
rect 707475 733298 708475 733438
rect 709076 733299 710076 733461
rect 687623 726386 687629 726834
rect 696682 726255 696686 727460
rect 687623 723314 687629 723788
rect 711444 721915 711460 734096
rect 714591 733040 714617 733074
rect 712274 721915 712296 729026
rect 707475 721134 708475 721175
rect 709076 721134 710076 721175
rect 699187 720503 700187 720658
rect 700787 720503 701787 720658
rect 707475 720403 708475 720613
rect 709076 720403 710076 720613
rect 699187 720178 700187 720333
rect 700787 720178 701787 720333
rect 711444 720090 711470 721872
rect 711444 720080 711484 720090
rect 711444 720066 712328 720080
rect 5000 704124 5884 704138
rect 5844 704114 5884 704124
rect 5858 702332 5884 704114
rect 15541 703871 16541 704026
rect 17141 703871 18141 704026
rect 7252 703591 8252 703801
rect 8853 703591 9853 703801
rect 15541 703546 16541 703701
rect 17141 703546 18141 703701
rect 7252 703029 8252 703070
rect 8853 703029 9853 703070
rect 5032 695178 5054 702289
rect 2711 691130 2737 691164
rect 5868 690108 5884 702289
rect 29699 700416 29705 700890
rect 20642 696744 20646 697949
rect 29699 697370 29705 697818
rect 7252 690743 8252 690905
rect 8853 690766 9853 690906
rect 15541 690378 16541 690480
rect 17141 690378 18141 690480
rect 15541 690307 16541 690333
rect 17141 690307 18141 690333
rect 2711 689896 2737 689930
rect 19379 689816 19410 696740
rect 29815 695542 29818 701095
rect 29878 696361 29890 702084
rect 38809 701030 38817 701055
rect 38809 697820 38817 697846
rect 29878 696351 30584 696361
rect 29878 696335 30581 696351
rect 31686 693747 31924 693779
rect 31344 693727 31660 693745
rect 35934 693312 35961 693802
rect 31344 692527 31660 692539
rect 31344 692523 31924 692527
rect 31686 692489 31924 692523
rect 20672 690525 20684 690581
rect 14607 689642 19353 689790
rect 697975 687814 702721 687962
rect 696644 687023 696656 687079
rect 685404 685081 685642 685115
rect 685404 685077 685984 685081
rect 685668 685065 685984 685077
rect 681367 683802 681394 684292
rect 685668 683859 685984 683877
rect 685404 683825 685642 683857
rect 686747 681253 687450 681269
rect 686744 681243 687450 681253
rect 678511 679758 678519 679784
rect 678511 676549 678519 676574
rect 687438 675520 687450 681243
rect 687510 676509 687513 682062
rect 697918 680864 697949 687788
rect 714591 687674 714617 687708
rect 699187 687271 700187 687297
rect 700787 687271 701787 687297
rect 699187 687124 700187 687226
rect 700787 687124 701787 687226
rect 707475 686698 708475 686838
rect 709076 686699 710076 686861
rect 687623 679786 687629 680234
rect 696682 679655 696686 680860
rect 687623 676714 687629 677188
rect 711444 675315 711460 687496
rect 714591 686440 714617 686474
rect 712274 675315 712296 682426
rect 707475 674534 708475 674575
rect 709076 674534 710076 674575
rect 699187 673903 700187 674058
rect 700787 673903 701787 674058
rect 707475 673803 708475 674013
rect 709076 673803 710076 674013
rect 699187 673578 700187 673733
rect 700787 673578 701787 673733
rect 711444 673490 711470 675272
rect 711444 673480 711484 673490
rect 711444 673466 712328 673480
rect 5000 659524 5884 659538
rect 5844 659514 5884 659524
rect 5858 657732 5884 659514
rect 15541 659271 16541 659426
rect 17141 659271 18141 659426
rect 7252 658991 8252 659201
rect 8853 658991 9853 659201
rect 15541 658946 16541 659101
rect 17141 658946 18141 659101
rect 7252 658429 8252 658470
rect 8853 658429 9853 658470
rect 5032 650578 5054 657689
rect 2711 646530 2737 646564
rect 5868 645508 5884 657689
rect 29699 655816 29705 656290
rect 20642 652144 20646 653349
rect 29699 652770 29705 653218
rect 7252 646143 8252 646305
rect 8853 646166 9853 646306
rect 15541 645778 16541 645880
rect 17141 645778 18141 645880
rect 15541 645707 16541 645733
rect 17141 645707 18141 645733
rect 2711 645296 2737 645330
rect 19379 645216 19410 652140
rect 29815 650942 29818 656495
rect 29878 651761 29890 657484
rect 38809 656430 38817 656455
rect 38809 653220 38817 653246
rect 29878 651751 30584 651761
rect 29878 651735 30581 651751
rect 31686 649147 31924 649179
rect 31344 649127 31660 649145
rect 35934 648712 35961 649202
rect 31344 647927 31660 647939
rect 31344 647923 31924 647927
rect 31686 647889 31924 647923
rect 20672 645925 20684 645981
rect 14607 645042 19353 645190
rect 697975 641214 702721 641362
rect 696644 640423 696656 640479
rect 685404 638481 685642 638515
rect 685404 638477 685984 638481
rect 685668 638465 685984 638477
rect 681367 637202 681394 637692
rect 685668 637259 685984 637277
rect 685404 637225 685642 637257
rect 686747 634653 687450 634669
rect 686744 634643 687450 634653
rect 678511 633158 678519 633184
rect 678511 629949 678519 629974
rect 687438 628920 687450 634643
rect 687510 629909 687513 635462
rect 697918 634264 697949 641188
rect 714591 641074 714617 641108
rect 699187 640671 700187 640697
rect 700787 640671 701787 640697
rect 699187 640524 700187 640626
rect 700787 640524 701787 640626
rect 707475 640098 708475 640238
rect 709076 640099 710076 640261
rect 687623 633186 687629 633634
rect 696682 633055 696686 634260
rect 687623 630114 687629 630588
rect 711444 628715 711460 640896
rect 714591 639840 714617 639874
rect 712274 628715 712296 635826
rect 707475 627934 708475 627975
rect 709076 627934 710076 627975
rect 699187 627303 700187 627458
rect 700787 627303 701787 627458
rect 707475 627203 708475 627413
rect 709076 627203 710076 627413
rect 699187 626978 700187 627133
rect 700787 626978 701787 627133
rect 711444 626890 711470 628672
rect 711444 626880 711484 626890
rect 711444 626866 712328 626880
rect 5000 614924 5884 614938
rect 5844 614914 5884 614924
rect 5858 613132 5884 614914
rect 15541 614671 16541 614826
rect 17141 614671 18141 614826
rect 7252 614391 8252 614601
rect 8853 614391 9853 614601
rect 15541 614346 16541 614501
rect 17141 614346 18141 614501
rect 7252 613829 8252 613870
rect 8853 613829 9853 613870
rect 5032 605978 5054 613089
rect 2711 601930 2737 601964
rect 5868 600908 5884 613089
rect 29699 611216 29705 611690
rect 20642 607544 20646 608749
rect 29699 608170 29705 608618
rect 7252 601543 8252 601705
rect 8853 601566 9853 601706
rect 15541 601178 16541 601280
rect 17141 601178 18141 601280
rect 15541 601107 16541 601133
rect 17141 601107 18141 601133
rect 2711 600696 2737 600730
rect 19379 600616 19410 607540
rect 29815 606342 29818 611895
rect 29878 607161 29890 612884
rect 38809 611830 38817 611855
rect 38809 608620 38817 608646
rect 29878 607151 30584 607161
rect 29878 607135 30581 607151
rect 31686 604547 31924 604579
rect 31344 604527 31660 604545
rect 35934 604112 35961 604602
rect 31344 603327 31660 603339
rect 31344 603323 31924 603327
rect 31686 603289 31924 603323
rect 20672 601325 20684 601381
rect 14607 600442 19353 600590
rect 697975 594614 702721 594762
rect 696644 593823 696656 593879
rect 685404 591881 685642 591915
rect 685404 591877 685984 591881
rect 685668 591865 685984 591877
rect 681367 590602 681394 591092
rect 685668 590659 685984 590677
rect 685404 590625 685642 590657
rect 686747 588053 687450 588069
rect 686744 588043 687450 588053
rect 678511 586558 678519 586584
rect 678511 583349 678519 583374
rect 687438 582320 687450 588043
rect 687510 583309 687513 588862
rect 697918 587664 697949 594588
rect 714591 594474 714617 594508
rect 699187 594071 700187 594097
rect 700787 594071 701787 594097
rect 699187 593924 700187 594026
rect 700787 593924 701787 594026
rect 707475 593498 708475 593638
rect 709076 593499 710076 593661
rect 687623 586586 687629 587034
rect 696682 586455 696686 587660
rect 687623 583514 687629 583988
rect 711444 582115 711460 594296
rect 714591 593240 714617 593274
rect 712274 582115 712296 589226
rect 707475 581334 708475 581375
rect 709076 581334 710076 581375
rect 699187 580703 700187 580858
rect 700787 580703 701787 580858
rect 707475 580603 708475 580813
rect 709076 580603 710076 580813
rect 699187 580378 700187 580533
rect 700787 580378 701787 580533
rect 711444 580290 711470 582072
rect 711444 580280 711484 580290
rect 711444 580266 712328 580280
rect 5000 570524 5884 570538
rect 5844 570514 5884 570524
rect 5858 568732 5884 570514
rect 15541 570271 16541 570426
rect 17141 570271 18141 570426
rect 7252 569991 8252 570201
rect 8853 569991 9853 570201
rect 15541 569946 16541 570101
rect 17141 569946 18141 570101
rect 7252 569429 8252 569470
rect 8853 569429 9853 569470
rect 5032 561578 5054 568689
rect 2711 557530 2737 557564
rect 5868 556508 5884 568689
rect 29699 566816 29705 567290
rect 20642 563144 20646 564349
rect 29699 563770 29705 564218
rect 7252 557143 8252 557305
rect 8853 557166 9853 557306
rect 15541 556778 16541 556880
rect 17141 556778 18141 556880
rect 15541 556707 16541 556733
rect 17141 556707 18141 556733
rect 2711 556296 2737 556330
rect 19379 556216 19410 563140
rect 29815 561942 29818 567495
rect 29878 562761 29890 568484
rect 38809 567430 38817 567455
rect 38809 564220 38817 564246
rect 29878 562751 30584 562761
rect 29878 562735 30581 562751
rect 31686 560147 31924 560179
rect 31344 560127 31660 560145
rect 35934 559712 35961 560202
rect 31344 558927 31660 558939
rect 31344 558923 31924 558927
rect 31686 558889 31924 558923
rect 20672 556925 20684 556981
rect 14607 556042 19353 556190
rect 697975 548014 702721 548162
rect 696644 547223 696656 547279
rect 685404 545281 685642 545315
rect 685404 545277 685984 545281
rect 685668 545265 685984 545277
rect 681367 544002 681394 544492
rect 685668 544059 685984 544077
rect 685404 544025 685642 544057
rect 686747 541453 687450 541469
rect 686744 541443 687450 541453
rect 678511 539958 678519 539984
rect 678511 536749 678519 536774
rect 687438 535720 687450 541443
rect 687510 536709 687513 542262
rect 697918 541064 697949 547988
rect 714591 547874 714617 547908
rect 699187 547471 700187 547497
rect 700787 547471 701787 547497
rect 699187 547324 700187 547426
rect 700787 547324 701787 547426
rect 707475 546898 708475 547038
rect 709076 546899 710076 547061
rect 687623 539986 687629 540434
rect 696682 539855 696686 541060
rect 687623 536914 687629 537388
rect 711444 535515 711460 547696
rect 714591 546640 714617 546674
rect 712274 535515 712296 542626
rect 707475 534734 708475 534775
rect 709076 534734 710076 534775
rect 699187 534103 700187 534258
rect 700787 534103 701787 534258
rect 707475 534003 708475 534213
rect 709076 534003 710076 534213
rect 699187 533778 700187 533933
rect 700787 533778 701787 533933
rect 711444 533690 711470 535472
rect 711444 533680 711484 533690
rect 711444 533666 712328 533680
rect 5000 525924 5884 525938
rect 5844 525914 5884 525924
rect 5858 524132 5884 525914
rect 15541 525671 16541 525826
rect 17141 525671 18141 525826
rect 7252 525391 8252 525601
rect 8853 525391 9853 525601
rect 15541 525346 16541 525501
rect 17141 525346 18141 525501
rect 7252 524829 8252 524870
rect 8853 524829 9853 524870
rect 5032 516978 5054 524089
rect 2711 512930 2737 512964
rect 5868 511908 5884 524089
rect 29699 522216 29705 522690
rect 20642 518544 20646 519749
rect 29699 519170 29705 519618
rect 7252 512543 8252 512705
rect 8853 512566 9853 512706
rect 15541 512178 16541 512280
rect 17141 512178 18141 512280
rect 15541 512107 16541 512133
rect 17141 512107 18141 512133
rect 2711 511696 2737 511730
rect 19379 511616 19410 518540
rect 29815 517342 29818 522895
rect 29878 518161 29890 523884
rect 38809 522830 38817 522855
rect 38809 519620 38817 519646
rect 29878 518151 30584 518161
rect 29878 518135 30581 518151
rect 31686 515547 31924 515579
rect 31344 515527 31660 515545
rect 35934 515112 35961 515602
rect 31344 514327 31660 514339
rect 31344 514323 31924 514327
rect 31686 514289 31924 514323
rect 20672 512325 20684 512381
rect 14607 511442 19353 511590
rect 678146 453589 681534 453647
rect 678146 449673 681534 449687
rect 35794 430917 39182 430931
rect 35794 426957 39182 427015
rect 5000 394324 5884 394338
rect 5844 394314 5884 394324
rect 5858 392532 5884 394314
rect 15541 394071 16541 394226
rect 17141 394071 18141 394226
rect 7252 393791 8252 394001
rect 8853 393791 9853 394001
rect 15541 393746 16541 393901
rect 17141 393746 18141 393901
rect 7252 393229 8252 393270
rect 8853 393229 9853 393270
rect 5032 385378 5054 392489
rect 2711 381330 2737 381364
rect 5868 380308 5884 392489
rect 29699 390616 29705 391090
rect 20642 386944 20646 388149
rect 29699 387570 29705 388018
rect 7252 380943 8252 381105
rect 8853 380966 9853 381106
rect 15541 380578 16541 380680
rect 17141 380578 18141 380680
rect 15541 380507 16541 380533
rect 17141 380507 18141 380533
rect 2711 380096 2737 380130
rect 19379 380016 19410 386940
rect 29815 385742 29818 391295
rect 29878 386561 29890 392284
rect 38809 391230 38817 391255
rect 38809 388020 38817 388046
rect 29878 386551 30584 386561
rect 29878 386535 30581 386551
rect 31686 383947 31924 383979
rect 31344 383927 31660 383945
rect 35934 383512 35961 384002
rect 31344 382727 31660 382739
rect 31344 382723 31924 382727
rect 31686 382689 31924 382723
rect 20672 380725 20684 380781
rect 14607 379842 19353 379990
rect 697975 364814 702721 364962
rect 696644 364023 696656 364079
rect 685404 362081 685642 362115
rect 685404 362077 685984 362081
rect 685668 362065 685984 362077
rect 681367 360802 681394 361292
rect 685668 360859 685984 360877
rect 685404 360825 685642 360857
rect 686747 358253 687450 358269
rect 686744 358243 687450 358253
rect 678511 356758 678519 356784
rect 678511 353549 678519 353574
rect 687438 352520 687450 358243
rect 687510 353509 687513 359062
rect 697918 357864 697949 364788
rect 714591 364674 714617 364708
rect 699187 364271 700187 364297
rect 700787 364271 701787 364297
rect 699187 364124 700187 364226
rect 700787 364124 701787 364226
rect 707475 363698 708475 363838
rect 709076 363699 710076 363861
rect 687623 356786 687629 357234
rect 696682 356655 696686 357860
rect 687623 353714 687629 354188
rect 711444 352315 711460 364496
rect 714591 363440 714617 363474
rect 712274 352315 712296 359426
rect 707475 351534 708475 351575
rect 709076 351534 710076 351575
rect 699187 350903 700187 351058
rect 700787 350903 701787 351058
rect 707475 350803 708475 351013
rect 709076 350803 710076 351013
rect 699187 350578 700187 350733
rect 700787 350578 701787 350733
rect 711444 350490 711470 352272
rect 711444 350480 711484 350490
rect 711444 350466 712328 350480
rect 5000 349724 5884 349738
rect 5844 349714 5884 349724
rect 5858 347932 5884 349714
rect 15541 349471 16541 349626
rect 17141 349471 18141 349626
rect 7252 349191 8252 349401
rect 8853 349191 9853 349401
rect 15541 349146 16541 349301
rect 17141 349146 18141 349301
rect 7252 348629 8252 348670
rect 8853 348629 9853 348670
rect 5032 340778 5054 347889
rect 2711 336730 2737 336764
rect 5868 335708 5884 347889
rect 29699 346016 29705 346490
rect 20642 342344 20646 343549
rect 29699 342970 29705 343418
rect 7252 336343 8252 336505
rect 8853 336366 9853 336506
rect 15541 335978 16541 336080
rect 17141 335978 18141 336080
rect 15541 335907 16541 335933
rect 17141 335907 18141 335933
rect 2711 335496 2737 335530
rect 19379 335416 19410 342340
rect 29815 341142 29818 346695
rect 29878 341961 29890 347684
rect 38809 346630 38817 346655
rect 38809 343420 38817 343446
rect 29878 341951 30584 341961
rect 29878 341935 30581 341951
rect 31686 339347 31924 339379
rect 31344 339327 31660 339345
rect 35934 338912 35961 339402
rect 31344 338127 31660 338139
rect 31344 338123 31924 338127
rect 31686 338089 31924 338123
rect 20672 336125 20684 336181
rect 14607 335242 19353 335390
rect 697975 318214 702721 318362
rect 696644 317423 696656 317479
rect 685404 315481 685642 315515
rect 685404 315477 685984 315481
rect 685668 315465 685984 315477
rect 681367 314202 681394 314692
rect 685668 314259 685984 314277
rect 685404 314225 685642 314257
rect 686747 311653 687450 311669
rect 686744 311643 687450 311653
rect 678511 310158 678519 310184
rect 678511 306949 678519 306974
rect 687438 305920 687450 311643
rect 687510 306909 687513 312462
rect 697918 311264 697949 318188
rect 714591 318074 714617 318108
rect 699187 317671 700187 317697
rect 700787 317671 701787 317697
rect 699187 317524 700187 317626
rect 700787 317524 701787 317626
rect 707475 317098 708475 317238
rect 709076 317099 710076 317261
rect 687623 310186 687629 310634
rect 696682 310055 696686 311260
rect 687623 307114 687629 307588
rect 711444 305715 711460 317896
rect 714591 316840 714617 316874
rect 712274 305715 712296 312826
rect 5000 305324 5884 305338
rect 5844 305314 5884 305324
rect 5858 303532 5884 305314
rect 15541 305071 16541 305226
rect 17141 305071 18141 305226
rect 7252 304791 8252 305001
rect 8853 304791 9853 305001
rect 707475 304934 708475 304975
rect 709076 304934 710076 304975
rect 15541 304746 16541 304901
rect 17141 304746 18141 304901
rect 699187 304303 700187 304458
rect 700787 304303 701787 304458
rect 7252 304229 8252 304270
rect 8853 304229 9853 304270
rect 707475 304203 708475 304413
rect 709076 304203 710076 304413
rect 699187 303978 700187 304133
rect 700787 303978 701787 304133
rect 711444 303890 711470 305672
rect 711444 303880 711484 303890
rect 711444 303866 712328 303880
rect 5032 296378 5054 303489
rect 2711 292330 2737 292364
rect 5868 291308 5884 303489
rect 29699 301616 29705 302090
rect 20642 297944 20646 299149
rect 29699 298570 29705 299018
rect 7252 291943 8252 292105
rect 8853 291966 9853 292106
rect 15541 291578 16541 291680
rect 17141 291578 18141 291680
rect 15541 291507 16541 291533
rect 17141 291507 18141 291533
rect 2711 291096 2737 291130
rect 19379 291016 19410 297940
rect 29815 296742 29818 302295
rect 29878 297561 29890 303284
rect 38809 302230 38817 302255
rect 38809 299020 38817 299046
rect 29878 297551 30584 297561
rect 29878 297535 30581 297551
rect 31686 294947 31924 294979
rect 31344 294927 31660 294945
rect 35934 294512 35961 295002
rect 31344 293727 31660 293739
rect 31344 293723 31924 293727
rect 31686 293689 31924 293723
rect 20672 291725 20684 291781
rect 14607 290842 19353 290990
rect 697975 271814 702721 271962
rect 696644 271023 696656 271079
rect 685404 269081 685642 269115
rect 685404 269077 685984 269081
rect 685668 269065 685984 269077
rect 681367 267802 681394 268292
rect 685668 267859 685984 267877
rect 685404 267825 685642 267857
rect 686747 265253 687450 265269
rect 686744 265243 687450 265253
rect 678511 263758 678519 263784
rect 5000 260724 5884 260738
rect 5844 260714 5884 260724
rect 5858 258932 5884 260714
rect 15541 260471 16541 260626
rect 17141 260471 18141 260626
rect 678511 260549 678519 260574
rect 7252 260191 8252 260401
rect 8853 260191 9853 260401
rect 15541 260146 16541 260301
rect 17141 260146 18141 260301
rect 7252 259629 8252 259670
rect 8853 259629 9853 259670
rect 687438 259520 687450 265243
rect 687510 260509 687513 266062
rect 697918 264864 697949 271788
rect 714591 271674 714617 271708
rect 699187 271271 700187 271297
rect 700787 271271 701787 271297
rect 699187 271124 700187 271226
rect 700787 271124 701787 271226
rect 707475 270698 708475 270838
rect 709076 270699 710076 270861
rect 687623 263786 687629 264234
rect 696682 263655 696686 264860
rect 687623 260714 687629 261188
rect 711444 259315 711460 271496
rect 714591 270440 714617 270474
rect 712274 259315 712296 266426
rect 5032 251778 5054 258889
rect 2711 247730 2737 247764
rect 5868 246708 5884 258889
rect 29699 257016 29705 257490
rect 20642 253344 20646 254549
rect 29699 253970 29705 254418
rect 7252 247343 8252 247505
rect 8853 247366 9853 247506
rect 15541 246978 16541 247080
rect 17141 246978 18141 247080
rect 15541 246907 16541 246933
rect 17141 246907 18141 246933
rect 2711 246496 2737 246530
rect 19379 246416 19410 253340
rect 29815 252142 29818 257695
rect 29878 252961 29890 258684
rect 707475 258534 708475 258575
rect 709076 258534 710076 258575
rect 699187 257903 700187 258058
rect 700787 257903 701787 258058
rect 707475 257803 708475 258013
rect 709076 257803 710076 258013
rect 38809 257630 38817 257655
rect 699187 257578 700187 257733
rect 700787 257578 701787 257733
rect 711444 257490 711470 259272
rect 711444 257480 711484 257490
rect 711444 257466 712328 257480
rect 38809 254420 38817 254446
rect 29878 252951 30584 252961
rect 29878 252935 30581 252951
rect 31686 250347 31924 250379
rect 31344 250327 31660 250345
rect 35934 249912 35961 250402
rect 31344 249127 31660 249139
rect 31344 249123 31924 249127
rect 31686 249089 31924 249123
rect 20672 247125 20684 247181
rect 14607 246242 19353 246390
rect 697975 225214 702721 225362
rect 696644 224423 696656 224479
rect 685404 222481 685642 222515
rect 685404 222477 685984 222481
rect 685668 222465 685984 222477
rect 681367 221202 681394 221692
rect 685668 221259 685984 221277
rect 685404 221225 685642 221257
rect 686747 218653 687450 218669
rect 686744 218643 687450 218653
rect 678511 217158 678519 217184
rect 5000 216124 5884 216138
rect 5844 216114 5884 216124
rect 5858 214332 5884 216114
rect 15541 215871 16541 216026
rect 17141 215871 18141 216026
rect 7252 215591 8252 215801
rect 8853 215591 9853 215801
rect 15541 215546 16541 215701
rect 17141 215546 18141 215701
rect 7252 215029 8252 215070
rect 8853 215029 9853 215070
rect 5032 207178 5054 214289
rect 2711 203130 2737 203164
rect 5868 202108 5884 214289
rect 29699 212416 29705 212890
rect 20642 208744 20646 209949
rect 29699 209370 29705 209818
rect 7252 202743 8252 202905
rect 8853 202766 9853 202906
rect 15541 202378 16541 202480
rect 17141 202378 18141 202480
rect 15541 202307 16541 202333
rect 17141 202307 18141 202333
rect 2711 201896 2737 201930
rect 19379 201816 19410 208740
rect 29815 207542 29818 213095
rect 29878 208361 29890 214084
rect 678511 213949 678519 213974
rect 38809 213030 38817 213055
rect 687438 212920 687450 218643
rect 687510 213909 687513 219462
rect 697918 218264 697949 225188
rect 714591 225074 714617 225108
rect 699187 224671 700187 224697
rect 700787 224671 701787 224697
rect 699187 224524 700187 224626
rect 700787 224524 701787 224626
rect 707475 224098 708475 224238
rect 709076 224099 710076 224261
rect 687623 217186 687629 217634
rect 696682 217055 696686 218260
rect 687623 214114 687629 214588
rect 711444 212715 711460 224896
rect 714591 223840 714617 223874
rect 712274 212715 712296 219826
rect 707475 211934 708475 211975
rect 709076 211934 710076 211975
rect 699187 211303 700187 211458
rect 700787 211303 701787 211458
rect 707475 211203 708475 211413
rect 709076 211203 710076 211413
rect 699187 210978 700187 211133
rect 700787 210978 701787 211133
rect 711444 210890 711470 212672
rect 711444 210880 711484 210890
rect 711444 210866 712328 210880
rect 38809 209820 38817 209846
rect 29878 208351 30584 208361
rect 29878 208335 30581 208351
rect 31686 205747 31924 205779
rect 31344 205727 31660 205745
rect 35934 205312 35961 205802
rect 31344 204527 31660 204539
rect 31344 204523 31924 204527
rect 31686 204489 31924 204523
rect 20672 202525 20684 202581
rect 14607 201642 19353 201790
rect 697975 178614 702721 178762
rect 696644 177823 696656 177879
rect 685404 175881 685642 175915
rect 685404 175877 685984 175881
rect 685668 175865 685984 175877
rect 681367 174602 681394 175092
rect 685668 174659 685984 174677
rect 685404 174625 685642 174657
rect 686747 172053 687450 172069
rect 686744 172043 687450 172053
rect 5000 171724 5884 171738
rect 5844 171714 5884 171724
rect 5858 169932 5884 171714
rect 15541 171471 16541 171626
rect 17141 171471 18141 171626
rect 7252 171191 8252 171401
rect 8853 171191 9853 171401
rect 15541 171146 16541 171301
rect 17141 171146 18141 171301
rect 7252 170629 8252 170670
rect 8853 170629 9853 170670
rect 678511 170558 678519 170584
rect 5032 162778 5054 169889
rect 2711 158730 2737 158764
rect 5868 157708 5884 169889
rect 29699 168016 29705 168490
rect 20642 164344 20646 165549
rect 29699 164970 29705 165418
rect 7252 158343 8252 158505
rect 8853 158366 9853 158506
rect 15541 157978 16541 158080
rect 17141 157978 18141 158080
rect 15541 157907 16541 157933
rect 17141 157907 18141 157933
rect 2711 157496 2737 157530
rect 19379 157416 19410 164340
rect 29815 163142 29818 168695
rect 29878 163961 29890 169684
rect 38809 168630 38817 168655
rect 678511 167349 678519 167374
rect 687438 166320 687450 172043
rect 687510 167309 687513 172862
rect 697918 171664 697949 178588
rect 714591 178474 714617 178508
rect 699187 178071 700187 178097
rect 700787 178071 701787 178097
rect 699187 177924 700187 178026
rect 700787 177924 701787 178026
rect 707475 177498 708475 177638
rect 709076 177499 710076 177661
rect 687623 170586 687629 171034
rect 696682 170455 696686 171660
rect 687623 167514 687629 167988
rect 711444 166115 711460 178296
rect 714591 177240 714617 177274
rect 712274 166115 712296 173226
rect 38809 165420 38817 165446
rect 707475 165334 708475 165375
rect 709076 165334 710076 165375
rect 699187 164703 700187 164858
rect 700787 164703 701787 164858
rect 707475 164603 708475 164813
rect 709076 164603 710076 164813
rect 699187 164378 700187 164533
rect 700787 164378 701787 164533
rect 711444 164290 711470 166072
rect 711444 164280 711484 164290
rect 711444 164266 712328 164280
rect 29878 163951 30584 163961
rect 29878 163935 30581 163951
rect 31686 161347 31924 161379
rect 31344 161327 31660 161345
rect 35934 160912 35961 161402
rect 31344 160127 31660 160139
rect 31344 160123 31924 160127
rect 31686 160089 31924 160123
rect 20672 158125 20684 158181
rect 14607 157242 19353 157390
rect 697975 132014 702721 132162
rect 696644 131223 696656 131279
rect 685404 129281 685642 129315
rect 685404 129277 685984 129281
rect 685668 129265 685984 129277
rect 681367 128002 681394 128492
rect 685668 128059 685984 128077
rect 685404 128025 685642 128057
rect 686747 125453 687450 125469
rect 686744 125443 687450 125453
rect 678511 123958 678519 123984
rect 678511 120749 678519 120774
rect 687438 119720 687450 125443
rect 687510 120709 687513 126262
rect 697918 125064 697949 131988
rect 714591 131874 714617 131908
rect 699187 131471 700187 131497
rect 700787 131471 701787 131497
rect 699187 131324 700187 131426
rect 700787 131324 701787 131426
rect 707475 130898 708475 131038
rect 709076 130899 710076 131061
rect 687623 123986 687629 124434
rect 696682 123855 696686 125060
rect 687623 120914 687629 121388
rect 711444 119515 711460 131696
rect 714591 130640 714617 130674
rect 712274 119515 712296 126626
rect 707475 118734 708475 118775
rect 709076 118734 710076 118775
rect 699187 118103 700187 118258
rect 700787 118103 701787 118258
rect 707475 118003 708475 118213
rect 709076 118003 710076 118213
rect 699187 117778 700187 117933
rect 700787 117778 701787 117933
rect 711444 117690 711470 119472
rect 711444 117680 711484 117690
rect 711444 117666 712328 117680
rect 697975 85414 702721 85562
rect 696644 84623 696656 84679
rect 685404 82681 685642 82715
rect 685404 82677 685984 82681
rect 685668 82665 685984 82677
rect 681367 81402 681394 81892
rect 685668 81459 685984 81477
rect 685404 81425 685642 81457
rect 686747 78853 687450 78869
rect 686744 78843 687450 78853
rect 678511 77358 678519 77384
rect 35794 76517 39182 76531
rect 678511 74149 678519 74174
rect 687438 73120 687450 78843
rect 687510 74109 687513 79662
rect 697918 78464 697949 85388
rect 714591 85274 714617 85308
rect 699187 84871 700187 84897
rect 700787 84871 701787 84897
rect 699187 84724 700187 84826
rect 700787 84724 701787 84826
rect 707475 84298 708475 84438
rect 709076 84299 710076 84461
rect 687623 77386 687629 77834
rect 696682 77255 696686 78460
rect 687623 74314 687629 74788
rect 711444 72915 711460 85096
rect 714591 84040 714617 84074
rect 712274 72915 712296 80026
rect 35794 72557 39182 72615
rect 707475 72134 708475 72175
rect 709076 72134 710076 72175
rect 699187 71503 700187 71658
rect 700787 71503 701787 71658
rect 707475 71403 708475 71613
rect 709076 71403 710076 71613
rect 699187 71178 700187 71333
rect 700787 71178 701787 71333
rect 711444 71090 711470 72872
rect 711444 71080 711484 71090
rect 711444 71066 712328 71080
rect 190011 38947 190036 38955
rect 193220 38947 193246 38955
rect 146051 38282 146317 38293
rect 144582 36868 144602 37392
rect 197264 36072 197754 36099
rect 248735 35932 248749 39320
rect 252651 35932 252709 39320
rect 298611 38947 298636 38955
rect 301820 38947 301846 38955
rect 353411 38947 353436 38955
rect 356620 38947 356646 38955
rect 408211 38947 408236 38955
rect 411420 38947 411446 38955
rect 463011 38947 463036 38955
rect 466220 38947 466246 38955
rect 517811 38947 517836 38955
rect 521020 38947 521046 38955
rect 305864 36072 306354 36099
rect 360664 36072 361154 36099
rect 415464 36072 415954 36099
rect 470264 36072 470754 36099
rect 525064 36072 525554 36099
rect 143271 35904 143327 35925
rect 143271 35795 143293 35904
rect 197287 31824 197319 32062
rect 198539 31824 198577 32062
rect 305887 31824 305919 32062
rect 307139 31824 307177 32062
rect 360687 31824 360719 32062
rect 361939 31824 361977 32062
rect 415487 31824 415519 32062
rect 416739 31824 416777 32062
rect 470287 31824 470319 32062
rect 471539 31824 471577 32062
rect 525087 31824 525119 32062
rect 526339 31824 526377 32062
rect 198539 31798 198543 31824
rect 307139 31798 307143 31824
rect 361939 31798 361943 31824
rect 416739 31798 416743 31824
rect 471539 31798 471543 31824
rect 526339 31798 526343 31824
rect 197321 31482 197339 31798
rect 198527 31482 198543 31798
rect 305921 31482 305939 31798
rect 307127 31482 307143 31798
rect 360721 31482 360739 31798
rect 361927 31482 361943 31798
rect 415521 31482 415539 31798
rect 416727 31482 416743 31798
rect 470321 31482 470339 31798
rect 471527 31482 471543 31798
rect 525121 31482 525139 31798
rect 526327 31482 526343 31798
rect 194705 30719 194715 30722
rect 303305 30719 303315 30722
rect 358105 30719 358115 30722
rect 412905 30719 412915 30722
rect 467705 30719 467715 30722
rect 522505 30719 522515 30722
rect 194705 30028 194731 30719
rect 303305 30028 303331 30719
rect 358105 30028 358131 30719
rect 412905 30028 412931 30719
rect 467705 30028 467731 30719
rect 522505 30028 522531 30719
rect 188982 30016 194731 30028
rect 297582 30016 303331 30028
rect 352382 30016 358131 30028
rect 407182 30016 412931 30028
rect 461982 30016 467731 30028
rect 516782 30016 522531 30028
rect 189971 29953 195524 29956
rect 298571 29953 304124 29956
rect 353371 29953 358924 29956
rect 408171 29953 413724 29956
rect 462971 29953 468524 29956
rect 517771 29953 523324 29956
rect 190176 29837 190650 29843
rect 193248 29837 193696 29843
rect 298776 29837 299250 29843
rect 301848 29837 302296 29843
rect 353576 29837 354050 29843
rect 356648 29837 357096 29843
rect 408376 29837 408850 29843
rect 411448 29837 411896 29843
rect 463176 29837 463650 29843
rect 466248 29837 466696 29843
rect 517976 29837 518450 29843
rect 521048 29837 521496 29843
rect 200485 20810 200541 20822
rect 309085 20810 309141 20822
rect 363885 20810 363941 20822
rect 418685 20810 418741 20822
rect 473485 20810 473541 20822
rect 528285 20810 528341 20822
rect 193117 20780 194322 20784
rect 301717 20780 302922 20784
rect 356517 20780 357722 20784
rect 411317 20780 412522 20784
rect 466117 20780 467322 20784
rect 520917 20780 522122 20784
rect 147373 19549 147437 19620
rect 194326 19517 201250 19548
rect 302926 19517 309850 19548
rect 357726 19517 364650 19548
rect 412526 19517 419450 19548
rect 467326 19517 474250 19548
rect 522126 19517 529050 19548
rect 133105 17480 133260 18480
rect 133430 17480 133585 18480
rect 146651 17480 146753 18480
rect 146798 17480 146824 18480
rect 187040 17279 187195 18279
rect 187365 17279 187520 18279
rect 200586 17279 200688 18279
rect 200733 17279 200759 18279
rect 133105 15880 133260 16880
rect 133430 15880 133585 16880
rect 146651 15880 146753 16880
rect 146798 15880 146824 16880
rect 187040 15679 187195 16679
rect 187365 15679 187520 16679
rect 200586 15679 200688 16679
rect 200733 15679 200759 16679
rect 201276 14745 201424 19491
rect 295640 17279 295795 18279
rect 295965 17279 296120 18279
rect 309186 17279 309288 18279
rect 309333 17279 309359 18279
rect 295640 15679 295795 16679
rect 295965 15679 296120 16679
rect 309186 15679 309288 16679
rect 309333 15679 309359 16679
rect 309876 14745 310024 19491
rect 350440 17279 350595 18279
rect 350765 17279 350920 18279
rect 363986 17279 364088 18279
rect 364133 17279 364159 18279
rect 350440 15679 350595 16679
rect 350765 15679 350920 16679
rect 363986 15679 364088 16679
rect 364133 15679 364159 16679
rect 364676 14745 364824 19491
rect 405240 17279 405395 18279
rect 405565 17279 405720 18279
rect 418786 17279 418888 18279
rect 418933 17279 418959 18279
rect 405240 15679 405395 16679
rect 405565 15679 405720 16679
rect 418786 15679 418888 16679
rect 418933 15679 418959 16679
rect 419476 14745 419624 19491
rect 460040 17279 460195 18279
rect 460365 17279 460520 18279
rect 473586 17279 473688 18279
rect 473733 17279 473759 18279
rect 460040 15679 460195 16679
rect 460365 15679 460520 16679
rect 473586 15679 473688 16679
rect 473733 15679 473759 16679
rect 474276 14745 474424 19491
rect 514840 17279 514995 18279
rect 515165 17279 515320 18279
rect 528386 17279 528488 18279
rect 528533 17279 528559 18279
rect 514840 15679 514995 16679
rect 515165 15679 515320 16679
rect 528386 15679 528488 16679
rect 528533 15679 528559 16679
rect 529076 14745 529224 19491
rect 133470 8992 133680 9992
rect 134201 8992 134242 9992
rect 146365 8992 146505 9992
rect 187265 8991 187475 9991
rect 187996 8991 188037 9991
rect 200160 8991 200300 9991
rect 295865 8991 296075 9991
rect 296596 8991 296637 9991
rect 308760 8991 308900 9991
rect 350665 8991 350875 9991
rect 351396 8991 351437 9991
rect 363560 8991 363700 9991
rect 405465 8991 405675 9991
rect 406196 8991 406237 9991
rect 418360 8991 418500 9991
rect 460265 8991 460475 9991
rect 460996 8991 461037 9991
rect 473160 8991 473300 9991
rect 515065 8991 515275 9991
rect 515796 8991 515837 9991
rect 527960 8991 528100 9991
rect 133470 7391 133680 8391
rect 134201 7391 134242 8391
rect 146366 7391 146528 8391
rect 187265 7390 187475 8390
rect 187996 7390 188037 8390
rect 200161 7390 200323 8390
rect 295865 7390 296075 8390
rect 296596 7390 296637 8390
rect 308761 7390 308923 8390
rect 350665 7390 350875 8390
rect 351396 7390 351437 8390
rect 363561 7390 363723 8390
rect 405465 7390 405675 8390
rect 406196 7390 406237 8390
rect 418361 7390 418523 8390
rect 460265 7390 460475 8390
rect 460996 7390 461037 8390
rect 473161 7390 473323 8390
rect 515065 7390 515275 8390
rect 515796 7390 515837 8390
rect 527961 7390 528123 8390
rect 186928 5996 188734 6022
rect 188777 6006 200958 6022
rect 295528 5996 297334 6022
rect 297377 6006 309558 6022
rect 350328 5996 352134 6022
rect 352177 6006 364358 6022
rect 405128 5996 406934 6022
rect 406977 6006 419158 6022
rect 459928 5996 461734 6022
rect 461777 6006 473958 6022
rect 514728 5996 516534 6022
rect 516577 6006 528758 6022
rect 186928 5982 186952 5996
rect 295528 5982 295552 5996
rect 350328 5982 350352 5996
rect 405128 5982 405152 5996
rect 459928 5982 459952 5996
rect 514728 5982 514752 5996
rect 186928 5138 186942 5982
rect 188777 5170 195888 5192
rect 295528 5138 295542 5982
rect 297377 5170 304488 5192
rect 350328 5138 350342 5982
rect 352177 5170 359288 5192
rect 405128 5138 405142 5982
rect 406977 5170 414088 5192
rect 459928 5138 459942 5982
rect 461777 5170 468888 5192
rect 514728 5138 514742 5982
rect 516577 5170 523688 5192
rect 199902 2849 199936 2875
rect 201136 2849 201170 2875
rect 308502 2849 308536 2875
rect 309736 2849 309770 2875
rect 363302 2849 363336 2875
rect 364536 2849 364570 2875
rect 418102 2849 418136 2875
rect 419336 2849 419370 2875
rect 472902 2849 472936 2875
rect 474136 2849 474170 2875
rect 527702 2849 527736 2875
rect 528936 2849 528970 2875
<< metal1 >>
rect 311390 995462 311396 995514
rect 311448 995502 311454 995514
rect 312770 995502 312776 995514
rect 311448 995474 312776 995502
rect 311448 995462 311454 995474
rect 312770 995462 312776 995474
rect 312828 995462 312834 995514
rect 466962 995462 466968 995514
rect 467020 995502 467026 995514
rect 473770 995502 473776 995514
rect 467020 995474 473776 995502
rect 467020 995462 467026 995474
rect 473770 995462 473776 995474
rect 473828 995462 473834 995514
rect 467698 995258 467704 995310
rect 467756 995298 467762 995310
rect 475610 995298 475616 995310
rect 467756 995270 475616 995298
rect 467756 995258 467762 995270
rect 475610 995258 475616 995270
rect 475668 995258 475674 995310
rect 250394 994170 250400 994222
rect 250452 994210 250458 994222
rect 256650 994210 256656 994222
rect 250452 994182 256656 994210
rect 250452 994170 250458 994182
rect 256650 994170 256656 994182
rect 256708 994210 256714 994222
rect 259042 994210 259048 994222
rect 256708 994182 259048 994210
rect 256708 994170 256714 994182
rect 259042 994170 259048 994182
rect 259100 994170 259106 994222
rect 82402 993558 82408 993610
rect 82460 993598 82466 993610
rect 136958 993598 136964 993610
rect 82460 993570 136964 993598
rect 82460 993558 82466 993570
rect 136958 993558 136964 993570
rect 137016 993598 137022 993610
rect 191606 993598 191612 993610
rect 137016 993570 191612 993598
rect 137016 993558 137022 993570
rect 191606 993558 191612 993570
rect 191664 993558 191670 993610
rect 195930 993558 195936 993610
rect 195988 993598 195994 993610
rect 203934 993598 203940 993610
rect 195988 993570 203940 993598
rect 195988 993558 195994 993570
rect 203934 993558 203940 993570
rect 203992 993558 203998 993610
rect 250394 993598 250400 993610
rect 204044 993570 250400 993598
rect 86726 993490 86732 993542
rect 86784 993530 86790 993542
rect 94730 993530 94736 993542
rect 86784 993502 94736 993530
rect 86784 993490 86790 993502
rect 94730 993490 94736 993502
rect 94788 993490 94794 993542
rect 100066 993490 100072 993542
rect 100124 993530 100130 993542
rect 102918 993530 102924 993542
rect 100124 993502 102924 993530
rect 100124 993490 100130 993502
rect 102918 993490 102924 993502
rect 102976 993490 102982 993542
rect 136314 993530 136320 993542
rect 132284 993502 136320 993530
rect 81758 993422 81764 993474
rect 81816 993462 81822 993474
rect 93718 993462 93724 993474
rect 81816 993434 93724 993462
rect 81816 993422 81822 993434
rect 93718 993422 93724 993434
rect 93776 993422 93782 993474
rect 115706 993422 115712 993474
rect 115764 993462 115770 993474
rect 132284 993462 132312 993502
rect 136314 993490 136320 993502
rect 136372 993490 136378 993542
rect 202094 993490 202100 993542
rect 202152 993530 202158 993542
rect 204044 993530 204072 993570
rect 250394 993558 250400 993570
rect 250452 993558 250458 993610
rect 250486 993558 250492 993610
rect 250544 993598 250550 993610
rect 258490 993598 258496 993610
rect 250544 993570 258496 993598
rect 250544 993558 250550 993570
rect 258490 993558 258496 993570
rect 258548 993558 258554 993610
rect 259042 993558 259048 993610
rect 259100 993598 259106 993610
rect 312770 993598 312776 993610
rect 259100 993570 312776 993598
rect 259100 993558 259106 993570
rect 312770 993558 312776 993570
rect 312828 993558 312834 993610
rect 437798 993558 437804 993610
rect 437856 993598 437862 993610
rect 450586 993598 450592 993610
rect 437856 993570 450592 993598
rect 437856 993558 437862 993570
rect 450586 993558 450592 993570
rect 450644 993558 450650 993610
rect 517286 993558 517292 993610
rect 517344 993598 517350 993610
rect 518022 993598 518028 993610
rect 517344 993570 518028 993598
rect 517344 993558 517350 993570
rect 518022 993558 518028 993570
rect 518080 993598 518086 993610
rect 625754 993598 625760 993610
rect 518080 993570 625760 993598
rect 518080 993558 518086 993570
rect 625754 993558 625760 993570
rect 625812 993598 625818 993610
rect 626214 993598 626220 993610
rect 625812 993570 626220 993598
rect 625812 993558 625818 993570
rect 626214 993558 626220 993570
rect 626272 993558 626278 993610
rect 630538 993558 630544 993610
rect 630596 993598 630602 993610
rect 638542 993598 638548 993610
rect 630596 993570 638548 993598
rect 630596 993558 630602 993570
rect 638542 993558 638548 993570
rect 638600 993558 638606 993610
rect 202152 993502 204072 993530
rect 202152 993490 202158 993502
rect 222610 993490 222616 993542
rect 222668 993530 222674 993542
rect 222668 993502 232960 993530
rect 222668 993490 222674 993502
rect 115764 993434 119432 993462
rect 115764 993422 115770 993434
rect 119404 993394 119432 993434
rect 119496 993434 132312 993462
rect 119496 993394 119524 993434
rect 141282 993422 141288 993474
rect 141340 993462 141346 993474
rect 149286 993462 149292 993474
rect 141340 993434 149292 993462
rect 141340 993422 141346 993434
rect 149286 993422 149292 993434
rect 149344 993422 149350 993474
rect 157934 993462 157940 993474
rect 151604 993434 157940 993462
rect 119404 993366 119524 993394
rect 136314 993354 136320 993406
rect 136372 993394 136378 993406
rect 151604 993394 151632 993434
rect 157934 993422 157940 993434
rect 157992 993422 157998 993474
rect 158118 993422 158124 993474
rect 158176 993462 158182 993474
rect 170906 993462 170912 993474
rect 158176 993434 170912 993462
rect 158176 993422 158182 993434
rect 170906 993422 170912 993434
rect 170964 993422 170970 993474
rect 170998 993422 171004 993474
rect 171056 993462 171062 993474
rect 178358 993462 178364 993474
rect 171056 993434 178364 993462
rect 171056 993422 171062 993434
rect 178358 993422 178364 993434
rect 178416 993422 178422 993474
rect 209822 993422 209828 993474
rect 209880 993462 209886 993474
rect 209880 993434 218792 993462
rect 209880 993422 209886 993434
rect 136372 993366 151632 993394
rect 218764 993394 218792 993434
rect 222426 993394 222432 993406
rect 218764 993366 222432 993394
rect 136372 993354 136378 993366
rect 222426 993354 222432 993366
rect 222484 993354 222490 993406
rect 232932 993394 232960 993502
rect 248370 993490 248376 993542
rect 248428 993530 248434 993542
rect 261158 993530 261164 993542
rect 248428 993502 261164 993530
rect 248428 993490 248434 993502
rect 261158 993490 261164 993502
rect 261216 993490 261222 993542
rect 273964 993502 274084 993530
rect 273964 993474 273992 993502
rect 274056 993474 274084 993502
rect 312586 993490 312592 993542
rect 312644 993530 312650 993542
rect 408082 993530 408088 993542
rect 312644 993502 408088 993530
rect 312644 993490 312650 993502
rect 408082 993490 408088 993502
rect 408140 993530 408146 993542
rect 462730 993530 462736 993542
rect 408140 993502 462736 993530
rect 408140 993490 408146 993502
rect 462730 993490 462736 993502
rect 462788 993530 462794 993542
rect 462788 993502 517424 993530
rect 462788 993490 462794 993502
rect 517396 993474 517424 993502
rect 528510 993490 528516 993542
rect 528568 993530 528574 993542
rect 636702 993530 636708 993542
rect 528568 993502 636708 993530
rect 528568 993490 528574 993502
rect 636702 993490 636708 993502
rect 636760 993490 636766 993542
rect 273946 993422 273952 993474
rect 274004 993422 274010 993474
rect 274038 993422 274044 993474
rect 274096 993422 274102 993474
rect 287010 993422 287016 993474
rect 287068 993462 287074 993474
rect 287068 993434 299752 993462
rect 287068 993422 287074 993434
rect 245518 993394 245524 993406
rect 232932 993366 245524 993394
rect 245518 993354 245524 993366
rect 245576 993394 245582 993406
rect 248278 993394 248284 993406
rect 245576 993366 248284 993394
rect 245576 993354 245582 993366
rect 248278 993354 248284 993366
rect 248336 993354 248342 993406
rect 92706 993286 92712 993338
rect 92764 993326 92770 993338
rect 92890 993326 92896 993338
rect 92764 993298 92896 993326
rect 92764 993286 92770 993298
rect 92890 993286 92896 993298
rect 92948 993326 92954 993338
rect 147446 993326 147452 993338
rect 92948 993298 147452 993326
rect 92948 993286 92954 993298
rect 147446 993286 147452 993298
rect 147504 993326 147510 993338
rect 202094 993326 202100 993338
rect 147504 993298 150252 993326
rect 147504 993286 147510 993298
rect 93718 993218 93724 993270
rect 93776 993258 93782 993270
rect 100066 993258 100072 993270
rect 93776 993230 100072 993258
rect 93776 993218 93782 993230
rect 100066 993218 100072 993230
rect 100124 993218 100130 993270
rect 150224 993258 150252 993298
rect 151696 993298 202100 993326
rect 151696 993258 151724 993298
rect 202094 993286 202100 993298
rect 202152 993286 202158 993338
rect 209730 993286 209736 993338
rect 209788 993326 209794 993338
rect 209788 993298 225232 993326
rect 209788 993286 209794 993298
rect 150224 993230 151724 993258
rect 191606 993150 191612 993202
rect 191664 993190 191670 993202
rect 209546 993190 209552 993202
rect 191664 993162 209552 993190
rect 191664 993150 191670 993162
rect 209546 993150 209552 993162
rect 209604 993150 209610 993202
rect 178542 993082 178548 993134
rect 178600 993122 178606 993134
rect 190962 993122 190968 993134
rect 178600 993094 190968 993122
rect 178600 993082 178606 993094
rect 190962 993082 190968 993094
rect 191020 993122 191026 993134
rect 209822 993122 209828 993134
rect 191020 993094 209828 993122
rect 191020 993082 191026 993094
rect 209822 993082 209828 993094
rect 209880 993082 209886 993134
rect 225204 993054 225232 993298
rect 261084 993298 261204 993326
rect 261084 993054 261112 993298
rect 261176 993258 261204 993298
rect 274038 993286 274044 993338
rect 274096 993326 274102 993338
rect 286826 993326 286832 993338
rect 274096 993298 286832 993326
rect 274096 993286 274102 993298
rect 286826 993286 286832 993298
rect 286884 993286 286890 993338
rect 261176 993230 273992 993258
rect 273964 993122 273992 993230
rect 295842 993190 295848 993202
rect 283256 993162 295848 993190
rect 283256 993122 283284 993162
rect 295842 993150 295848 993162
rect 295900 993150 295906 993202
rect 299724 993190 299752 993434
rect 299798 993422 299804 993474
rect 299856 993462 299862 993474
rect 300810 993462 300816 993474
rect 299856 993434 300816 993462
rect 299856 993422 299862 993434
rect 300810 993422 300816 993434
rect 300868 993462 300874 993474
rect 353158 993462 353164 993474
rect 300868 993434 353164 993462
rect 300868 993422 300874 993434
rect 353158 993422 353164 993434
rect 353216 993462 353222 993474
rect 406610 993462 406616 993474
rect 353216 993434 406616 993462
rect 353216 993422 353222 993434
rect 406610 993422 406616 993434
rect 406668 993462 406674 993474
rect 463374 993462 463380 993474
rect 406668 993434 463380 993462
rect 406668 993422 406674 993434
rect 463374 993422 463380 993434
rect 463432 993462 463438 993474
rect 517286 993462 517292 993474
rect 463432 993434 517292 993462
rect 463432 993422 463438 993434
rect 517286 993422 517292 993434
rect 517344 993422 517350 993474
rect 517378 993422 517384 993474
rect 517436 993462 517442 993474
rect 625570 993462 625576 993474
rect 517436 993434 625576 993462
rect 517436 993422 517442 993434
rect 625570 993422 625576 993434
rect 625628 993422 625634 993474
rect 305134 993354 305140 993406
rect 305192 993394 305198 993406
rect 313138 993394 313144 993406
rect 305192 993366 313144 993394
rect 305192 993354 305198 993366
rect 313138 993354 313144 993366
rect 313196 993354 313202 993406
rect 419122 993394 419128 993406
rect 411964 993366 419128 993394
rect 411964 993326 411992 993366
rect 419122 993354 419128 993366
rect 419180 993354 419186 993406
rect 528510 993394 528516 993406
rect 492924 993366 528516 993394
rect 437798 993326 437804 993338
rect 399176 993298 411992 993326
rect 428616 993298 437804 993326
rect 334666 993218 334672 993270
rect 334724 993258 334730 993270
rect 338346 993258 338352 993270
rect 334724 993230 338352 993258
rect 334724 993218 334730 993230
rect 338346 993218 338352 993230
rect 338404 993218 338410 993270
rect 338438 993218 338444 993270
rect 338496 993258 338502 993270
rect 338496 993230 341152 993258
rect 338496 993218 338502 993230
rect 300166 993190 300172 993202
rect 299724 993162 300172 993190
rect 300166 993150 300172 993162
rect 300224 993190 300230 993202
rect 300224 993162 304536 993190
rect 300224 993150 300230 993162
rect 273964 993094 283284 993122
rect 304508 993122 304536 993162
rect 312770 993150 312776 993202
rect 312828 993190 312834 993202
rect 321878 993190 321884 993202
rect 312828 993162 321884 993190
rect 312828 993150 312834 993162
rect 321878 993150 321884 993162
rect 321936 993150 321942 993202
rect 341124 993190 341152 993230
rect 360426 993218 360432 993270
rect 360484 993258 360490 993270
rect 364106 993258 364112 993270
rect 360484 993230 364112 993258
rect 360484 993218 360490 993230
rect 364106 993218 364112 993230
rect 364164 993218 364170 993270
rect 364198 993218 364204 993270
rect 364256 993258 364262 993270
rect 364256 993230 366912 993258
rect 364256 993218 364262 993230
rect 347638 993190 347644 993202
rect 341124 993162 347644 993190
rect 347638 993150 347644 993162
rect 347696 993150 347702 993202
rect 366884 993190 366912 993230
rect 386186 993218 386192 993270
rect 386244 993258 386250 993270
rect 389866 993258 389872 993270
rect 386244 993230 389872 993258
rect 386244 993218 386250 993230
rect 389866 993218 389872 993230
rect 389924 993218 389930 993270
rect 389958 993218 389964 993270
rect 390016 993258 390022 993270
rect 390016 993230 392672 993258
rect 390016 993218 390022 993230
rect 373398 993190 373404 993202
rect 366884 993162 373404 993190
rect 373398 993150 373404 993162
rect 373456 993150 373462 993202
rect 392644 993190 392672 993230
rect 399176 993190 399204 993298
rect 419122 993218 419128 993270
rect 419180 993258 419186 993270
rect 428616 993258 428644 993298
rect 437798 993286 437804 993298
rect 437856 993286 437862 993338
rect 450586 993286 450592 993338
rect 450644 993326 450650 993338
rect 466962 993326 466968 993338
rect 450644 993298 454312 993326
rect 450644 993286 450650 993298
rect 419180 993230 428644 993258
rect 454284 993258 454312 993298
rect 454376 993298 466968 993326
rect 454376 993258 454404 993298
rect 466962 993286 466968 993298
rect 467020 993286 467026 993338
rect 492924 993326 492952 993366
rect 528510 993354 528516 993366
rect 528568 993354 528574 993406
rect 480136 993298 492952 993326
rect 454284 993230 454404 993258
rect 419180 993218 419186 993230
rect 473862 993218 473868 993270
rect 473920 993258 473926 993270
rect 480136 993258 480164 993298
rect 522346 993286 522352 993338
rect 522404 993326 522410 993338
rect 530350 993326 530356 993338
rect 522404 993298 530356 993326
rect 522404 993286 522410 993298
rect 530350 993286 530356 993298
rect 530408 993286 530414 993338
rect 473920 993230 480164 993258
rect 473920 993218 473926 993230
rect 392644 993162 399204 993190
rect 312586 993122 312592 993134
rect 304508 993094 312592 993122
rect 312586 993082 312592 993094
rect 312644 993082 312650 993134
rect 225204 993026 231764 993054
rect 231736 992986 231764 993026
rect 257404 993026 261112 993054
rect 257404 992998 257432 993026
rect 231736 992958 231856 992986
rect 231828 992850 231856 992958
rect 257386 992946 257392 992998
rect 257444 992946 257450 992998
rect 296026 992946 296032 992998
rect 296084 992986 296090 992998
rect 299706 992986 299712 992998
rect 296084 992958 299712 992986
rect 296084 992946 296090 992958
rect 299706 992946 299712 992958
rect 299764 992946 299770 992998
rect 244598 992850 244604 992862
rect 231828 992822 244604 992850
rect 244598 992810 244604 992822
rect 244656 992810 244662 992862
rect 636702 992810 636708 992862
rect 636760 992850 636766 992862
rect 675158 992850 675164 992862
rect 636760 992822 675164 992850
rect 636760 992810 636766 992822
rect 675158 992810 675164 992822
rect 675216 992810 675222 992862
rect 625754 992742 625760 992794
rect 625812 992782 625818 992794
rect 675342 992782 675348 992794
rect 625812 992754 675348 992782
rect 625812 992742 625818 992754
rect 675342 992742 675348 992754
rect 675400 992742 675406 992794
rect 244598 992674 244604 992726
rect 244656 992714 244662 992726
rect 246162 992714 246168 992726
rect 244656 992686 246168 992714
rect 244656 992674 244662 992686
rect 246162 992674 246168 992686
rect 246220 992714 246226 992726
rect 257386 992714 257392 992726
rect 246220 992686 257392 992714
rect 246220 992674 246226 992686
rect 257386 992674 257392 992686
rect 257444 992674 257450 992726
rect 625570 992674 625576 992726
rect 625628 992714 625634 992726
rect 675250 992714 675256 992726
rect 625628 992686 675256 992714
rect 625628 992674 625634 992686
rect 675250 992674 675256 992686
rect 675308 992674 675314 992726
rect 81666 992334 81672 992386
rect 81724 992374 81730 992386
rect 82402 992374 82408 992386
rect 81724 992346 82408 992374
rect 81724 992334 81730 992346
rect 82402 992334 82408 992346
rect 82460 992334 82466 992386
rect 364198 975198 364204 975250
rect 364256 975238 364262 975250
rect 364382 975238 364388 975250
rect 364256 975210 364388 975238
rect 364256 975198 364262 975210
rect 364382 975198 364388 975210
rect 364440 975198 364446 975250
rect 581318 975198 581324 975250
rect 581376 975238 581382 975250
rect 581502 975238 581508 975250
rect 581376 975210 581508 975238
rect 581376 975198 581382 975210
rect 581502 975198 581508 975210
rect 581560 975198 581566 975250
rect 42106 970574 42112 970626
rect 42164 970614 42170 970626
rect 92706 970614 92712 970626
rect 42164 970586 92712 970614
rect 42164 970574 42170 970586
rect 92706 970574 92712 970586
rect 92764 970574 92770 970626
rect 41646 968126 41652 968178
rect 41704 968166 41710 968178
rect 42290 968166 42296 968178
rect 41704 968138 42296 968166
rect 41704 968126 41710 968138
rect 42290 968126 42296 968138
rect 42348 968126 42354 968178
rect 41646 967242 41652 967294
rect 41704 967282 41710 967294
rect 42198 967282 42204 967294
rect 41704 967254 42204 967282
rect 41704 967242 41710 967254
rect 42198 967242 42204 967254
rect 42256 967242 42262 967294
rect 674974 966018 674980 966070
rect 675032 966058 675038 966070
rect 675342 966058 675348 966070
rect 675032 966030 675348 966058
rect 675032 966018 675038 966030
rect 675342 966018 675348 966030
rect 675400 966018 675406 966070
rect 675066 965950 675072 966002
rect 675124 965990 675130 966002
rect 675250 965990 675256 966002
rect 675124 965962 675256 965990
rect 675124 965950 675130 965962
rect 675250 965950 675256 965962
rect 675308 965950 675314 966002
rect 675158 963978 675164 964030
rect 675216 963978 675222 964030
rect 675176 963826 675204 963978
rect 675158 963774 675164 963826
rect 675216 963774 675222 963826
rect 674974 962958 674980 963010
rect 675032 962998 675038 963010
rect 675250 962998 675256 963010
rect 675032 962970 675256 962998
rect 675032 962958 675038 962970
rect 675250 962958 675256 962970
rect 675308 962958 675314 963010
rect 42014 962414 42020 962466
rect 42072 962454 42078 962466
rect 42198 962454 42204 962466
rect 42072 962426 42204 962454
rect 42072 962414 42078 962426
rect 42198 962414 42204 962426
rect 42256 962414 42262 962466
rect 675158 962346 675164 962398
rect 675216 962346 675222 962398
rect 675176 962194 675204 962346
rect 675158 962142 675164 962194
rect 675216 962142 675222 962194
rect 42106 961870 42112 961922
rect 42164 961910 42170 961922
rect 42290 961910 42296 961922
rect 42164 961882 42296 961910
rect 42164 961870 42170 961882
rect 42290 961870 42296 961882
rect 42348 961870 42354 961922
rect 43026 960102 43032 960154
rect 43084 960142 43090 960154
rect 364382 960142 364388 960154
rect 43084 960114 364388 960142
rect 43084 960102 43090 960114
rect 364382 960102 364388 960114
rect 364440 960102 364446 960154
rect 99606 960034 99612 960086
rect 99664 960074 99670 960086
rect 632930 960074 632936 960086
rect 99664 960046 632936 960074
rect 99664 960034 99670 960046
rect 632930 960034 632936 960046
rect 632988 960034 632994 960086
rect 674790 958606 674796 958658
rect 674848 958646 674854 958658
rect 675158 958646 675164 958658
rect 674848 958618 675164 958646
rect 674848 958606 674854 958618
rect 675158 958606 675164 958618
rect 675216 958606 675222 958658
rect 41646 955818 41652 955870
rect 41704 955858 41710 955870
rect 42382 955858 42388 955870
rect 41704 955830 42388 955858
rect 41704 955818 41710 955830
rect 42382 955818 42388 955830
rect 42440 955818 42446 955870
rect 41646 955274 41652 955326
rect 41704 955314 41710 955326
rect 42198 955314 42204 955326
rect 41704 955286 42204 955314
rect 41704 955274 41710 955286
rect 42198 955274 42204 955286
rect 42256 955274 42262 955326
rect 632930 954934 632936 954986
rect 632988 954974 632994 954986
rect 641026 954974 641032 954986
rect 632988 954946 641032 954974
rect 632988 954934 632994 954946
rect 641026 954934 641032 954946
rect 641084 954934 641090 954986
rect 93902 953778 93908 953830
rect 93960 953818 93966 953830
rect 99606 953818 99612 953830
rect 93960 953790 99612 953818
rect 93960 953778 93966 953790
rect 99606 953778 99612 953790
rect 99664 953778 99670 953830
rect 41646 953030 41652 953082
rect 41704 953070 41710 953082
rect 42382 953070 42388 953082
rect 41704 953042 42388 953070
rect 41704 953030 41710 953042
rect 42382 953030 42388 953042
rect 42440 953070 42446 953082
rect 81666 953070 81672 953082
rect 42440 953042 81672 953070
rect 42440 953030 42446 953042
rect 81666 953030 81672 953042
rect 81724 953030 81730 953082
rect 42198 952962 42204 953014
rect 42256 953002 42262 953014
rect 81758 953002 81764 953014
rect 42256 952974 81764 953002
rect 42256 952962 42262 952974
rect 81758 952962 81764 952974
rect 81816 952962 81822 953014
rect 674790 951874 674796 951926
rect 674848 951914 674854 951926
rect 675250 951914 675256 951926
rect 674848 951886 675256 951914
rect 674848 951874 674854 951886
rect 675250 951874 675256 951886
rect 675308 951874 675314 951926
rect 92430 951330 92436 951382
rect 92488 951370 92494 951382
rect 93902 951370 93908 951382
rect 92488 951342 93908 951370
rect 92488 951330 92494 951342
rect 93902 951330 93908 951342
rect 93960 951330 93966 951382
rect 581318 949426 581324 949478
rect 581376 949466 581382 949478
rect 581502 949466 581508 949478
rect 581376 949438 581508 949466
rect 581376 949426 581382 949438
rect 581502 949426 581508 949438
rect 581560 949426 581566 949478
rect 674790 948542 674796 948594
rect 674848 948582 674854 948594
rect 675158 948582 675164 948594
rect 674848 948554 675164 948582
rect 674848 948542 674854 948554
rect 675158 948542 675164 948554
rect 675216 948542 675222 948594
rect 641026 947590 641032 947642
rect 641084 947630 641090 947642
rect 641084 947602 642084 947630
rect 641084 947590 641090 947602
rect 642056 947562 642084 947602
rect 646638 947562 646644 947574
rect 642056 947534 646644 947562
rect 646638 947522 646644 947534
rect 646696 947522 646702 947574
rect 646638 943374 646644 943426
rect 646696 943414 646702 943426
rect 653906 943414 653912 943426
rect 646696 943386 653912 943414
rect 646696 943374 646702 943386
rect 653906 943374 653912 943386
rect 653964 943374 653970 943426
rect 90038 941130 90044 941182
rect 90096 941170 90102 941182
rect 92430 941170 92436 941182
rect 90096 941142 92436 941170
rect 90096 941130 90102 941142
rect 92430 941130 92436 941142
rect 92488 941130 92494 941182
rect 88198 937458 88204 937510
rect 88256 937498 88262 937510
rect 90038 937498 90044 937510
rect 88256 937470 90044 937498
rect 88256 937458 88262 937470
rect 90038 937458 90044 937470
rect 90096 937458 90102 937510
rect 87002 934738 87008 934790
rect 87060 934778 87066 934790
rect 88198 934778 88204 934790
rect 87060 934750 88204 934778
rect 87060 934738 87066 934750
rect 88198 934738 88204 934750
rect 88256 934738 88262 934790
rect 653906 934738 653912 934790
rect 653964 934778 653970 934790
rect 655746 934778 655752 934790
rect 653964 934750 655752 934778
rect 653964 934738 653970 934750
rect 655746 934738 655752 934750
rect 655804 934738 655810 934790
rect 80838 931882 80844 931934
rect 80896 931922 80902 931934
rect 87002 931922 87008 931934
rect 80896 931894 87008 931922
rect 80896 931882 80902 931894
rect 87002 931882 87008 931894
rect 87060 931882 87066 931934
rect 44038 926442 44044 926494
rect 44096 926482 44102 926494
rect 80838 926482 80844 926494
rect 44096 926454 80844 926482
rect 44096 926442 44102 926454
rect 80838 926442 80844 926454
rect 80896 926442 80902 926494
rect 39254 925558 39260 925610
rect 39312 925598 39318 925610
rect 44038 925598 44044 925610
rect 39312 925570 44044 925598
rect 39312 925558 39318 925570
rect 44038 925558 44044 925570
rect 44096 925558 44102 925610
rect 581318 923722 581324 923774
rect 581376 923762 581382 923774
rect 581502 923762 581508 923774
rect 581376 923734 581508 923762
rect 581376 923722 581382 923734
rect 581502 923722 581508 923734
rect 581560 923722 581566 923774
rect 655746 919982 655752 920034
rect 655804 920022 655810 920034
rect 655804 919994 656804 920022
rect 655804 919982 655810 919994
rect 656776 919954 656804 919994
rect 661266 919954 661272 919966
rect 656776 919926 661272 919954
rect 661266 919914 661272 919926
rect 661324 919914 661330 919966
rect 39622 913250 39628 913302
rect 39680 913290 39686 913302
rect 40450 913290 40456 913302
rect 39680 913262 40456 913290
rect 39680 913250 39686 913262
rect 40450 913250 40456 913262
rect 40508 913290 40514 913302
rect 41646 913290 41652 913302
rect 40508 913262 41652 913290
rect 40508 913250 40514 913262
rect 41646 913250 41652 913262
rect 41704 913250 41710 913302
rect 661266 908898 661272 908950
rect 661324 908938 661330 908950
rect 669454 908938 669460 908950
rect 661324 908910 669460 908938
rect 661324 908898 661330 908910
rect 669454 908898 669460 908910
rect 669512 908898 669518 908950
rect 675342 908898 675348 908950
rect 675400 908938 675406 908950
rect 677550 908938 677556 908950
rect 675400 908910 677556 908938
rect 675400 908898 675406 908910
rect 677550 908898 677556 908910
rect 677608 908898 677614 908950
rect 669454 905294 669460 905346
rect 669512 905334 669518 905346
rect 669512 905306 671524 905334
rect 669512 905294 669518 905306
rect 671496 905266 671524 905306
rect 677550 905266 677556 905278
rect 671496 905238 677556 905266
rect 677550 905226 677556 905238
rect 677608 905226 677614 905278
rect 674514 875306 674520 875358
rect 674572 875346 674578 875358
rect 675066 875346 675072 875358
rect 674572 875318 675072 875346
rect 674572 875306 674578 875318
rect 675066 875306 675072 875318
rect 675124 875306 675130 875358
rect 675158 875034 675164 875086
rect 675216 875074 675222 875086
rect 675342 875074 675348 875086
rect 675216 875046 675348 875074
rect 675216 875034 675222 875046
rect 675342 875034 675348 875046
rect 675400 875034 675406 875086
rect 674974 873742 674980 873794
rect 675032 873782 675038 873794
rect 675250 873782 675256 873794
rect 675032 873754 675256 873782
rect 675032 873742 675038 873754
rect 675250 873742 675256 873754
rect 675308 873742 675314 873794
rect 41922 872178 41928 872230
rect 41980 872218 41986 872230
rect 42106 872218 42112 872230
rect 41980 872190 42112 872218
rect 41980 872178 41986 872190
rect 42106 872178 42112 872190
rect 42164 872178 42170 872230
rect 581318 872178 581324 872230
rect 581376 872218 581382 872230
rect 581502 872218 581508 872230
rect 581376 872190 581508 872218
rect 581376 872178 581382 872190
rect 581502 872178 581508 872190
rect 581560 872178 581566 872230
rect 674974 871702 674980 871754
rect 675032 871742 675038 871754
rect 675250 871742 675256 871754
rect 675032 871714 675256 871742
rect 675032 871702 675038 871714
rect 675250 871702 675256 871714
rect 675308 871702 675314 871754
rect 675158 870138 675164 870190
rect 675216 870138 675222 870190
rect 675176 869986 675204 870138
rect 675158 869934 675164 869986
rect 675216 869934 675222 869986
rect 674882 866738 674888 866790
rect 674940 866778 674946 866790
rect 675158 866778 675164 866790
rect 674940 866750 675164 866778
rect 674940 866738 674946 866750
rect 675158 866738 675164 866750
rect 675216 866738 675222 866790
rect 39714 865786 39720 865838
rect 39772 865826 39778 865838
rect 40450 865826 40456 865838
rect 39772 865798 40456 865826
rect 39772 865786 39778 865798
rect 40450 865786 40456 865798
rect 40508 865826 40514 865838
rect 41646 865826 41652 865838
rect 40508 865798 41652 865826
rect 40508 865786 40514 865798
rect 41646 865786 41652 865798
rect 41704 865786 41710 865838
rect 674514 862998 674520 863050
rect 674572 863038 674578 863050
rect 674606 863038 674612 863050
rect 674572 863010 674612 863038
rect 674572 862998 674578 863010
rect 674606 862998 674612 863010
rect 674664 862998 674670 863050
rect 674882 860618 674888 860670
rect 674940 860658 674946 860670
rect 675250 860658 675256 860670
rect 674940 860630 675256 860658
rect 674940 860618 674946 860630
rect 675250 860618 675256 860630
rect 675308 860618 675314 860670
rect 674606 853682 674612 853734
rect 674664 853722 674670 853734
rect 674974 853722 674980 853734
rect 674664 853694 674980 853722
rect 674664 853682 674670 853694
rect 674974 853682 674980 853694
rect 675032 853682 675038 853734
rect 675250 850010 675256 850062
rect 675308 850050 675314 850062
rect 675342 850050 675348 850062
rect 675308 850022 675348 850050
rect 675308 850010 675314 850022
rect 675342 850010 675348 850022
rect 675400 850010 675406 850062
rect 41738 846474 41744 846526
rect 41796 846514 41802 846526
rect 41922 846514 41928 846526
rect 41796 846486 41928 846514
rect 41796 846474 41802 846486
rect 41922 846474 41928 846486
rect 41980 846474 41986 846526
rect 581318 846406 581324 846458
rect 581376 846446 581382 846458
rect 581502 846446 581508 846458
rect 581376 846418 581508 846446
rect 581376 846406 581382 846418
rect 581502 846406 581508 846418
rect 581560 846406 581566 846458
rect 674882 840898 674888 840950
rect 674940 840898 674946 840950
rect 674900 840870 674928 840898
rect 674974 840870 674980 840882
rect 674900 840842 674980 840870
rect 674974 840830 674980 840842
rect 675032 840830 675038 840882
rect 41738 837226 41744 837278
rect 41796 837266 41802 837278
rect 42014 837266 42020 837278
rect 41796 837238 42020 837266
rect 41796 837226 41802 837238
rect 42014 837226 42020 837238
rect 42072 837226 42078 837278
rect 674882 837226 674888 837278
rect 674940 837266 674946 837278
rect 674974 837266 674980 837278
rect 674940 837238 674980 837266
rect 674940 837226 674946 837238
rect 674974 837226 674980 837238
rect 675032 837226 675038 837278
rect 675250 837226 675256 837278
rect 675308 837266 675314 837278
rect 675526 837266 675532 837278
rect 675308 837238 675532 837266
rect 675308 837226 675314 837238
rect 675526 837226 675532 837238
rect 675584 837226 675590 837278
rect 675158 836138 675164 836190
rect 675216 836178 675222 836190
rect 675434 836178 675440 836190
rect 675216 836150 675440 836178
rect 675216 836138 675222 836150
rect 675434 836138 675440 836150
rect 675492 836138 675498 836190
rect 42014 828086 42020 828098
rect 41940 828058 42020 828086
rect 41940 827962 41968 828058
rect 42014 828046 42020 828058
rect 42072 828046 42078 828098
rect 675250 827978 675256 828030
rect 675308 828018 675314 828030
rect 675526 828018 675532 828030
rect 675308 827990 675532 828018
rect 675308 827978 675314 827990
rect 675526 827978 675532 827990
rect 675584 827978 675590 828030
rect 41922 827910 41928 827962
rect 41980 827910 41986 827962
rect 573958 821518 573964 821570
rect 574016 821558 574022 821570
rect 674974 821558 674980 821570
rect 574016 821530 674980 821558
rect 574016 821518 574022 821530
rect 674974 821518 674980 821530
rect 675032 821518 675038 821570
rect 675158 821518 675164 821570
rect 675216 821558 675222 821570
rect 675434 821558 675440 821570
rect 675216 821530 675440 821558
rect 675216 821518 675222 821530
rect 675434 821518 675440 821530
rect 675492 821518 675498 821570
rect 581318 820634 581324 820686
rect 581376 820674 581382 820686
rect 581502 820674 581508 820686
rect 581376 820646 581508 820674
rect 581376 820634 581382 820646
rect 581502 820634 581508 820646
rect 581560 820634 581566 820686
rect 581318 817846 581324 817898
rect 581376 817886 581382 817898
rect 674882 817886 674888 817898
rect 581376 817858 674888 817886
rect 581376 817846 581382 817858
rect 674882 817846 674888 817858
rect 674940 817846 674946 817898
rect 675250 811386 675256 811438
rect 675308 811426 675314 811438
rect 675342 811426 675348 811438
rect 675308 811398 675348 811426
rect 675308 811386 675314 811398
rect 675342 811386 675348 811398
rect 675400 811386 675406 811438
rect 674698 809550 674704 809602
rect 674756 809590 674762 809602
rect 674882 809590 674888 809602
rect 674756 809562 674888 809590
rect 674756 809550 674762 809562
rect 674882 809550 674888 809562
rect 674940 809550 674946 809602
rect 675158 808258 675164 808310
rect 675216 808298 675222 808310
rect 675434 808298 675440 808310
rect 675216 808270 675440 808298
rect 675216 808258 675222 808270
rect 675434 808258 675440 808270
rect 675492 808258 675498 808310
rect 675342 798602 675348 798654
rect 675400 798642 675406 798654
rect 675526 798642 675532 798654
rect 675400 798614 675532 798642
rect 675400 798602 675406 798614
rect 675526 798602 675532 798614
rect 675584 798602 675590 798654
rect 674698 796698 674704 796750
rect 674756 796738 674762 796750
rect 674882 796738 674888 796750
rect 674756 796710 674888 796738
rect 674756 796698 674762 796710
rect 674882 796698 674888 796710
rect 674940 796698 674946 796750
rect 675158 795746 675164 795798
rect 675216 795786 675222 795798
rect 675434 795786 675440 795798
rect 675216 795758 675440 795786
rect 675216 795746 675222 795758
rect 675434 795746 675440 795758
rect 675492 795746 675498 795798
rect 41922 793910 41928 793962
rect 41980 793950 41986 793962
rect 42566 793950 42572 793962
rect 41980 793922 42572 793950
rect 41980 793910 41986 793922
rect 42566 793910 42572 793922
rect 42624 793910 42630 793962
rect 41646 791122 41652 791174
rect 41704 791162 41710 791174
rect 42566 791162 42572 791174
rect 41704 791134 42572 791162
rect 41704 791122 41710 791134
rect 42566 791122 42572 791134
rect 42624 791122 42630 791174
rect 674790 790442 674796 790494
rect 674848 790482 674854 790494
rect 675066 790482 675072 790494
rect 674848 790454 675072 790482
rect 674848 790442 674854 790454
rect 675066 790442 675072 790454
rect 675124 790442 675130 790494
rect 674790 782894 674796 782946
rect 674848 782934 674854 782946
rect 675066 782934 675072 782946
rect 674848 782906 675072 782934
rect 674848 782894 674854 782906
rect 675066 782894 675072 782906
rect 675124 782894 675130 782946
rect 42106 782078 42112 782130
rect 42164 782118 42170 782130
rect 42566 782118 42572 782130
rect 42164 782090 42572 782118
rect 42164 782078 42170 782090
rect 42566 782078 42572 782090
rect 42624 782078 42630 782130
rect 41646 781874 41652 781926
rect 41704 781874 41710 781926
rect 41664 781722 41692 781874
rect 41646 781670 41652 781722
rect 41704 781670 41710 781722
rect 674514 781534 674520 781586
rect 674572 781574 674578 781586
rect 675526 781574 675532 781586
rect 674572 781546 675532 781574
rect 674572 781534 674578 781546
rect 675526 781534 675532 781546
rect 675584 781534 675590 781586
rect 674514 778950 674520 779002
rect 674572 778990 674578 779002
rect 675250 778990 675256 779002
rect 674572 778962 675256 778990
rect 674572 778950 674578 778962
rect 675250 778950 675256 778962
rect 675308 778950 675314 779002
rect 674698 778542 674704 778594
rect 674756 778582 674762 778594
rect 675158 778582 675164 778594
rect 674756 778554 675164 778582
rect 674756 778542 674762 778554
rect 675158 778542 675164 778554
rect 675216 778542 675222 778594
rect 674790 774190 674796 774242
rect 674848 774230 674854 774242
rect 675158 774230 675164 774242
rect 674848 774202 675164 774230
rect 674848 774190 674854 774202
rect 675158 774190 675164 774202
rect 675216 774190 675222 774242
rect 674606 770042 674612 770094
rect 674664 770082 674670 770094
rect 675066 770082 675072 770094
rect 674664 770054 675072 770082
rect 674664 770042 674670 770054
rect 675066 770042 675072 770054
rect 675124 770042 675130 770094
rect 674698 768478 674704 768530
rect 674756 768518 674762 768530
rect 675250 768518 675256 768530
rect 674756 768490 675256 768518
rect 674756 768478 674762 768490
rect 675250 768478 675256 768490
rect 675308 768478 675314 768530
rect 675158 767594 675164 767646
rect 675216 767594 675222 767646
rect 675176 767442 675204 767594
rect 675158 767390 675164 767442
rect 675216 767390 675222 767442
rect 674790 765962 674796 766014
rect 674848 766002 674854 766014
rect 675526 766002 675532 766014
rect 674848 765974 675532 766002
rect 674848 765962 674854 765974
rect 675526 765962 675532 765974
rect 675584 765962 675590 766014
rect 674514 765894 674520 765946
rect 674572 765934 674578 765946
rect 675250 765934 675256 765946
rect 674572 765906 675256 765934
rect 674572 765894 674578 765906
rect 675250 765894 675256 765906
rect 675308 765894 675314 765946
rect 674422 759978 674428 760030
rect 674480 760018 674486 760030
rect 674882 760018 674888 760030
rect 674480 759990 674888 760018
rect 674480 759978 674486 759990
rect 674882 759978 674888 759990
rect 674940 759978 674946 760030
rect 674698 758006 674704 758058
rect 674756 758046 674762 758058
rect 674882 758046 674888 758058
rect 674756 758018 674888 758046
rect 674756 758006 674762 758018
rect 674882 758006 674888 758018
rect 674940 758006 674946 758058
rect 675526 758006 675532 758058
rect 675584 758046 675590 758058
rect 675710 758046 675716 758058
rect 675584 758018 675716 758046
rect 675584 758006 675590 758018
rect 675710 758006 675716 758018
rect 675768 758006 675774 758058
rect 674606 757122 674612 757174
rect 674664 757162 674670 757174
rect 675066 757162 675072 757174
rect 674664 757134 675072 757162
rect 674664 757122 674670 757134
rect 675066 757122 675072 757134
rect 675124 757122 675130 757174
rect 42106 749778 42112 749830
rect 42164 749818 42170 749830
rect 42566 749818 42572 749830
rect 42164 749790 42572 749818
rect 42164 749778 42170 749790
rect 42566 749778 42572 749790
rect 42624 749778 42630 749830
rect 41646 748350 41652 748402
rect 41704 748390 41710 748402
rect 42658 748390 42664 748402
rect 41704 748362 42664 748390
rect 41704 748350 41710 748362
rect 42658 748350 42664 748362
rect 42716 748350 42722 748402
rect 41830 747126 41836 747178
rect 41888 747166 41894 747178
rect 42566 747166 42572 747178
rect 41888 747138 42572 747166
rect 41888 747126 41894 747138
rect 42566 747126 42572 747138
rect 42624 747126 42630 747178
rect 41830 746514 41836 746566
rect 41888 746554 41894 746566
rect 42566 746554 42572 746566
rect 41888 746526 42572 746554
rect 41888 746514 41894 746526
rect 42566 746514 42572 746526
rect 42624 746514 42630 746566
rect 674790 744270 674796 744322
rect 674848 744310 674854 744322
rect 674974 744310 674980 744322
rect 674848 744282 674980 744310
rect 674848 744270 674854 744282
rect 674974 744270 674980 744282
rect 675032 744270 675038 744322
rect 42106 743386 42112 743438
rect 42164 743426 42170 743438
rect 42658 743426 42664 743438
rect 42164 743398 42664 743426
rect 42164 743386 42170 743398
rect 42658 743386 42664 743398
rect 42716 743386 42722 743438
rect 41646 741414 41652 741466
rect 41704 741454 41710 741466
rect 42106 741454 42112 741466
rect 41704 741426 42112 741454
rect 41704 741414 41710 741426
rect 42106 741414 42112 741426
rect 42164 741414 42170 741466
rect 674606 735294 674612 735346
rect 674664 735334 674670 735346
rect 675066 735334 675072 735346
rect 674664 735306 675072 735334
rect 674664 735294 674670 735306
rect 675066 735294 675072 735306
rect 675124 735294 675130 735346
rect 674698 735226 674704 735278
rect 674756 735266 674762 735278
rect 675158 735266 675164 735278
rect 674756 735238 675164 735266
rect 674756 735226 674762 735238
rect 675158 735226 675164 735238
rect 675216 735226 675222 735278
rect 674882 734342 674888 734394
rect 674940 734342 674946 734394
rect 674900 734258 674928 734342
rect 674882 734206 674888 734258
rect 674940 734206 674946 734258
rect 42106 733254 42112 733306
rect 42164 733294 42170 733306
rect 42566 733294 42572 733306
rect 42164 733266 42572 733294
rect 42164 733254 42170 733266
rect 42566 733254 42572 733266
rect 42624 733254 42630 733306
rect 675158 725298 675164 725350
rect 675216 725298 675222 725350
rect 675066 725026 675072 725078
rect 675124 725066 675130 725078
rect 675176 725066 675204 725298
rect 675124 725038 675204 725066
rect 675124 725026 675130 725038
rect 674606 724958 674612 725010
rect 674664 724998 674670 725010
rect 674974 724998 674980 725010
rect 674664 724970 674980 724998
rect 674664 724958 674670 724970
rect 674974 724958 674980 724970
rect 675032 724958 675038 725010
rect 674698 722034 674704 722086
rect 674756 722074 674762 722086
rect 675250 722074 675256 722086
rect 674756 722046 675256 722074
rect 674756 722034 674762 722046
rect 675250 722034 675256 722046
rect 675308 722034 675314 722086
rect 674422 721898 674428 721950
rect 674480 721938 674486 721950
rect 674698 721938 674704 721950
rect 674480 721910 674704 721938
rect 674480 721898 674486 721910
rect 674698 721898 674704 721910
rect 674756 721898 674762 721950
rect 41738 721286 41744 721338
rect 41796 721326 41802 721338
rect 42014 721326 42020 721338
rect 41796 721298 42020 721326
rect 41796 721286 41802 721298
rect 42014 721286 42020 721298
rect 42072 721286 42078 721338
rect 675066 720198 675072 720250
rect 675124 720238 675130 720250
rect 675250 720238 675256 720250
rect 675124 720210 675256 720238
rect 675124 720198 675130 720210
rect 675250 720198 675256 720210
rect 675308 720198 675314 720250
rect 674606 714894 674612 714946
rect 674664 714934 674670 714946
rect 674974 714934 674980 714946
rect 674664 714906 674980 714934
rect 674664 714894 674670 714906
rect 674974 714894 674980 714906
rect 675032 714894 675038 714946
rect 674698 708502 674704 708554
rect 674756 708542 674762 708554
rect 674882 708542 674888 708554
rect 674756 708514 674888 708542
rect 674756 708502 674762 708514
rect 674882 708502 674888 708514
rect 674940 708502 674946 708554
rect 674606 708366 674612 708418
rect 674664 708406 674670 708418
rect 675066 708406 675072 708418
rect 674664 708378 675072 708406
rect 674664 708366 674670 708378
rect 675066 708366 675072 708378
rect 675124 708366 675130 708418
rect 675158 708366 675164 708418
rect 675216 708406 675222 708418
rect 675342 708406 675348 708418
rect 675216 708378 675348 708406
rect 675216 708366 675222 708378
rect 675342 708366 675348 708378
rect 675400 708366 675406 708418
rect 674698 706530 674704 706582
rect 674756 706570 674762 706582
rect 674882 706570 674888 706582
rect 674756 706542 674888 706570
rect 674756 706530 674762 706542
rect 674882 706530 674888 706542
rect 674940 706530 674946 706582
rect 675158 705646 675164 705698
rect 675216 705686 675222 705698
rect 675434 705686 675440 705698
rect 675216 705658 675440 705686
rect 675216 705646 675222 705658
rect 675434 705646 675440 705658
rect 675492 705646 675498 705698
rect 41646 702178 41652 702230
rect 41704 702218 41710 702230
rect 42106 702218 42112 702230
rect 41704 702190 42112 702218
rect 41704 702178 41710 702190
rect 42106 702178 42112 702190
rect 42164 702218 42170 702230
rect 42566 702218 42572 702230
rect 42164 702190 42572 702218
rect 42164 702178 42170 702190
rect 42566 702178 42572 702190
rect 42624 702178 42630 702230
rect 675342 699186 675348 699238
rect 675400 699226 675406 699238
rect 675400 699198 675664 699226
rect 675400 699186 675406 699198
rect 675636 699170 675664 699198
rect 675618 699118 675624 699170
rect 675676 699118 675682 699170
rect 674698 693678 674704 693730
rect 674756 693718 674762 693730
rect 674882 693718 674888 693730
rect 674756 693690 674888 693718
rect 674756 693678 674762 693690
rect 674882 693678 674888 693690
rect 674940 693678 674946 693730
rect 674790 692182 674796 692234
rect 674848 692222 674854 692234
rect 674974 692222 674980 692234
rect 674848 692194 674980 692222
rect 674848 692182 674854 692194
rect 674974 692182 674980 692194
rect 675032 692182 675038 692234
rect 41646 691094 41652 691146
rect 41704 691134 41710 691146
rect 42106 691134 42112 691146
rect 41704 691106 42112 691134
rect 41704 691094 41710 691106
rect 42106 691094 42112 691106
rect 42164 691094 42170 691146
rect 41646 688986 41652 689038
rect 41704 689026 41710 689038
rect 42106 689026 42112 689038
rect 41704 688998 42112 689026
rect 41704 688986 41710 688998
rect 42106 688986 42112 688998
rect 42164 688986 42170 689038
rect 674698 688714 674704 688766
rect 674756 688754 674762 688766
rect 675158 688754 675164 688766
rect 674756 688726 675164 688754
rect 674756 688714 674762 688726
rect 675158 688714 675164 688726
rect 675216 688714 675222 688766
rect 675158 688578 675164 688630
rect 675216 688618 675222 688630
rect 675618 688618 675624 688630
rect 675216 688590 675624 688618
rect 675216 688578 675222 688590
rect 675618 688578 675624 688590
rect 675676 688578 675682 688630
rect 674882 686442 674888 686454
rect 674808 686414 674888 686442
rect 674808 686318 674836 686414
rect 674882 686402 674888 686414
rect 674940 686402 674946 686454
rect 674790 686266 674796 686318
rect 674848 686266 674854 686318
rect 674514 682594 674520 682646
rect 674572 682634 674578 682646
rect 674790 682634 674796 682646
rect 674572 682606 674796 682634
rect 674572 682594 674578 682606
rect 674790 682594 674796 682606
rect 674848 682594 674854 682646
rect 674882 681166 674888 681218
rect 674940 681206 674946 681218
rect 675158 681206 675164 681218
rect 674940 681178 675164 681206
rect 674940 681166 674946 681178
rect 675158 681166 675164 681178
rect 675216 681166 675222 681218
rect 674514 680010 674520 680062
rect 674572 680050 674578 680062
rect 674790 680050 674796 680062
rect 674572 680022 674796 680050
rect 674572 680010 674578 680022
rect 674790 680010 674796 680022
rect 674848 680010 674854 680062
rect 674514 679874 674520 679926
rect 674572 679914 674578 679926
rect 674974 679914 674980 679926
rect 674572 679886 674980 679914
rect 674572 679874 674578 679886
rect 674974 679874 674980 679886
rect 675032 679874 675038 679926
rect 674422 675454 674428 675506
rect 674480 675494 674486 675506
rect 675250 675494 675256 675506
rect 674480 675466 675256 675494
rect 674480 675454 674486 675466
rect 675250 675454 675256 675466
rect 675308 675454 675314 675506
rect 41922 673590 41928 673602
rect 41848 673562 41928 673590
rect 41848 673398 41876 673562
rect 41922 673550 41928 673562
rect 41980 673550 41986 673602
rect 41830 673346 41836 673398
rect 41888 673346 41894 673398
rect 674974 672938 674980 672990
rect 675032 672978 675038 672990
rect 675250 672978 675256 672990
rect 675032 672950 675256 672978
rect 675032 672938 675038 672950
rect 675250 672938 675256 672950
rect 675308 672938 675314 672990
rect 674790 672870 674796 672922
rect 674848 672910 674854 672922
rect 675618 672910 675624 672922
rect 674848 672882 675624 672910
rect 674848 672870 674854 672882
rect 675618 672870 675624 672882
rect 675676 672870 675682 672922
rect 674422 672802 674428 672854
rect 674480 672842 674486 672854
rect 675342 672842 675348 672854
rect 674480 672814 675348 672842
rect 674480 672802 674486 672814
rect 675342 672802 675348 672814
rect 675400 672802 675406 672854
rect 674514 666954 674520 667006
rect 674572 666994 674578 667006
rect 674974 666994 674980 667006
rect 674572 666966 674980 666994
rect 674572 666954 674578 666966
rect 674974 666954 674980 666966
rect 675032 666954 675038 667006
rect 42106 660154 42112 660206
rect 42164 660194 42170 660206
rect 42566 660194 42572 660206
rect 42164 660166 42572 660194
rect 42164 660154 42170 660166
rect 42566 660154 42572 660166
rect 42624 660154 42630 660206
rect 41646 660018 41652 660070
rect 41704 660058 41710 660070
rect 42106 660058 42112 660070
rect 41704 660030 42112 660058
rect 41704 660018 41710 660030
rect 42106 660018 42112 660030
rect 42164 660018 42170 660070
rect 42014 653218 42020 653270
rect 42072 653258 42078 653270
rect 42658 653258 42664 653270
rect 42072 653230 42664 653258
rect 42072 653218 42078 653230
rect 42658 653218 42664 653230
rect 42716 653218 42722 653270
rect 41646 648050 41652 648102
rect 41704 648090 41710 648102
rect 42566 648090 42572 648102
rect 41704 648062 42572 648090
rect 41704 648050 41710 648062
rect 42566 648050 42572 648062
rect 42624 648050 42630 648102
rect 42014 647642 42020 647694
rect 42072 647642 42078 647694
rect 42032 647490 42060 647642
rect 41646 647438 41652 647490
rect 41704 647478 41710 647490
rect 42014 647478 42020 647490
rect 41704 647450 42020 647478
rect 41704 647438 41710 647450
rect 42014 647438 42020 647450
rect 42072 647438 42078 647490
rect 42106 644486 42112 644498
rect 41664 644458 42112 644486
rect 41664 644430 41692 644458
rect 42106 644446 42112 644458
rect 42164 644446 42170 644498
rect 41646 644378 41652 644430
rect 41704 644378 41710 644430
rect 42106 644310 42112 644362
rect 42164 644350 42170 644362
rect 42566 644350 42572 644362
rect 42164 644322 42572 644350
rect 42164 644310 42170 644322
rect 42566 644310 42572 644322
rect 42624 644310 42630 644362
rect 674790 641998 674796 642050
rect 674848 642038 674854 642050
rect 675250 642038 675256 642050
rect 674848 642010 675256 642038
rect 674848 641998 674854 642010
rect 675250 641998 675256 642010
rect 675308 641998 675314 642050
rect 674698 641182 674704 641234
rect 674756 641222 674762 641234
rect 674974 641222 674980 641234
rect 674756 641194 674980 641222
rect 674756 641182 674762 641194
rect 674974 641182 674980 641194
rect 675032 641182 675038 641234
rect 674790 638938 674796 638990
rect 674848 638978 674854 638990
rect 675250 638978 675256 638990
rect 674848 638950 675256 638978
rect 674848 638938 674854 638950
rect 675250 638938 675256 638950
rect 675308 638938 675314 638990
rect 674698 628330 674704 628382
rect 674756 628370 674762 628382
rect 674974 628370 674980 628382
rect 674756 628342 674980 628370
rect 674756 628330 674762 628342
rect 674974 628330 674980 628342
rect 675032 628330 675038 628382
rect 41554 627378 41560 627430
rect 41612 627418 41618 627430
rect 41738 627418 41744 627430
rect 41612 627390 41744 627418
rect 41612 627378 41618 627390
rect 41738 627378 41744 627390
rect 41796 627378 41802 627430
rect 674790 626358 674796 626410
rect 674848 626398 674854 626410
rect 675250 626398 675256 626410
rect 674848 626370 675256 626398
rect 674848 626358 674854 626370
rect 675250 626358 675256 626370
rect 675308 626358 675314 626410
rect 674790 615478 674796 615530
rect 674848 615518 674854 615530
rect 674974 615518 674980 615530
rect 674848 615490 674980 615518
rect 674848 615478 674854 615490
rect 674974 615478 674980 615490
rect 675032 615478 675038 615530
rect 42106 615410 42112 615462
rect 42164 615450 42170 615462
rect 42566 615450 42572 615462
rect 42164 615422 42572 615450
rect 42164 615410 42170 615422
rect 42566 615410 42572 615422
rect 42624 615410 42630 615462
rect 41646 612894 41652 612946
rect 41704 612934 41710 612946
rect 42566 612934 42572 612946
rect 41704 612906 42572 612934
rect 41704 612894 41710 612906
rect 42566 612894 42572 612906
rect 42624 612894 42630 612946
rect 675342 609018 675348 609070
rect 675400 609058 675406 609070
rect 675526 609058 675532 609070
rect 675400 609030 675532 609058
rect 675400 609018 675406 609030
rect 675526 609018 675532 609030
rect 675584 609018 675590 609070
rect 42106 608950 42112 609002
rect 42164 608990 42170 609002
rect 42566 608990 42572 609002
rect 42164 608962 42572 608990
rect 42164 608950 42170 608962
rect 42566 608950 42572 608962
rect 42624 608950 42630 609002
rect 674790 602558 674796 602610
rect 674848 602598 674854 602610
rect 674974 602598 674980 602610
rect 674848 602570 674980 602598
rect 674848 602558 674854 602570
rect 674974 602558 674980 602570
rect 675032 602558 675038 602610
rect 42106 599810 42112 599822
rect 41664 599782 42112 599810
rect 41554 599498 41560 599550
rect 41612 599538 41618 599550
rect 41664 599538 41692 599782
rect 42106 599770 42112 599782
rect 42164 599770 42170 599822
rect 41612 599510 41692 599538
rect 41612 599498 41618 599510
rect 674790 595486 674796 595538
rect 674848 595526 674854 595538
rect 675250 595526 675256 595538
rect 674848 595498 675256 595526
rect 674848 595486 674854 595498
rect 675250 595486 675256 595498
rect 675308 595486 675314 595538
rect 674422 595418 674428 595470
rect 674480 595458 674486 595470
rect 675158 595458 675164 595470
rect 674480 595430 675164 595458
rect 674480 595418 674486 595430
rect 675158 595418 675164 595430
rect 675216 595418 675222 595470
rect 674790 592358 674796 592410
rect 674848 592398 674854 592410
rect 675250 592398 675256 592410
rect 674848 592370 675256 592398
rect 674848 592358 674854 592370
rect 675250 592358 675256 592370
rect 675308 592358 675314 592410
rect 674698 587394 674704 587446
rect 674756 587434 674762 587446
rect 675250 587434 675256 587446
rect 674756 587406 675256 587434
rect 674756 587394 674762 587406
rect 675250 587394 675256 587406
rect 675308 587394 675314 587446
rect 674790 583450 674796 583502
rect 674848 583450 674854 583502
rect 674808 583354 674836 583450
rect 675250 583354 675256 583366
rect 674808 583326 675256 583354
rect 675250 583314 675256 583326
rect 675308 583314 675314 583366
rect 674790 580390 674796 580442
rect 674848 580430 674854 580442
rect 675250 580430 675256 580442
rect 674848 580402 675256 580430
rect 674848 580390 674854 580402
rect 675250 580390 675256 580402
rect 675308 580390 675314 580442
rect 674422 579778 674428 579830
rect 674480 579818 674486 579830
rect 675250 579818 675256 579830
rect 674480 579790 675256 579818
rect 674480 579778 674486 579790
rect 675250 579778 675256 579790
rect 675308 579778 675314 579830
rect 41554 579642 41560 579694
rect 41612 579682 41618 579694
rect 41830 579682 41836 579694
rect 41612 579654 41836 579682
rect 41612 579642 41618 579654
rect 41830 579642 41836 579654
rect 41888 579642 41894 579694
rect 41646 576786 41652 576838
rect 41704 576826 41710 576838
rect 42014 576826 42020 576838
rect 41704 576798 42020 576826
rect 41704 576786 41710 576798
rect 42014 576786 42020 576798
rect 42072 576786 42078 576838
rect 42106 571074 42112 571126
rect 42164 571114 42170 571126
rect 42566 571114 42572 571126
rect 42164 571086 42572 571114
rect 42164 571074 42170 571086
rect 42566 571074 42572 571086
rect 42624 571074 42630 571126
rect 677458 566722 677464 566774
rect 677516 566762 677522 566774
rect 677734 566762 677740 566774
rect 677516 566734 677740 566762
rect 677516 566722 677522 566734
rect 677734 566722 677740 566734
rect 677792 566722 677798 566774
rect 41646 559038 41652 559090
rect 41704 559078 41710 559090
rect 42566 559078 42572 559090
rect 41704 559050 42572 559078
rect 41704 559038 41710 559050
rect 42566 559038 42572 559050
rect 42624 559038 42630 559090
rect 675158 557406 675164 557458
rect 675216 557446 675222 557458
rect 675434 557446 675440 557458
rect 675216 557418 675440 557446
rect 675216 557406 675222 557418
rect 675434 557406 675440 557418
rect 675492 557406 675498 557458
rect 41738 551218 41744 551270
rect 41796 551258 41802 551270
rect 42106 551258 42112 551270
rect 41796 551230 42112 551258
rect 41796 551218 41802 551230
rect 42106 551218 42112 551230
rect 42164 551218 42170 551270
rect 674514 551082 674520 551134
rect 674572 551122 674578 551134
rect 674974 551122 674980 551134
rect 674572 551094 674980 551122
rect 674572 551082 674578 551094
rect 674974 551082 674980 551094
rect 675032 551082 675038 551134
rect 675158 551082 675164 551134
rect 675216 551122 675222 551134
rect 675342 551122 675348 551134
rect 675216 551094 675348 551122
rect 675216 551082 675222 551094
rect 675342 551082 675348 551094
rect 675400 551082 675406 551134
rect 674790 548838 674796 548890
rect 674848 548878 674854 548890
rect 675434 548878 675440 548890
rect 674848 548850 675440 548878
rect 674848 548838 674854 548850
rect 675434 548838 675440 548850
rect 675492 548838 675498 548890
rect 674974 548770 674980 548822
rect 675032 548810 675038 548822
rect 675250 548810 675256 548822
rect 675032 548782 675256 548810
rect 675032 548770 675038 548782
rect 675250 548770 675256 548782
rect 675308 548770 675314 548822
rect 674790 546662 674796 546714
rect 674848 546702 674854 546714
rect 675250 546702 675256 546714
rect 674848 546674 675256 546702
rect 674848 546662 674854 546674
rect 675250 546662 675256 546674
rect 675308 546662 675314 546714
rect 674974 546118 674980 546170
rect 675032 546158 675038 546170
rect 675342 546158 675348 546170
rect 675032 546130 675348 546158
rect 675032 546118 675038 546130
rect 675342 546118 675348 546130
rect 675400 546118 675406 546170
rect 674606 545098 674612 545150
rect 674664 545138 674670 545150
rect 675250 545138 675256 545150
rect 674664 545110 675256 545138
rect 674664 545098 674670 545110
rect 675250 545098 675256 545110
rect 675308 545098 675314 545150
rect 674974 541426 674980 541478
rect 675032 541466 675038 541478
rect 675158 541466 675164 541478
rect 675032 541438 675164 541466
rect 675032 541426 675038 541438
rect 675158 541426 675164 541438
rect 675216 541426 675222 541478
rect 674974 535646 674980 535698
rect 675032 535686 675038 535698
rect 675250 535686 675256 535698
rect 675032 535658 675256 535686
rect 675032 535646 675038 535658
rect 675250 535646 675256 535658
rect 675308 535646 675314 535698
rect 674514 535510 674520 535562
rect 674572 535550 674578 535562
rect 674974 535550 674980 535562
rect 674572 535522 674980 535550
rect 674572 535510 674578 535522
rect 674974 535510 674980 535522
rect 675032 535510 675038 535562
rect 674790 533198 674796 533250
rect 674848 533238 674854 533250
rect 675158 533238 675164 533250
rect 674848 533210 675164 533238
rect 674848 533198 674854 533210
rect 675158 533198 675164 533210
rect 675216 533198 675222 533250
rect 674606 533062 674612 533114
rect 674664 533102 674670 533114
rect 675250 533102 675256 533114
rect 674664 533074 675256 533102
rect 674664 533062 674670 533074
rect 675250 533062 675256 533074
rect 675308 533062 675314 533114
rect 674790 530818 674796 530870
rect 674848 530858 674854 530870
rect 674974 530858 674980 530870
rect 674848 530830 674980 530858
rect 674848 530818 674854 530830
rect 674974 530818 674980 530830
rect 675032 530818 675038 530870
rect 41738 526398 41744 526450
rect 41796 526438 41802 526450
rect 42566 526438 42572 526450
rect 41796 526410 42572 526438
rect 41796 526398 41802 526410
rect 42566 526398 42572 526410
rect 42624 526398 42630 526450
rect 41646 523882 41652 523934
rect 41704 523922 41710 523934
rect 42566 523922 42572 523934
rect 41704 523894 42572 523922
rect 41704 523882 41710 523894
rect 42566 523882 42572 523894
rect 42624 523882 42630 523934
rect 42106 518238 42112 518290
rect 42164 518278 42170 518290
rect 42566 518278 42572 518290
rect 42164 518250 42572 518278
rect 42164 518238 42170 518250
rect 42566 518238 42572 518250
rect 42624 518238 42630 518290
rect 674790 511506 674796 511558
rect 674848 511546 674854 511558
rect 674974 511546 674980 511558
rect 674848 511518 674980 511546
rect 674848 511506 674854 511518
rect 674974 511506 674980 511518
rect 675032 511506 675038 511558
rect 41646 499538 41652 499590
rect 41704 499578 41710 499590
rect 42106 499578 42112 499590
rect 41704 499550 42112 499578
rect 41704 499538 41710 499550
rect 42106 499538 42112 499550
rect 42164 499538 42170 499590
rect 674606 498586 674612 498638
rect 674664 498626 674670 498638
rect 674882 498626 674888 498638
rect 674664 498598 674888 498626
rect 674664 498586 674670 498598
rect 674882 498586 674888 498598
rect 674940 498586 674946 498638
rect 674790 498518 674796 498570
rect 674848 498558 674854 498570
rect 674974 498558 674980 498570
rect 674848 498530 674980 498558
rect 674848 498518 674854 498530
rect 674974 498518 674980 498530
rect 675032 498518 675038 498570
rect 674698 472814 674704 472866
rect 674756 472854 674762 472866
rect 674974 472854 674980 472866
rect 674756 472826 674980 472854
rect 674756 472814 674762 472826
rect 674974 472814 674980 472826
rect 675032 472814 675038 472866
rect 674698 454454 674704 454506
rect 674756 454494 674762 454506
rect 674882 454494 674888 454506
rect 674756 454466 674888 454494
rect 674756 454454 674762 454466
rect 674882 454454 674888 454466
rect 674940 454454 674946 454506
rect 675250 447042 675256 447094
rect 675308 447082 675314 447094
rect 677550 447082 677556 447094
rect 675308 447054 677556 447082
rect 675308 447042 675314 447054
rect 677550 447042 677556 447054
rect 677608 447042 677614 447094
rect 41830 441602 41836 441654
rect 41888 441642 41894 441654
rect 42014 441642 42020 441654
rect 41888 441614 42020 441642
rect 41888 441602 41894 441614
rect 42014 441602 42020 441614
rect 42072 441602 42078 441654
rect 39254 439766 39260 439818
rect 39312 439806 39318 439818
rect 44038 439806 44044 439818
rect 39312 439778 44044 439806
rect 39312 439766 39318 439778
rect 44038 439766 44044 439778
rect 44096 439806 44102 439818
rect 44866 439806 44872 439818
rect 44096 439778 44872 439806
rect 44096 439766 44102 439778
rect 44866 439766 44872 439778
rect 44924 439766 44930 439818
rect 675342 437930 675348 437982
rect 675400 437970 675406 437982
rect 677918 437970 677924 437982
rect 675400 437942 677924 437970
rect 675400 437930 675406 437942
rect 677918 437930 677924 437942
rect 677976 437930 677982 437982
rect 675342 430586 675348 430638
rect 675400 430586 675406 430638
rect 672398 430518 672404 430570
rect 672456 430558 672462 430570
rect 675360 430558 675388 430586
rect 672456 430530 675388 430558
rect 672456 430518 672462 430530
rect 39622 428546 39628 428598
rect 39680 428586 39686 428598
rect 41830 428586 41836 428598
rect 39680 428558 41836 428586
rect 39680 428546 39686 428558
rect 41830 428546 41836 428558
rect 41888 428586 41894 428598
rect 42014 428586 42020 428598
rect 41888 428558 42020 428586
rect 41888 428546 41894 428558
rect 42014 428546 42020 428558
rect 42072 428546 42078 428598
rect 41554 425010 41560 425062
rect 41612 425050 41618 425062
rect 42014 425050 42020 425062
rect 41612 425022 42020 425050
rect 41612 425010 41618 425022
rect 42014 425010 42020 425022
rect 42072 425010 42078 425062
rect 674882 425010 674888 425062
rect 674940 425050 674946 425062
rect 675066 425050 675072 425062
rect 674940 425022 675072 425050
rect 674940 425010 674946 425022
rect 675066 425010 675072 425022
rect 675124 425010 675130 425062
rect 672398 423282 672404 423294
rect 669656 423254 672404 423282
rect 668626 423174 668632 423226
rect 668684 423214 668690 423226
rect 669656 423214 669684 423254
rect 672398 423242 672404 423254
rect 672456 423242 672462 423294
rect 668684 423186 669684 423214
rect 668684 423174 668690 423186
rect 41554 412158 41560 412210
rect 41612 412198 41618 412210
rect 41830 412198 41836 412210
rect 41612 412170 41836 412198
rect 41612 412158 41618 412170
rect 41830 412158 41836 412170
rect 41888 412158 41894 412210
rect 664670 408486 664676 408538
rect 664728 408526 664734 408538
rect 668626 408526 668632 408538
rect 664728 408498 668632 408526
rect 664728 408486 664734 408498
rect 668626 408486 668632 408498
rect 668684 408486 668690 408538
rect 663106 404814 663112 404866
rect 663164 404854 663170 404866
rect 664670 404854 664676 404866
rect 663164 404826 664676 404854
rect 663164 404814 663170 404826
rect 664670 404814 664676 404826
rect 664728 404814 664734 404866
rect 41830 399238 41836 399290
rect 41888 399278 41894 399290
rect 42290 399278 42296 399290
rect 41888 399250 42296 399278
rect 41888 399238 41894 399250
rect 42290 399238 42296 399250
rect 42348 399238 42354 399290
rect 41646 394886 41652 394938
rect 41704 394926 41710 394938
rect 42382 394926 42388 394938
rect 41704 394898 42388 394926
rect 41704 394886 41710 394898
rect 42382 394886 42388 394898
rect 42440 394886 42446 394938
rect 41738 394818 41744 394870
rect 41796 394858 41802 394870
rect 42474 394858 42480 394870
rect 41796 394830 42480 394858
rect 41796 394818 41802 394830
rect 42474 394818 42480 394830
rect 42532 394818 42538 394870
rect 41646 394138 41652 394190
rect 41704 394178 41710 394190
rect 42106 394178 42112 394190
rect 41704 394150 42112 394178
rect 41704 394138 41710 394150
rect 42106 394138 42112 394150
rect 42164 394138 42170 394190
rect 41646 392710 41652 392762
rect 41704 392750 41710 392762
rect 42382 392750 42388 392762
rect 41704 392722 42388 392750
rect 41704 392710 41710 392722
rect 42382 392710 42388 392722
rect 42440 392710 42446 392762
rect 41646 387202 41652 387254
rect 41704 387242 41710 387254
rect 42106 387242 42112 387254
rect 41704 387214 42112 387242
rect 41704 387202 41710 387214
rect 42106 387202 42112 387214
rect 42164 387202 42170 387254
rect 42106 386726 42112 386778
rect 42164 386766 42170 386778
rect 42474 386766 42480 386778
rect 42164 386738 42480 386766
rect 42164 386726 42170 386738
rect 42474 386726 42480 386738
rect 42532 386726 42538 386778
rect 41646 381830 41652 381882
rect 41704 381870 41710 381882
rect 42106 381870 42112 381882
rect 41704 381842 42112 381870
rect 41704 381830 41710 381842
rect 42106 381830 42112 381842
rect 42164 381870 42170 381882
rect 42290 381870 42296 381882
rect 42164 381842 42296 381870
rect 42164 381830 42170 381842
rect 42290 381830 42296 381842
rect 42348 381830 42354 381882
rect 41646 379178 41652 379230
rect 41704 379218 41710 379230
rect 42106 379218 42112 379230
rect 41704 379190 42112 379218
rect 41704 379178 41710 379190
rect 42106 379178 42112 379190
rect 42164 379178 42170 379230
rect 42014 374350 42020 374402
rect 42072 374390 42078 374402
rect 42382 374390 42388 374402
rect 42072 374362 42388 374390
rect 42072 374350 42078 374362
rect 42382 374350 42388 374362
rect 42440 374350 42446 374402
rect 675158 365714 675164 365766
rect 675216 365714 675222 365766
rect 675176 365562 675204 365714
rect 675158 365510 675164 365562
rect 675216 365510 675222 365562
rect 42014 364354 42020 364406
rect 42072 364354 42078 364406
rect 42032 364270 42060 364354
rect 42014 364218 42020 364270
rect 42072 364218 42078 364270
rect 675066 362926 675072 362978
rect 675124 362966 675130 362978
rect 675250 362966 675256 362978
rect 675124 362938 675256 362966
rect 675124 362926 675130 362938
rect 675250 362926 675256 362938
rect 675308 362926 675314 362978
rect 675158 362042 675164 362094
rect 675216 362042 675222 362094
rect 675176 361890 675204 362042
rect 675158 361838 675164 361890
rect 675216 361838 675222 361890
rect 660438 358982 660444 359034
rect 660496 359022 660502 359034
rect 663106 359022 663112 359034
rect 660496 358994 663112 359022
rect 660496 358982 660502 358994
rect 663106 358982 663112 358994
rect 663164 358982 663170 359034
rect 674882 357554 674888 357606
rect 674940 357594 674946 357606
rect 675250 357594 675256 357606
rect 674940 357566 675256 357594
rect 674940 357554 674946 357566
rect 675250 357554 675256 357566
rect 675308 357554 675314 357606
rect 675066 357146 675072 357198
rect 675124 357146 675130 357198
rect 675084 356982 675112 357146
rect 675158 356982 675164 356994
rect 675084 356954 675164 356982
rect 675158 356942 675164 356954
rect 675216 356942 675222 356994
rect 674790 356874 674796 356926
rect 674848 356914 674854 356926
rect 675066 356914 675072 356926
rect 674848 356886 675072 356914
rect 674848 356874 674854 356886
rect 675066 356874 675072 356886
rect 675124 356874 675130 356926
rect 42014 352182 42020 352234
rect 42072 352222 42078 352234
rect 42382 352222 42388 352234
rect 42072 352194 42388 352222
rect 42072 352182 42078 352194
rect 42382 352182 42388 352194
rect 42440 352182 42446 352234
rect 41646 350278 41652 350330
rect 41704 350318 41710 350330
rect 42106 350318 42112 350330
rect 41704 350290 42112 350318
rect 41704 350278 41710 350290
rect 42106 350278 42112 350290
rect 42164 350278 42170 350330
rect 41738 350210 41744 350262
rect 41796 350250 41802 350262
rect 42566 350250 42572 350262
rect 41796 350222 42572 350250
rect 41796 350210 41802 350222
rect 42566 350210 42572 350222
rect 42624 350210 42630 350262
rect 657126 350006 657132 350058
rect 657184 350046 657190 350058
rect 660346 350046 660352 350058
rect 657184 350018 660352 350046
rect 657184 350006 657190 350018
rect 660346 350006 660352 350018
rect 660404 350006 660410 350058
rect 674974 349938 674980 349990
rect 675032 349978 675038 349990
rect 675342 349978 675348 349990
rect 675032 349950 675348 349978
rect 675032 349938 675038 349950
rect 675342 349938 675348 349950
rect 675400 349938 675406 349990
rect 674790 349870 674796 349922
rect 674848 349910 674854 349922
rect 675250 349910 675256 349922
rect 674848 349882 675256 349910
rect 674848 349870 674854 349882
rect 675250 349870 675256 349882
rect 675308 349870 675314 349922
rect 41646 349530 41652 349582
rect 41704 349570 41710 349582
rect 42290 349570 42296 349582
rect 41704 349542 42296 349570
rect 41704 349530 41710 349542
rect 42290 349530 42296 349542
rect 42348 349530 42354 349582
rect 41830 348646 41836 348698
rect 41888 348686 41894 348698
rect 42382 348686 42388 348698
rect 41888 348658 42388 348686
rect 41888 348646 41894 348658
rect 42382 348646 42388 348658
rect 42440 348646 42446 348698
rect 41830 347694 41836 347746
rect 41888 347734 41894 347746
rect 42382 347734 42388 347746
rect 41888 347706 42388 347734
rect 41888 347694 41894 347706
rect 42382 347694 42388 347706
rect 42440 347694 42446 347746
rect 655746 344770 655752 344822
rect 655804 344810 655810 344822
rect 657126 344810 657132 344822
rect 655804 344782 657132 344810
rect 655804 344770 655810 344782
rect 657126 344770 657132 344782
rect 657184 344770 657190 344822
rect 42106 344566 42112 344618
rect 42164 344606 42170 344618
rect 42474 344606 42480 344618
rect 42164 344578 42480 344606
rect 42164 344566 42170 344578
rect 42474 344566 42480 344578
rect 42532 344566 42538 344618
rect 42106 344430 42112 344482
rect 42164 344470 42170 344482
rect 42290 344470 42296 344482
rect 42164 344442 42296 344470
rect 42164 344430 42170 344442
rect 42290 344430 42296 344442
rect 42348 344430 42354 344482
rect 42382 344198 42388 344210
rect 42124 344170 42388 344198
rect 42124 343994 42152 344170
rect 42382 344158 42388 344170
rect 42440 344158 42446 344210
rect 42382 343994 42388 344006
rect 42124 343966 42388 343994
rect 42382 343954 42388 343966
rect 42440 343954 42446 344006
rect 41646 338242 41652 338294
rect 41704 338282 41710 338294
rect 42106 338282 42112 338294
rect 41704 338254 42112 338282
rect 41704 338242 41710 338254
rect 42106 338242 42112 338254
rect 42164 338282 42170 338294
rect 42474 338282 42480 338294
rect 42164 338254 42480 338282
rect 42164 338242 42170 338254
rect 42474 338242 42480 338254
rect 42532 338242 42538 338294
rect 41646 337630 41652 337682
rect 41704 337670 41710 337682
rect 42566 337670 42572 337682
rect 41704 337642 42572 337670
rect 41704 337630 41710 337642
rect 42566 337630 42572 337642
rect 42624 337630 42630 337682
rect 41830 335114 41836 335166
rect 41888 335154 41894 335166
rect 42566 335154 42572 335166
rect 41888 335126 42572 335154
rect 41888 335114 41894 335126
rect 42566 335114 42572 335126
rect 42624 335114 42630 335166
rect 41830 334842 41836 334894
rect 41888 334842 41894 334894
rect 41646 334570 41652 334622
rect 41704 334610 41710 334622
rect 41848 334610 41876 334842
rect 41704 334582 41876 334610
rect 41704 334570 41710 334582
rect 42106 334366 42112 334418
rect 42164 334406 42170 334418
rect 42382 334406 42388 334418
rect 42164 334378 42388 334406
rect 42164 334366 42170 334378
rect 42382 334366 42388 334378
rect 42440 334366 42446 334418
rect 41646 333958 41652 334010
rect 41704 333998 41710 334010
rect 42014 333998 42020 334010
rect 41704 333970 42020 333998
rect 41704 333958 41710 333970
rect 42014 333958 42020 333970
rect 42072 333958 42078 334010
rect 655746 331278 655752 331290
rect 653096 331250 655752 331278
rect 651238 331170 651244 331222
rect 651296 331210 651302 331222
rect 653096 331210 653124 331250
rect 655746 331238 655752 331250
rect 655804 331238 655810 331290
rect 651296 331182 653124 331210
rect 651296 331170 651302 331182
rect 649398 319338 649404 319390
rect 649456 319378 649462 319390
rect 651238 319378 651244 319390
rect 649456 319350 651244 319378
rect 649456 319338 649462 319350
rect 651238 319338 651244 319350
rect 651296 319338 651302 319390
rect 675158 319066 675164 319118
rect 675216 319066 675222 319118
rect 675176 318914 675204 319066
rect 675158 318862 675164 318914
rect 675216 318862 675222 318914
rect 675066 316346 675072 316398
rect 675124 316386 675130 316398
rect 675250 316386 675256 316398
rect 675124 316358 675256 316386
rect 675124 316346 675130 316358
rect 675250 316346 675256 316358
rect 675308 316346 675314 316398
rect 640842 313830 640848 313882
rect 640900 313870 640906 313882
rect 649398 313870 649404 313882
rect 640900 313842 649404 313870
rect 640900 313830 640906 313842
rect 649398 313830 649404 313842
rect 649456 313830 649462 313882
rect 41554 312810 41560 312862
rect 41612 312850 41618 312862
rect 41738 312850 41744 312862
rect 41612 312822 41744 312850
rect 41612 312810 41618 312822
rect 41738 312810 41744 312822
rect 41796 312810 41802 312862
rect 41922 312810 41928 312862
rect 41980 312810 41986 312862
rect 41940 312782 41968 312810
rect 42014 312782 42020 312794
rect 41940 312754 42020 312782
rect 42014 312742 42020 312754
rect 42072 312742 42078 312794
rect 636886 310226 636892 310278
rect 636944 310266 636950 310278
rect 640842 310266 640848 310278
rect 636944 310238 640848 310266
rect 636944 310226 636950 310238
rect 640842 310226 640848 310238
rect 640900 310226 640906 310278
rect 41922 309138 41928 309190
rect 41980 309178 41986 309190
rect 42014 309178 42020 309190
rect 41980 309150 42020 309178
rect 41980 309138 41986 309150
rect 42014 309138 42020 309150
rect 42072 309138 42078 309190
rect 674882 309070 674888 309122
rect 674940 309110 674946 309122
rect 675066 309110 675072 309122
rect 674940 309082 675072 309110
rect 674940 309070 674946 309082
rect 675066 309070 675072 309082
rect 675124 309070 675130 309122
rect 634678 306418 634684 306470
rect 634736 306458 634742 306470
rect 636886 306458 636892 306470
rect 634736 306430 636892 306458
rect 634736 306418 634742 306430
rect 636886 306418 636892 306430
rect 636944 306418 636950 306470
rect 41922 305874 41928 305926
rect 41980 305914 41986 305926
rect 42382 305914 42388 305926
rect 41980 305886 42388 305914
rect 41980 305874 41986 305886
rect 42382 305874 42388 305886
rect 42440 305874 42446 305926
rect 42106 305330 42112 305382
rect 42164 305370 42170 305382
rect 42290 305370 42296 305382
rect 42164 305342 42296 305370
rect 42164 305330 42170 305342
rect 42290 305330 42296 305342
rect 42348 305330 42354 305382
rect 41830 305126 41836 305178
rect 41888 305166 41894 305178
rect 42106 305166 42112 305178
rect 41888 305138 42112 305166
rect 41888 305126 41894 305138
rect 42106 305126 42112 305138
rect 42164 305126 42170 305178
rect 674974 304922 674980 304974
rect 675032 304962 675038 304974
rect 675250 304962 675256 304974
rect 675032 304934 675256 304962
rect 675032 304922 675038 304934
rect 675250 304922 675256 304934
rect 675308 304922 675314 304974
rect 674974 303358 674980 303410
rect 675032 303398 675038 303410
rect 675434 303398 675440 303410
rect 675032 303370 675440 303398
rect 675032 303358 675038 303370
rect 675434 303358 675440 303370
rect 675492 303358 675498 303410
rect 41646 303290 41652 303342
rect 41704 303330 41710 303342
rect 42382 303330 42388 303342
rect 41704 303302 42388 303330
rect 41704 303290 41710 303302
rect 42382 303290 42388 303302
rect 42440 303290 42446 303342
rect 634678 299998 634684 300010
rect 632856 299970 634684 299998
rect 630354 299890 630360 299942
rect 630412 299930 630418 299942
rect 632856 299930 632884 299970
rect 634678 299958 634684 299970
rect 634736 299958 634742 300010
rect 630412 299902 632884 299930
rect 630412 299890 630418 299902
rect 674882 296218 674888 296270
rect 674940 296258 674946 296270
rect 675342 296258 675348 296270
rect 674940 296230 675348 296258
rect 674940 296218 674946 296230
rect 675342 296218 675348 296230
rect 675400 296218 675406 296270
rect 630354 294422 630360 294434
rect 625496 294394 630360 294422
rect 620694 294246 620700 294298
rect 620752 294286 620758 294298
rect 625496 294286 625524 294394
rect 630354 294382 630360 294394
rect 630412 294382 630418 294434
rect 620752 294258 625524 294286
rect 620752 294246 620758 294258
rect 41646 293566 41652 293618
rect 41704 293606 41710 293618
rect 42106 293606 42112 293618
rect 41704 293578 42112 293606
rect 41704 293566 41710 293578
rect 42106 293566 42112 293578
rect 42164 293566 42170 293618
rect 42106 293430 42112 293482
rect 42164 293470 42170 293482
rect 42382 293470 42388 293482
rect 42164 293442 42388 293470
rect 42164 293430 42170 293442
rect 42382 293430 42388 293442
rect 42440 293430 42446 293482
rect 41922 287378 41928 287430
rect 41980 287418 41986 287430
rect 42106 287418 42112 287430
rect 41980 287390 42112 287418
rect 41980 287378 41986 287390
rect 42106 287378 42112 287390
rect 42164 287378 42170 287430
rect 615542 286290 615548 286342
rect 615600 286330 615606 286342
rect 620694 286330 620700 286342
rect 615600 286302 620700 286330
rect 615600 286290 615606 286302
rect 620694 286290 620700 286302
rect 620752 286290 620758 286342
rect 613426 284114 613432 284166
rect 613484 284154 613490 284166
rect 615542 284154 615548 284166
rect 613484 284126 615548 284154
rect 613484 284114 613490 284126
rect 615542 284114 615548 284126
rect 615600 284114 615606 284166
rect 613426 276062 613432 276074
rect 610776 276034 613432 276062
rect 609746 275954 609752 276006
rect 609804 275994 609810 276006
rect 610776 275994 610804 276034
rect 613426 276022 613432 276034
rect 613484 276022 613490 276074
rect 609804 275966 610804 275994
rect 609804 275954 609810 275966
rect 674790 274118 674796 274170
rect 674848 274158 674854 274170
rect 675158 274158 675164 274170
rect 674848 274130 675164 274158
rect 674848 274118 674854 274130
rect 675158 274118 675164 274130
rect 675216 274118 675222 274170
rect 675158 272554 675164 272606
rect 675216 272594 675222 272606
rect 675434 272594 675440 272606
rect 675216 272566 675440 272594
rect 675216 272554 675222 272566
rect 675434 272554 675440 272566
rect 675492 272554 675498 272606
rect 675526 270718 675532 270770
rect 675584 270718 675590 270770
rect 675434 270514 675440 270566
rect 675492 270554 675498 270566
rect 675544 270554 675572 270718
rect 675492 270526 675572 270554
rect 675492 270514 675498 270526
rect 674974 269562 674980 269614
rect 675032 269602 675038 269614
rect 675250 269602 675256 269614
rect 675032 269574 675256 269602
rect 675032 269562 675038 269574
rect 675250 269562 675256 269574
rect 675308 269562 675314 269614
rect 674790 268882 674796 268934
rect 674848 268922 674854 268934
rect 675250 268922 675256 268934
rect 674848 268894 675256 268922
rect 674848 268882 674854 268894
rect 675250 268882 675256 268894
rect 675308 268882 675314 268934
rect 42106 266706 42112 266758
rect 42164 266746 42170 266758
rect 42382 266746 42388 266758
rect 42164 266718 42388 266746
rect 42164 266706 42170 266718
rect 42382 266706 42388 266718
rect 42440 266706 42446 266758
rect 41646 266570 41652 266622
rect 41704 266610 41710 266622
rect 42106 266610 42112 266622
rect 41704 266582 42112 266610
rect 41704 266570 41710 266582
rect 42106 266570 42112 266582
rect 42164 266570 42170 266622
rect 605330 264938 605336 264990
rect 605388 264978 605394 264990
rect 609746 264978 609752 264990
rect 605388 264950 609752 264978
rect 605388 264938 605394 264950
rect 609746 264938 609752 264950
rect 609804 264938 609810 264990
rect 674882 264666 674888 264718
rect 674940 264706 674946 264718
rect 675158 264706 675164 264718
rect 674940 264678 675164 264706
rect 674940 264666 674946 264678
rect 675158 264666 675164 264678
rect 675216 264666 675222 264718
rect 600546 262150 600552 262202
rect 600604 262190 600610 262202
rect 605330 262190 605336 262202
rect 600604 262162 605336 262190
rect 600604 262150 600610 262162
rect 605330 262150 605336 262162
rect 605388 262150 605394 262202
rect 41738 261266 41744 261318
rect 41796 261306 41802 261318
rect 42658 261306 42664 261318
rect 41796 261278 42664 261306
rect 41796 261266 41802 261278
rect 42658 261266 42664 261278
rect 42716 261266 42722 261318
rect 41646 260518 41652 260570
rect 41704 260558 41710 260570
rect 42290 260558 42296 260570
rect 41704 260530 42296 260558
rect 41704 260518 41710 260530
rect 42290 260518 42296 260530
rect 42348 260518 42354 260570
rect 41646 259634 41652 259686
rect 41704 259674 41710 259686
rect 42382 259674 42388 259686
rect 41704 259646 42388 259674
rect 41704 259634 41710 259646
rect 42382 259634 42388 259646
rect 42440 259634 42446 259686
rect 675158 259498 675164 259550
rect 675216 259498 675222 259550
rect 675176 259346 675204 259498
rect 675158 259294 675164 259346
rect 675216 259294 675222 259346
rect 674882 259226 674888 259278
rect 674940 259266 674946 259278
rect 675250 259266 675256 259278
rect 674940 259238 675256 259266
rect 674940 259226 674946 259238
rect 675250 259226 675256 259238
rect 675308 259226 675314 259278
rect 674882 257594 674888 257646
rect 674940 257634 674946 257646
rect 675342 257634 675348 257646
rect 674940 257606 675348 257634
rect 674940 257594 674946 257606
rect 675342 257594 675348 257606
rect 675400 257594 675406 257646
rect 675342 257186 675348 257238
rect 675400 257226 675406 257238
rect 675400 257198 675572 257226
rect 675400 257186 675406 257198
rect 674974 257050 674980 257102
rect 675032 257050 675038 257102
rect 674992 257022 675020 257050
rect 675544 257034 675572 257198
rect 675342 257022 675348 257034
rect 674992 256994 675348 257022
rect 675342 256982 675348 256994
rect 675400 256982 675406 257034
rect 675526 256982 675532 257034
rect 675584 256982 675590 257034
rect 42290 254166 42296 254178
rect 41664 254138 42296 254166
rect 41664 253634 41692 254138
rect 42290 254126 42296 254138
rect 42348 254126 42354 254178
rect 42382 254098 42388 254110
rect 42124 254070 42388 254098
rect 42124 253894 42152 254070
rect 42382 254058 42388 254070
rect 42440 254058 42446 254110
rect 42290 253922 42296 253974
rect 42348 253962 42354 253974
rect 42658 253962 42664 253974
rect 42348 253934 42664 253962
rect 42348 253922 42354 253934
rect 42658 253922 42664 253934
rect 42716 253922 42722 253974
rect 42382 253894 42388 253906
rect 42124 253866 42388 253894
rect 42382 253854 42388 253866
rect 42440 253854 42446 253906
rect 41646 253582 41652 253634
rect 41704 253582 41710 253634
rect 600546 248454 600552 248466
rect 597896 248426 600552 248454
rect 594106 248346 594112 248398
rect 594164 248386 594170 248398
rect 597896 248386 597924 248426
rect 600546 248414 600552 248426
rect 600604 248414 600610 248466
rect 594164 248358 597924 248386
rect 594164 248346 594170 248358
rect 41922 245558 41928 245610
rect 41980 245598 41986 245610
rect 42382 245598 42388 245610
rect 41980 245570 42388 245598
rect 41980 245558 41986 245570
rect 42382 245558 42388 245570
rect 42440 245558 42446 245610
rect 41646 245490 41652 245542
rect 41704 245530 41710 245542
rect 42106 245530 42112 245542
rect 41704 245502 42112 245530
rect 41704 245490 41710 245502
rect 42106 245490 42112 245502
rect 42164 245490 42170 245542
rect 594106 242946 594112 242958
rect 590536 242918 594112 242946
rect 590426 242838 590432 242890
rect 590484 242878 590490 242890
rect 590536 242878 590564 242918
rect 594106 242906 594112 242918
rect 594164 242906 594170 242958
rect 590484 242850 590564 242878
rect 590484 242838 590490 242850
rect 675158 241002 675164 241054
rect 675216 241042 675222 241054
rect 675434 241042 675440 241054
rect 675216 241014 675440 241042
rect 675216 241002 675222 241014
rect 675434 241002 675440 241014
rect 675492 241002 675498 241054
rect 587666 234882 587672 234934
rect 587724 234922 587730 234934
rect 590426 234922 590432 234934
rect 587724 234894 590432 234922
rect 587724 234882 587730 234894
rect 590426 234882 590432 234894
rect 590484 234882 590490 234934
rect 41922 228150 41928 228202
rect 41980 228190 41986 228202
rect 42106 228190 42112 228202
rect 41980 228162 42112 228190
rect 41980 228150 41986 228162
rect 42106 228150 42112 228162
rect 42164 228150 42170 228202
rect 674974 226042 674980 226094
rect 675032 226082 675038 226094
rect 675434 226082 675440 226094
rect 675032 226054 675440 226082
rect 675032 226042 675038 226054
rect 675434 226042 675440 226054
rect 675492 226042 675498 226094
rect 674882 225974 674888 226026
rect 674940 226014 674946 226026
rect 675526 226014 675532 226026
rect 674940 225986 675532 226014
rect 674940 225974 674946 225986
rect 675526 225974 675532 225986
rect 675584 225974 675590 226026
rect 674974 223322 674980 223374
rect 675032 223362 675038 223374
rect 675342 223362 675348 223374
rect 675032 223334 675348 223362
rect 675032 223322 675038 223334
rect 675342 223322 675348 223334
rect 675400 223322 675406 223374
rect 675250 222954 675256 222966
rect 675176 222926 675256 222954
rect 675176 222694 675204 222926
rect 675250 222914 675256 222926
rect 675308 222914 675314 222966
rect 675158 222642 675164 222694
rect 675216 222642 675222 222694
rect 585826 221418 585832 221470
rect 585884 221458 585890 221470
rect 587666 221458 587672 221470
rect 585884 221430 587672 221458
rect 585884 221418 585890 221430
rect 587666 221418 587672 221430
rect 587724 221418 587730 221470
rect 42106 216658 42112 216710
rect 42164 216698 42170 216710
rect 42474 216698 42480 216710
rect 42164 216670 42480 216698
rect 42164 216658 42170 216670
rect 42474 216658 42480 216670
rect 42532 216658 42538 216710
rect 41646 215978 41652 216030
rect 41704 216018 41710 216030
rect 42290 216018 42296 216030
rect 41704 215990 42296 216018
rect 41704 215978 41710 215990
rect 42290 215978 42296 215990
rect 42348 215978 42354 216030
rect 42474 215270 42480 215282
rect 41664 215242 42480 215270
rect 41664 215146 41692 215242
rect 42474 215230 42480 215242
rect 42532 215230 42538 215282
rect 42106 215162 42112 215214
rect 42164 215202 42170 215214
rect 42382 215202 42388 215214
rect 42164 215174 42388 215202
rect 42164 215162 42170 215174
rect 42382 215162 42388 215174
rect 42440 215162 42446 215214
rect 41646 215094 41652 215146
rect 41704 215094 41710 215146
rect 674882 210334 674888 210386
rect 674940 210374 674946 210386
rect 675250 210374 675256 210386
rect 674940 210346 675256 210374
rect 674940 210334 674946 210346
rect 675250 210334 675256 210346
rect 675308 210334 675314 210386
rect 674974 210198 674980 210250
rect 675032 210238 675038 210250
rect 675342 210238 675348 210250
rect 675032 210210 675348 210238
rect 675032 210198 675038 210210
rect 675342 210198 675348 210210
rect 675400 210198 675406 210250
rect 42106 209762 42112 209774
rect 41664 209734 42112 209762
rect 41664 209570 41692 209734
rect 42106 209722 42112 209734
rect 42164 209722 42170 209774
rect 41646 209518 41652 209570
rect 41704 209518 41710 209570
rect 41646 208974 41652 209026
rect 41704 209014 41710 209026
rect 42290 209014 42296 209026
rect 41704 208986 42296 209014
rect 41704 208974 41710 208986
rect 42290 208974 42296 208986
rect 42348 208974 42354 209026
rect 585826 206158 585832 206170
rect 583636 206130 585832 206158
rect 581502 206050 581508 206102
rect 581560 206090 581566 206102
rect 583636 206090 583664 206130
rect 585826 206118 585832 206130
rect 585884 206118 585890 206170
rect 581560 206062 583664 206090
rect 581560 206050 581566 206062
rect 41646 203058 41652 203110
rect 41704 203098 41710 203110
rect 42382 203098 42388 203110
rect 41704 203070 42388 203098
rect 41704 203058 41710 203070
rect 42382 203058 42388 203070
rect 42440 203058 42446 203110
rect 578098 200610 578104 200662
rect 578156 200650 578162 200662
rect 581502 200650 581508 200662
rect 578156 200622 581508 200650
rect 578156 200610 578162 200622
rect 581502 200610 581508 200622
rect 581560 200610 581566 200662
rect 573958 198706 573964 198758
rect 574016 198746 574022 198758
rect 578098 198746 578104 198758
rect 574016 198718 578104 198746
rect 574016 198706 574022 198718
rect 578098 198706 578104 198718
rect 578156 198706 578162 198758
rect 41830 193198 41836 193250
rect 41888 193238 41894 193250
rect 42382 193238 42388 193250
rect 41888 193210 42388 193238
rect 41888 193198 41894 193210
rect 42382 193198 42388 193210
rect 42440 193198 42446 193250
rect 570646 191906 570652 191958
rect 570704 191946 570710 191958
rect 573958 191946 573964 191958
rect 570704 191918 573964 191946
rect 570704 191906 570710 191918
rect 573958 191906 573964 191918
rect 574016 191906 574022 191958
rect 675158 189390 675164 189442
rect 675216 189430 675222 189442
rect 675342 189430 675348 189442
rect 675216 189402 675348 189430
rect 675216 189390 675222 189402
rect 675342 189390 675348 189402
rect 675400 189390 675406 189442
rect 566598 187690 566604 187742
rect 566656 187730 566662 187742
rect 570646 187730 570652 187742
rect 566656 187702 570652 187730
rect 566656 187690 566662 187702
rect 570646 187690 570652 187702
rect 570704 187690 570710 187742
rect 41830 184018 41836 184070
rect 41888 184018 41894 184070
rect 41848 183922 41876 184018
rect 41922 183922 41928 183934
rect 41848 183894 41928 183922
rect 41922 183882 41928 183894
rect 41980 183882 41986 183934
rect 674974 179802 674980 179854
rect 675032 179842 675038 179854
rect 675618 179842 675624 179854
rect 675032 179814 675624 179842
rect 675032 179802 675038 179814
rect 675618 179802 675624 179814
rect 675676 179802 675682 179854
rect 675158 179666 675164 179718
rect 675216 179706 675222 179718
rect 675710 179706 675716 179718
rect 675216 179678 675716 179706
rect 675216 179666 675222 179678
rect 675710 179666 675716 179678
rect 675768 179666 675774 179718
rect 555006 178510 555012 178562
rect 555064 178550 555070 178562
rect 566506 178550 566512 178562
rect 555064 178522 566512 178550
rect 555064 178510 555070 178522
rect 566506 178510 566512 178522
rect 566564 178510 566570 178562
rect 675066 176742 675072 176794
rect 675124 176782 675130 176794
rect 675342 176782 675348 176794
rect 675124 176754 675348 176782
rect 675124 176742 675130 176754
rect 675342 176742 675348 176754
rect 675400 176742 675406 176794
rect 674882 175654 674888 175706
rect 674940 175694 674946 175706
rect 675250 175694 675256 175706
rect 674940 175666 675256 175694
rect 674940 175654 674946 175666
rect 675250 175654 675256 175666
rect 675308 175654 675314 175706
rect 41922 172254 41928 172306
rect 41980 172294 41986 172306
rect 42382 172294 42388 172306
rect 41980 172266 42388 172294
rect 41980 172254 41986 172266
rect 42382 172254 42388 172266
rect 42440 172254 42446 172306
rect 41646 172186 41652 172238
rect 41704 172226 41710 172238
rect 42290 172226 42296 172238
rect 41704 172198 42296 172226
rect 41704 172186 41710 172198
rect 42290 172186 42296 172198
rect 42348 172186 42354 172238
rect 552154 167562 552160 167614
rect 552212 167602 552218 167614
rect 555006 167602 555012 167614
rect 552212 167574 555012 167602
rect 552212 167562 552218 167574
rect 555006 167562 555012 167574
rect 555064 167562 555070 167614
rect 674790 167358 674796 167410
rect 674848 167398 674854 167410
rect 674974 167398 674980 167410
rect 674848 167370 674980 167398
rect 674848 167358 674854 167370
rect 674974 167358 674980 167370
rect 675032 167358 675038 167410
rect 674790 165318 674796 165370
rect 674848 165358 674854 165370
rect 675250 165358 675256 165370
rect 674848 165330 675256 165358
rect 674848 165318 674854 165330
rect 675250 165318 675256 165330
rect 675308 165318 675314 165370
rect 550038 164842 550044 164894
rect 550096 164882 550102 164894
rect 552154 164882 552160 164894
rect 550096 164854 552160 164882
rect 550096 164842 550102 164854
rect 552154 164842 552160 164854
rect 552212 164842 552218 164894
rect 42290 164134 42296 164146
rect 42124 164106 42296 164134
rect 42124 164066 42152 164106
rect 42290 164094 42296 164106
rect 42348 164094 42354 164146
rect 42032 164038 42152 164066
rect 42032 164010 42060 164038
rect 42014 163958 42020 164010
rect 42072 163958 42078 164010
rect 674882 163754 674888 163806
rect 674940 163794 674946 163806
rect 675342 163794 675348 163806
rect 674940 163766 675348 163794
rect 674940 163754 674946 163766
rect 675342 163754 675348 163766
rect 675400 163754 675406 163806
rect 41646 158994 41652 159046
rect 41704 159034 41710 159046
rect 42290 159034 42296 159046
rect 41704 159006 42296 159034
rect 41704 158994 41710 159006
rect 42290 158994 42296 159006
rect 42348 158994 42354 159046
rect 675158 157294 675164 157346
rect 675216 157334 675222 157346
rect 675434 157334 675440 157346
rect 675216 157306 675440 157334
rect 675216 157294 675222 157306
rect 675434 157294 675440 157306
rect 675492 157294 675498 157346
rect 674790 157158 674796 157210
rect 674848 157198 674854 157210
rect 675158 157198 675164 157210
rect 674848 157170 675164 157198
rect 674848 157158 674854 157170
rect 675158 157158 675164 157170
rect 675216 157158 675222 157210
rect 546358 155730 546364 155782
rect 546416 155770 546422 155782
rect 550038 155770 550044 155782
rect 546416 155742 550044 155770
rect 546416 155730 546422 155742
rect 550038 155730 550044 155742
rect 550096 155730 550102 155782
rect 42290 155458 42296 155510
rect 42348 155498 42354 155510
rect 87186 155498 87192 155510
rect 42348 155470 87192 155498
rect 42348 155458 42354 155470
rect 87186 155458 87192 155470
rect 87244 155458 87250 155510
rect 42474 154574 42480 154626
rect 42532 154614 42538 154626
rect 42566 154614 42572 154626
rect 42532 154586 42572 154614
rect 42532 154574 42538 154586
rect 42566 154574 42572 154586
rect 42624 154574 42630 154626
rect 42290 154438 42296 154490
rect 42348 154478 42354 154490
rect 42474 154478 42480 154490
rect 42348 154450 42480 154478
rect 42348 154438 42354 154450
rect 42474 154438 42480 154450
rect 42532 154438 42538 154490
rect 542678 151786 542684 151838
rect 542736 151826 542742 151838
rect 546358 151826 546364 151838
rect 542736 151798 546364 151826
rect 542736 151786 542742 151798
rect 546358 151786 546364 151798
rect 546416 151786 546422 151838
rect 542678 143598 542684 143610
rect 540856 143570 542684 143598
rect 540010 143490 540016 143542
rect 540068 143530 540074 143542
rect 540856 143530 540884 143570
rect 542678 143558 542684 143570
rect 542736 143558 542742 143610
rect 540068 143502 540884 143530
rect 540068 143490 540074 143502
rect 42290 141722 42296 141774
rect 42348 141762 42354 141774
rect 42566 141762 42572 141774
rect 42348 141734 42572 141762
rect 42348 141722 42354 141734
rect 42566 141722 42572 141734
rect 42624 141722 42630 141774
rect 87186 141654 87192 141706
rect 87244 141694 87250 141706
rect 88658 141694 88664 141706
rect 87244 141666 88664 141694
rect 87244 141654 87250 141666
rect 88658 141654 88664 141666
rect 88716 141654 88722 141706
rect 675158 137914 675164 137966
rect 675216 137954 675222 137966
rect 675526 137954 675532 137966
rect 675216 137926 675532 137954
rect 675216 137914 675222 137926
rect 675526 137914 675532 137926
rect 675584 137914 675590 137966
rect 88658 134310 88664 134362
rect 88716 134350 88722 134362
rect 90866 134350 90872 134362
rect 88716 134322 90872 134350
rect 88716 134310 88722 134322
rect 90866 134310 90872 134322
rect 90924 134310 90930 134362
rect 674882 132814 674888 132866
rect 674940 132854 674946 132866
rect 675526 132854 675532 132866
rect 674940 132826 675532 132854
rect 674940 132814 674946 132826
rect 675526 132814 675532 132826
rect 675584 132814 675590 132866
rect 675342 132786 675348 132798
rect 675084 132758 675348 132786
rect 675084 132730 675112 132758
rect 675342 132746 675348 132758
rect 675400 132746 675406 132798
rect 675434 132746 675440 132798
rect 675492 132746 675498 132798
rect 675066 132678 675072 132730
rect 675124 132678 675130 132730
rect 675452 132582 675480 132746
rect 675526 132582 675532 132594
rect 675452 132554 675532 132582
rect 675526 132542 675532 132554
rect 675584 132542 675590 132594
rect 42382 132474 42388 132526
rect 42440 132514 42446 132526
rect 42566 132514 42572 132526
rect 42440 132486 42572 132514
rect 42440 132474 42446 132486
rect 42566 132474 42572 132486
rect 42624 132474 42630 132526
rect 674974 129074 674980 129126
rect 675032 129114 675038 129126
rect 675250 129114 675256 129126
rect 675032 129086 675256 129114
rect 675032 129074 675038 129086
rect 675250 129074 675256 129086
rect 675308 129074 675314 129126
rect 42382 128734 42388 128786
rect 42440 128774 42446 128786
rect 42474 128774 42480 128786
rect 42440 128746 42480 128774
rect 42440 128734 42446 128746
rect 42474 128734 42480 128746
rect 42532 128734 42538 128786
rect 675158 124858 675164 124910
rect 675216 124858 675222 124910
rect 675176 124706 675204 124858
rect 675158 124654 675164 124706
rect 675216 124654 675222 124706
rect 674882 119894 674888 119946
rect 674940 119934 674946 119946
rect 675158 119934 675164 119946
rect 674940 119906 675164 119934
rect 674940 119894 674946 119906
rect 675158 119894 675164 119906
rect 675216 119894 675222 119946
rect 675066 119826 675072 119878
rect 675124 119826 675130 119878
rect 42474 119622 42480 119674
rect 42532 119622 42538 119674
rect 675084 119662 675112 119826
rect 675158 119662 675164 119674
rect 675084 119634 675164 119662
rect 675158 119622 675164 119634
rect 675216 119622 675222 119674
rect 42382 119554 42388 119606
rect 42440 119594 42446 119606
rect 42492 119594 42520 119622
rect 42440 119566 42520 119594
rect 42440 119554 42446 119566
rect 90866 118738 90872 118790
rect 90924 118778 90930 118790
rect 92522 118778 92528 118790
rect 90924 118750 92528 118778
rect 90924 118738 90930 118750
rect 92522 118738 92528 118750
rect 92580 118738 92586 118790
rect 674882 118670 674888 118722
rect 674940 118710 674946 118722
rect 675250 118710 675256 118722
rect 674940 118682 675256 118710
rect 674940 118670 674946 118682
rect 675250 118670 675256 118682
rect 675308 118670 675314 118722
rect 675066 117242 675072 117294
rect 675124 117242 675130 117294
rect 675084 117214 675112 117242
rect 675526 117214 675532 117226
rect 675084 117186 675532 117214
rect 675526 117174 675532 117186
rect 675584 117174 675590 117226
rect 39898 115950 39904 116002
rect 39956 115990 39962 116002
rect 40358 115990 40364 116002
rect 39956 115962 40364 115990
rect 39956 115950 39962 115962
rect 40358 115950 40364 115962
rect 40416 115990 40422 116002
rect 42106 115990 42112 116002
rect 40416 115962 42112 115990
rect 40416 115950 40422 115962
rect 42106 115950 42112 115962
rect 42164 115950 42170 116002
rect 92522 115882 92528 115934
rect 92580 115922 92586 115934
rect 93994 115922 94000 115934
rect 92580 115894 94000 115922
rect 92580 115882 92586 115894
rect 93994 115882 94000 115894
rect 94052 115882 94058 115934
rect 42198 109422 42204 109474
rect 42256 109462 42262 109474
rect 42474 109462 42480 109474
rect 42256 109434 42480 109462
rect 42256 109422 42262 109434
rect 42474 109422 42480 109434
rect 42532 109422 42538 109474
rect 93994 108538 94000 108590
rect 94052 108578 94058 108590
rect 94052 108550 95604 108578
rect 94052 108538 94058 108550
rect 95576 108510 95604 108550
rect 97398 108510 97404 108522
rect 95576 108482 97404 108510
rect 97398 108470 97404 108482
rect 97456 108470 97462 108522
rect 97398 102486 97404 102538
rect 97456 102526 97462 102538
rect 99698 102526 99704 102538
rect 97456 102498 99704 102526
rect 97456 102486 97462 102498
rect 99698 102486 99704 102498
rect 99756 102486 99762 102538
rect 44866 100106 44872 100158
rect 44924 100146 44930 100158
rect 45786 100146 45792 100158
rect 44924 100118 45792 100146
rect 44924 100106 44930 100118
rect 45786 100106 45792 100118
rect 45844 100106 45850 100158
rect 45786 99902 45792 99954
rect 45844 99942 45850 99954
rect 540102 99942 540108 99954
rect 45844 99914 540108 99942
rect 45844 99902 45850 99914
rect 540102 99902 540108 99914
rect 540160 99902 540166 99954
rect 99698 99834 99704 99886
rect 99756 99874 99762 99886
rect 126838 99874 126844 99886
rect 99756 99846 126844 99874
rect 99756 99834 99762 99846
rect 126838 99834 126844 99846
rect 126896 99834 126902 99886
rect 126838 95686 126844 95738
rect 126896 95726 126902 95738
rect 126896 95698 128724 95726
rect 126896 95686 126902 95698
rect 128696 95658 128724 95698
rect 130978 95658 130984 95670
rect 128696 95630 130984 95658
rect 130978 95618 130984 95630
rect 131036 95618 131042 95670
rect 42198 93782 42204 93834
rect 42256 93822 42262 93834
rect 42382 93822 42388 93834
rect 42256 93794 42388 93822
rect 42256 93782 42262 93794
rect 42382 93782 42388 93794
rect 42440 93782 42446 93834
rect 130978 91946 130984 91998
rect 131036 91986 131042 91998
rect 135026 91986 135032 91998
rect 131036 91958 135032 91986
rect 131036 91946 131042 91958
rect 135026 91946 135032 91958
rect 135084 91946 135090 91998
rect 42106 90110 42112 90162
rect 42164 90150 42170 90162
rect 42382 90150 42388 90162
rect 42164 90122 42388 90150
rect 42164 90110 42170 90122
rect 42382 90110 42388 90122
rect 42440 90110 42446 90162
rect 674790 86302 674796 86354
rect 674848 86342 674854 86354
rect 675526 86342 675532 86354
rect 674848 86314 675532 86342
rect 674848 86302 674854 86314
rect 675526 86302 675532 86314
rect 675584 86302 675590 86354
rect 675158 86234 675164 86286
rect 675216 86234 675222 86286
rect 675176 86082 675204 86234
rect 675158 86030 675164 86082
rect 675216 86030 675222 86082
rect 45142 85554 45148 85606
rect 45200 85594 45206 85606
rect 45786 85594 45792 85606
rect 45200 85566 45792 85594
rect 45200 85554 45206 85566
rect 45786 85554 45792 85566
rect 45844 85594 45850 85606
rect 465490 85594 465496 85606
rect 45844 85566 465496 85594
rect 45844 85554 45850 85566
rect 465490 85554 465496 85566
rect 465548 85554 465554 85606
rect 39254 84670 39260 84722
rect 39312 84710 39318 84722
rect 45142 84710 45148 84722
rect 39312 84682 45148 84710
rect 39312 84670 39318 84682
rect 45142 84670 45148 84682
rect 45200 84670 45206 84722
rect 674790 83786 674796 83838
rect 674848 83826 674854 83838
rect 675250 83826 675256 83838
rect 674848 83798 675256 83826
rect 674848 83786 674854 83798
rect 675250 83786 675256 83798
rect 675308 83786 675314 83838
rect 135026 83582 135032 83634
rect 135084 83622 135090 83634
rect 136038 83622 136044 83634
rect 135084 83594 136044 83622
rect 135084 83582 135090 83594
rect 136038 83582 136044 83594
rect 136096 83582 136102 83634
rect 675066 83514 675072 83566
rect 675124 83554 675130 83566
rect 675250 83554 675256 83566
rect 675124 83526 675256 83554
rect 675124 83514 675130 83526
rect 675250 83514 675256 83526
rect 675308 83514 675314 83566
rect 674882 82494 674888 82546
rect 674940 82534 674946 82546
rect 675250 82534 675256 82546
rect 674940 82506 675256 82534
rect 674940 82494 674946 82506
rect 675250 82494 675256 82506
rect 675308 82494 675314 82546
rect 42106 77258 42112 77310
rect 42164 77298 42170 77310
rect 42290 77298 42296 77310
rect 42164 77270 42296 77298
rect 42164 77258 42170 77270
rect 42290 77258 42296 77270
rect 42348 77258 42354 77310
rect 43946 76306 43952 76358
rect 44004 76346 44010 76358
rect 149746 76346 149752 76358
rect 44004 76318 149752 76346
rect 44004 76306 44010 76318
rect 149746 76306 149752 76318
rect 149804 76306 149810 76358
rect 136038 74606 136044 74658
rect 136096 74646 136102 74658
rect 138798 74646 138804 74658
rect 136096 74618 138804 74646
rect 136096 74606 136102 74618
rect 138798 74606 138804 74618
rect 138856 74606 138862 74658
rect 674882 73994 674888 74046
rect 674940 74034 674946 74046
rect 674940 74006 675020 74034
rect 674940 73994 674946 74006
rect 674992 73842 675020 74006
rect 674974 73790 674980 73842
rect 675032 73790 675038 73842
rect 674790 73654 674796 73706
rect 674848 73694 674854 73706
rect 675158 73694 675164 73706
rect 674848 73666 675164 73694
rect 674848 73654 674854 73666
rect 675158 73654 675164 73666
rect 675216 73654 675222 73706
rect 675158 73558 675164 73570
rect 675084 73530 675164 73558
rect 675084 73298 675112 73530
rect 675158 73518 675164 73530
rect 675216 73518 675222 73570
rect 675066 73246 675072 73298
rect 675124 73246 675130 73298
rect 39714 72634 39720 72686
rect 39772 72674 39778 72686
rect 90866 72674 90872 72686
rect 39772 72646 90872 72674
rect 39772 72634 39778 72646
rect 90866 72634 90872 72646
rect 90924 72634 90930 72686
rect 674882 72090 674888 72142
rect 674940 72130 674946 72142
rect 675250 72130 675256 72142
rect 674940 72102 675256 72130
rect 674940 72090 674946 72102
rect 675250 72090 675256 72102
rect 675308 72090 675314 72142
rect 39530 67126 39536 67178
rect 39588 67166 39594 67178
rect 140546 67166 140552 67178
rect 39588 67138 140552 67166
rect 39588 67126 39594 67138
rect 140546 67126 140552 67138
rect 140604 67126 140610 67178
rect 138798 66174 138804 66226
rect 138856 66214 138862 66226
rect 140638 66214 140644 66226
rect 138856 66186 140644 66214
rect 138856 66174 138862 66186
rect 140638 66174 140644 66186
rect 140696 66174 140702 66226
rect 140638 62502 140644 62554
rect 140696 62542 140702 62554
rect 142386 62542 142392 62554
rect 140696 62514 142392 62542
rect 140696 62502 140702 62514
rect 142386 62502 142392 62514
rect 142444 62502 142450 62554
rect 670282 45910 670288 45962
rect 670340 45950 670346 45962
rect 675158 45950 675164 45962
rect 670340 45922 675164 45950
rect 670340 45910 670346 45922
rect 675158 45910 675164 45922
rect 675216 45910 675222 45962
rect 183786 45134 183792 45146
rect 180216 45106 183792 45134
rect 43026 45026 43032 45078
rect 43084 45066 43090 45078
rect 180216 45066 180244 45106
rect 183786 45094 183792 45106
rect 183844 45094 183850 45146
rect 195838 45134 195844 45146
rect 193004 45106 195844 45134
rect 43084 45038 180244 45066
rect 43084 45026 43090 45038
rect 183878 45026 183884 45078
rect 183936 45066 183942 45078
rect 193004 45066 193032 45106
rect 195838 45094 195844 45106
rect 195896 45134 195902 45146
rect 196666 45134 196672 45146
rect 195896 45106 196672 45134
rect 195896 45094 195902 45106
rect 196666 45094 196672 45106
rect 196724 45094 196730 45146
rect 515078 45094 515084 45146
rect 515136 45134 515142 45146
rect 516182 45134 516188 45146
rect 515136 45106 516188 45134
rect 515136 45094 515142 45106
rect 516182 45094 516188 45106
rect 516240 45134 516246 45146
rect 516240 45106 525060 45134
rect 516240 45094 516246 45106
rect 183936 45038 193032 45066
rect 525032 45066 525060 45106
rect 527314 45094 527320 45146
rect 527372 45134 527378 45146
rect 675342 45134 675348 45146
rect 527372 45106 675348 45134
rect 527372 45094 527378 45106
rect 675342 45094 675348 45106
rect 675400 45094 675406 45146
rect 540838 45066 540844 45078
rect 525032 45038 540844 45066
rect 183936 45026 183942 45038
rect 540838 45026 540844 45038
rect 540896 45026 540902 45078
rect 553626 44958 553632 45010
rect 553684 44998 553690 45010
rect 553684 44970 557352 44998
rect 553684 44958 553690 44970
rect 218838 44794 218844 44806
rect 212324 44766 218844 44794
rect 196666 44686 196672 44738
rect 196724 44726 196730 44738
rect 209546 44726 209552 44738
rect 196724 44698 209552 44726
rect 196724 44686 196730 44698
rect 209546 44686 209552 44698
rect 209604 44686 209610 44738
rect 209638 44686 209644 44738
rect 209696 44726 209702 44738
rect 212324 44726 212352 44766
rect 218838 44754 218844 44766
rect 218896 44754 218902 44806
rect 244598 44794 244604 44806
rect 238084 44766 244604 44794
rect 209696 44698 212352 44726
rect 209696 44686 209702 44698
rect 231626 44686 231632 44738
rect 231684 44726 231690 44738
rect 235306 44726 235312 44738
rect 231684 44698 235312 44726
rect 231684 44686 231690 44698
rect 235306 44686 235312 44698
rect 235364 44686 235370 44738
rect 235398 44686 235404 44738
rect 235456 44726 235462 44738
rect 238084 44726 238112 44766
rect 244598 44754 244604 44766
rect 244656 44754 244662 44806
rect 273946 44794 273952 44806
rect 263844 44766 273952 44794
rect 235456 44698 238112 44726
rect 235456 44686 235462 44698
rect 257386 44686 257392 44738
rect 257444 44726 257450 44738
rect 261066 44726 261072 44738
rect 257444 44698 261072 44726
rect 257444 44686 257450 44698
rect 261066 44686 261072 44698
rect 261124 44686 261130 44738
rect 261158 44686 261164 44738
rect 261216 44726 261222 44738
rect 263844 44726 263872 44766
rect 273946 44754 273952 44766
rect 274004 44754 274010 44806
rect 417466 44754 417472 44806
rect 417524 44794 417530 44806
rect 424918 44794 424924 44806
rect 417524 44766 424924 44794
rect 417524 44754 417530 44766
rect 424918 44754 424924 44766
rect 424976 44754 424982 44806
rect 515078 44794 515084 44806
rect 505804 44766 515084 44794
rect 261216 44698 263872 44726
rect 261216 44686 261222 44698
rect 274130 44686 274136 44738
rect 274188 44726 274194 44738
rect 274188 44698 281444 44726
rect 274188 44686 274194 44698
rect 281416 44658 281444 44698
rect 307434 44686 307440 44738
rect 307492 44726 307498 44738
rect 318106 44726 318112 44738
rect 307492 44698 318112 44726
rect 307492 44686 307498 44698
rect 318106 44686 318112 44698
rect 318164 44686 318170 44738
rect 344786 44686 344792 44738
rect 344844 44726 344850 44738
rect 351778 44726 351784 44738
rect 344844 44698 351784 44726
rect 344844 44686 344850 44698
rect 351778 44686 351784 44698
rect 351836 44686 351842 44738
rect 359230 44686 359236 44738
rect 359288 44726 359294 44738
rect 359288 44698 412912 44726
rect 359288 44686 359294 44698
rect 283146 44658 283152 44670
rect 281416 44630 283152 44658
rect 283146 44618 283152 44630
rect 283204 44618 283210 44670
rect 299614 44658 299620 44670
rect 296044 44630 299620 44658
rect 283330 44550 283336 44602
rect 283388 44590 283394 44602
rect 296044 44590 296072 44630
rect 299614 44618 299620 44630
rect 299672 44618 299678 44670
rect 412884 44658 412912 44698
rect 437706 44686 437712 44738
rect 437764 44726 437770 44738
rect 441386 44726 441392 44738
rect 437764 44698 441392 44726
rect 437764 44686 437770 44698
rect 441386 44686 441392 44698
rect 441444 44686 441450 44738
rect 505804 44726 505832 44766
rect 515078 44754 515084 44766
rect 515136 44754 515142 44806
rect 557324 44794 557352 44970
rect 570186 44794 570192 44806
rect 557324 44766 570192 44794
rect 570186 44754 570192 44766
rect 570244 44754 570250 44806
rect 570278 44754 570284 44806
rect 570336 44794 570342 44806
rect 570336 44766 572992 44794
rect 570336 44754 570342 44766
rect 493016 44698 505832 44726
rect 572964 44726 572992 44766
rect 592266 44754 592272 44806
rect 592324 44794 592330 44806
rect 595946 44794 595952 44806
rect 592324 44766 595952 44794
rect 592324 44754 592330 44766
rect 595946 44754 595952 44766
rect 596004 44754 596010 44806
rect 596038 44754 596044 44806
rect 596096 44794 596102 44806
rect 596096 44766 598752 44794
rect 596096 44754 596102 44766
rect 579478 44726 579484 44738
rect 572964 44698 579484 44726
rect 413878 44658 413884 44670
rect 389884 44630 410428 44658
rect 412884 44630 413884 44658
rect 283388 44562 296072 44590
rect 283388 44550 283394 44562
rect 308078 44550 308084 44602
rect 308136 44590 308142 44602
rect 358586 44590 358592 44602
rect 308136 44562 358592 44590
rect 308136 44550 308142 44562
rect 358586 44550 358592 44562
rect 358644 44550 358650 44602
rect 376986 44590 376992 44602
rect 364216 44562 376992 44590
rect 195194 44482 195200 44534
rect 195252 44522 195258 44534
rect 199518 44522 199524 44534
rect 195252 44494 199524 44522
rect 195252 44482 195258 44494
rect 199518 44482 199524 44494
rect 199576 44522 199582 44534
rect 303754 44522 303760 44534
rect 199576 44494 303760 44522
rect 199576 44482 199582 44494
rect 303754 44482 303760 44494
rect 303812 44482 303818 44534
rect 318106 44482 318112 44534
rect 318164 44522 318170 44534
rect 331078 44522 331084 44534
rect 318164 44494 331084 44522
rect 318164 44482 318170 44494
rect 331078 44482 331084 44494
rect 331136 44482 331142 44534
rect 362818 44482 362824 44534
rect 362876 44522 362882 44534
rect 364216 44522 364244 44562
rect 376986 44550 376992 44562
rect 377044 44550 377050 44602
rect 377170 44550 377176 44602
rect 377228 44590 377234 44602
rect 389884 44590 389912 44630
rect 377228 44562 389912 44590
rect 377228 44550 377234 44562
rect 362876 44494 364244 44522
rect 362876 44482 362882 44494
rect 200714 44414 200720 44466
rect 200772 44454 200778 44466
rect 242758 44454 242764 44466
rect 200772 44426 242764 44454
rect 200772 44414 200778 44426
rect 242758 44414 242764 44426
rect 242816 44414 242822 44466
rect 306238 44414 306244 44466
rect 306296 44454 306302 44466
rect 309274 44454 309280 44466
rect 306296 44426 309280 44454
rect 306296 44414 306302 44426
rect 309274 44414 309280 44426
rect 309332 44454 309338 44466
rect 352422 44454 352428 44466
rect 309332 44426 352428 44454
rect 309332 44414 309338 44426
rect 352422 44414 352428 44426
rect 352480 44454 352486 44466
rect 355458 44454 355464 44466
rect 352480 44426 355464 44454
rect 352480 44414 352486 44426
rect 355458 44414 355464 44426
rect 355516 44454 355522 44466
rect 361070 44454 361076 44466
rect 355516 44426 361076 44454
rect 355516 44414 355522 44426
rect 361070 44414 361076 44426
rect 361128 44454 361134 44466
rect 364106 44454 364112 44466
rect 361128 44426 364112 44454
rect 361128 44414 361134 44426
rect 364106 44414 364112 44426
rect 364164 44454 364170 44466
rect 407254 44454 407260 44466
rect 364164 44426 407260 44454
rect 364164 44414 364170 44426
rect 407254 44414 407260 44426
rect 407312 44454 407318 44466
rect 410290 44454 410296 44466
rect 407312 44426 410296 44454
rect 407312 44414 407318 44426
rect 410290 44414 410296 44426
rect 410348 44414 410354 44466
rect 410400 44454 410428 44630
rect 413878 44618 413884 44630
rect 413936 44618 413942 44670
rect 441570 44618 441576 44670
rect 441628 44658 441634 44670
rect 450678 44658 450684 44670
rect 441628 44630 450684 44658
rect 441628 44618 441634 44630
rect 450678 44618 450684 44630
rect 450736 44618 450742 44670
rect 459510 44618 459516 44670
rect 459568 44658 459574 44670
rect 467514 44658 467520 44670
rect 459568 44630 467520 44658
rect 459568 44618 459574 44630
rect 467514 44618 467520 44630
rect 467572 44618 467578 44670
rect 471838 44618 471844 44670
rect 471896 44658 471902 44670
rect 473770 44658 473776 44670
rect 471896 44630 473776 44658
rect 471896 44618 471902 44630
rect 473770 44618 473776 44630
rect 473828 44618 473834 44670
rect 473862 44618 473868 44670
rect 473920 44658 473926 44670
rect 480118 44658 480124 44670
rect 473920 44630 480124 44658
rect 473920 44618 473926 44630
rect 480118 44618 480124 44630
rect 480176 44618 480182 44670
rect 489226 44618 489232 44670
rect 489284 44658 489290 44670
rect 493016 44658 493044 44698
rect 579478 44686 579484 44698
rect 579536 44686 579542 44738
rect 598724 44726 598752 44766
rect 618026 44754 618032 44806
rect 618084 44794 618090 44806
rect 621706 44794 621712 44806
rect 618084 44766 621712 44794
rect 618084 44754 618090 44766
rect 621706 44754 621712 44766
rect 621764 44754 621770 44806
rect 621798 44754 621804 44806
rect 621856 44794 621862 44806
rect 621856 44766 624512 44794
rect 621856 44754 621862 44766
rect 605238 44726 605244 44738
rect 598724 44698 605244 44726
rect 605238 44686 605244 44698
rect 605296 44686 605302 44738
rect 624484 44726 624512 44766
rect 643786 44754 643792 44806
rect 643844 44794 643850 44806
rect 647466 44794 647472 44806
rect 643844 44766 647472 44794
rect 643844 44754 643850 44766
rect 647466 44754 647472 44766
rect 647524 44754 647530 44806
rect 647558 44754 647564 44806
rect 647616 44794 647622 44806
rect 647616 44766 650272 44794
rect 647616 44754 647622 44766
rect 630998 44726 631004 44738
rect 624484 44698 631004 44726
rect 630998 44686 631004 44698
rect 631056 44686 631062 44738
rect 650244 44726 650272 44766
rect 669546 44754 669552 44806
rect 669604 44794 669610 44806
rect 670282 44794 670288 44806
rect 669604 44766 670288 44794
rect 669604 44754 669610 44766
rect 670282 44754 670288 44766
rect 670340 44754 670346 44806
rect 656758 44726 656764 44738
rect 650244 44698 656764 44726
rect 656758 44686 656764 44698
rect 656816 44686 656822 44738
rect 489284 44630 493044 44658
rect 489284 44618 489290 44630
rect 463466 44550 463472 44602
rect 463524 44590 463530 44602
rect 471856 44590 471884 44618
rect 463524 44562 471884 44590
rect 463524 44550 463530 44562
rect 413878 44482 413884 44534
rect 413936 44522 413942 44534
rect 414062 44522 414068 44534
rect 413936 44494 414068 44522
rect 413936 44482 413942 44494
rect 414062 44482 414068 44494
rect 414120 44522 414126 44534
rect 468802 44522 468808 44534
rect 414120 44494 468808 44522
rect 414120 44482 414126 44494
rect 468802 44482 468808 44494
rect 468860 44482 468866 44534
rect 476346 44482 476352 44534
rect 476404 44522 476410 44534
rect 515078 44522 515084 44534
rect 476404 44494 515084 44522
rect 476404 44482 476410 44494
rect 515078 44482 515084 44494
rect 515136 44482 515142 44534
rect 412958 44454 412964 44466
rect 410400 44426 412964 44454
rect 412958 44414 412964 44426
rect 413016 44414 413022 44466
rect 419030 44414 419036 44466
rect 419088 44454 419094 44466
rect 461994 44454 462000 44466
rect 419088 44426 462000 44454
rect 419088 44414 419094 44426
rect 461994 44414 462000 44426
rect 462052 44454 462058 44466
rect 465030 44454 465036 44466
rect 462052 44426 465036 44454
rect 462052 44414 462058 44426
rect 465030 44414 465036 44426
rect 465088 44454 465094 44466
rect 465490 44454 465496 44466
rect 465088 44426 465496 44454
rect 465088 44414 465094 44426
rect 465490 44414 465496 44426
rect 465548 44414 465554 44466
rect 473586 44414 473592 44466
rect 473644 44454 473650 44466
rect 516826 44454 516832 44466
rect 473644 44426 516832 44454
rect 473644 44414 473650 44426
rect 516826 44414 516832 44426
rect 516884 44454 516890 44466
rect 519862 44454 519868 44466
rect 516884 44426 519868 44454
rect 516884 44414 516890 44426
rect 519862 44414 519868 44426
rect 519920 44414 519926 44466
rect 201358 44346 201364 44398
rect 201416 44386 201422 44398
rect 244506 44386 244512 44398
rect 201416 44358 244512 44386
rect 201416 44346 201422 44358
rect 244506 44346 244512 44358
rect 244564 44346 244570 44398
rect 296946 44346 296952 44398
rect 297004 44386 297010 44398
rect 299430 44386 299436 44398
rect 297004 44358 299436 44386
rect 297004 44346 297010 44358
rect 299430 44346 299436 44358
rect 299488 44386 299494 44398
rect 305594 44386 305600 44398
rect 299488 44358 305600 44386
rect 299488 44346 299494 44358
rect 305594 44346 305600 44358
rect 305652 44386 305658 44398
rect 344786 44386 344792 44398
rect 305652 44358 344792 44386
rect 305652 44346 305658 44358
rect 344786 44346 344792 44358
rect 344844 44346 344850 44398
rect 344878 44346 344884 44398
rect 344936 44386 344942 44398
rect 362266 44386 362272 44398
rect 344936 44358 362272 44386
rect 344936 44346 344942 44358
rect 362266 44346 362272 44358
rect 362324 44386 362330 44398
rect 362818 44386 362824 44398
rect 362324 44358 362824 44386
rect 362324 44346 362330 44358
rect 362818 44346 362824 44358
rect 362876 44346 362882 44398
rect 362910 44346 362916 44398
rect 362968 44386 362974 44398
rect 413418 44386 413424 44398
rect 362968 44358 413424 44386
rect 362968 44346 362974 44358
rect 413418 44346 413424 44358
rect 413476 44386 413482 44398
rect 417742 44386 417748 44398
rect 413476 44358 417748 44386
rect 413476 44346 413482 44358
rect 417742 44346 417748 44358
rect 417800 44386 417806 44398
rect 468158 44386 468164 44398
rect 417800 44358 468164 44386
rect 417800 44346 417806 44358
rect 468158 44346 468164 44358
rect 468216 44346 468222 44398
rect 472482 44346 472488 44398
rect 472540 44386 472546 44398
rect 522990 44386 522996 44398
rect 472540 44358 522996 44386
rect 472540 44346 472546 44358
rect 522990 44346 522996 44358
rect 523048 44346 523054 44398
rect 90866 44278 90872 44330
rect 90924 44318 90930 44330
rect 198874 44318 198880 44330
rect 90924 44290 198880 44318
rect 90924 44278 90930 44290
rect 198874 44278 198880 44290
rect 198932 44318 198938 44330
rect 247082 44318 247088 44330
rect 198932 44290 247088 44318
rect 198932 44278 198938 44290
rect 247082 44278 247088 44290
rect 247140 44318 247146 44330
rect 307434 44318 307440 44330
rect 247140 44290 307440 44318
rect 247140 44278 247146 44290
rect 307434 44278 307440 44290
rect 307492 44278 307498 44330
rect 331078 44278 331084 44330
rect 331136 44318 331142 44330
rect 334758 44318 334764 44330
rect 331136 44290 334764 44318
rect 331136 44278 331142 44290
rect 334758 44278 334764 44290
rect 334816 44278 334822 44330
rect 351778 44278 351784 44330
rect 351836 44318 351842 44330
rect 354262 44318 354268 44330
rect 351836 44290 354268 44318
rect 351836 44278 351842 44290
rect 354262 44278 354268 44290
rect 354320 44318 354326 44330
rect 360426 44318 360432 44330
rect 354320 44290 360432 44318
rect 354320 44278 354326 44290
rect 360426 44278 360432 44290
rect 360484 44318 360490 44330
rect 406610 44318 406616 44330
rect 360484 44290 406616 44318
rect 360484 44278 360490 44290
rect 406610 44278 406616 44290
rect 406668 44318 406674 44330
rect 461350 44318 461356 44330
rect 406668 44290 461356 44318
rect 406668 44278 406674 44290
rect 461350 44278 461356 44290
rect 461408 44318 461414 44330
rect 473862 44318 473868 44330
rect 461408 44290 473868 44318
rect 461408 44278 461414 44290
rect 473862 44278 473868 44290
rect 473920 44278 473926 44330
rect 518666 44278 518672 44330
rect 518724 44318 518730 44330
rect 524830 44318 524836 44330
rect 518724 44290 524836 44318
rect 518724 44278 518730 44290
rect 524830 44278 524836 44290
rect 524888 44278 524894 44330
rect 525934 44278 525940 44330
rect 525992 44318 525998 44330
rect 568990 44318 568996 44330
rect 525992 44290 568996 44318
rect 525992 44278 525998 44290
rect 568990 44278 568996 44290
rect 569048 44278 569054 44330
rect 148918 44210 148924 44262
rect 148976 44250 148982 44262
rect 149746 44250 149752 44262
rect 148976 44222 149752 44250
rect 148976 44210 148982 44222
rect 149746 44210 149752 44222
rect 149804 44250 149810 44262
rect 188386 44250 188392 44262
rect 149804 44222 188392 44250
rect 149804 44210 149810 44222
rect 188386 44210 188392 44222
rect 188444 44250 188450 44262
rect 192710 44250 192716 44262
rect 188444 44222 192716 44250
rect 188444 44210 188450 44222
rect 192710 44210 192716 44222
rect 192768 44250 192774 44262
rect 201358 44250 201364 44262
rect 192768 44222 201364 44250
rect 192768 44210 192774 44222
rect 201358 44210 201364 44222
rect 201416 44210 201422 44262
rect 304398 44210 304404 44262
rect 304456 44250 304462 44262
rect 338346 44250 338352 44262
rect 304456 44222 338352 44250
rect 304456 44210 304462 44222
rect 338346 44210 338352 44222
rect 338404 44210 338410 44262
rect 338530 44210 338536 44262
rect 338588 44250 338594 44262
rect 359230 44250 359236 44262
rect 338588 44222 359236 44250
rect 338588 44210 338594 44222
rect 359230 44210 359236 44222
rect 359288 44210 359294 44262
rect 410934 44210 410940 44262
rect 410992 44250 410998 44262
rect 410992 44222 412912 44250
rect 410992 44210 410998 44222
rect 186546 44142 186552 44194
rect 186604 44182 186610 44194
rect 194550 44182 194556 44194
rect 186604 44154 194556 44182
rect 186604 44142 186610 44154
rect 194550 44142 194556 44154
rect 194608 44142 194614 44194
rect 295106 44142 295112 44194
rect 295164 44182 295170 44194
rect 303110 44182 303116 44194
rect 295164 44154 303116 44182
rect 295164 44142 295170 44154
rect 303110 44142 303116 44154
rect 303168 44142 303174 44194
rect 349938 44142 349944 44194
rect 349996 44182 350002 44194
rect 357942 44182 357948 44194
rect 349996 44154 357948 44182
rect 349996 44142 350002 44154
rect 357942 44142 357948 44154
rect 358000 44142 358006 44194
rect 358586 44142 358592 44194
rect 358644 44182 358650 44194
rect 362910 44182 362916 44194
rect 358644 44154 362916 44182
rect 358644 44142 358650 44154
rect 362910 44142 362916 44154
rect 362968 44142 362974 44194
rect 404770 44142 404776 44194
rect 404828 44182 404834 44194
rect 412774 44182 412780 44194
rect 404828 44154 412780 44182
rect 404828 44142 404834 44154
rect 412774 44142 412780 44154
rect 412832 44142 412838 44194
rect 412884 44182 412912 44222
rect 412958 44210 412964 44262
rect 413016 44250 413022 44262
rect 417098 44250 417104 44262
rect 413016 44222 417104 44250
rect 413016 44210 413022 44222
rect 417098 44210 417104 44222
rect 417156 44250 417162 44262
rect 417466 44250 417472 44262
rect 417156 44222 417472 44250
rect 417156 44210 417162 44222
rect 417466 44210 417472 44222
rect 417524 44210 417530 44262
rect 473770 44210 473776 44262
rect 473828 44250 473834 44262
rect 526670 44250 526676 44262
rect 473828 44222 526676 44250
rect 473828 44210 473834 44222
rect 526670 44210 526676 44222
rect 526728 44250 526734 44262
rect 630262 44250 630268 44262
rect 526728 44222 630268 44250
rect 526728 44210 526734 44222
rect 630262 44210 630268 44222
rect 630320 44210 630326 44262
rect 419582 44182 419588 44194
rect 412884 44154 419588 44182
rect 419582 44142 419588 44154
rect 419640 44142 419646 44194
rect 465674 44142 465680 44194
rect 465732 44182 465738 44194
rect 474322 44182 474328 44194
rect 465732 44154 474328 44182
rect 465732 44142 465738 44154
rect 474322 44142 474328 44154
rect 474380 44142 474386 44194
rect 514342 44142 514348 44194
rect 514400 44182 514406 44194
rect 522346 44182 522352 44194
rect 514400 44154 522352 44182
rect 514400 44142 514406 44154
rect 522346 44142 522352 44154
rect 522404 44142 522410 44194
rect 522990 44142 522996 44194
rect 523048 44182 523054 44194
rect 527314 44182 527320 44194
rect 523048 44154 527320 44182
rect 523048 44142 523054 44154
rect 527314 44142 527320 44154
rect 527372 44142 527378 44194
rect 515078 43530 515084 43582
rect 515136 43570 515142 43582
rect 523634 43570 523640 43582
rect 515136 43542 523640 43570
rect 515136 43530 515142 43542
rect 523634 43530 523640 43542
rect 523692 43570 523698 43582
rect 525934 43570 525940 43582
rect 523692 43542 525940 43570
rect 523692 43530 523698 43542
rect 525934 43530 525940 43542
rect 525992 43530 525998 43582
rect 142386 43326 142392 43378
rect 142444 43366 142450 43378
rect 144962 43366 144968 43378
rect 142444 43338 144968 43366
rect 142444 43326 142450 43338
rect 144962 43326 144968 43338
rect 145020 43326 145026 43378
rect 251314 43190 251320 43242
rect 251372 43230 251378 43242
rect 297590 43230 297596 43242
rect 251372 43202 297596 43230
rect 251372 43190 251378 43202
rect 297590 43190 297596 43202
rect 297648 43190 297654 43242
rect 579478 43190 579484 43242
rect 579536 43230 579542 43242
rect 675250 43230 675256 43242
rect 579536 43202 675256 43230
rect 579536 43190 579542 43202
rect 675250 43190 675256 43202
rect 675308 43190 675314 43242
rect 299614 42442 299620 42494
rect 299672 42482 299678 42494
rect 304398 42482 304404 42494
rect 299672 42454 304404 42482
rect 299672 42442 299678 42454
rect 304398 42442 304404 42454
rect 304456 42442 304462 42494
rect 144962 42374 144968 42426
rect 145020 42414 145026 42426
rect 195194 42414 195200 42426
rect 145020 42386 195200 42414
rect 145020 42374 145026 42386
rect 195194 42374 195200 42386
rect 195252 42374 195258 42426
rect 242758 42374 242764 42426
rect 242816 42414 242822 42426
rect 251314 42414 251320 42426
rect 242816 42386 251320 42414
rect 242816 42374 242822 42386
rect 251314 42374 251320 42386
rect 251372 42374 251378 42426
rect 297590 42374 297596 42426
rect 297648 42414 297654 42426
rect 300626 42414 300632 42426
rect 297648 42386 300632 42414
rect 297648 42374 297654 42386
rect 300626 42374 300632 42386
rect 300684 42374 300690 42426
rect 144410 42306 144416 42358
rect 144468 42346 144474 42358
rect 253798 42346 253804 42358
rect 144468 42318 253804 42346
rect 144468 42306 144474 42318
rect 253798 42306 253804 42318
rect 253856 42346 253862 42358
rect 569082 42346 569088 42358
rect 253856 42318 569088 42346
rect 253856 42306 253862 42318
rect 569082 42306 569088 42318
rect 569140 42346 569146 42358
rect 579478 42346 579484 42358
rect 569140 42318 579484 42346
rect 569140 42306 569146 42318
rect 579478 42306 579484 42318
rect 579536 42306 579542 42358
rect 303754 42238 303760 42290
rect 303812 42278 303818 42290
rect 308078 42278 308084 42290
rect 303812 42250 308084 42278
rect 303812 42238 303818 42250
rect 308078 42238 308084 42250
rect 308136 42238 308142 42290
rect 468158 42238 468164 42290
rect 468216 42278 468222 42290
rect 472482 42278 472488 42290
rect 468216 42250 472488 42278
rect 468216 42238 468222 42250
rect 472482 42238 472488 42250
rect 472540 42238 472546 42290
rect 189122 41898 189128 41950
rect 189180 41938 189186 41950
rect 306146 41938 306152 41950
rect 189180 41910 191008 41938
rect 189180 41898 189186 41910
rect 190980 41814 191008 41910
rect 304876 41910 306152 41938
rect 198322 41830 198328 41882
rect 198380 41870 198386 41882
rect 199978 41870 199984 41882
rect 198380 41842 199984 41870
rect 198380 41830 198386 41842
rect 199978 41830 199984 41842
rect 200036 41830 200042 41882
rect 304876 41814 304904 41910
rect 306146 41898 306152 41910
rect 306204 41898 306210 41950
rect 409186 41830 409192 41882
rect 409244 41870 409250 41882
rect 412222 41870 412228 41882
rect 409244 41842 412228 41870
rect 409244 41830 409250 41842
rect 412222 41830 412228 41842
rect 412280 41870 412286 41882
rect 415074 41870 415080 41882
rect 412280 41842 415080 41870
rect 412280 41830 412286 41842
rect 415074 41830 415080 41842
rect 415132 41830 415138 41882
rect 464018 41830 464024 41882
rect 464076 41870 464082 41882
rect 467054 41870 467060 41882
rect 464076 41842 467060 41870
rect 464076 41830 464082 41842
rect 467054 41830 467060 41842
rect 467112 41870 467118 41882
rect 469906 41870 469912 41882
rect 467112 41842 469912 41870
rect 467112 41830 467118 41842
rect 469906 41830 469912 41842
rect 469964 41830 469970 41882
rect 519954 41830 519960 41882
rect 520012 41870 520018 41882
rect 521242 41870 521248 41882
rect 520012 41842 521248 41870
rect 520012 41830 520018 41842
rect 521242 41830 521248 41842
rect 521300 41870 521306 41882
rect 524278 41870 524284 41882
rect 521300 41842 524284 41870
rect 521300 41830 521306 41842
rect 524278 41830 524284 41842
rect 524336 41870 524342 41882
rect 525566 41870 525572 41882
rect 524336 41842 525572 41870
rect 524336 41830 524342 41842
rect 525566 41830 525572 41842
rect 525624 41870 525630 41882
rect 527774 41870 527780 41882
rect 525624 41842 527780 41870
rect 525624 41830 525630 41842
rect 527774 41830 527780 41842
rect 527832 41830 527838 41882
rect 190962 41762 190968 41814
rect 191020 41802 191026 41814
rect 192158 41802 192164 41814
rect 191020 41774 192164 41802
rect 191020 41762 191026 41774
rect 192158 41762 192164 41774
rect 192216 41802 192222 41814
rect 193446 41802 193452 41814
rect 192216 41774 193452 41802
rect 192216 41762 192222 41774
rect 193446 41762 193452 41774
rect 193504 41802 193510 41814
rect 196298 41802 196304 41814
rect 193504 41774 196304 41802
rect 193504 41762 193510 41774
rect 196298 41762 196304 41774
rect 196356 41762 196362 41814
rect 297130 41762 297136 41814
rect 297188 41762 297194 41814
rect 302098 41762 302104 41814
rect 302156 41802 302162 41814
rect 304858 41802 304864 41814
rect 302156 41774 304864 41802
rect 302156 41762 302162 41774
rect 304858 41762 304864 41774
rect 304916 41762 304922 41814
rect 359874 41762 359880 41814
rect 359932 41802 359938 41814
rect 360978 41802 360984 41814
rect 359932 41774 360984 41802
rect 359932 41762 359938 41774
rect 360978 41762 360984 41774
rect 361036 41762 361042 41814
rect 410382 41762 410388 41814
rect 410440 41802 410446 41814
rect 411394 41802 411400 41814
rect 410440 41774 411400 41802
rect 410440 41762 410446 41774
rect 411394 41762 411400 41774
rect 411452 41802 411458 41814
rect 414430 41802 414436 41814
rect 411452 41774 414436 41802
rect 411452 41762 411458 41774
rect 414430 41762 414436 41774
rect 414488 41802 414494 41814
rect 415718 41802 415724 41814
rect 414488 41774 415724 41802
rect 414488 41762 414494 41774
rect 415718 41762 415724 41774
rect 415776 41802 415782 41814
rect 418110 41802 418116 41814
rect 415776 41774 418116 41802
rect 415776 41762 415782 41774
rect 418110 41762 418116 41774
rect 418168 41802 418174 41814
rect 419030 41802 419036 41814
rect 418168 41774 419036 41802
rect 418168 41762 418174 41774
rect 419030 41762 419036 41774
rect 419088 41762 419094 41814
rect 251958 41558 251964 41610
rect 252016 41598 252022 41610
rect 252016 41570 261204 41598
rect 252016 41558 252022 41570
rect 261176 41530 261204 41570
rect 286918 41558 286924 41610
rect 286976 41598 286982 41610
rect 297148 41598 297176 41762
rect 286976 41570 297176 41598
rect 286976 41558 286982 41570
rect 261176 41502 273992 41530
rect 273964 41394 273992 41502
rect 286918 41394 286924 41406
rect 273964 41366 286924 41394
rect 286918 41354 286924 41366
rect 286976 41354 286982 41406
rect 134106 40130 134112 40182
rect 134164 40170 134170 40182
rect 143398 40170 143404 40182
rect 134164 40142 143404 40170
rect 134164 40130 134170 40142
rect 143398 40130 143404 40142
rect 143456 40130 143462 40182
rect 140854 40062 140860 40114
rect 140912 40102 140918 40114
rect 142930 40102 142936 40114
rect 140912 40074 142936 40102
rect 140912 40062 140918 40074
rect 142450 39952 142478 40074
rect 142930 40062 142936 40074
rect 142988 40102 142994 40114
rect 144410 40102 144416 40114
rect 142988 40074 144416 40102
rect 142988 40062 142994 40074
rect 144410 40062 144416 40074
rect 144468 40062 144474 40114
rect 241102 39654 241108 39706
rect 241160 39694 241166 39706
rect 242758 39694 242764 39706
rect 241160 39666 242764 39694
rect 241160 39654 241166 39666
rect 242758 39654 242764 39666
rect 242816 39654 242822 39706
rect 251958 39654 251964 39706
rect 252016 39694 252022 39706
rect 253798 39694 253804 39706
rect 252016 39666 253804 39694
rect 252016 39654 252022 39666
rect 253798 39654 253804 39666
rect 253856 39654 253862 39706
<< via1 >>
rect 311396 995462 311448 995514
rect 312776 995462 312828 995514
rect 466968 995462 467020 995514
rect 473776 995462 473828 995514
rect 467704 995258 467756 995310
rect 475616 995258 475668 995310
rect 250400 994170 250452 994222
rect 256656 994170 256708 994222
rect 259048 994170 259100 994222
rect 82408 993558 82460 993610
rect 136964 993558 137016 993610
rect 191612 993558 191664 993610
rect 195936 993558 195988 993610
rect 203940 993558 203992 993610
rect 86732 993490 86784 993542
rect 94736 993490 94788 993542
rect 100072 993490 100124 993542
rect 102924 993490 102976 993542
rect 81764 993422 81816 993474
rect 93724 993422 93776 993474
rect 115712 993422 115764 993474
rect 136320 993490 136372 993542
rect 202100 993490 202152 993542
rect 250400 993558 250452 993610
rect 250492 993558 250544 993610
rect 258496 993558 258548 993610
rect 259048 993558 259100 993610
rect 312776 993558 312828 993610
rect 437804 993558 437856 993610
rect 450592 993558 450644 993610
rect 517292 993558 517344 993610
rect 518028 993558 518080 993610
rect 625760 993558 625812 993610
rect 626220 993558 626272 993610
rect 630544 993558 630596 993610
rect 638548 993558 638600 993610
rect 222616 993490 222668 993542
rect 141288 993422 141340 993474
rect 149292 993422 149344 993474
rect 136320 993354 136372 993406
rect 157940 993422 157992 993474
rect 158124 993422 158176 993474
rect 170912 993422 170964 993474
rect 171004 993422 171056 993474
rect 178364 993422 178416 993474
rect 209828 993422 209880 993474
rect 222432 993354 222484 993406
rect 248376 993490 248428 993542
rect 261164 993490 261216 993542
rect 312592 993490 312644 993542
rect 408088 993490 408140 993542
rect 462736 993490 462788 993542
rect 528516 993490 528568 993542
rect 636708 993490 636760 993542
rect 273952 993422 274004 993474
rect 274044 993422 274096 993474
rect 287016 993422 287068 993474
rect 245524 993354 245576 993406
rect 248284 993354 248336 993406
rect 92712 993286 92764 993338
rect 92896 993286 92948 993338
rect 147452 993286 147504 993338
rect 93724 993218 93776 993270
rect 100072 993218 100124 993270
rect 202100 993286 202152 993338
rect 209736 993286 209788 993338
rect 191612 993150 191664 993202
rect 209552 993150 209604 993202
rect 178548 993082 178600 993134
rect 190968 993082 191020 993134
rect 209828 993082 209880 993134
rect 274044 993286 274096 993338
rect 286832 993286 286884 993338
rect 295848 993150 295900 993202
rect 299804 993422 299856 993474
rect 300816 993422 300868 993474
rect 353164 993422 353216 993474
rect 406616 993422 406668 993474
rect 463380 993422 463432 993474
rect 517292 993422 517344 993474
rect 517384 993422 517436 993474
rect 625576 993422 625628 993474
rect 305140 993354 305192 993406
rect 313144 993354 313196 993406
rect 419128 993354 419180 993406
rect 334672 993218 334724 993270
rect 338352 993218 338404 993270
rect 338444 993218 338496 993270
rect 300172 993150 300224 993202
rect 312776 993150 312828 993202
rect 321884 993150 321936 993202
rect 360432 993218 360484 993270
rect 364112 993218 364164 993270
rect 364204 993218 364256 993270
rect 347644 993150 347696 993202
rect 386192 993218 386244 993270
rect 389872 993218 389924 993270
rect 389964 993218 390016 993270
rect 373404 993150 373456 993202
rect 419128 993218 419180 993270
rect 437804 993286 437856 993338
rect 450592 993286 450644 993338
rect 466968 993286 467020 993338
rect 528516 993354 528568 993406
rect 473868 993218 473920 993270
rect 522352 993286 522404 993338
rect 530356 993286 530408 993338
rect 312592 993082 312644 993134
rect 257392 992946 257444 992998
rect 296032 992946 296084 992998
rect 299712 992946 299764 992998
rect 244604 992810 244656 992862
rect 636708 992810 636760 992862
rect 675164 992810 675216 992862
rect 625760 992742 625812 992794
rect 675348 992742 675400 992794
rect 244604 992674 244656 992726
rect 246168 992674 246220 992726
rect 257392 992674 257444 992726
rect 625576 992674 625628 992726
rect 675256 992674 675308 992726
rect 81672 992334 81724 992386
rect 82408 992334 82460 992386
rect 364204 975198 364256 975250
rect 364388 975198 364440 975250
rect 581324 975198 581376 975250
rect 581508 975198 581560 975250
rect 42112 970574 42164 970626
rect 92712 970574 92764 970626
rect 41652 968126 41704 968178
rect 42296 968126 42348 968178
rect 41652 967242 41704 967294
rect 42204 967242 42256 967294
rect 674980 966018 675032 966070
rect 675348 966018 675400 966070
rect 675072 965950 675124 966002
rect 675256 965950 675308 966002
rect 675164 963978 675216 964030
rect 675164 963774 675216 963826
rect 674980 962958 675032 963010
rect 675256 962958 675308 963010
rect 42020 962414 42072 962466
rect 42204 962414 42256 962466
rect 675164 962346 675216 962398
rect 675164 962142 675216 962194
rect 42112 961870 42164 961922
rect 42296 961870 42348 961922
rect 43032 960102 43084 960154
rect 364388 960102 364440 960154
rect 99612 960034 99664 960086
rect 632936 960034 632988 960086
rect 674796 958606 674848 958658
rect 675164 958606 675216 958658
rect 41652 955818 41704 955870
rect 42388 955818 42440 955870
rect 41652 955274 41704 955326
rect 42204 955274 42256 955326
rect 632936 954934 632988 954986
rect 641032 954934 641084 954986
rect 93908 953778 93960 953830
rect 99612 953778 99664 953830
rect 41652 953030 41704 953082
rect 42388 953030 42440 953082
rect 81672 953030 81724 953082
rect 42204 952962 42256 953014
rect 81764 952962 81816 953014
rect 674796 951874 674848 951926
rect 675256 951874 675308 951926
rect 92436 951330 92488 951382
rect 93908 951330 93960 951382
rect 581324 949426 581376 949478
rect 581508 949426 581560 949478
rect 674796 948542 674848 948594
rect 675164 948542 675216 948594
rect 641032 947590 641084 947642
rect 646644 947522 646696 947574
rect 646644 943374 646696 943426
rect 653912 943374 653964 943426
rect 90044 941130 90096 941182
rect 92436 941130 92488 941182
rect 88204 937458 88256 937510
rect 90044 937458 90096 937510
rect 87008 934738 87060 934790
rect 88204 934738 88256 934790
rect 653912 934738 653964 934790
rect 655752 934738 655804 934790
rect 80844 931882 80896 931934
rect 87008 931882 87060 931934
rect 44044 926442 44096 926494
rect 80844 926442 80896 926494
rect 39260 925558 39312 925610
rect 44044 925558 44096 925610
rect 581324 923722 581376 923774
rect 581508 923722 581560 923774
rect 655752 919982 655804 920034
rect 661272 919914 661324 919966
rect 39628 913250 39680 913302
rect 40456 913250 40508 913302
rect 41652 913250 41704 913302
rect 661272 908898 661324 908950
rect 669460 908898 669512 908950
rect 675348 908898 675400 908950
rect 677556 908898 677608 908950
rect 669460 905294 669512 905346
rect 677556 905226 677608 905278
rect 674520 875306 674572 875358
rect 675072 875306 675124 875358
rect 675164 875034 675216 875086
rect 675348 875034 675400 875086
rect 674980 873742 675032 873794
rect 675256 873742 675308 873794
rect 41928 872178 41980 872230
rect 42112 872178 42164 872230
rect 581324 872178 581376 872230
rect 581508 872178 581560 872230
rect 674980 871702 675032 871754
rect 675256 871702 675308 871754
rect 675164 870138 675216 870190
rect 675164 869934 675216 869986
rect 674888 866738 674940 866790
rect 675164 866738 675216 866790
rect 39720 865786 39772 865838
rect 40456 865786 40508 865838
rect 41652 865786 41704 865838
rect 674520 862998 674572 863050
rect 674612 862998 674664 863050
rect 674888 860618 674940 860670
rect 675256 860618 675308 860670
rect 674612 853682 674664 853734
rect 674980 853682 675032 853734
rect 675256 850010 675308 850062
rect 675348 850010 675400 850062
rect 41744 846474 41796 846526
rect 41928 846474 41980 846526
rect 581324 846406 581376 846458
rect 581508 846406 581560 846458
rect 674888 840898 674940 840950
rect 674980 840830 675032 840882
rect 41744 837226 41796 837278
rect 42020 837226 42072 837278
rect 674888 837226 674940 837278
rect 674980 837226 675032 837278
rect 675256 837226 675308 837278
rect 675532 837226 675584 837278
rect 675164 836138 675216 836190
rect 675440 836138 675492 836190
rect 42020 828046 42072 828098
rect 675256 827978 675308 828030
rect 675532 827978 675584 828030
rect 41928 827910 41980 827962
rect 573964 821518 574016 821570
rect 674980 821518 675032 821570
rect 675164 821518 675216 821570
rect 675440 821518 675492 821570
rect 581324 820634 581376 820686
rect 581508 820634 581560 820686
rect 581324 817846 581376 817898
rect 674888 817846 674940 817898
rect 675256 811386 675308 811438
rect 675348 811386 675400 811438
rect 674704 809550 674756 809602
rect 674888 809550 674940 809602
rect 675164 808258 675216 808310
rect 675440 808258 675492 808310
rect 675348 798602 675400 798654
rect 675532 798602 675584 798654
rect 674704 796698 674756 796750
rect 674888 796698 674940 796750
rect 675164 795746 675216 795798
rect 675440 795746 675492 795798
rect 41928 793910 41980 793962
rect 42572 793910 42624 793962
rect 41652 791122 41704 791174
rect 42572 791122 42624 791174
rect 674796 790442 674848 790494
rect 675072 790442 675124 790494
rect 674796 782894 674848 782946
rect 675072 782894 675124 782946
rect 42112 782078 42164 782130
rect 42572 782078 42624 782130
rect 41652 781874 41704 781926
rect 41652 781670 41704 781722
rect 674520 781534 674572 781586
rect 675532 781534 675584 781586
rect 674520 778950 674572 779002
rect 675256 778950 675308 779002
rect 674704 778542 674756 778594
rect 675164 778542 675216 778594
rect 674796 774190 674848 774242
rect 675164 774190 675216 774242
rect 674612 770042 674664 770094
rect 675072 770042 675124 770094
rect 674704 768478 674756 768530
rect 675256 768478 675308 768530
rect 675164 767594 675216 767646
rect 675164 767390 675216 767442
rect 674796 765962 674848 766014
rect 675532 765962 675584 766014
rect 674520 765894 674572 765946
rect 675256 765894 675308 765946
rect 674428 759978 674480 760030
rect 674888 759978 674940 760030
rect 674704 758006 674756 758058
rect 674888 758006 674940 758058
rect 675532 758006 675584 758058
rect 675716 758006 675768 758058
rect 674612 757122 674664 757174
rect 675072 757122 675124 757174
rect 42112 749778 42164 749830
rect 42572 749778 42624 749830
rect 41652 748350 41704 748402
rect 42664 748350 42716 748402
rect 41836 747126 41888 747178
rect 42572 747126 42624 747178
rect 41836 746514 41888 746566
rect 42572 746514 42624 746566
rect 674796 744270 674848 744322
rect 674980 744270 675032 744322
rect 42112 743386 42164 743438
rect 42664 743386 42716 743438
rect 41652 741414 41704 741466
rect 42112 741414 42164 741466
rect 674612 735294 674664 735346
rect 675072 735294 675124 735346
rect 674704 735226 674756 735278
rect 675164 735226 675216 735278
rect 674888 734342 674940 734394
rect 674888 734206 674940 734258
rect 42112 733254 42164 733306
rect 42572 733254 42624 733306
rect 675164 725298 675216 725350
rect 675072 725026 675124 725078
rect 674612 724958 674664 725010
rect 674980 724958 675032 725010
rect 674704 722034 674756 722086
rect 675256 722034 675308 722086
rect 674428 721898 674480 721950
rect 674704 721898 674756 721950
rect 41744 721286 41796 721338
rect 42020 721286 42072 721338
rect 675072 720198 675124 720250
rect 675256 720198 675308 720250
rect 674612 714894 674664 714946
rect 674980 714894 675032 714946
rect 674704 708502 674756 708554
rect 674888 708502 674940 708554
rect 674612 708366 674664 708418
rect 675072 708366 675124 708418
rect 675164 708366 675216 708418
rect 675348 708366 675400 708418
rect 674704 706530 674756 706582
rect 674888 706530 674940 706582
rect 675164 705646 675216 705698
rect 675440 705646 675492 705698
rect 41652 702178 41704 702230
rect 42112 702178 42164 702230
rect 42572 702178 42624 702230
rect 675348 699186 675400 699238
rect 675624 699118 675676 699170
rect 674704 693678 674756 693730
rect 674888 693678 674940 693730
rect 674796 692182 674848 692234
rect 674980 692182 675032 692234
rect 41652 691094 41704 691146
rect 42112 691094 42164 691146
rect 41652 688986 41704 689038
rect 42112 688986 42164 689038
rect 674704 688714 674756 688766
rect 675164 688714 675216 688766
rect 675164 688578 675216 688630
rect 675624 688578 675676 688630
rect 674888 686402 674940 686454
rect 674796 686266 674848 686318
rect 674520 682594 674572 682646
rect 674796 682594 674848 682646
rect 674888 681166 674940 681218
rect 675164 681166 675216 681218
rect 674520 680010 674572 680062
rect 674796 680010 674848 680062
rect 674520 679874 674572 679926
rect 674980 679874 675032 679926
rect 674428 675454 674480 675506
rect 675256 675454 675308 675506
rect 41928 673550 41980 673602
rect 41836 673346 41888 673398
rect 674980 672938 675032 672990
rect 675256 672938 675308 672990
rect 674796 672870 674848 672922
rect 675624 672870 675676 672922
rect 674428 672802 674480 672854
rect 675348 672802 675400 672854
rect 674520 666954 674572 667006
rect 674980 666954 675032 667006
rect 42112 660154 42164 660206
rect 42572 660154 42624 660206
rect 41652 660018 41704 660070
rect 42112 660018 42164 660070
rect 42020 653218 42072 653270
rect 42664 653218 42716 653270
rect 41652 648050 41704 648102
rect 42572 648050 42624 648102
rect 42020 647642 42072 647694
rect 41652 647438 41704 647490
rect 42020 647438 42072 647490
rect 42112 644446 42164 644498
rect 41652 644378 41704 644430
rect 42112 644310 42164 644362
rect 42572 644310 42624 644362
rect 674796 641998 674848 642050
rect 675256 641998 675308 642050
rect 674704 641182 674756 641234
rect 674980 641182 675032 641234
rect 674796 638938 674848 638990
rect 675256 638938 675308 638990
rect 674704 628330 674756 628382
rect 674980 628330 675032 628382
rect 41560 627378 41612 627430
rect 41744 627378 41796 627430
rect 674796 626358 674848 626410
rect 675256 626358 675308 626410
rect 674796 615478 674848 615530
rect 674980 615478 675032 615530
rect 42112 615410 42164 615462
rect 42572 615410 42624 615462
rect 41652 612894 41704 612946
rect 42572 612894 42624 612946
rect 675348 609018 675400 609070
rect 675532 609018 675584 609070
rect 42112 608950 42164 609002
rect 42572 608950 42624 609002
rect 674796 602558 674848 602610
rect 674980 602558 675032 602610
rect 41560 599498 41612 599550
rect 42112 599770 42164 599822
rect 674796 595486 674848 595538
rect 675256 595486 675308 595538
rect 674428 595418 674480 595470
rect 675164 595418 675216 595470
rect 674796 592358 674848 592410
rect 675256 592358 675308 592410
rect 674704 587394 674756 587446
rect 675256 587394 675308 587446
rect 674796 583450 674848 583502
rect 675256 583314 675308 583366
rect 674796 580390 674848 580442
rect 675256 580390 675308 580442
rect 674428 579778 674480 579830
rect 675256 579778 675308 579830
rect 41560 579642 41612 579694
rect 41836 579642 41888 579694
rect 41652 576786 41704 576838
rect 42020 576786 42072 576838
rect 42112 571074 42164 571126
rect 42572 571074 42624 571126
rect 677464 566722 677516 566774
rect 677740 566722 677792 566774
rect 41652 559038 41704 559090
rect 42572 559038 42624 559090
rect 675164 557406 675216 557458
rect 675440 557406 675492 557458
rect 41744 551218 41796 551270
rect 42112 551218 42164 551270
rect 674520 551082 674572 551134
rect 674980 551082 675032 551134
rect 675164 551082 675216 551134
rect 675348 551082 675400 551134
rect 674796 548838 674848 548890
rect 675440 548838 675492 548890
rect 674980 548770 675032 548822
rect 675256 548770 675308 548822
rect 674796 546662 674848 546714
rect 675256 546662 675308 546714
rect 674980 546118 675032 546170
rect 675348 546118 675400 546170
rect 674612 545098 674664 545150
rect 675256 545098 675308 545150
rect 674980 541426 675032 541478
rect 675164 541426 675216 541478
rect 674980 535646 675032 535698
rect 675256 535646 675308 535698
rect 674520 535510 674572 535562
rect 674980 535510 675032 535562
rect 674796 533198 674848 533250
rect 675164 533198 675216 533250
rect 674612 533062 674664 533114
rect 675256 533062 675308 533114
rect 674796 530818 674848 530870
rect 674980 530818 675032 530870
rect 41744 526398 41796 526450
rect 42572 526398 42624 526450
rect 41652 523882 41704 523934
rect 42572 523882 42624 523934
rect 42112 518238 42164 518290
rect 42572 518238 42624 518290
rect 674796 511506 674848 511558
rect 674980 511506 675032 511558
rect 41652 499538 41704 499590
rect 42112 499538 42164 499590
rect 674612 498586 674664 498638
rect 674888 498586 674940 498638
rect 674796 498518 674848 498570
rect 674980 498518 675032 498570
rect 674704 472814 674756 472866
rect 674980 472814 675032 472866
rect 674704 454454 674756 454506
rect 674888 454454 674940 454506
rect 675256 447042 675308 447094
rect 677556 447042 677608 447094
rect 41836 441602 41888 441654
rect 42020 441602 42072 441654
rect 39260 439766 39312 439818
rect 44044 439766 44096 439818
rect 44872 439766 44924 439818
rect 675348 437930 675400 437982
rect 677924 437930 677976 437982
rect 675348 430586 675400 430638
rect 672404 430518 672456 430570
rect 39628 428546 39680 428598
rect 41836 428546 41888 428598
rect 42020 428546 42072 428598
rect 41560 425010 41612 425062
rect 42020 425010 42072 425062
rect 674888 425010 674940 425062
rect 675072 425010 675124 425062
rect 668632 423174 668684 423226
rect 672404 423242 672456 423294
rect 41560 412158 41612 412210
rect 41836 412158 41888 412210
rect 664676 408486 664728 408538
rect 668632 408486 668684 408538
rect 663112 404814 663164 404866
rect 664676 404814 664728 404866
rect 41836 399238 41888 399290
rect 42296 399238 42348 399290
rect 41652 394886 41704 394938
rect 42388 394886 42440 394938
rect 41744 394818 41796 394870
rect 42480 394818 42532 394870
rect 41652 394138 41704 394190
rect 42112 394138 42164 394190
rect 41652 392710 41704 392762
rect 42388 392710 42440 392762
rect 41652 387202 41704 387254
rect 42112 387202 42164 387254
rect 42112 386726 42164 386778
rect 42480 386726 42532 386778
rect 41652 381830 41704 381882
rect 42112 381830 42164 381882
rect 42296 381830 42348 381882
rect 41652 379178 41704 379230
rect 42112 379178 42164 379230
rect 42020 374350 42072 374402
rect 42388 374350 42440 374402
rect 675164 365714 675216 365766
rect 675164 365510 675216 365562
rect 42020 364354 42072 364406
rect 42020 364218 42072 364270
rect 675072 362926 675124 362978
rect 675256 362926 675308 362978
rect 675164 362042 675216 362094
rect 675164 361838 675216 361890
rect 660444 358982 660496 359034
rect 663112 358982 663164 359034
rect 674888 357554 674940 357606
rect 675256 357554 675308 357606
rect 675072 357146 675124 357198
rect 675164 356942 675216 356994
rect 674796 356874 674848 356926
rect 675072 356874 675124 356926
rect 42020 352182 42072 352234
rect 42388 352182 42440 352234
rect 41652 350278 41704 350330
rect 42112 350278 42164 350330
rect 41744 350210 41796 350262
rect 42572 350210 42624 350262
rect 657132 350006 657184 350058
rect 660352 350006 660404 350058
rect 674980 349938 675032 349990
rect 675348 349938 675400 349990
rect 674796 349870 674848 349922
rect 675256 349870 675308 349922
rect 41652 349530 41704 349582
rect 42296 349530 42348 349582
rect 41836 348646 41888 348698
rect 42388 348646 42440 348698
rect 41836 347694 41888 347746
rect 42388 347694 42440 347746
rect 655752 344770 655804 344822
rect 657132 344770 657184 344822
rect 42112 344566 42164 344618
rect 42480 344566 42532 344618
rect 42112 344430 42164 344482
rect 42296 344430 42348 344482
rect 42388 344158 42440 344210
rect 42388 343954 42440 344006
rect 41652 338242 41704 338294
rect 42112 338242 42164 338294
rect 42480 338242 42532 338294
rect 41652 337630 41704 337682
rect 42572 337630 42624 337682
rect 41836 335114 41888 335166
rect 42572 335114 42624 335166
rect 41836 334842 41888 334894
rect 41652 334570 41704 334622
rect 42112 334366 42164 334418
rect 42388 334366 42440 334418
rect 41652 333958 41704 334010
rect 42020 333958 42072 334010
rect 651244 331170 651296 331222
rect 655752 331238 655804 331290
rect 649404 319338 649456 319390
rect 651244 319338 651296 319390
rect 675164 319066 675216 319118
rect 675164 318862 675216 318914
rect 675072 316346 675124 316398
rect 675256 316346 675308 316398
rect 640848 313830 640900 313882
rect 649404 313830 649456 313882
rect 41560 312810 41612 312862
rect 41744 312810 41796 312862
rect 41928 312810 41980 312862
rect 42020 312742 42072 312794
rect 636892 310226 636944 310278
rect 640848 310226 640900 310278
rect 41928 309138 41980 309190
rect 42020 309138 42072 309190
rect 674888 309070 674940 309122
rect 675072 309070 675124 309122
rect 634684 306418 634736 306470
rect 636892 306418 636944 306470
rect 41928 305874 41980 305926
rect 42388 305874 42440 305926
rect 42112 305330 42164 305382
rect 42296 305330 42348 305382
rect 41836 305126 41888 305178
rect 42112 305126 42164 305178
rect 674980 304922 675032 304974
rect 675256 304922 675308 304974
rect 674980 303358 675032 303410
rect 675440 303358 675492 303410
rect 41652 303290 41704 303342
rect 42388 303290 42440 303342
rect 630360 299890 630412 299942
rect 634684 299958 634736 300010
rect 674888 296218 674940 296270
rect 675348 296218 675400 296270
rect 620700 294246 620752 294298
rect 630360 294382 630412 294434
rect 41652 293566 41704 293618
rect 42112 293566 42164 293618
rect 42112 293430 42164 293482
rect 42388 293430 42440 293482
rect 41928 287378 41980 287430
rect 42112 287378 42164 287430
rect 615548 286290 615600 286342
rect 620700 286290 620752 286342
rect 613432 284114 613484 284166
rect 615548 284114 615600 284166
rect 609752 275954 609804 276006
rect 613432 276022 613484 276074
rect 674796 274118 674848 274170
rect 675164 274118 675216 274170
rect 675164 272554 675216 272606
rect 675440 272554 675492 272606
rect 675532 270718 675584 270770
rect 675440 270514 675492 270566
rect 674980 269562 675032 269614
rect 675256 269562 675308 269614
rect 674796 268882 674848 268934
rect 675256 268882 675308 268934
rect 42112 266706 42164 266758
rect 42388 266706 42440 266758
rect 41652 266570 41704 266622
rect 42112 266570 42164 266622
rect 605336 264938 605388 264990
rect 609752 264938 609804 264990
rect 674888 264666 674940 264718
rect 675164 264666 675216 264718
rect 600552 262150 600604 262202
rect 605336 262150 605388 262202
rect 41744 261266 41796 261318
rect 42664 261266 42716 261318
rect 41652 260518 41704 260570
rect 42296 260518 42348 260570
rect 41652 259634 41704 259686
rect 42388 259634 42440 259686
rect 675164 259498 675216 259550
rect 675164 259294 675216 259346
rect 674888 259226 674940 259278
rect 675256 259226 675308 259278
rect 674888 257594 674940 257646
rect 675348 257594 675400 257646
rect 675348 257186 675400 257238
rect 674980 257050 675032 257102
rect 675348 256982 675400 257034
rect 675532 256982 675584 257034
rect 42296 254126 42348 254178
rect 42388 254058 42440 254110
rect 42296 253922 42348 253974
rect 42664 253922 42716 253974
rect 42388 253854 42440 253906
rect 41652 253582 41704 253634
rect 594112 248346 594164 248398
rect 600552 248414 600604 248466
rect 41928 245558 41980 245610
rect 42388 245558 42440 245610
rect 41652 245490 41704 245542
rect 42112 245490 42164 245542
rect 590432 242838 590484 242890
rect 594112 242906 594164 242958
rect 675164 241002 675216 241054
rect 675440 241002 675492 241054
rect 587672 234882 587724 234934
rect 590432 234882 590484 234934
rect 41928 228150 41980 228202
rect 42112 228150 42164 228202
rect 674980 226042 675032 226094
rect 675440 226042 675492 226094
rect 674888 225974 674940 226026
rect 675532 225974 675584 226026
rect 674980 223322 675032 223374
rect 675348 223322 675400 223374
rect 675256 222914 675308 222966
rect 675164 222642 675216 222694
rect 585832 221418 585884 221470
rect 587672 221418 587724 221470
rect 42112 216658 42164 216710
rect 42480 216658 42532 216710
rect 41652 215978 41704 216030
rect 42296 215978 42348 216030
rect 42480 215230 42532 215282
rect 42112 215162 42164 215214
rect 42388 215162 42440 215214
rect 41652 215094 41704 215146
rect 674888 210334 674940 210386
rect 675256 210334 675308 210386
rect 674980 210198 675032 210250
rect 675348 210198 675400 210250
rect 42112 209722 42164 209774
rect 41652 209518 41704 209570
rect 41652 208974 41704 209026
rect 42296 208974 42348 209026
rect 581508 206050 581560 206102
rect 585832 206118 585884 206170
rect 41652 203058 41704 203110
rect 42388 203058 42440 203110
rect 578104 200610 578156 200662
rect 581508 200610 581560 200662
rect 573964 198706 574016 198758
rect 578104 198706 578156 198758
rect 41836 193198 41888 193250
rect 42388 193198 42440 193250
rect 570652 191906 570704 191958
rect 573964 191906 574016 191958
rect 675164 189390 675216 189442
rect 675348 189390 675400 189442
rect 566604 187690 566656 187742
rect 570652 187690 570704 187742
rect 41836 184018 41888 184070
rect 41928 183882 41980 183934
rect 674980 179802 675032 179854
rect 675624 179802 675676 179854
rect 675164 179666 675216 179718
rect 675716 179666 675768 179718
rect 555012 178510 555064 178562
rect 566512 178510 566564 178562
rect 675072 176742 675124 176794
rect 675348 176742 675400 176794
rect 674888 175654 674940 175706
rect 675256 175654 675308 175706
rect 41928 172254 41980 172306
rect 42388 172254 42440 172306
rect 41652 172186 41704 172238
rect 42296 172186 42348 172238
rect 552160 167562 552212 167614
rect 555012 167562 555064 167614
rect 674796 167358 674848 167410
rect 674980 167358 675032 167410
rect 674796 165318 674848 165370
rect 675256 165318 675308 165370
rect 550044 164842 550096 164894
rect 552160 164842 552212 164894
rect 42296 164094 42348 164146
rect 42020 163958 42072 164010
rect 674888 163754 674940 163806
rect 675348 163754 675400 163806
rect 41652 158994 41704 159046
rect 42296 158994 42348 159046
rect 675164 157294 675216 157346
rect 675440 157294 675492 157346
rect 674796 157158 674848 157210
rect 675164 157158 675216 157210
rect 546364 155730 546416 155782
rect 550044 155730 550096 155782
rect 42296 155458 42348 155510
rect 87192 155458 87244 155510
rect 42480 154574 42532 154626
rect 42572 154574 42624 154626
rect 42296 154438 42348 154490
rect 42480 154438 42532 154490
rect 542684 151786 542736 151838
rect 546364 151786 546416 151838
rect 540016 143490 540068 143542
rect 542684 143558 542736 143610
rect 42296 141722 42348 141774
rect 42572 141722 42624 141774
rect 87192 141654 87244 141706
rect 88664 141654 88716 141706
rect 675164 137914 675216 137966
rect 675532 137914 675584 137966
rect 88664 134310 88716 134362
rect 90872 134310 90924 134362
rect 674888 132814 674940 132866
rect 675532 132814 675584 132866
rect 675348 132746 675400 132798
rect 675440 132746 675492 132798
rect 675072 132678 675124 132730
rect 675532 132542 675584 132594
rect 42388 132474 42440 132526
rect 42572 132474 42624 132526
rect 674980 129074 675032 129126
rect 675256 129074 675308 129126
rect 42388 128734 42440 128786
rect 42480 128734 42532 128786
rect 675164 124858 675216 124910
rect 675164 124654 675216 124706
rect 674888 119894 674940 119946
rect 675164 119894 675216 119946
rect 675072 119826 675124 119878
rect 42480 119622 42532 119674
rect 675164 119622 675216 119674
rect 42388 119554 42440 119606
rect 90872 118738 90924 118790
rect 92528 118738 92580 118790
rect 674888 118670 674940 118722
rect 675256 118670 675308 118722
rect 675072 117242 675124 117294
rect 675532 117174 675584 117226
rect 39904 115950 39956 116002
rect 40364 115950 40416 116002
rect 42112 115950 42164 116002
rect 92528 115882 92580 115934
rect 94000 115882 94052 115934
rect 42204 109422 42256 109474
rect 42480 109422 42532 109474
rect 94000 108538 94052 108590
rect 97404 108470 97456 108522
rect 97404 102486 97456 102538
rect 99704 102486 99756 102538
rect 44872 100106 44924 100158
rect 45792 100106 45844 100158
rect 45792 99902 45844 99954
rect 540108 99902 540160 99954
rect 99704 99834 99756 99886
rect 126844 99834 126896 99886
rect 126844 95686 126896 95738
rect 130984 95618 131036 95670
rect 42204 93782 42256 93834
rect 42388 93782 42440 93834
rect 130984 91946 131036 91998
rect 135032 91946 135084 91998
rect 42112 90110 42164 90162
rect 42388 90110 42440 90162
rect 674796 86302 674848 86354
rect 675532 86302 675584 86354
rect 675164 86234 675216 86286
rect 675164 86030 675216 86082
rect 45148 85554 45200 85606
rect 45792 85554 45844 85606
rect 465496 85554 465548 85606
rect 39260 84670 39312 84722
rect 45148 84670 45200 84722
rect 674796 83786 674848 83838
rect 675256 83786 675308 83838
rect 135032 83582 135084 83634
rect 136044 83582 136096 83634
rect 675072 83514 675124 83566
rect 675256 83514 675308 83566
rect 674888 82494 674940 82546
rect 675256 82494 675308 82546
rect 42112 77258 42164 77310
rect 42296 77258 42348 77310
rect 43952 76306 44004 76358
rect 149752 76306 149804 76358
rect 136044 74606 136096 74658
rect 138804 74606 138856 74658
rect 674888 73994 674940 74046
rect 674980 73790 675032 73842
rect 674796 73654 674848 73706
rect 675164 73654 675216 73706
rect 675164 73518 675216 73570
rect 675072 73246 675124 73298
rect 39720 72634 39772 72686
rect 90872 72634 90924 72686
rect 674888 72090 674940 72142
rect 675256 72090 675308 72142
rect 39536 67126 39588 67178
rect 140552 67126 140604 67178
rect 138804 66174 138856 66226
rect 140644 66174 140696 66226
rect 140644 62502 140696 62554
rect 142392 62502 142444 62554
rect 670288 45910 670340 45962
rect 675164 45910 675216 45962
rect 43032 45026 43084 45078
rect 183792 45094 183844 45146
rect 183884 45026 183936 45078
rect 195844 45094 195896 45146
rect 196672 45094 196724 45146
rect 515084 45094 515136 45146
rect 516188 45094 516240 45146
rect 527320 45094 527372 45146
rect 675348 45094 675400 45146
rect 540844 45026 540896 45078
rect 553632 44958 553684 45010
rect 196672 44686 196724 44738
rect 209552 44686 209604 44738
rect 209644 44686 209696 44738
rect 218844 44754 218896 44806
rect 231632 44686 231684 44738
rect 235312 44686 235364 44738
rect 235404 44686 235456 44738
rect 244604 44754 244656 44806
rect 257392 44686 257444 44738
rect 261072 44686 261124 44738
rect 261164 44686 261216 44738
rect 273952 44754 274004 44806
rect 417472 44754 417524 44806
rect 424924 44754 424976 44806
rect 274136 44686 274188 44738
rect 307440 44686 307492 44738
rect 318112 44686 318164 44738
rect 344792 44686 344844 44738
rect 351784 44686 351836 44738
rect 359236 44686 359288 44738
rect 283152 44618 283204 44670
rect 283336 44550 283388 44602
rect 299620 44618 299672 44670
rect 437712 44686 437764 44738
rect 441392 44686 441444 44738
rect 515084 44754 515136 44806
rect 570192 44754 570244 44806
rect 570284 44754 570336 44806
rect 592272 44754 592324 44806
rect 595952 44754 596004 44806
rect 596044 44754 596096 44806
rect 308084 44550 308136 44602
rect 358592 44550 358644 44602
rect 195200 44482 195252 44534
rect 199524 44482 199576 44534
rect 303760 44482 303812 44534
rect 318112 44482 318164 44534
rect 331084 44482 331136 44534
rect 362824 44482 362876 44534
rect 376992 44550 377044 44602
rect 377176 44550 377228 44602
rect 200720 44414 200772 44466
rect 242764 44414 242816 44466
rect 306244 44414 306296 44466
rect 309280 44414 309332 44466
rect 352428 44414 352480 44466
rect 355464 44414 355516 44466
rect 361076 44414 361128 44466
rect 364112 44414 364164 44466
rect 407260 44414 407312 44466
rect 410296 44414 410348 44466
rect 413884 44618 413936 44670
rect 441576 44618 441628 44670
rect 450684 44618 450736 44670
rect 459516 44618 459568 44670
rect 467520 44618 467572 44670
rect 471844 44618 471896 44670
rect 473776 44618 473828 44670
rect 473868 44618 473920 44670
rect 480124 44618 480176 44670
rect 489232 44618 489284 44670
rect 579484 44686 579536 44738
rect 618032 44754 618084 44806
rect 621712 44754 621764 44806
rect 621804 44754 621856 44806
rect 605244 44686 605296 44738
rect 643792 44754 643844 44806
rect 647472 44754 647524 44806
rect 647564 44754 647616 44806
rect 631004 44686 631056 44738
rect 669552 44754 669604 44806
rect 670288 44754 670340 44806
rect 656764 44686 656816 44738
rect 463472 44550 463524 44602
rect 413884 44482 413936 44534
rect 414068 44482 414120 44534
rect 468808 44482 468860 44534
rect 476352 44482 476404 44534
rect 515084 44482 515136 44534
rect 412964 44414 413016 44466
rect 419036 44414 419088 44466
rect 462000 44414 462052 44466
rect 465036 44414 465088 44466
rect 465496 44414 465548 44466
rect 473592 44414 473644 44466
rect 516832 44414 516884 44466
rect 519868 44414 519920 44466
rect 201364 44346 201416 44398
rect 244512 44346 244564 44398
rect 296952 44346 297004 44398
rect 299436 44346 299488 44398
rect 305600 44346 305652 44398
rect 344792 44346 344844 44398
rect 344884 44346 344936 44398
rect 362272 44346 362324 44398
rect 362824 44346 362876 44398
rect 362916 44346 362968 44398
rect 413424 44346 413476 44398
rect 417748 44346 417800 44398
rect 468164 44346 468216 44398
rect 472488 44346 472540 44398
rect 522996 44346 523048 44398
rect 90872 44278 90924 44330
rect 198880 44278 198932 44330
rect 247088 44278 247140 44330
rect 307440 44278 307492 44330
rect 331084 44278 331136 44330
rect 334764 44278 334816 44330
rect 351784 44278 351836 44330
rect 354268 44278 354320 44330
rect 360432 44278 360484 44330
rect 406616 44278 406668 44330
rect 461356 44278 461408 44330
rect 473868 44278 473920 44330
rect 518672 44278 518724 44330
rect 524836 44278 524888 44330
rect 525940 44278 525992 44330
rect 568996 44278 569048 44330
rect 148924 44210 148976 44262
rect 149752 44210 149804 44262
rect 188392 44210 188444 44262
rect 192716 44210 192768 44262
rect 201364 44210 201416 44262
rect 304404 44210 304456 44262
rect 338352 44210 338404 44262
rect 338536 44210 338588 44262
rect 359236 44210 359288 44262
rect 410940 44210 410992 44262
rect 186552 44142 186604 44194
rect 194556 44142 194608 44194
rect 295112 44142 295164 44194
rect 303116 44142 303168 44194
rect 349944 44142 349996 44194
rect 357948 44142 358000 44194
rect 358592 44142 358644 44194
rect 362916 44142 362968 44194
rect 404776 44142 404828 44194
rect 412780 44142 412832 44194
rect 412964 44210 413016 44262
rect 417104 44210 417156 44262
rect 417472 44210 417524 44262
rect 473776 44210 473828 44262
rect 526676 44210 526728 44262
rect 630268 44210 630320 44262
rect 419588 44142 419640 44194
rect 465680 44142 465732 44194
rect 474328 44142 474380 44194
rect 514348 44142 514400 44194
rect 522352 44142 522404 44194
rect 522996 44142 523048 44194
rect 527320 44142 527372 44194
rect 515084 43530 515136 43582
rect 523640 43530 523692 43582
rect 525940 43530 525992 43582
rect 142392 43326 142444 43378
rect 144968 43326 145020 43378
rect 251320 43190 251372 43242
rect 297596 43190 297648 43242
rect 579484 43190 579536 43242
rect 675256 43190 675308 43242
rect 299620 42442 299672 42494
rect 304404 42442 304456 42494
rect 144968 42374 145020 42426
rect 195200 42374 195252 42426
rect 242764 42374 242816 42426
rect 251320 42374 251372 42426
rect 297596 42374 297648 42426
rect 300632 42374 300684 42426
rect 144416 42306 144468 42358
rect 253804 42306 253856 42358
rect 569088 42306 569140 42358
rect 579484 42306 579536 42358
rect 303760 42238 303812 42290
rect 308084 42238 308136 42290
rect 468164 42238 468216 42290
rect 472488 42238 472540 42290
rect 189128 41898 189180 41950
rect 198328 41830 198380 41882
rect 199984 41830 200036 41882
rect 306152 41898 306204 41950
rect 409192 41830 409244 41882
rect 412228 41830 412280 41882
rect 415080 41830 415132 41882
rect 464024 41830 464076 41882
rect 467060 41830 467112 41882
rect 469912 41830 469964 41882
rect 519960 41830 520012 41882
rect 521248 41830 521300 41882
rect 524284 41830 524336 41882
rect 525572 41830 525624 41882
rect 527780 41830 527832 41882
rect 190968 41762 191020 41814
rect 192164 41762 192216 41814
rect 193452 41762 193504 41814
rect 196304 41762 196356 41814
rect 297136 41762 297188 41814
rect 302104 41762 302156 41814
rect 304864 41762 304916 41814
rect 359880 41762 359932 41814
rect 360984 41762 361036 41814
rect 410388 41762 410440 41814
rect 411400 41762 411452 41814
rect 414436 41762 414488 41814
rect 415724 41762 415776 41814
rect 418116 41762 418168 41814
rect 419036 41762 419088 41814
rect 251964 41558 252016 41610
rect 286924 41558 286976 41610
rect 286924 41354 286976 41406
rect 134112 40130 134164 40182
rect 143404 40130 143456 40182
rect 140860 40062 140912 40114
rect 142936 40062 142988 40114
rect 144416 40062 144468 40114
rect 241108 39654 241160 39706
rect 242764 39654 242816 39706
rect 251964 39654 252016 39706
rect 253804 39654 253856 39706
<< metal2 >>
rect 352150 997658 352206 997667
rect 352150 997593 352206 997602
rect 362192 997531 362220 997630
rect 579404 997531 579432 997630
rect 353162 997522 353218 997531
rect 353162 997457 353218 997466
rect 362178 997522 362234 997531
rect 362178 997457 362234 997466
rect 364386 997522 364442 997531
rect 364386 997457 364442 997466
rect 579390 997522 579446 997531
rect 579390 997457 579446 997466
rect 581506 997522 581562 997531
rect 581506 997457 581562 997466
rect 256668 995636 256718 995664
rect 258508 995636 258558 995664
rect 81776 993480 81804 995454
rect 82420 993616 82448 995454
rect 82408 993610 82460 993616
rect 82408 993552 82460 993558
rect 81764 993474 81816 993480
rect 81764 993416 81816 993422
rect 81672 992386 81724 992392
rect 81672 992328 81724 992334
rect 42112 970626 42164 970632
rect 42112 970568 42164 970574
rect 42124 968812 42152 970568
rect 42124 968784 42244 968812
rect 41586 968682 41692 968710
rect 41664 968184 41692 968682
rect 41652 968178 41704 968184
rect 41652 968120 41704 968126
rect 42216 967300 42244 968784
rect 42296 968178 42348 968184
rect 42296 968120 42348 968126
rect 41652 967294 41704 967300
rect 41652 967236 41704 967242
rect 42204 967294 42256 967300
rect 42204 967236 42256 967242
rect 41664 966870 41692 967236
rect 41586 966842 41692 966870
rect 42216 962472 42244 967236
rect 42020 962466 42072 962472
rect 42020 962408 42072 962414
rect 42204 962466 42256 962472
rect 42204 962408 42256 962414
rect 42032 962012 42060 962408
rect 42032 961984 42244 962012
rect 42112 961922 42164 961928
rect 42112 961864 42164 961870
rect 42124 960788 42152 961864
rect 41664 960760 42152 960788
rect 41664 960706 41692 960760
rect 42216 960706 42244 961984
rect 42308 961928 42336 968120
rect 42296 961922 42348 961928
rect 42296 961864 42348 961870
rect 41586 960678 41692 960706
rect 42124 960678 42244 960706
rect 41586 956354 41692 956382
rect 41664 955876 41692 956354
rect 41652 955870 41704 955876
rect 41652 955812 41704 955818
rect 41586 955728 41692 955756
rect 41664 955332 41692 955728
rect 41652 955326 41704 955332
rect 41652 955268 41704 955274
rect 41652 953082 41704 953088
rect 41652 953024 41704 953030
rect 39260 925610 39312 925616
rect 39260 925552 39312 925558
rect 39272 920396 39300 925552
rect 39194 920368 39300 920396
rect 39718 917146 39774 917155
rect 39718 917081 39774 917090
rect 39417 916424 39668 916452
rect 39417 916302 39445 916424
rect 39640 913308 39668 916424
rect 39732 915251 39760 917081
rect 39718 915242 39774 915251
rect 39718 915177 39774 915186
rect 41664 913308 41692 953024
rect 42124 949364 42152 960678
rect 43032 960154 43084 960160
rect 43032 960096 43084 960102
rect 42388 955870 42440 955876
rect 42388 955812 42440 955818
rect 42204 955326 42256 955332
rect 42204 955268 42256 955274
rect 42216 953020 42244 955268
rect 42400 953088 42428 955812
rect 42388 953082 42440 953088
rect 42388 953024 42440 953030
rect 42204 953014 42256 953020
rect 42204 952956 42256 952962
rect 42032 949336 42152 949364
rect 42032 918220 42060 949336
rect 42032 918192 42152 918220
rect 39628 913302 39680 913308
rect 39628 913244 39680 913250
rect 40456 913302 40508 913308
rect 40456 913244 40508 913250
rect 41652 913302 41704 913308
rect 41652 913244 41704 913250
rect 39180 909624 39392 909652
rect 39180 909502 39208 909624
rect 39364 903691 39392 909624
rect 39350 903682 39406 903691
rect 39350 903617 39406 903626
rect 39470 875896 39944 875924
rect 39916 875811 39944 875896
rect 39902 875802 39958 875811
rect 39902 875737 39958 875746
rect 39470 865968 39760 865996
rect 39732 865844 39760 865968
rect 40468 865844 40496 913244
rect 42124 885036 42152 918192
rect 42294 914698 42350 914707
rect 42294 914633 42350 914642
rect 42308 910899 42336 914633
rect 42294 910890 42350 910899
rect 42294 910825 42350 910834
rect 41940 885008 42152 885036
rect 41940 872236 41968 885008
rect 42202 875802 42258 875811
rect 42202 875737 42258 875746
rect 41928 872230 41980 872236
rect 41928 872172 41980 872178
rect 42112 872230 42164 872236
rect 42112 872172 42164 872178
rect 42124 872116 42152 872172
rect 41940 872088 42152 872116
rect 39720 865838 39772 865844
rect 39720 865780 39772 865786
rect 40456 865838 40508 865844
rect 40456 865780 40508 865786
rect 41652 865838 41704 865844
rect 41652 865780 41704 865786
rect 39994 822762 40050 822771
rect 39994 822697 40050 822706
rect 40008 822612 40036 822697
rect 39470 822584 40036 822612
rect 40008 822363 40036 822584
rect 39994 822354 40050 822363
rect 39994 822289 40050 822298
rect 41664 793667 41692 865780
rect 41940 846532 41968 872088
rect 41744 846526 41796 846532
rect 41744 846468 41796 846474
rect 41928 846526 41980 846532
rect 41928 846468 41980 846474
rect 41756 837284 41784 846468
rect 41744 837278 41796 837284
rect 41744 837220 41796 837226
rect 42020 837278 42072 837284
rect 42020 837220 42072 837226
rect 42032 828104 42060 837220
rect 42020 828098 42072 828104
rect 42020 828040 42072 828046
rect 41928 827962 41980 827968
rect 41928 827904 41980 827910
rect 41940 793968 41968 827904
rect 41928 793962 41980 793968
rect 41928 793904 41980 793910
rect 41650 793658 41706 793667
rect 41650 793593 41706 793602
rect 41586 793480 42152 793508
rect 41586 791642 41692 791670
rect 41664 791180 41692 791642
rect 41652 791174 41704 791180
rect 41652 791116 41704 791122
rect 41926 789714 41982 789723
rect 41926 789649 41982 789658
rect 41940 789428 41968 789649
rect 42124 789587 42152 793480
rect 42110 789578 42166 789587
rect 42110 789513 42166 789522
rect 41940 789400 42152 789428
rect 41650 786042 41706 786051
rect 41650 785977 41706 785986
rect 41664 785484 41692 785977
rect 41586 785456 41692 785484
rect 42124 782220 42152 789400
rect 41664 782192 42152 782220
rect 41664 781932 41692 782192
rect 42112 782130 42164 782136
rect 42112 782072 42164 782078
rect 41652 781926 41704 781932
rect 41652 781868 41704 781874
rect 41652 781722 41704 781728
rect 41652 781664 41704 781670
rect 41664 781182 41692 781664
rect 41586 781154 41692 781182
rect 41664 780747 41692 781154
rect 41650 780738 41706 780747
rect 41650 780673 41706 780682
rect 41558 780552 41614 780561
rect 41558 780487 41614 780496
rect 41650 778018 41706 778027
rect 41650 777953 41706 777962
rect 41664 749036 41692 777953
rect 42124 749836 42152 782072
rect 42112 749830 42164 749836
rect 42112 749772 42164 749778
rect 41664 749008 42152 749036
rect 41586 748872 41692 748900
rect 41664 748408 41692 748872
rect 41652 748402 41704 748408
rect 41652 748344 41704 748350
rect 41836 747178 41888 747184
rect 41836 747120 41888 747126
rect 41848 747077 41876 747120
rect 41586 747049 41876 747077
rect 41848 746572 41876 747049
rect 41836 746566 41888 746572
rect 41836 746508 41888 746514
rect 42124 743619 42152 749008
rect 42110 743610 42166 743619
rect 42110 743545 42166 743554
rect 42112 743438 42164 743444
rect 42112 743380 42164 743386
rect 42124 741472 42152 743380
rect 41652 741466 41704 741472
rect 41652 741408 41704 741414
rect 42112 741466 42164 741472
rect 42112 741408 42164 741414
rect 41664 740906 41692 741408
rect 41586 740878 41692 740906
rect 41558 736596 41614 736605
rect 41558 736531 41614 736540
rect 41558 735952 41614 735961
rect 41558 735887 41614 735896
rect 42110 735952 42166 735961
rect 42110 735887 42166 735896
rect 41650 733410 41706 733419
rect 42124 733396 42152 735887
rect 41650 733345 41706 733354
rect 42032 733368 42152 733396
rect 41664 704723 41692 733345
rect 42032 721344 42060 733368
rect 42112 733306 42164 733312
rect 42112 733248 42164 733254
rect 41744 721338 41796 721344
rect 41744 721280 41796 721286
rect 42020 721338 42072 721344
rect 42020 721280 42072 721286
rect 41756 704859 41784 721280
rect 41742 704850 41798 704859
rect 41742 704785 41798 704794
rect 41650 704714 41706 704723
rect 41650 704649 41706 704658
rect 41558 704524 41614 704533
rect 41558 704459 41614 704468
rect 41586 702632 41692 702660
rect 41664 702236 41692 702632
rect 42124 702236 42152 733248
rect 41652 702230 41704 702236
rect 41652 702172 41704 702178
rect 42112 702230 42164 702236
rect 42112 702172 42164 702178
rect 41558 696520 41614 696529
rect 41558 696455 41614 696464
rect 42110 696418 42166 696427
rect 42110 696353 42166 696362
rect 41650 692746 41706 692755
rect 41650 692681 41706 692690
rect 41664 692188 41692 692681
rect 41586 692160 41692 692188
rect 41586 691510 41692 691538
rect 41664 691152 41692 691510
rect 42124 691152 42152 696353
rect 41652 691146 41704 691152
rect 41652 691088 41704 691094
rect 42112 691146 42164 691152
rect 42112 691088 42164 691094
rect 42124 689044 42152 691088
rect 41652 689038 41704 689044
rect 41652 688980 41704 688986
rect 42112 689038 42164 689044
rect 42112 688980 42164 688986
rect 41664 660076 41692 688980
rect 42110 688938 42166 688947
rect 42110 688873 42166 688882
rect 41926 682682 41982 682691
rect 41926 682617 41982 682626
rect 41940 673608 41968 682617
rect 41928 673602 41980 673608
rect 41928 673544 41980 673550
rect 41836 673398 41888 673404
rect 41836 673340 41888 673346
rect 41848 660115 41876 673340
rect 42124 660212 42152 688873
rect 42112 660206 42164 660212
rect 42112 660148 42164 660154
rect 41834 660106 41890 660115
rect 41652 660070 41704 660076
rect 41834 660041 41890 660050
rect 42112 660070 42164 660076
rect 41652 660012 41704 660018
rect 42112 660012 42164 660018
rect 41558 659924 41614 659933
rect 41558 659859 41614 659868
rect 41558 658066 41614 658075
rect 41558 658001 41614 658010
rect 42018 653306 42074 653315
rect 42018 653241 42020 653250
rect 42072 653241 42074 653250
rect 42020 653212 42072 653218
rect 41650 652354 41706 652363
rect 41650 652289 41706 652298
rect 41664 651932 41692 652289
rect 41586 651904 41692 651932
rect 41652 648102 41704 648108
rect 42124 648090 42152 660012
rect 41652 648044 41704 648050
rect 42032 648062 42152 648090
rect 41664 647580 41692 648044
rect 42032 647700 42060 648062
rect 42110 648002 42166 648011
rect 42110 647937 42166 647946
rect 42020 647694 42072 647700
rect 42020 647636 42072 647642
rect 41586 647552 41692 647580
rect 41652 647490 41704 647496
rect 41652 647432 41704 647438
rect 42020 647490 42072 647496
rect 42020 647432 42072 647438
rect 41664 646938 41692 647432
rect 41586 646910 41692 646938
rect 42032 646492 42060 647432
rect 42124 647059 42152 647937
rect 42110 647050 42166 647059
rect 42110 646985 42166 646994
rect 42032 646464 42152 646492
rect 42124 644504 42152 646464
rect 42112 644498 42164 644504
rect 42112 644440 42164 644446
rect 41652 644430 41704 644436
rect 41652 644372 41704 644378
rect 41560 627430 41612 627436
rect 41560 627372 41612 627378
rect 41572 615779 41600 627372
rect 41558 615770 41614 615779
rect 41558 615705 41614 615714
rect 41664 615507 41692 644372
rect 42112 644362 42164 644368
rect 42112 644304 42164 644310
rect 41742 644194 41798 644203
rect 41742 644129 41798 644138
rect 41756 627436 41784 644129
rect 41744 627430 41796 627436
rect 41744 627372 41796 627378
rect 41650 615498 41706 615507
rect 42124 615468 42152 644304
rect 41650 615433 41706 615442
rect 42112 615462 42164 615468
rect 42112 615404 42164 615410
rect 41558 615324 41614 615333
rect 41558 615259 41614 615268
rect 41650 613866 41706 613875
rect 41650 613801 41706 613810
rect 41664 613444 41692 613801
rect 41586 613416 41692 613444
rect 41664 612952 41692 613416
rect 41652 612946 41704 612952
rect 41652 612888 41704 612894
rect 42112 609002 42164 609008
rect 42112 608944 42164 608950
rect 41558 607338 41614 607347
rect 41558 607273 41614 607282
rect 41558 602986 41614 602995
rect 41558 602921 41614 602930
rect 41558 602352 41614 602361
rect 41558 602287 41614 602296
rect 41650 599858 41706 599867
rect 42124 599828 42152 608944
rect 41650 599793 41706 599802
rect 42112 599822 42164 599828
rect 41560 599550 41612 599556
rect 41560 599492 41612 599498
rect 41572 579700 41600 599492
rect 41560 579694 41612 579700
rect 41560 579636 41612 579642
rect 41664 576844 41692 599793
rect 42112 599764 42164 599770
rect 42110 599722 42166 599731
rect 42110 599657 42166 599666
rect 41836 579694 41888 579700
rect 41836 579636 41888 579642
rect 41652 576838 41704 576844
rect 41652 576780 41704 576786
rect 41848 571035 41876 579636
rect 42020 576838 42072 576844
rect 42020 576780 42072 576786
rect 41834 571026 41890 571035
rect 42032 571012 42060 576780
rect 42124 571132 42152 599657
rect 42112 571126 42164 571132
rect 42112 571068 42164 571074
rect 42032 570984 42152 571012
rect 41834 570961 41890 570970
rect 41586 570882 41692 570910
rect 41664 570491 41692 570882
rect 41650 570482 41706 570491
rect 41650 570417 41706 570426
rect 41558 569084 41614 569093
rect 41558 569019 41614 569028
rect 41650 563410 41706 563419
rect 41650 563345 41706 563354
rect 41664 562906 41692 563345
rect 41586 562878 41692 562906
rect 41652 559090 41704 559096
rect 41652 559032 41704 559038
rect 41664 558582 41692 559032
rect 41586 558554 41692 558582
rect 41664 558115 41692 558554
rect 41650 558106 41706 558115
rect 41650 558041 41706 558050
rect 42124 557979 42152 570984
rect 41558 557970 41614 557979
rect 41558 557905 41614 557914
rect 42110 557970 42166 557979
rect 42110 557905 42166 557914
rect 42110 557834 42166 557843
rect 42110 557769 42166 557778
rect 41834 555386 41890 555395
rect 41834 555321 41890 555330
rect 41744 551270 41796 551276
rect 41744 551212 41796 551218
rect 41756 526456 41784 551212
rect 41744 526450 41796 526456
rect 41744 526392 41796 526398
rect 41848 526404 41876 555321
rect 41926 555250 41982 555259
rect 41926 555185 41982 555194
rect 41940 551156 41968 555185
rect 42124 551276 42152 557769
rect 42112 551270 42164 551276
rect 42112 551212 42164 551218
rect 41940 551128 42152 551156
rect 42124 526563 42152 551128
rect 42110 526554 42166 526563
rect 42110 526489 42166 526498
rect 41848 526376 42152 526404
rect 41558 526324 41614 526333
rect 41558 526259 41614 526268
rect 41586 524442 41692 524470
rect 41664 523940 41692 524442
rect 41652 523934 41704 523940
rect 41652 523876 41704 523882
rect 42124 519083 42152 526376
rect 42110 519074 42166 519083
rect 42110 519009 42166 519018
rect 41558 518320 41614 518329
rect 41558 518255 41614 518264
rect 42112 518290 42164 518296
rect 42112 518232 42164 518238
rect 41558 513996 41614 514005
rect 41558 513931 41614 513940
rect 41558 513362 41614 513371
rect 41558 513297 41614 513306
rect 41650 510778 41706 510787
rect 41650 510713 41706 510722
rect 41926 510778 41982 510787
rect 41926 510713 41982 510722
rect 41664 499884 41692 510713
rect 41664 499856 41784 499884
rect 41652 499590 41704 499596
rect 41652 499532 41704 499538
rect 39260 439818 39312 439824
rect 39260 439760 39312 439766
rect 39272 434604 39300 439760
rect 39718 437882 39774 437891
rect 39718 437817 39774 437826
rect 39194 434576 39300 434604
rect 39431 430496 39668 430524
rect 39640 428604 39668 430496
rect 39628 428598 39680 428604
rect 39628 428540 39680 428546
rect 39180 423832 39392 423860
rect 39180 423710 39208 423832
rect 39364 423724 39392 423832
rect 39732 423747 39760 437817
rect 41560 425062 41612 425068
rect 41560 425004 41612 425010
rect 39534 423738 39590 423747
rect 39364 423696 39534 423724
rect 39534 423673 39590 423682
rect 39718 423738 39774 423747
rect 39718 423673 39774 423682
rect 41572 412216 41600 425004
rect 41560 412210 41612 412216
rect 41560 412152 41612 412158
rect 41664 394944 41692 499532
rect 41652 394938 41704 394944
rect 41652 394880 41704 394886
rect 41756 394876 41784 499856
rect 41940 493220 41968 510713
rect 42124 499596 42152 518232
rect 42112 499590 42164 499596
rect 42112 499532 42164 499538
rect 41848 493192 41968 493220
rect 41848 454460 41876 493192
rect 41848 454432 42060 454460
rect 42032 441660 42060 454432
rect 41836 441654 41888 441660
rect 41836 441596 41888 441602
rect 42020 441654 42072 441660
rect 42020 441596 42072 441602
rect 41848 428604 41876 441596
rect 41836 428598 41888 428604
rect 41836 428540 41888 428546
rect 42020 428598 42072 428604
rect 42020 428540 42072 428546
rect 42032 425068 42060 428540
rect 42020 425062 42072 425068
rect 42020 425004 42072 425010
rect 41836 412210 41888 412216
rect 41836 412152 41888 412158
rect 41848 399296 41876 412152
rect 41836 399290 41888 399296
rect 41836 399232 41888 399238
rect 41744 394870 41796 394876
rect 41744 394812 41796 394818
rect 41586 394682 41692 394710
rect 41664 394196 41692 394682
rect 41652 394190 41704 394196
rect 41652 394132 41704 394138
rect 42112 394190 42164 394196
rect 42112 394132 42164 394138
rect 41586 392824 41692 392852
rect 41664 392768 41692 392824
rect 41652 392762 41704 392768
rect 41652 392704 41704 392710
rect 42124 387260 42152 394132
rect 41652 387254 41704 387260
rect 41652 387196 41704 387202
rect 42112 387254 42164 387260
rect 42112 387196 42164 387202
rect 41664 386732 41692 387196
rect 41586 386704 41692 386732
rect 42112 386778 42164 386784
rect 42112 386720 42164 386726
rect 41586 382352 41692 382380
rect 41664 381888 41692 382352
rect 42124 381995 42152 386720
rect 42110 381986 42166 381995
rect 42110 381921 42166 381930
rect 41652 381882 41704 381888
rect 41652 381824 41704 381830
rect 42112 381882 42164 381888
rect 42112 381824 42164 381830
rect 41558 381752 41614 381761
rect 41558 381687 41614 381696
rect 41742 379266 41798 379275
rect 41652 379230 41704 379236
rect 42124 379236 42152 381824
rect 41742 379201 41798 379210
rect 42112 379230 42164 379236
rect 41652 379172 41704 379178
rect 41664 350336 41692 379172
rect 41652 350330 41704 350336
rect 41652 350272 41704 350278
rect 41756 350268 41784 379201
rect 42112 379172 42164 379178
rect 42020 374402 42072 374408
rect 42020 374344 42072 374350
rect 42032 364412 42060 374344
rect 42020 364406 42072 364412
rect 42020 364348 42072 364354
rect 42020 364270 42072 364276
rect 42020 364212 42072 364218
rect 42032 352240 42060 364212
rect 42020 352234 42072 352240
rect 42020 352176 42072 352182
rect 42112 350330 42164 350336
rect 42112 350272 42164 350278
rect 41744 350262 41796 350268
rect 41744 350204 41796 350210
rect 41586 350082 41692 350110
rect 41664 349588 41692 350082
rect 41652 349582 41704 349588
rect 41652 349524 41704 349530
rect 41836 348698 41888 348704
rect 41836 348640 41888 348646
rect 41848 348244 41876 348640
rect 41586 348216 41876 348244
rect 41848 347752 41876 348216
rect 41836 347746 41888 347752
rect 41836 347688 41888 347694
rect 42124 344624 42152 350272
rect 42112 344618 42164 344624
rect 42112 344560 42164 344566
rect 42112 344482 42164 344488
rect 42112 344424 42164 344430
rect 42124 342260 42152 344424
rect 41664 342232 42152 342260
rect 41664 342124 41692 342232
rect 41586 342096 41692 342124
rect 41652 338294 41704 338300
rect 41652 338236 41704 338242
rect 42112 338294 42164 338300
rect 42112 338236 42164 338242
rect 41664 337772 41692 338236
rect 41586 337744 41692 337772
rect 41652 337682 41704 337688
rect 41652 337624 41704 337630
rect 41664 337138 41692 337624
rect 41586 337110 41692 337138
rect 41836 335166 41888 335172
rect 41836 335108 41888 335114
rect 41848 334900 41876 335108
rect 41836 334894 41888 334900
rect 41836 334836 41888 334842
rect 42124 334644 42152 338236
rect 41652 334622 41704 334628
rect 41652 334564 41704 334570
rect 42032 334616 42152 334644
rect 41664 334100 41692 334564
rect 41572 334072 41692 334100
rect 41572 312868 41600 334072
rect 42032 334016 42060 334616
rect 42112 334418 42164 334424
rect 42112 334360 42164 334366
rect 41652 334010 41704 334016
rect 41652 333952 41704 333958
rect 42020 334010 42072 334016
rect 42020 333952 42072 333958
rect 41560 312862 41612 312868
rect 41560 312804 41612 312810
rect 41664 305835 41692 333952
rect 42124 325668 42152 334360
rect 42032 325640 42152 325668
rect 42032 321996 42060 325640
rect 41940 321968 42060 321996
rect 41940 312868 41968 321968
rect 41744 312862 41796 312868
rect 41744 312804 41796 312810
rect 41928 312862 41980 312868
rect 41928 312804 41980 312810
rect 41650 305826 41706 305835
rect 41756 305812 41784 312804
rect 42020 312794 42072 312800
rect 42020 312736 42072 312742
rect 42032 309196 42060 312736
rect 41928 309190 41980 309196
rect 41928 309132 41980 309138
rect 42020 309190 42072 309196
rect 42020 309132 42072 309138
rect 41940 305932 41968 309132
rect 41928 305926 41980 305932
rect 41928 305868 41980 305874
rect 41756 305784 42152 305812
rect 41650 305761 41706 305770
rect 41586 305682 41876 305710
rect 41848 305184 41876 305682
rect 42124 305388 42152 305784
rect 42112 305382 42164 305388
rect 42112 305324 42164 305330
rect 41836 305178 41888 305184
rect 41836 305120 41888 305126
rect 42112 305178 42164 305184
rect 42112 305120 42164 305126
rect 41586 303842 41692 303870
rect 41664 303348 41692 303842
rect 41652 303342 41704 303348
rect 41652 303284 41704 303290
rect 42124 297788 42152 305120
rect 41664 297760 42152 297788
rect 41664 297706 41692 297760
rect 41586 297678 41692 297706
rect 42110 297666 42166 297675
rect 42110 297601 42166 297610
rect 42124 293624 42152 297601
rect 41652 293618 41704 293624
rect 41652 293560 41704 293566
rect 42112 293618 42164 293624
rect 42112 293560 42164 293566
rect 41558 293396 41614 293405
rect 41664 293382 41692 293560
rect 42112 293482 42164 293488
rect 42112 293424 42164 293430
rect 41614 293354 41692 293382
rect 41558 293331 41614 293340
rect 41558 292770 41614 292779
rect 41558 292705 41614 292714
rect 41742 290186 41798 290195
rect 41742 290121 41798 290130
rect 41650 287194 41706 287203
rect 41650 287129 41706 287138
rect 41664 266628 41692 287129
rect 41652 266622 41704 266628
rect 41652 266564 41704 266570
rect 41756 261324 41784 290121
rect 42124 287436 42152 293424
rect 42216 292484 42244 875737
rect 42308 431363 42336 910825
rect 43044 879483 43072 960096
rect 81684 953088 81712 992328
rect 81672 953082 81724 953088
rect 81672 953024 81724 953030
rect 81776 953020 81804 993416
rect 82420 992392 82448 993552
rect 86744 993548 86772 995454
rect 86732 993542 86784 993548
rect 86732 993484 86784 993490
rect 92908 993344 92936 995454
rect 94748 993548 94776 995454
rect 136332 995440 136386 995468
rect 136976 995440 137030 995468
rect 141300 995440 141354 995468
rect 147464 995440 147518 995468
rect 149304 995440 149358 995468
rect 102922 993578 102978 993587
rect 94736 993542 94788 993548
rect 94736 993484 94788 993490
rect 100072 993542 100124 993548
rect 102922 993513 102924 993522
rect 100072 993484 100124 993490
rect 102976 993513 102978 993522
rect 115710 993578 115766 993587
rect 136332 993548 136360 995440
rect 136976 993616 137004 995440
rect 136964 993610 137016 993616
rect 136964 993552 137016 993558
rect 115710 993513 115766 993522
rect 136320 993542 136372 993548
rect 102924 993484 102976 993490
rect 93724 993474 93776 993480
rect 93724 993416 93776 993422
rect 92712 993338 92764 993344
rect 92712 993280 92764 993286
rect 92896 993338 92948 993344
rect 92896 993280 92948 993286
rect 82408 992386 82460 992392
rect 82408 992328 82460 992334
rect 92724 970632 92752 993280
rect 93736 993276 93764 993416
rect 100084 993276 100112 993484
rect 115724 993480 115752 993513
rect 136320 993484 136372 993490
rect 115712 993474 115764 993480
rect 115712 993416 115764 993422
rect 136332 993412 136360 993484
rect 141300 993480 141328 995440
rect 141288 993474 141340 993480
rect 141288 993416 141340 993422
rect 136320 993406 136372 993412
rect 136320 993348 136372 993354
rect 147464 993344 147492 995440
rect 149304 993480 149332 995440
rect 178376 993536 178588 993564
rect 178376 993480 178404 993536
rect 149292 993474 149344 993480
rect 149292 993416 149344 993422
rect 157940 993474 157992 993480
rect 158124 993474 158176 993480
rect 157992 993422 158124 993428
rect 157940 993416 158176 993422
rect 170912 993474 170964 993480
rect 171004 993474 171056 993480
rect 170964 993422 171004 993428
rect 170912 993416 171056 993422
rect 178364 993474 178416 993480
rect 178364 993416 178416 993422
rect 157952 993400 158164 993416
rect 170924 993400 171044 993416
rect 147452 993338 147504 993344
rect 147452 993280 147504 993286
rect 93724 993270 93776 993276
rect 93724 993212 93776 993218
rect 100072 993270 100124 993276
rect 100072 993212 100124 993218
rect 178560 993140 178588 993536
rect 190980 993140 191008 995454
rect 191624 993616 191652 995454
rect 195948 993616 195976 995454
rect 191612 993610 191664 993616
rect 191612 993552 191664 993558
rect 195936 993610 195988 993616
rect 195936 993552 195988 993558
rect 191624 993208 191652 993552
rect 202112 993548 202140 995454
rect 203952 993616 203980 995454
rect 245536 995440 245586 995468
rect 246180 995440 246230 995468
rect 250504 995440 250554 995468
rect 203940 993610 203992 993616
rect 203940 993552 203992 993558
rect 202100 993542 202152 993548
rect 202100 993484 202152 993490
rect 222616 993542 222668 993548
rect 222616 993484 222668 993490
rect 202112 993344 202140 993484
rect 209828 993474 209880 993480
rect 222628 993428 222656 993484
rect 209828 993416 209880 993422
rect 202100 993338 202152 993344
rect 209736 993338 209788 993344
rect 202100 993280 202152 993286
rect 209564 993286 209736 993292
rect 209564 993280 209788 993286
rect 209564 993264 209776 993280
rect 209564 993208 209592 993264
rect 191612 993202 191664 993208
rect 191612 993144 191664 993150
rect 209552 993202 209604 993208
rect 209552 993144 209604 993150
rect 209840 993140 209868 993416
rect 222444 993412 222656 993428
rect 245536 993412 245564 995440
rect 222432 993406 222656 993412
rect 222484 993400 222656 993406
rect 245524 993406 245576 993412
rect 222432 993348 222484 993354
rect 245524 993348 245576 993354
rect 178548 993134 178600 993140
rect 178548 993076 178600 993082
rect 190968 993134 191020 993140
rect 190968 993076 191020 993082
rect 209828 993134 209880 993140
rect 209828 993076 209880 993082
rect 244604 992862 244656 992868
rect 244604 992804 244656 992810
rect 244616 992732 244644 992804
rect 246180 992732 246208 995440
rect 250400 994222 250452 994228
rect 250400 994164 250452 994170
rect 250412 993616 250440 994164
rect 250504 993616 250532 995440
rect 256668 994228 256696 995636
rect 256656 994222 256708 994228
rect 256656 994164 256708 994170
rect 258508 993616 258536 995636
rect 311396 995514 311448 995520
rect 311330 995462 311396 995468
rect 311330 995456 311448 995462
rect 312776 995514 312828 995520
rect 312776 995456 312828 995462
rect 259048 994222 259100 994228
rect 259048 994164 259100 994170
rect 259060 993616 259088 994164
rect 250400 993610 250452 993616
rect 250400 993552 250452 993558
rect 250492 993610 250544 993616
rect 250492 993552 250544 993558
rect 258496 993610 258548 993616
rect 258496 993552 258548 993558
rect 259048 993610 259100 993616
rect 259048 993552 259100 993558
rect 261162 993578 261218 993587
rect 248376 993542 248428 993548
rect 261162 993513 261164 993522
rect 248376 993484 248428 993490
rect 261216 993513 261218 993522
rect 261164 993484 261216 993490
rect 248284 993406 248336 993412
rect 248388 993394 248416 993484
rect 273952 993474 274004 993480
rect 248336 993366 248416 993394
rect 273950 993442 273952 993451
rect 274044 993474 274096 993480
rect 274004 993442 274006 993451
rect 287016 993474 287068 993480
rect 274044 993416 274096 993422
rect 286844 993422 287016 993428
rect 286844 993416 287068 993422
rect 299804 993474 299856 993480
rect 299804 993416 299856 993422
rect 273950 993377 274006 993386
rect 248284 993348 248336 993354
rect 274056 993344 274084 993416
rect 286844 993400 287056 993416
rect 286844 993344 286872 993400
rect 274044 993338 274096 993344
rect 274044 993280 274096 993286
rect 286832 993338 286884 993344
rect 286832 993280 286884 993286
rect 295848 993202 295900 993208
rect 295848 993144 295900 993150
rect 257392 992998 257444 993004
rect 257392 992940 257444 992946
rect 257404 992732 257432 992940
rect 295860 992884 295888 993144
rect 296032 992998 296084 993004
rect 296032 992940 296084 992946
rect 299712 992998 299764 993004
rect 299816 992986 299844 993416
rect 300184 993208 300212 995454
rect 300828 993480 300856 995454
rect 300816 993474 300868 993480
rect 300816 993416 300868 993422
rect 305152 993412 305180 995454
rect 311330 995440 311436 995456
rect 312788 993616 312816 995456
rect 312776 993610 312828 993616
rect 312776 993552 312828 993558
rect 312592 993542 312644 993548
rect 312592 993484 312644 993490
rect 305140 993406 305192 993412
rect 305140 993348 305192 993354
rect 300172 993202 300224 993208
rect 300172 993144 300224 993150
rect 312604 993140 312632 993484
rect 312788 993208 312816 993552
rect 313156 993412 313184 995454
rect 353176 993480 353204 997457
rect 353164 993474 353216 993480
rect 353164 993416 353216 993422
rect 313144 993406 313196 993412
rect 313144 993348 313196 993354
rect 338364 993276 338484 993292
rect 364124 993276 364244 993292
rect 334672 993270 334724 993276
rect 334672 993212 334724 993218
rect 338352 993270 338496 993276
rect 338404 993264 338444 993270
rect 338352 993212 338404 993218
rect 338444 993212 338496 993218
rect 360432 993270 360484 993276
rect 360432 993212 360484 993218
rect 364112 993270 364256 993276
rect 364164 993264 364204 993270
rect 364112 993212 364164 993218
rect 364204 993212 364256 993218
rect 312776 993202 312828 993208
rect 321884 993202 321936 993208
rect 312776 993144 312828 993150
rect 321882 993170 321884 993179
rect 334684 993179 334712 993212
rect 347644 993202 347696 993208
rect 321936 993170 321938 993179
rect 312592 993134 312644 993140
rect 321882 993105 321938 993114
rect 334670 993170 334726 993179
rect 334670 993105 334726 993114
rect 347642 993170 347644 993179
rect 360444 993179 360472 993212
rect 347696 993170 347698 993179
rect 347642 993105 347698 993114
rect 360430 993170 360486 993179
rect 360430 993105 360486 993114
rect 312592 993076 312644 993082
rect 299764 992958 299844 992986
rect 299712 992940 299764 992946
rect 296044 992884 296072 992940
rect 295860 992856 296072 992884
rect 244604 992726 244656 992732
rect 244604 992668 244656 992674
rect 246168 992726 246220 992732
rect 246168 992668 246220 992674
rect 257392 992726 257444 992732
rect 257392 992668 257444 992674
rect 364400 975256 364428 997457
rect 573962 997386 574018 997395
rect 573962 997321 574018 997330
rect 408100 995576 408220 995604
rect 406614 995482 406670 995491
rect 406614 995417 406670 995426
rect 406628 993480 406656 995417
rect 408100 993548 408128 995576
rect 408192 995454 408220 995576
rect 466968 995514 467020 995520
rect 408822 995482 408878 995491
rect 408822 995417 408878 995426
rect 413146 995482 413202 995491
rect 421150 995482 421206 995491
rect 413146 995417 413202 995426
rect 419140 995440 419338 995468
rect 408088 993542 408140 993548
rect 408088 993484 408140 993490
rect 406616 993474 406668 993480
rect 406616 993416 406668 993422
rect 419140 993412 419168 995440
rect 466968 995456 467020 995462
rect 473776 995514 473828 995520
rect 473828 995462 473894 995468
rect 473776 995456 473894 995462
rect 421150 995417 421206 995426
rect 437804 993610 437856 993616
rect 437804 993552 437856 993558
rect 450592 993610 450644 993616
rect 450592 993552 450644 993558
rect 419128 993406 419180 993412
rect 419128 993348 419180 993354
rect 389884 993276 390004 993292
rect 419140 993276 419168 993348
rect 437816 993344 437844 993552
rect 450604 993344 450632 993552
rect 462748 993548 462776 995454
rect 462736 993542 462788 993548
rect 462736 993484 462788 993490
rect 463392 993480 463420 995454
rect 463380 993474 463432 993480
rect 463380 993416 463432 993422
rect 466980 993344 467008 995456
rect 473788 995454 473894 995456
rect 467716 995316 467744 995454
rect 473788 995440 473908 995454
rect 467704 995310 467756 995316
rect 467704 995252 467756 995258
rect 437804 993338 437856 993344
rect 437804 993280 437856 993286
rect 450592 993338 450644 993344
rect 450592 993280 450644 993286
rect 466968 993338 467020 993344
rect 466968 993280 467020 993286
rect 473880 993276 473908 995440
rect 475628 995440 475734 995468
rect 475628 995316 475656 995440
rect 475616 995310 475668 995316
rect 475616 995252 475668 995258
rect 517292 993610 517344 993616
rect 517292 993552 517344 993558
rect 517304 993480 517332 993552
rect 517396 993480 517424 995454
rect 518040 993616 518068 995454
rect 518028 993610 518080 993616
rect 518028 993552 518080 993558
rect 517292 993474 517344 993480
rect 517292 993416 517344 993422
rect 517384 993474 517436 993480
rect 517384 993416 517436 993422
rect 522364 993344 522392 995454
rect 528528 993548 528556 995454
rect 528516 993542 528568 993548
rect 528516 993484 528568 993490
rect 528528 993412 528556 993484
rect 528516 993406 528568 993412
rect 528516 993348 528568 993354
rect 530368 993344 530396 995454
rect 522352 993338 522404 993344
rect 522352 993280 522404 993286
rect 530356 993338 530408 993344
rect 530356 993280 530408 993286
rect 386192 993270 386244 993276
rect 386192 993212 386244 993218
rect 389872 993270 390016 993276
rect 389924 993264 389964 993270
rect 389872 993212 389924 993218
rect 389964 993212 390016 993218
rect 419128 993270 419180 993276
rect 419128 993212 419180 993218
rect 473868 993270 473920 993276
rect 473868 993212 473920 993218
rect 373404 993202 373456 993208
rect 373402 993170 373404 993179
rect 386204 993179 386232 993212
rect 373456 993170 373458 993179
rect 373402 993105 373458 993114
rect 386190 993170 386246 993179
rect 386190 993105 386246 993114
rect 364204 975250 364256 975256
rect 364388 975250 364440 975256
rect 364256 975198 364336 975204
rect 364204 975192 364336 975198
rect 364388 975192 364440 975198
rect 364216 975176 364336 975192
rect 92712 970626 92764 970632
rect 92712 970568 92764 970574
rect 364308 962420 364336 975176
rect 364308 962392 364428 962420
rect 364400 960160 364428 962392
rect 364388 960154 364440 960160
rect 364388 960096 364440 960102
rect 99612 960086 99664 960092
rect 99612 960028 99664 960034
rect 99624 953836 99652 960028
rect 93908 953830 93960 953836
rect 93908 953772 93960 953778
rect 99612 953830 99664 953836
rect 99612 953772 99664 953778
rect 81764 953014 81816 953020
rect 81764 952956 81816 952962
rect 93920 951388 93948 953772
rect 92436 951382 92488 951388
rect 92436 951324 92488 951330
rect 93908 951382 93960 951388
rect 93908 951324 93960 951330
rect 92448 941188 92476 951324
rect 90044 941182 90096 941188
rect 90044 941124 90096 941130
rect 92436 941182 92488 941188
rect 92436 941124 92488 941130
rect 90056 937516 90084 941124
rect 88204 937510 88256 937516
rect 88204 937452 88256 937458
rect 90044 937510 90096 937516
rect 90044 937452 90096 937458
rect 88216 934796 88244 937452
rect 87008 934790 87060 934796
rect 87008 934732 87060 934738
rect 88204 934790 88256 934796
rect 88204 934732 88256 934738
rect 87020 931940 87048 934732
rect 80844 931934 80896 931940
rect 80844 931876 80896 931882
rect 87008 931934 87060 931940
rect 87008 931876 87060 931882
rect 80856 926500 80884 931876
rect 44044 926494 44096 926500
rect 44044 926436 44096 926442
rect 80844 926494 80896 926500
rect 80844 926436 80896 926442
rect 44056 925616 44084 926436
rect 44044 925610 44096 925616
rect 44044 925552 44096 925558
rect 43030 879474 43086 879483
rect 43030 879409 43086 879418
rect 42478 830106 42534 830115
rect 42478 830041 42534 830050
rect 42386 822354 42442 822363
rect 42386 822289 42442 822298
rect 42400 472979 42428 822289
rect 42492 476515 42520 830041
rect 42572 793962 42624 793968
rect 42572 793904 42624 793910
rect 42584 791180 42612 793904
rect 42572 791174 42624 791180
rect 42572 791116 42624 791122
rect 42584 782136 42612 791116
rect 42572 782130 42624 782136
rect 42572 782072 42624 782078
rect 42572 749830 42624 749836
rect 42572 749772 42624 749778
rect 42584 747184 42612 749772
rect 42664 748402 42716 748408
rect 42664 748344 42716 748350
rect 42572 747178 42624 747184
rect 42572 747120 42624 747126
rect 42572 746566 42624 746572
rect 42572 746508 42624 746514
rect 42584 733312 42612 746508
rect 42676 743444 42704 748344
rect 42664 743438 42716 743444
rect 42664 743380 42716 743386
rect 42572 733306 42624 733312
rect 42572 733248 42624 733254
rect 42572 702230 42624 702236
rect 42572 702172 42624 702178
rect 42584 682691 42612 702172
rect 42570 682682 42626 682691
rect 42570 682617 42626 682626
rect 42572 660206 42624 660212
rect 42572 660148 42624 660154
rect 42584 648108 42612 660148
rect 42662 658066 42718 658075
rect 42662 658001 42718 658010
rect 42676 653276 42704 658001
rect 42664 653270 42716 653276
rect 42664 653212 42716 653218
rect 42572 648102 42624 648108
rect 42572 648044 42624 648050
rect 42584 644368 42612 648044
rect 42572 644362 42624 644368
rect 42572 644304 42624 644310
rect 42572 615462 42624 615468
rect 42572 615404 42624 615410
rect 42584 614532 42612 615404
rect 42584 614504 42796 614532
rect 42572 612946 42624 612952
rect 42572 612888 42624 612894
rect 42584 609008 42612 612888
rect 42572 609002 42624 609008
rect 42572 608944 42624 608950
rect 42768 602995 42796 614504
rect 42754 602986 42810 602995
rect 42754 602921 42810 602930
rect 42572 571126 42624 571132
rect 42572 571068 42624 571074
rect 42584 559096 42612 571068
rect 42572 559090 42624 559096
rect 42572 559032 42624 559038
rect 42572 526450 42624 526456
rect 42572 526392 42624 526398
rect 42584 523940 42612 526392
rect 42572 523934 42624 523940
rect 42572 523876 42624 523882
rect 42584 518296 42612 523876
rect 42572 518290 42624 518296
rect 42572 518232 42624 518238
rect 42478 476506 42534 476515
rect 42478 476441 42534 476450
rect 42492 474883 42520 476441
rect 42478 474874 42534 474883
rect 42478 474809 42534 474818
rect 42386 472970 42442 472979
rect 42386 472905 42442 472914
rect 44056 439824 44084 925552
rect 573976 821576 574004 997321
rect 581520 975256 581548 997457
rect 625588 993480 625616 995454
rect 626232 993616 626260 995454
rect 630556 993616 630584 995454
rect 625760 993610 625812 993616
rect 625760 993552 625812 993558
rect 626220 993610 626272 993616
rect 626220 993552 626272 993558
rect 630544 993610 630596 993616
rect 630544 993552 630596 993558
rect 625576 993474 625628 993480
rect 625576 993416 625628 993422
rect 625588 992732 625616 993416
rect 625772 992800 625800 993552
rect 636720 993548 636748 995454
rect 638560 993616 638588 995454
rect 638548 993610 638600 993616
rect 638548 993552 638600 993558
rect 636708 993542 636760 993548
rect 636708 993484 636760 993490
rect 636720 992868 636748 993484
rect 636708 992862 636760 992868
rect 636708 992804 636760 992810
rect 675164 992862 675216 992868
rect 675164 992804 675216 992810
rect 625760 992794 625812 992800
rect 625760 992736 625812 992742
rect 625576 992726 625628 992732
rect 625576 992668 625628 992674
rect 581324 975250 581376 975256
rect 581508 975250 581560 975256
rect 581376 975198 581456 975204
rect 581324 975192 581456 975198
rect 581508 975192 581560 975198
rect 581336 975176 581456 975192
rect 581428 962420 581456 975176
rect 674980 966070 675032 966076
rect 674980 966012 675032 966018
rect 674992 963372 675020 966012
rect 675072 966002 675124 966008
rect 675072 965944 675124 965950
rect 675084 963916 675112 965944
rect 675176 964036 675204 992804
rect 675348 992794 675400 992800
rect 675348 992736 675400 992742
rect 675256 992726 675308 992732
rect 675256 992668 675308 992674
rect 675268 966008 675296 992668
rect 675360 966076 675388 992736
rect 675348 966070 675400 966076
rect 675348 966012 675400 966018
rect 675256 966002 675308 966008
rect 675256 965944 675308 965950
rect 675164 964030 675216 964036
rect 675164 963972 675216 963978
rect 675084 963888 675296 963916
rect 675164 963826 675216 963832
rect 675164 963768 675216 963774
rect 674992 963344 675112 963372
rect 674980 963010 675032 963016
rect 674980 962952 675032 962958
rect 581428 962392 581548 962420
rect 581520 949484 581548 962392
rect 632936 960086 632988 960092
rect 632936 960028 632988 960034
rect 632948 954992 632976 960028
rect 674796 958658 674848 958664
rect 674796 958600 674848 958606
rect 632936 954986 632988 954992
rect 632936 954928 632988 954934
rect 641032 954986 641084 954992
rect 641032 954928 641084 954934
rect 581324 949478 581376 949484
rect 581324 949420 581376 949426
rect 581508 949478 581560 949484
rect 581508 949420 581560 949426
rect 581336 949364 581364 949420
rect 581336 949336 581456 949364
rect 581428 936580 581456 949336
rect 641044 947648 641072 954928
rect 674808 951932 674836 958600
rect 674796 951926 674848 951932
rect 674796 951868 674848 951874
rect 674808 948600 674836 951868
rect 674992 950316 675020 962952
rect 675084 962851 675112 963344
rect 675070 962842 675126 962851
rect 675070 962777 675126 962786
rect 675084 950860 675112 962777
rect 675176 962404 675204 963768
rect 675268 963016 675296 963888
rect 675256 963010 675308 963016
rect 675256 962952 675308 962958
rect 675254 962842 675310 962851
rect 675254 962777 675310 962786
rect 675164 962398 675216 962404
rect 675164 962340 675216 962346
rect 675164 962194 675216 962200
rect 675164 962136 675216 962142
rect 675176 958664 675204 962136
rect 675164 958658 675216 958664
rect 675164 958600 675216 958606
rect 675176 958498 675282 958526
rect 675176 950996 675204 958498
rect 675268 951932 675296 952342
rect 675256 951926 675308 951932
rect 675256 951868 675308 951874
rect 675176 950968 675296 950996
rect 675084 950832 675204 950860
rect 675176 950452 675204 950832
rect 675268 950508 675296 950968
rect 675176 950424 675388 950452
rect 674992 950288 675296 950316
rect 674796 948594 674848 948600
rect 674796 948536 674848 948542
rect 675164 948594 675216 948600
rect 675164 948536 675216 948542
rect 641032 947642 641084 947648
rect 641032 947584 641084 947590
rect 646644 947574 646696 947580
rect 646644 947516 646696 947522
rect 646656 943432 646684 947516
rect 646644 943426 646696 943432
rect 646644 943368 646696 943374
rect 653912 943426 653964 943432
rect 653912 943368 653964 943374
rect 581428 936552 581548 936580
rect 581520 923780 581548 936552
rect 653924 934796 653952 943368
rect 653912 934790 653964 934796
rect 653912 934732 653964 934738
rect 655752 934790 655804 934796
rect 655752 934732 655804 934738
rect 581324 923774 581376 923780
rect 581324 923716 581376 923722
rect 581508 923774 581560 923780
rect 581508 923716 581560 923722
rect 581336 923660 581364 923716
rect 581336 923632 581456 923660
rect 581428 910876 581456 923632
rect 655764 920040 655792 934732
rect 655752 920034 655804 920040
rect 655752 919976 655804 919982
rect 661272 919966 661324 919972
rect 661272 919908 661324 919914
rect 581428 910848 581548 910876
rect 581520 897956 581548 910848
rect 661284 908956 661312 919908
rect 675070 911026 675126 911035
rect 675070 910961 675126 910970
rect 661272 908950 661324 908956
rect 661272 908892 661324 908898
rect 669460 908950 669512 908956
rect 669460 908892 669512 908898
rect 669472 905352 669500 908892
rect 669460 905346 669512 905352
rect 675084 905323 675112 910961
rect 669460 905288 669512 905294
rect 675070 905314 675126 905323
rect 675070 905249 675126 905258
rect 581336 897928 581548 897956
rect 581336 885036 581364 897928
rect 581336 885008 581548 885036
rect 581520 872236 581548 885008
rect 675084 875364 675112 905249
rect 674520 875358 674572 875364
rect 674520 875300 674572 875306
rect 675072 875358 675124 875364
rect 675072 875300 675124 875306
rect 581324 872230 581376 872236
rect 581324 872172 581376 872178
rect 581508 872230 581560 872236
rect 581508 872172 581560 872178
rect 581336 872116 581364 872172
rect 581336 872088 581548 872116
rect 581520 846464 581548 872088
rect 674532 863056 674560 875300
rect 675176 875244 675204 948536
rect 675084 875216 675204 875244
rect 674980 873794 675032 873800
rect 674980 873736 675032 873742
rect 674992 871760 675020 873736
rect 674980 871754 675032 871760
rect 674980 871696 675032 871702
rect 674888 866790 674940 866796
rect 674888 866732 674940 866738
rect 674520 863050 674572 863056
rect 674520 862992 674572 862998
rect 674612 863050 674664 863056
rect 674612 862992 674664 862998
rect 674624 853740 674652 862992
rect 674900 860676 674928 866732
rect 674992 866676 675020 871696
rect 675084 870484 675112 875216
rect 675164 875086 675216 875092
rect 675164 875028 675216 875034
rect 675176 870650 675204 875028
rect 675268 873800 675296 950288
rect 675360 908956 675388 950424
rect 677738 915650 677794 915659
rect 677794 915608 677950 915636
rect 677738 915585 677794 915594
rect 677568 910848 677896 910876
rect 677568 908956 677596 910848
rect 675348 908950 675400 908956
rect 675348 908892 675400 908898
rect 677556 908950 677608 908956
rect 677556 908892 677608 908898
rect 675360 875092 675388 908892
rect 677556 905278 677608 905284
rect 677556 905220 677608 905226
rect 677568 904756 677596 905220
rect 677568 904728 677950 904756
rect 675348 875086 675400 875092
rect 675348 875028 675400 875034
rect 675256 873794 675308 873800
rect 675256 873736 675308 873742
rect 675256 871754 675308 871760
rect 675256 871696 675308 871702
rect 675268 871286 675296 871696
rect 675176 870622 675282 870650
rect 675084 870456 675204 870484
rect 675176 870196 675204 870456
rect 675164 870190 675216 870196
rect 675164 870132 675216 870138
rect 675164 869986 675216 869992
rect 675164 869928 675216 869934
rect 675176 866796 675204 869928
rect 675164 866790 675216 866796
rect 675164 866732 675216 866738
rect 674992 866648 675204 866676
rect 675176 866404 675204 866648
rect 675084 866376 675204 866404
rect 674888 860670 674940 860676
rect 674888 860612 674940 860618
rect 674900 858108 674928 860612
rect 675084 858244 675112 866376
rect 675176 866298 675282 866326
rect 675176 858322 675204 866298
rect 675256 860670 675308 860676
rect 675256 860612 675308 860618
rect 675268 860134 675296 860612
rect 675176 858294 675282 858322
rect 675084 858216 675388 858244
rect 674900 858080 675204 858108
rect 674612 853734 674664 853740
rect 674612 853676 674664 853682
rect 674980 853734 675032 853740
rect 674980 853676 675032 853682
rect 674992 850084 675020 853676
rect 674900 850056 675020 850084
rect 581324 846458 581376 846464
rect 581324 846400 581376 846406
rect 581508 846458 581560 846464
rect 581508 846400 581560 846406
rect 581336 833492 581364 846400
rect 674900 840956 674928 850056
rect 674888 840950 674940 840956
rect 674888 840892 674940 840898
rect 674980 840882 675032 840888
rect 674980 840824 675032 840830
rect 674992 837284 675020 840824
rect 674888 837278 674940 837284
rect 674888 837220 674940 837226
rect 674980 837278 675032 837284
rect 674980 837220 675032 837226
rect 581336 833464 581548 833492
rect 573964 821570 574016 821576
rect 573964 821512 574016 821518
rect 581520 820692 581548 833464
rect 674900 828052 674928 837220
rect 675176 836196 675204 858080
rect 675360 850068 675388 858216
rect 675256 850062 675308 850068
rect 675256 850004 675308 850010
rect 675348 850062 675400 850068
rect 675348 850004 675400 850010
rect 675268 837284 675296 850004
rect 675256 837278 675308 837284
rect 675256 837220 675308 837226
rect 675532 837278 675584 837284
rect 675532 837220 675584 837226
rect 675164 836190 675216 836196
rect 675164 836132 675216 836138
rect 675440 836190 675492 836196
rect 675440 836132 675492 836138
rect 674900 828024 675112 828052
rect 674978 822490 675034 822499
rect 674978 822425 675034 822434
rect 674992 821576 675020 822425
rect 674980 821570 675032 821576
rect 674980 821512 675032 821518
rect 581324 820686 581376 820692
rect 581324 820628 581376 820634
rect 581508 820686 581560 820692
rect 581508 820628 581560 820634
rect 581336 817904 581364 820628
rect 581324 817898 581376 817904
rect 581324 817840 581376 817846
rect 674888 817898 674940 817904
rect 674888 817840 674940 817846
rect 674900 817739 674928 817840
rect 674886 817730 674942 817739
rect 674886 817665 674942 817674
rect 674900 813387 674928 817665
rect 674886 813378 674942 813387
rect 674886 813313 674942 813322
rect 674900 809608 674928 813313
rect 674704 809602 674756 809608
rect 674704 809544 674756 809550
rect 674888 809602 674940 809608
rect 674888 809544 674940 809550
rect 674716 796756 674744 809544
rect 674704 796750 674756 796756
rect 674704 796692 674756 796698
rect 674888 796750 674940 796756
rect 674888 796692 674940 796698
rect 674796 790494 674848 790500
rect 674796 790436 674848 790442
rect 674426 783866 674482 783875
rect 674426 783801 674482 783810
rect 674440 760036 674468 783801
rect 674808 782952 674836 790436
rect 674900 783875 674928 796692
rect 674886 783866 674942 783875
rect 674886 783801 674942 783810
rect 674796 782946 674848 782952
rect 674796 782888 674848 782894
rect 674520 781586 674572 781592
rect 674520 781528 674572 781534
rect 674532 779008 674560 781528
rect 674520 779002 674572 779008
rect 674520 778944 674572 778950
rect 674532 765952 674560 778944
rect 674704 778594 674756 778600
rect 674704 778536 674756 778542
rect 674612 770094 674664 770100
rect 674612 770036 674664 770042
rect 674520 765946 674572 765952
rect 674520 765888 674572 765894
rect 674428 760030 674480 760036
rect 674428 759972 674480 759978
rect 674624 757180 674652 770036
rect 674716 768536 674744 778536
rect 674796 774242 674848 774248
rect 674796 774184 674848 774190
rect 674704 768530 674756 768536
rect 674704 768472 674756 768478
rect 674808 766020 674836 774184
rect 674796 766014 674848 766020
rect 674796 765956 674848 765962
rect 674888 760030 674940 760036
rect 674888 759972 674940 759978
rect 674900 758064 674928 759972
rect 674704 758058 674756 758064
rect 674704 758000 674756 758006
rect 674888 758058 674940 758064
rect 674888 758000 674940 758006
rect 674612 757174 674664 757180
rect 674612 757116 674664 757122
rect 674716 745251 674744 758000
rect 674702 745242 674758 745251
rect 674702 745177 674758 745186
rect 674886 745242 674942 745251
rect 674886 745177 674942 745186
rect 674796 744322 674848 744328
rect 674796 744264 674848 744270
rect 674612 735346 674664 735352
rect 674612 735288 674664 735294
rect 674426 732322 674482 732331
rect 674426 732257 674482 732266
rect 674440 721956 674468 732257
rect 674624 725016 674652 735288
rect 674704 735278 674756 735284
rect 674704 735220 674756 735226
rect 674612 725010 674664 725016
rect 674612 724952 674664 724958
rect 674716 722092 674744 735220
rect 674704 722086 674756 722092
rect 674704 722028 674756 722034
rect 674428 721950 674480 721956
rect 674428 721892 674480 721898
rect 674704 721950 674756 721956
rect 674704 721892 674756 721898
rect 674612 714946 674664 714952
rect 674612 714888 674664 714894
rect 674624 708424 674652 714888
rect 674716 708560 674744 721892
rect 674704 708554 674756 708560
rect 674704 708496 674756 708502
rect 674612 708418 674664 708424
rect 674612 708360 674664 708366
rect 674704 706582 674756 706588
rect 674704 706524 674756 706530
rect 674716 693736 674744 706524
rect 674704 693730 674756 693736
rect 674704 693672 674756 693678
rect 674808 692240 674836 744264
rect 674900 734400 674928 745177
rect 674992 744328 675020 821512
rect 675084 790500 675112 828024
rect 675256 828030 675308 828036
rect 675256 827972 675308 827978
rect 675164 821570 675216 821576
rect 675164 821512 675216 821518
rect 675176 808316 675204 821512
rect 675268 811444 675296 827972
rect 675452 821576 675480 836132
rect 675544 828036 675572 837220
rect 675532 828030 675584 828036
rect 675532 827972 675584 827978
rect 677292 822584 677490 822612
rect 677292 822499 677320 822584
rect 677278 822490 677334 822499
rect 677278 822425 677334 822434
rect 675440 821570 675492 821576
rect 675440 821512 675492 821518
rect 675256 811438 675308 811444
rect 675256 811380 675308 811386
rect 675348 811438 675400 811444
rect 675348 811380 675400 811386
rect 675164 808310 675216 808316
rect 675164 808252 675216 808258
rect 675360 798660 675388 811380
rect 675440 808310 675492 808316
rect 675440 808252 675492 808258
rect 675348 798654 675400 798660
rect 675348 798596 675400 798602
rect 675452 795804 675480 808252
rect 675532 798654 675584 798660
rect 675532 798596 675584 798602
rect 675164 795798 675216 795804
rect 675164 795740 675216 795746
rect 675440 795798 675492 795804
rect 675440 795740 675492 795746
rect 675072 790494 675124 790500
rect 675072 790436 675124 790442
rect 675072 782946 675124 782952
rect 675072 782888 675124 782894
rect 675084 770100 675112 782888
rect 675176 778600 675204 795740
rect 675544 781592 675572 798596
rect 675532 781586 675584 781592
rect 675532 781528 675584 781534
rect 675268 779008 675296 779078
rect 675256 779002 675308 779008
rect 675256 778944 675308 778950
rect 675164 778594 675216 778600
rect 675164 778536 675216 778542
rect 675176 778422 675282 778450
rect 675176 774248 675204 778422
rect 675164 774242 675216 774248
rect 675164 774184 675216 774190
rect 675176 774098 675282 774126
rect 675072 770094 675124 770100
rect 675072 770036 675124 770042
rect 675176 767652 675204 774098
rect 675256 768530 675308 768536
rect 675256 768472 675308 768478
rect 675164 767646 675216 767652
rect 675164 767588 675216 767594
rect 675268 767532 675296 768472
rect 675084 767504 675296 767532
rect 675084 766036 675112 767504
rect 675164 767442 675216 767448
rect 675164 767384 675216 767390
rect 675176 766122 675204 767384
rect 675176 766094 675282 766122
rect 675084 766008 675204 766036
rect 675072 757174 675124 757180
rect 675072 757116 675124 757122
rect 674980 744322 675032 744328
rect 674980 744264 675032 744270
rect 675084 735352 675112 757116
rect 675072 735346 675124 735352
rect 675072 735288 675124 735294
rect 675176 735284 675204 766008
rect 675532 766014 675584 766020
rect 675532 765956 675584 765962
rect 675256 765946 675308 765952
rect 675256 765888 675308 765894
rect 675164 735278 675216 735284
rect 675164 735220 675216 735226
rect 675268 735164 675296 765888
rect 675544 758064 675572 765956
rect 675532 758058 675584 758064
rect 675532 758000 675584 758006
rect 675716 758058 675768 758064
rect 675716 758000 675768 758006
rect 675728 745251 675756 758000
rect 675438 745242 675494 745251
rect 675438 745177 675494 745186
rect 675714 745242 675770 745251
rect 675714 745177 675770 745186
rect 675452 744435 675480 745177
rect 675438 744426 675494 744435
rect 675438 744361 675494 744370
rect 675176 735136 675296 735164
rect 674888 734394 674940 734400
rect 674888 734336 674940 734342
rect 674888 734258 674940 734264
rect 674888 734200 674940 734206
rect 674900 732331 674928 734200
rect 675176 733124 675204 735136
rect 675176 733096 675296 733124
rect 675268 732580 675296 733096
rect 675268 732552 675388 732580
rect 674886 732322 674942 732331
rect 674886 732257 674942 732266
rect 675360 732172 675388 732552
rect 675176 732144 675388 732172
rect 675176 727820 675204 732144
rect 675254 732050 675310 732059
rect 675254 731985 675310 731994
rect 675084 727792 675204 727820
rect 675084 725236 675112 727792
rect 675176 727698 675282 727726
rect 675176 725356 675204 727698
rect 675164 725350 675216 725356
rect 675164 725292 675216 725298
rect 675084 725208 675204 725236
rect 675072 725078 675124 725084
rect 675072 725020 675124 725026
rect 674980 725010 675032 725016
rect 674980 724952 675032 724958
rect 674992 714952 675020 724952
rect 675084 720256 675112 725020
rect 675072 720250 675124 720256
rect 675072 720192 675124 720198
rect 674980 714946 675032 714952
rect 674980 714888 675032 714894
rect 674888 708554 674940 708560
rect 674888 708496 674940 708502
rect 674900 706588 674928 708496
rect 675176 708424 675204 725208
rect 675256 722086 675308 722092
rect 675256 722028 675308 722034
rect 675268 721179 675296 722028
rect 675254 721170 675310 721179
rect 675254 721105 675310 721114
rect 675256 720250 675308 720256
rect 675256 720192 675308 720198
rect 675268 719708 675296 720192
rect 675530 719538 675586 719547
rect 675530 719473 675586 719482
rect 675438 719266 675494 719275
rect 675438 719201 675494 719210
rect 675072 708418 675124 708424
rect 675072 708360 675124 708366
rect 675164 708418 675216 708424
rect 675164 708360 675216 708366
rect 675348 708418 675400 708424
rect 675348 708360 675400 708366
rect 674888 706582 674940 706588
rect 674888 706524 674940 706530
rect 674888 693730 674940 693736
rect 674888 693672 674940 693678
rect 674796 692234 674848 692240
rect 674796 692176 674848 692182
rect 674704 688766 674756 688772
rect 674704 688708 674756 688714
rect 674716 685660 674744 688708
rect 674900 686460 674928 693672
rect 674980 692234 675032 692240
rect 674980 692176 675032 692182
rect 674888 686454 674940 686460
rect 674888 686396 674940 686402
rect 674796 686318 674848 686324
rect 674796 686260 674848 686266
rect 674440 685632 674744 685660
rect 674440 675512 674468 685632
rect 674610 685402 674666 685411
rect 674610 685337 674666 685346
rect 674520 682646 674572 682652
rect 674520 682588 674572 682594
rect 674532 680068 674560 682588
rect 674520 680062 674572 680068
rect 674520 680004 674572 680010
rect 674520 679926 674572 679932
rect 674520 679868 674572 679874
rect 674428 675506 674480 675512
rect 674428 675448 674480 675454
rect 674440 672860 674468 675448
rect 674428 672854 674480 672860
rect 674428 672796 674480 672802
rect 674532 667012 674560 679868
rect 674624 678180 674652 685337
rect 674808 682652 674836 686260
rect 674796 682646 674848 682652
rect 674796 682588 674848 682594
rect 674888 681218 674940 681224
rect 674888 681160 674940 681166
rect 674796 680062 674848 680068
rect 674796 680004 674848 680010
rect 674808 678316 674836 680004
rect 674900 679812 674928 681160
rect 674992 679932 675020 692176
rect 674980 679926 675032 679932
rect 674980 679868 675032 679874
rect 674900 679784 675020 679812
rect 674808 678288 674928 678316
rect 674624 678152 674836 678180
rect 674808 672928 674836 678152
rect 674796 672922 674848 672928
rect 674796 672864 674848 672870
rect 674520 667006 674572 667012
rect 674520 666948 674572 666954
rect 674796 642050 674848 642056
rect 674796 641992 674848 641998
rect 674704 641234 674756 641240
rect 674704 641176 674756 641182
rect 674716 628388 674744 641176
rect 674808 638996 674836 641992
rect 674796 638990 674848 638996
rect 674796 638932 674848 638938
rect 674704 628382 674756 628388
rect 674704 628324 674756 628330
rect 674808 626416 674836 638932
rect 674796 626410 674848 626416
rect 674796 626352 674848 626358
rect 674796 615530 674848 615536
rect 674796 615472 674848 615478
rect 674808 602616 674836 615472
rect 674796 602610 674848 602616
rect 674796 602552 674848 602558
rect 674796 595538 674848 595544
rect 674796 595480 674848 595486
rect 674428 595470 674480 595476
rect 674428 595412 674480 595418
rect 674440 592251 674468 595412
rect 674808 592416 674836 595480
rect 674796 592410 674848 592416
rect 674796 592352 674848 592358
rect 674426 592242 674482 592251
rect 674426 592177 674482 592186
rect 674440 579836 674468 592177
rect 674704 587446 674756 587452
rect 674704 587388 674756 587394
rect 674716 583388 674744 587388
rect 674808 583508 674836 592352
rect 674796 583502 674848 583508
rect 674796 583444 674848 583450
rect 674716 583360 674836 583388
rect 674808 580448 674836 583360
rect 674796 580442 674848 580448
rect 674796 580384 674848 580390
rect 674428 579830 674480 579836
rect 674428 579772 674480 579778
rect 674520 551134 674572 551140
rect 674520 551076 674572 551082
rect 674532 535568 674560 551076
rect 674796 548890 674848 548896
rect 674796 548832 674848 548838
rect 674808 546720 674836 548832
rect 674796 546714 674848 546720
rect 674796 546656 674848 546662
rect 674612 545150 674664 545156
rect 674612 545092 674664 545098
rect 674520 535562 674572 535568
rect 674520 535504 674572 535510
rect 674624 533120 674652 545092
rect 674808 533256 674836 546656
rect 674796 533250 674848 533256
rect 674796 533192 674848 533198
rect 674612 533114 674664 533120
rect 674612 533056 674664 533062
rect 674796 530870 674848 530876
rect 674796 530812 674848 530818
rect 674808 511564 674836 530812
rect 674796 511558 674848 511564
rect 674796 511500 674848 511506
rect 674900 498683 674928 678288
rect 674992 672996 675020 679784
rect 674980 672990 675032 672996
rect 674980 672932 675032 672938
rect 674980 667006 675032 667012
rect 674980 666948 675032 666954
rect 674992 641240 675020 666948
rect 674980 641234 675032 641240
rect 674980 641176 675032 641182
rect 674980 628382 675032 628388
rect 674980 628324 675032 628330
rect 674992 615536 675020 628324
rect 674980 615530 675032 615536
rect 674980 615472 675032 615478
rect 674980 602610 675032 602616
rect 674980 602552 675032 602558
rect 674992 551140 675020 602552
rect 674980 551134 675032 551140
rect 674980 551076 675032 551082
rect 674980 548822 675032 548828
rect 674980 548764 675032 548770
rect 674992 546176 675020 548764
rect 674980 546170 675032 546176
rect 674980 546112 675032 546118
rect 674980 541478 675032 541484
rect 674980 541420 675032 541426
rect 674992 535704 675020 541420
rect 674980 535698 675032 535704
rect 674980 535640 675032 535646
rect 674980 535562 675032 535568
rect 674980 535504 675032 535510
rect 674992 530876 675020 535504
rect 674980 530870 675032 530876
rect 674980 530812 675032 530818
rect 674980 511558 675032 511564
rect 674980 511500 675032 511506
rect 674886 498674 674942 498683
rect 674612 498638 674664 498644
rect 674886 498609 674888 498618
rect 674612 498580 674664 498586
rect 674940 498609 674942 498618
rect 674888 498580 674940 498586
rect 674624 493243 674652 498580
rect 674992 498576 675020 511500
rect 674796 498570 674848 498576
rect 674796 498512 674848 498518
rect 674980 498570 675032 498576
rect 674980 498512 675032 498518
rect 674808 495283 674836 498512
rect 674794 495274 674850 495283
rect 674794 495209 674850 495218
rect 674610 493234 674666 493243
rect 674610 493169 674666 493178
rect 674704 472866 674756 472872
rect 674704 472808 674756 472814
rect 674716 454512 674744 472808
rect 674704 454506 674756 454512
rect 674704 454448 674756 454454
rect 44044 439818 44096 439824
rect 44044 439760 44096 439766
rect 44872 439818 44924 439824
rect 44872 439760 44924 439766
rect 42294 431354 42350 431363
rect 42294 431289 42350 431298
rect 42296 399290 42348 399296
rect 42296 399232 42348 399238
rect 42308 381888 42336 399232
rect 42388 394938 42440 394944
rect 42388 394880 42440 394886
rect 42400 392768 42428 394880
rect 42480 394870 42532 394876
rect 42480 394812 42532 394818
rect 42388 392762 42440 392768
rect 42388 392704 42440 392710
rect 42296 381882 42348 381888
rect 42296 381824 42348 381830
rect 42400 374408 42428 392704
rect 42492 386784 42520 394812
rect 42480 386778 42532 386784
rect 42480 386720 42532 386726
rect 42388 374402 42440 374408
rect 42388 374344 42440 374350
rect 42388 352234 42440 352240
rect 42388 352176 42440 352182
rect 42296 349582 42348 349588
rect 42296 349524 42348 349530
rect 42308 344488 42336 349524
rect 42400 348704 42428 352176
rect 42572 350262 42624 350268
rect 42572 350204 42624 350210
rect 42388 348698 42440 348704
rect 42388 348640 42440 348646
rect 42388 347746 42440 347752
rect 42388 347688 42440 347694
rect 42296 344482 42348 344488
rect 42296 344424 42348 344430
rect 42400 344216 42428 347688
rect 42480 344618 42532 344624
rect 42480 344560 42532 344566
rect 42388 344210 42440 344216
rect 42388 344152 42440 344158
rect 42388 344006 42440 344012
rect 42388 343948 42440 343954
rect 42400 334424 42428 343948
rect 42492 338300 42520 344560
rect 42480 338294 42532 338300
rect 42480 338236 42532 338242
rect 42584 337688 42612 350204
rect 42572 337682 42624 337688
rect 42572 337624 42624 337630
rect 42584 335172 42612 337624
rect 42572 335166 42624 335172
rect 42572 335108 42624 335114
rect 42388 334418 42440 334424
rect 42388 334360 42440 334366
rect 42388 305926 42440 305932
rect 42388 305868 42440 305874
rect 42296 305382 42348 305388
rect 42296 305324 42348 305330
rect 42308 292779 42336 305324
rect 42400 303348 42428 305868
rect 42388 303342 42440 303348
rect 42388 303284 42440 303290
rect 42400 293488 42428 303284
rect 42388 293482 42440 293488
rect 42388 293424 42440 293430
rect 42294 292770 42350 292779
rect 42294 292705 42350 292714
rect 42216 292456 42428 292484
rect 41928 287430 41980 287436
rect 41928 287372 41980 287378
rect 42112 287430 42164 287436
rect 42112 287372 42164 287378
rect 41940 285956 41968 287372
rect 41940 285928 42152 285956
rect 42124 266764 42152 285928
rect 42400 279700 42428 292456
rect 42216 279672 42428 279700
rect 42112 266758 42164 266764
rect 42112 266700 42164 266706
rect 42112 266622 42164 266628
rect 42112 266564 42164 266570
rect 41744 261318 41796 261324
rect 41744 261260 41796 261266
rect 41586 261082 41692 261110
rect 41664 260576 41692 261082
rect 41652 260570 41704 260576
rect 41652 260512 41704 260518
rect 41652 259686 41704 259692
rect 41652 259628 41704 259634
rect 41664 259270 41692 259628
rect 41586 259242 41692 259270
rect 41652 253634 41704 253640
rect 41652 253576 41704 253582
rect 41664 253106 41692 253576
rect 41586 253078 41692 253106
rect 42124 248782 42152 266564
rect 41586 248754 42152 248782
rect 41558 248162 41614 248171
rect 41558 248097 41614 248106
rect 41928 245610 41980 245616
rect 41742 245578 41798 245587
rect 41652 245542 41704 245548
rect 41928 245552 41980 245558
rect 41742 245513 41798 245522
rect 41652 245484 41704 245490
rect 41664 216755 41692 245484
rect 41650 216746 41706 216755
rect 41650 216681 41706 216690
rect 41756 216596 41784 245513
rect 41940 228208 41968 245552
rect 42124 245548 42152 248754
rect 42112 245542 42164 245548
rect 42112 245484 42164 245490
rect 41928 228202 41980 228208
rect 41928 228144 41980 228150
rect 42112 228202 42164 228208
rect 42112 228144 42164 228150
rect 42124 216716 42152 228144
rect 42112 216710 42164 216716
rect 42112 216652 42164 216658
rect 41756 216568 42152 216596
rect 41586 216482 41692 216510
rect 41664 216036 41692 216482
rect 41652 216030 41704 216036
rect 41652 215972 41704 215978
rect 42124 215220 42152 216568
rect 42112 215214 42164 215220
rect 42112 215156 42164 215162
rect 41652 215146 41704 215152
rect 41652 215088 41704 215094
rect 42110 215114 42166 215123
rect 41664 214692 41692 215088
rect 42110 215049 42166 215058
rect 41586 214664 41692 214692
rect 41664 214171 41692 214664
rect 41650 214162 41706 214171
rect 41650 214097 41706 214106
rect 42124 209780 42152 215049
rect 42112 209774 42164 209780
rect 42112 209716 42164 209722
rect 42110 209674 42166 209683
rect 42110 209609 42166 209618
rect 41652 209570 41704 209576
rect 41652 209512 41704 209518
rect 41664 209275 41692 209512
rect 41650 209266 41706 209275
rect 41650 209201 41706 209210
rect 41652 209026 41704 209032
rect 41652 208968 41704 208974
rect 41664 208506 41692 208968
rect 41586 208478 41692 208506
rect 41558 204196 41614 204205
rect 41558 204131 41614 204140
rect 41586 203512 41692 203540
rect 41664 203116 41692 203512
rect 41652 203110 41704 203116
rect 41652 203052 41704 203058
rect 41650 200970 41706 200979
rect 41650 200905 41706 200914
rect 41664 172244 41692 200905
rect 41836 193250 41888 193256
rect 41836 193192 41888 193198
rect 41848 184076 41876 193192
rect 41836 184070 41888 184076
rect 41836 184012 41888 184018
rect 41928 183934 41980 183940
rect 41928 183876 41980 183882
rect 41940 172312 41968 183876
rect 41928 172306 41980 172312
rect 42124 172283 42152 209609
rect 41928 172248 41980 172254
rect 42110 172274 42166 172283
rect 41652 172238 41704 172244
rect 42110 172209 42166 172218
rect 41652 172180 41704 172186
rect 41586 172096 42152 172124
rect 41558 170284 41614 170293
rect 41558 170219 41614 170228
rect 42124 164134 42152 172096
rect 41572 164106 42152 164134
rect 41572 164086 41600 164106
rect 42020 164010 42072 164016
rect 42020 163952 42072 163958
rect 42032 163556 42060 163952
rect 42032 163528 42152 163556
rect 42124 159884 42152 163528
rect 41756 159856 42152 159884
rect 41756 159782 41784 159856
rect 41586 159754 41784 159782
rect 41586 159110 41692 159138
rect 41664 159052 41692 159110
rect 41652 159046 41704 159052
rect 41652 158988 41704 158994
rect 42124 116008 42152 159856
rect 42216 120467 42244 279672
rect 42388 266758 42440 266764
rect 42388 266700 42440 266706
rect 42296 260570 42348 260576
rect 42296 260512 42348 260518
rect 42308 254184 42336 260512
rect 42400 259692 42428 266700
rect 42664 261318 42716 261324
rect 42664 261260 42716 261266
rect 42388 259686 42440 259692
rect 42388 259628 42440 259634
rect 42296 254178 42348 254184
rect 42296 254120 42348 254126
rect 42400 254116 42428 259628
rect 42388 254110 42440 254116
rect 42388 254052 42440 254058
rect 42676 253980 42704 261260
rect 42296 253974 42348 253980
rect 42296 253916 42348 253922
rect 42664 253974 42716 253980
rect 42664 253916 42716 253922
rect 42308 248171 42336 253916
rect 42388 253906 42440 253912
rect 42388 253848 42440 253854
rect 42294 248162 42350 248171
rect 42294 248097 42350 248106
rect 42400 245616 42428 253848
rect 42388 245610 42440 245616
rect 42388 245552 42440 245558
rect 42480 216710 42532 216716
rect 42480 216652 42532 216658
rect 42296 216030 42348 216036
rect 42296 215972 42348 215978
rect 42308 209032 42336 215972
rect 42492 215288 42520 216652
rect 42480 215282 42532 215288
rect 42480 215224 42532 215230
rect 42388 215214 42440 215220
rect 42388 215156 42440 215162
rect 42296 209026 42348 209032
rect 42296 208968 42348 208974
rect 42400 203116 42428 215156
rect 42388 203110 42440 203116
rect 42388 203052 42440 203058
rect 42400 193256 42428 203052
rect 42388 193250 42440 193256
rect 42388 193192 42440 193198
rect 42388 172306 42440 172312
rect 42388 172248 42440 172254
rect 42296 172238 42348 172244
rect 42296 172180 42348 172186
rect 42308 164152 42336 172180
rect 42296 164146 42348 164152
rect 42296 164088 42348 164094
rect 42400 160700 42428 172248
rect 42662 170234 42718 170243
rect 42662 170169 42718 170178
rect 42308 160672 42428 160700
rect 42308 159052 42336 160672
rect 42676 159340 42704 170169
rect 42584 159312 42704 159340
rect 42296 159046 42348 159052
rect 42296 158988 42348 158994
rect 42308 155516 42336 158988
rect 42296 155510 42348 155516
rect 42296 155452 42348 155458
rect 42584 154632 42612 159312
rect 42480 154626 42532 154632
rect 42480 154568 42532 154574
rect 42572 154626 42624 154632
rect 42572 154568 42624 154574
rect 42492 154496 42520 154568
rect 42296 154490 42348 154496
rect 42296 154432 42348 154438
rect 42480 154490 42532 154496
rect 42480 154432 42532 154438
rect 42308 141780 42336 154432
rect 42296 141774 42348 141780
rect 42296 141716 42348 141722
rect 42572 141774 42624 141780
rect 42572 141716 42624 141722
rect 42584 132532 42612 141716
rect 42388 132526 42440 132532
rect 42388 132468 42440 132474
rect 42572 132526 42624 132532
rect 42572 132468 42624 132474
rect 42400 128792 42428 132468
rect 42388 128786 42440 128792
rect 42388 128728 42440 128734
rect 42480 128786 42532 128792
rect 42480 128728 42532 128734
rect 42202 120458 42258 120467
rect 42202 120393 42258 120402
rect 39904 116002 39956 116008
rect 39470 115950 39904 115956
rect 39470 115944 39956 115950
rect 40364 116002 40416 116008
rect 40364 115944 40416 115950
rect 42112 116002 42164 116008
rect 42112 115944 42164 115950
rect 39470 115928 39944 115944
rect 39260 84722 39312 84728
rect 39260 84664 39312 84670
rect 39272 80188 39300 84664
rect 39194 80160 39300 80188
rect 39417 76352 39668 76380
rect 39417 76094 39445 76352
rect 39640 75972 39668 76352
rect 39640 75944 39760 75972
rect 39732 72692 39760 75944
rect 39720 72686 39772 72692
rect 39720 72628 39772 72634
rect 40376 69444 40404 115944
rect 42216 112987 42244 120393
rect 42492 119680 42520 128728
rect 42480 119674 42532 119680
rect 42480 119616 42532 119622
rect 42388 119606 42440 119612
rect 42388 119548 42440 119554
rect 42400 115956 42428 119548
rect 42400 115928 42520 115956
rect 42202 112978 42258 112987
rect 42202 112913 42258 112922
rect 42492 109480 42520 115928
rect 43030 112978 43086 112987
rect 43030 112913 43086 112922
rect 42204 109474 42256 109480
rect 42204 109416 42256 109422
rect 42480 109474 42532 109480
rect 42480 109416 42532 109422
rect 42216 93840 42244 109416
rect 42204 93834 42256 93840
rect 42204 93776 42256 93782
rect 42388 93834 42440 93840
rect 42388 93776 42440 93782
rect 42400 90168 42428 93776
rect 42112 90162 42164 90168
rect 42112 90104 42164 90110
rect 42388 90162 42440 90168
rect 42388 90104 42440 90110
rect 42124 77316 42152 90104
rect 42112 77310 42164 77316
rect 42112 77252 42164 77258
rect 42296 77310 42348 77316
rect 42296 77252 42348 77258
rect 42308 76947 42336 77252
rect 42294 76938 42350 76947
rect 42294 76873 42350 76882
rect 39194 69416 40404 69444
rect 39548 67184 39576 69416
rect 39536 67178 39588 67184
rect 39536 67120 39588 67126
rect 43044 45084 43072 112913
rect 44884 100164 44912 439760
rect 672404 430570 672456 430576
rect 672404 430512 672456 430518
rect 672416 423300 672444 430512
rect 672404 423294 672456 423300
rect 672404 423236 672456 423242
rect 668632 423226 668684 423232
rect 668632 423168 668684 423174
rect 668644 408544 668672 423168
rect 664676 408538 664728 408544
rect 664676 408480 664728 408486
rect 668632 408538 668684 408544
rect 668632 408480 668684 408486
rect 664688 404872 664716 408480
rect 674808 406611 674836 495209
rect 674978 493234 675034 493243
rect 674978 493169 675034 493178
rect 674992 472872 675020 493169
rect 674980 472866 675032 472872
rect 674980 472808 675032 472814
rect 674888 454506 674940 454512
rect 674888 454448 674940 454454
rect 674900 441676 674928 454448
rect 675084 449723 675112 708360
rect 675164 705698 675216 705704
rect 675164 705640 675216 705646
rect 675176 688772 675204 705640
rect 675360 699244 675388 708360
rect 675452 705704 675480 719201
rect 675440 705698 675492 705704
rect 675440 705640 675492 705646
rect 675544 699260 675572 719473
rect 675348 699238 675400 699244
rect 675544 699232 675756 699260
rect 675348 699180 675400 699186
rect 675624 699170 675676 699176
rect 675624 699112 675676 699118
rect 675164 688766 675216 688772
rect 675164 688708 675216 688714
rect 675636 688636 675664 699112
rect 675728 688947 675756 699232
rect 675714 688938 675770 688947
rect 675714 688873 675770 688882
rect 675164 688630 675216 688636
rect 675164 688572 675216 688578
rect 675624 688630 675676 688636
rect 675624 688572 675676 688578
rect 675176 686476 675204 688572
rect 675176 686448 675296 686476
rect 675268 686170 675296 686448
rect 675176 686142 675296 686170
rect 675176 681224 675204 686142
rect 675268 686054 675296 686142
rect 675254 685464 675310 685473
rect 675254 685399 675310 685408
rect 675164 681218 675216 681224
rect 675164 681160 675216 681166
rect 675176 681098 675282 681126
rect 675176 673692 675204 681098
rect 675256 675506 675308 675512
rect 675256 675448 675308 675454
rect 675268 674948 675296 675448
rect 675176 673664 675388 673692
rect 675360 673148 675388 673664
rect 675282 673120 675388 673148
rect 675256 672990 675308 672996
rect 675256 672932 675308 672938
rect 675268 642056 675296 672932
rect 675624 672922 675676 672928
rect 675624 672864 675676 672870
rect 675348 672854 675400 672860
rect 675348 672796 675400 672802
rect 675256 642050 675308 642056
rect 675360 642027 675388 672796
rect 675636 642163 675664 672864
rect 675622 642154 675678 642163
rect 675622 642089 675678 642098
rect 675256 641992 675308 641998
rect 675346 642018 675402 642027
rect 675346 641953 675402 641962
rect 675268 638996 675296 639480
rect 675256 638990 675308 638996
rect 675256 638932 675308 638938
rect 675254 638890 675310 638899
rect 675254 638825 675310 638834
rect 675176 634496 675282 634524
rect 675176 627044 675204 634496
rect 675254 628376 675310 628385
rect 675254 628311 675310 628320
rect 675176 627016 675296 627044
rect 675268 626486 675296 627016
rect 675256 626410 675308 626416
rect 675162 626378 675218 626387
rect 675256 626352 675308 626358
rect 675530 626378 675586 626387
rect 675162 626313 675218 626322
rect 675176 595476 675204 626313
rect 675268 595544 675296 626352
rect 675530 626313 675586 626322
rect 675544 609076 675572 626313
rect 675348 609070 675400 609076
rect 675348 609012 675400 609018
rect 675532 609070 675584 609076
rect 675532 609012 675584 609018
rect 675256 595538 675308 595544
rect 675256 595480 675308 595486
rect 675164 595470 675216 595476
rect 675164 595412 675216 595418
rect 675360 595356 675388 609012
rect 675176 595328 675388 595356
rect 675176 583411 675204 595328
rect 675268 592416 675296 592894
rect 675256 592410 675308 592416
rect 675256 592352 675308 592358
rect 675254 592242 675310 592251
rect 675254 592177 675310 592186
rect 675268 587452 675296 587912
rect 675256 587446 675308 587452
rect 675256 587388 675308 587394
rect 675162 583402 675218 583411
rect 675162 583337 675218 583346
rect 675256 583366 675308 583372
rect 675256 583308 675308 583314
rect 675268 583252 675296 583308
rect 675176 583224 675296 583252
rect 675176 557464 675204 583224
rect 675254 581770 675310 581779
rect 675254 581705 675310 581714
rect 675256 580442 675308 580448
rect 675256 580384 675308 580390
rect 675268 579908 675296 580384
rect 675256 579830 675308 579836
rect 675256 579772 675308 579778
rect 675164 557458 675216 557464
rect 675164 557400 675216 557406
rect 675164 551134 675216 551140
rect 675164 551076 675216 551082
rect 675176 541484 675204 551076
rect 675268 548828 675296 579772
rect 675346 579730 675402 579739
rect 675346 579665 675402 579674
rect 675360 551140 675388 579665
rect 677462 573202 677518 573211
rect 677462 573137 677518 573146
rect 677476 566780 677504 573137
rect 677464 566774 677516 566780
rect 677464 566716 677516 566722
rect 677740 566774 677792 566780
rect 677740 566716 677792 566722
rect 675440 557458 675492 557464
rect 675440 557400 675492 557406
rect 675348 551134 675400 551140
rect 675348 551076 675400 551082
rect 675452 548896 675480 557400
rect 677752 550091 677780 566716
rect 677738 550082 677794 550091
rect 677738 550017 677794 550026
rect 675440 548890 675492 548896
rect 675440 548832 675492 548838
rect 675256 548822 675308 548828
rect 675256 548764 675308 548770
rect 675256 546714 675308 546720
rect 675256 546656 675308 546662
rect 675268 546280 675296 546656
rect 675348 546170 675400 546176
rect 675348 546112 675400 546118
rect 675360 545650 675388 546112
rect 675282 545636 675388 545650
rect 675268 545622 675388 545636
rect 675268 545156 675296 545622
rect 675256 545150 675308 545156
rect 675256 545092 675308 545098
rect 675164 541478 675216 541484
rect 675164 541420 675216 541426
rect 675176 541298 675282 541326
rect 675176 533884 675204 541298
rect 675256 535698 675308 535704
rect 675256 535640 675308 535646
rect 675268 535148 675296 535640
rect 675176 533856 675388 533884
rect 675164 533250 675216 533256
rect 675268 533238 675296 533326
rect 675360 533238 675388 533856
rect 675268 533210 675388 533238
rect 675164 533192 675216 533198
rect 675070 449714 675126 449723
rect 675070 449649 675126 449658
rect 674900 441648 675020 441676
rect 674992 428915 675020 441648
rect 674978 428906 675034 428915
rect 674978 428841 675034 428850
rect 674886 425098 674942 425107
rect 674886 425033 674888 425042
rect 674940 425033 674942 425042
rect 675072 425062 675124 425068
rect 674888 425004 674940 425010
rect 675072 425004 675124 425010
rect 675084 415700 675112 425004
rect 674992 415672 675112 415700
rect 674794 406602 674850 406611
rect 674794 406537 674850 406546
rect 663112 404866 663164 404872
rect 663112 404808 663164 404814
rect 664676 404866 664728 404872
rect 664676 404808 664728 404814
rect 663124 359040 663152 404808
rect 674992 403052 675020 415672
rect 674992 403024 675112 403052
rect 675084 401715 675112 403024
rect 675070 401706 675126 401715
rect 675070 401641 675126 401650
rect 675176 365772 675204 533192
rect 675256 533114 675308 533120
rect 675256 533056 675308 533062
rect 675268 447100 675296 533056
rect 677922 459914 677978 459923
rect 677922 459849 677978 459858
rect 677936 452964 677964 459849
rect 677752 452950 677964 452964
rect 677752 452936 677950 452950
rect 677752 452171 677780 452936
rect 677738 452162 677794 452171
rect 677738 452097 677794 452106
rect 677568 448176 677896 448204
rect 677568 447100 677596 448176
rect 675256 447094 675308 447100
rect 675256 447036 675308 447042
rect 677556 447094 677608 447100
rect 677556 447036 677608 447042
rect 675164 365766 675216 365772
rect 675164 365708 675216 365714
rect 675268 365652 675296 447036
rect 677936 437988 677964 442070
rect 675348 437982 675400 437988
rect 675348 437924 675400 437930
rect 677924 437982 677976 437988
rect 677924 437924 677976 437930
rect 675360 430644 675388 437924
rect 675348 430638 675400 430644
rect 675348 430580 675400 430586
rect 677462 406602 677518 406611
rect 677462 406537 677518 406546
rect 675084 365624 675296 365652
rect 675084 362984 675112 365624
rect 675164 365562 675216 365568
rect 675164 365504 675216 365510
rect 675176 363340 675204 365504
rect 675176 363312 675296 363340
rect 675072 362978 675124 362984
rect 675072 362920 675124 362926
rect 675176 362100 675204 363312
rect 675268 363054 675296 363312
rect 675256 362978 675308 362984
rect 675256 362920 675308 362926
rect 675164 362094 675216 362100
rect 675164 362036 675216 362042
rect 675268 361980 675296 362920
rect 674992 361952 675296 361980
rect 660444 359034 660496 359040
rect 660444 358976 660496 358982
rect 663112 359034 663164 359040
rect 663112 358976 663164 358982
rect 660456 353412 660484 358976
rect 674888 357606 674940 357612
rect 674888 357548 674940 357554
rect 674796 356926 674848 356932
rect 674796 356868 674848 356874
rect 660364 353384 660484 353412
rect 660364 350064 660392 353384
rect 657132 350058 657184 350064
rect 657132 350000 657184 350006
rect 660352 350058 660404 350064
rect 660352 350000 660404 350006
rect 657144 344828 657172 350000
rect 674808 349928 674836 356868
rect 674900 350171 674928 357548
rect 674992 357084 675020 361952
rect 675164 361890 675216 361896
rect 675164 361832 675216 361838
rect 675176 358308 675204 361832
rect 675084 358280 675204 358308
rect 675084 357204 675112 358280
rect 675268 357612 675296 358112
rect 675256 357606 675308 357612
rect 675256 357548 675308 357554
rect 675072 357198 675124 357204
rect 675072 357140 675124 357146
rect 674992 357056 675112 357084
rect 675084 356932 675112 357056
rect 675164 356994 675216 357000
rect 675162 356962 675164 356971
rect 675216 356962 675218 356971
rect 675072 356926 675124 356932
rect 675162 356897 675218 356906
rect 675072 356868 675124 356874
rect 674978 356690 675034 356699
rect 674978 356625 675034 356634
rect 674886 350162 674942 350171
rect 674886 350097 674942 350106
rect 674992 349996 675020 356625
rect 675176 351934 675282 351962
rect 674980 349990 675032 349996
rect 674980 349932 675032 349938
rect 674796 349922 674848 349928
rect 674796 349864 674848 349870
rect 655752 344822 655804 344828
rect 655752 344764 655804 344770
rect 657132 344822 657184 344828
rect 657132 344764 657184 344770
rect 655764 331296 655792 344764
rect 655752 331290 655804 331296
rect 655752 331232 655804 331238
rect 651244 331222 651296 331228
rect 651244 331164 651296 331170
rect 651256 319396 651284 331164
rect 649404 319390 649456 319396
rect 649404 319332 649456 319338
rect 651244 319390 651296 319396
rect 651244 319332 651296 319338
rect 649416 313888 649444 319332
rect 675176 319124 675204 351934
rect 675254 350162 675310 350171
rect 675254 350097 675310 350106
rect 675348 349990 675400 349996
rect 675348 349932 675400 349938
rect 675256 349922 675308 349928
rect 675256 349864 675308 349870
rect 675164 319118 675216 319124
rect 675164 319060 675216 319066
rect 675268 319004 675296 349864
rect 675360 319027 675388 349932
rect 675084 318976 675296 319004
rect 675346 319018 675402 319027
rect 675084 316404 675112 318976
rect 675346 318953 675402 318962
rect 675164 318914 675216 318920
rect 675164 318856 675216 318862
rect 675072 316398 675124 316404
rect 675072 316340 675124 316346
rect 675176 315468 675204 318856
rect 675254 316508 675310 316517
rect 675254 316443 675310 316452
rect 675256 316398 675308 316404
rect 675256 316340 675308 316346
rect 674992 315440 675204 315468
rect 640848 313882 640900 313888
rect 640848 313824 640900 313830
rect 649404 313882 649456 313888
rect 649404 313824 649456 313830
rect 640860 310284 640888 313824
rect 636892 310278 636944 310284
rect 636892 310220 636944 310226
rect 640848 310278 640900 310284
rect 640848 310220 640900 310226
rect 636904 306476 636932 310220
rect 674888 309122 674940 309128
rect 674888 309064 674940 309070
rect 634684 306470 634736 306476
rect 634684 306412 634736 306418
rect 636892 306470 636944 306476
rect 636892 306412 636944 306418
rect 634696 300016 634724 306412
rect 634684 300010 634736 300016
rect 634684 299952 634736 299958
rect 630360 299942 630412 299948
rect 630360 299884 630412 299890
rect 630372 294440 630400 299884
rect 674900 296276 674928 309064
rect 674992 304980 675020 315440
rect 675268 315332 675296 316340
rect 675176 315304 675296 315332
rect 675176 311660 675204 315304
rect 675084 311632 675204 311660
rect 675084 309128 675112 311632
rect 675176 311496 675282 311524
rect 675072 309122 675124 309128
rect 675072 309064 675124 309070
rect 674980 304974 675032 304980
rect 674980 304916 675032 304922
rect 674992 303416 675020 304916
rect 675176 304044 675204 311496
rect 675268 304980 675296 305348
rect 675256 304974 675308 304980
rect 675256 304916 675308 304922
rect 675176 304016 675296 304044
rect 675268 303486 675296 304016
rect 674980 303410 675032 303416
rect 674980 303352 675032 303358
rect 675440 303410 675492 303416
rect 675440 303352 675492 303358
rect 674888 296270 674940 296276
rect 674888 296212 674940 296218
rect 675348 296270 675400 296276
rect 675348 296212 675400 296218
rect 675360 296156 675388 296212
rect 675176 296128 675388 296156
rect 630360 294434 630412 294440
rect 630360 294376 630412 294382
rect 620700 294298 620752 294304
rect 620700 294240 620752 294246
rect 620712 286348 620740 294240
rect 615548 286342 615600 286348
rect 615548 286284 615600 286290
rect 620700 286342 620752 286348
rect 620700 286284 620752 286290
rect 615560 284172 615588 286284
rect 613432 284166 613484 284172
rect 613432 284108 613484 284114
rect 615548 284166 615600 284172
rect 615548 284108 615600 284114
rect 613444 276080 613472 284108
rect 613432 276074 613484 276080
rect 613432 276016 613484 276022
rect 609752 276006 609804 276012
rect 609752 275948 609804 275954
rect 609764 264996 609792 275948
rect 675176 274176 675204 296128
rect 674796 274170 674848 274176
rect 674796 274112 674848 274118
rect 675164 274170 675216 274176
rect 675164 274112 675216 274118
rect 674808 268940 674836 274112
rect 675452 272612 675480 303352
rect 675164 272606 675216 272612
rect 675164 272548 675216 272554
rect 675440 272606 675492 272612
rect 675440 272548 675492 272554
rect 674980 269614 675032 269620
rect 674980 269556 675032 269562
rect 674796 268934 674848 268940
rect 674796 268876 674848 268882
rect 605336 264990 605388 264996
rect 605336 264932 605388 264938
rect 609752 264990 609804 264996
rect 609752 264932 609804 264938
rect 605348 262208 605376 264932
rect 600552 262202 600604 262208
rect 600552 262144 600604 262150
rect 605336 262202 605388 262208
rect 605336 262144 605388 262150
rect 600564 248472 600592 262144
rect 674808 256988 674836 268876
rect 674888 264718 674940 264724
rect 674888 264660 674940 264666
rect 674900 259284 674928 264660
rect 674888 259278 674940 259284
rect 674888 259220 674940 259226
rect 674900 257652 674928 259220
rect 674888 257646 674940 257652
rect 674888 257588 674940 257594
rect 674992 257108 675020 269556
rect 675176 264724 675204 272548
rect 675530 271146 675586 271155
rect 675530 271081 675586 271090
rect 675544 270776 675572 271081
rect 675532 270770 675584 270776
rect 675532 270712 675584 270718
rect 675440 270566 675492 270572
rect 675440 270508 675492 270514
rect 675452 270094 675480 270508
rect 675282 270080 675480 270094
rect 675268 270066 675480 270080
rect 675268 269620 675296 270066
rect 675256 269614 675308 269620
rect 675256 269556 675308 269562
rect 675268 268940 675296 269436
rect 675256 268934 675308 268940
rect 675256 268876 675308 268882
rect 675164 264718 675216 264724
rect 675164 264660 675216 264666
rect 675268 264604 675296 265134
rect 675176 264576 675296 264604
rect 675176 259556 675204 264576
rect 675164 259550 675216 259556
rect 675164 259492 675216 259498
rect 675164 259346 675216 259352
rect 675164 259288 675216 259294
rect 675176 257124 675204 259288
rect 675256 259278 675308 259284
rect 675256 259220 675308 259226
rect 675268 258948 675296 259220
rect 675348 257646 675400 257652
rect 675348 257588 675400 257594
rect 675360 257244 675388 257588
rect 675348 257238 675400 257244
rect 675348 257180 675400 257186
rect 674980 257102 675032 257108
rect 675176 257096 675282 257124
rect 674980 257044 675032 257050
rect 675348 257034 675400 257040
rect 674808 256960 675204 256988
rect 675348 256976 675400 256982
rect 675532 257034 675584 257040
rect 675532 256976 675584 256982
rect 600552 248466 600604 248472
rect 600552 248408 600604 248414
rect 594112 248398 594164 248404
rect 594112 248340 594164 248346
rect 594124 242964 594152 248340
rect 594112 242958 594164 242964
rect 594112 242900 594164 242906
rect 590432 242890 590484 242896
rect 590432 242832 590484 242838
rect 590444 234940 590472 242832
rect 675176 241060 675204 256960
rect 675164 241054 675216 241060
rect 675164 240996 675216 241002
rect 587672 234934 587724 234940
rect 587672 234876 587724 234882
rect 590432 234934 590484 234940
rect 590432 234876 590484 234882
rect 587684 221476 587712 234876
rect 674980 226094 675032 226100
rect 674980 226036 675032 226042
rect 674888 226026 674940 226032
rect 674888 225968 674940 225974
rect 585832 221470 585884 221476
rect 585832 221412 585884 221418
rect 587672 221470 587724 221476
rect 587672 221412 587724 221418
rect 585844 206176 585872 221412
rect 674900 212403 674928 225968
rect 674992 223380 675020 226036
rect 675360 225980 675388 256976
rect 675440 241054 675492 241060
rect 675440 240996 675492 241002
rect 675452 226100 675480 240996
rect 675440 226094 675492 226100
rect 675440 226036 675492 226042
rect 675544 226032 675572 256976
rect 675084 225952 675388 225980
rect 675532 226026 675584 226032
rect 675532 225968 675584 225974
rect 675084 223940 675112 225952
rect 675084 223912 675296 223940
rect 674980 223374 675032 223380
rect 674980 223316 675032 223322
rect 675268 222972 675296 223912
rect 675348 223374 675400 223380
rect 675348 223316 675400 223322
rect 675256 222966 675308 222972
rect 675256 222908 675308 222914
rect 675360 222852 675388 223316
rect 675282 222838 675388 222852
rect 675268 222824 675388 222838
rect 675164 222694 675216 222700
rect 675164 222636 675216 222642
rect 675176 222444 675204 222636
rect 675084 222416 675204 222444
rect 675084 222308 675112 222416
rect 675268 222308 675296 222824
rect 674992 222280 675112 222308
rect 675176 222280 675296 222308
rect 674886 212394 674942 212403
rect 674886 212329 674942 212338
rect 674900 210392 674928 212329
rect 674888 210386 674940 210392
rect 674888 210328 674940 210334
rect 674992 210256 675020 222280
rect 675176 218092 675204 222280
rect 675254 218514 675310 218523
rect 675254 218449 675310 218458
rect 675254 218378 675310 218387
rect 675254 218313 675310 218322
rect 675084 218064 675204 218092
rect 675084 210340 675112 218064
rect 675268 217956 675296 218313
rect 675176 217928 675296 217956
rect 675176 210522 675204 217928
rect 675254 212394 675310 212403
rect 675254 212329 675310 212338
rect 675176 210494 675282 210522
rect 675256 210386 675308 210392
rect 675084 210312 675204 210340
rect 675256 210328 675308 210334
rect 674980 210250 675032 210256
rect 674980 210192 675032 210198
rect 585832 206170 585884 206176
rect 585832 206112 585884 206118
rect 581508 206102 581560 206108
rect 581508 206044 581560 206050
rect 581520 200668 581548 206044
rect 578104 200662 578156 200668
rect 578104 200604 578156 200610
rect 581508 200662 581560 200668
rect 581508 200604 581560 200610
rect 578116 198764 578144 200604
rect 573964 198758 574016 198764
rect 573964 198700 574016 198706
rect 578104 198758 578156 198764
rect 578104 198700 578156 198706
rect 573976 191964 574004 198700
rect 570652 191958 570704 191964
rect 570652 191900 570704 191906
rect 573964 191958 574016 191964
rect 573964 191900 574016 191906
rect 570664 187748 570692 191900
rect 675176 189448 675204 210312
rect 675268 189555 675296 210328
rect 675348 210250 675400 210256
rect 675348 210192 675400 210198
rect 675254 189546 675310 189555
rect 675360 189532 675388 210192
rect 675360 189504 675756 189532
rect 675254 189481 675310 189490
rect 675164 189442 675216 189448
rect 675164 189384 675216 189390
rect 675348 189442 675400 189448
rect 675348 189384 675400 189390
rect 675622 189410 675678 189419
rect 566604 187742 566656 187748
rect 566604 187684 566656 187690
rect 570652 187742 570704 187748
rect 570652 187684 570704 187690
rect 566616 180420 566644 187684
rect 566524 180392 566644 180420
rect 566524 178568 566552 180392
rect 675360 179876 675388 189384
rect 675622 189345 675678 189354
rect 674980 179854 675032 179860
rect 674980 179796 675032 179802
rect 675084 179848 675388 179876
rect 675636 179860 675664 189345
rect 675624 179854 675676 179860
rect 555012 178562 555064 178568
rect 555012 178504 555064 178510
rect 566512 178562 566564 178568
rect 566512 178504 566564 178510
rect 555024 167620 555052 178504
rect 674888 175706 674940 175712
rect 674888 175648 674940 175654
rect 552160 167614 552212 167620
rect 552160 167556 552212 167562
rect 555012 167614 555064 167620
rect 555012 167556 555064 167562
rect 552172 164900 552200 167556
rect 674796 167410 674848 167416
rect 674796 167352 674848 167358
rect 674808 165376 674836 167352
rect 674796 165370 674848 165376
rect 674796 165312 674848 165318
rect 550044 164894 550096 164900
rect 550044 164836 550096 164842
rect 552160 164894 552212 164900
rect 552160 164836 552212 164842
rect 550056 155788 550084 164836
rect 674808 157216 674836 165312
rect 674900 163812 674928 175648
rect 674992 167416 675020 179796
rect 675084 176800 675112 179848
rect 675624 179796 675676 179802
rect 675728 179724 675756 189504
rect 675164 179718 675216 179724
rect 675164 179660 675216 179666
rect 675716 179718 675768 179724
rect 675716 179660 675768 179666
rect 675176 176884 675204 179660
rect 675176 176870 675282 176884
rect 675176 176856 675296 176870
rect 675072 176794 675124 176800
rect 675072 176736 675124 176742
rect 675268 176340 675296 176856
rect 675348 176794 675400 176800
rect 675348 176736 675400 176742
rect 675084 176312 675296 176340
rect 674980 167410 675032 167416
rect 674980 167352 675032 167358
rect 675084 163828 675112 176312
rect 675360 176250 675388 176736
rect 675282 176236 675388 176250
rect 675268 176222 675388 176236
rect 675268 175712 675296 176222
rect 675256 175706 675308 175712
rect 675256 175648 675308 175654
rect 675176 171898 675282 171926
rect 675176 163922 675204 171898
rect 675268 165376 675296 165748
rect 675256 165370 675308 165376
rect 675256 165312 675308 165318
rect 675176 163894 675282 163922
rect 674888 163806 674940 163812
rect 675084 163800 675204 163828
rect 674888 163748 674940 163754
rect 675176 157352 675204 163800
rect 675348 163806 675400 163812
rect 675348 163748 675400 163754
rect 675164 157346 675216 157352
rect 675164 157288 675216 157294
rect 674796 157210 674848 157216
rect 674796 157152 674848 157158
rect 675164 157210 675216 157216
rect 675164 157152 675216 157158
rect 546364 155782 546416 155788
rect 546364 155724 546416 155730
rect 550044 155782 550096 155788
rect 550044 155724 550096 155730
rect 87192 155510 87244 155516
rect 87192 155452 87244 155458
rect 87204 141712 87232 155452
rect 546376 151844 546404 155724
rect 542684 151838 542736 151844
rect 542684 151780 542736 151786
rect 546364 151838 546416 151844
rect 546364 151780 546416 151786
rect 542696 143616 542724 151780
rect 542684 143610 542736 143616
rect 542684 143552 542736 143558
rect 540016 143542 540068 143548
rect 540016 143484 540068 143490
rect 540028 143428 540056 143484
rect 539936 143400 540056 143428
rect 87192 141706 87244 141712
rect 87192 141648 87244 141654
rect 88664 141706 88716 141712
rect 88664 141648 88716 141654
rect 88676 134368 88704 141648
rect 539936 137988 539964 143400
rect 539936 137960 540148 137988
rect 675176 137972 675204 157152
rect 88664 134362 88716 134368
rect 88664 134304 88716 134310
rect 90872 134362 90924 134368
rect 90872 134304 90924 134310
rect 90884 118796 90912 134304
rect 90872 118790 90924 118796
rect 90872 118732 90924 118738
rect 92528 118790 92580 118796
rect 92528 118732 92580 118738
rect 92540 115940 92568 118732
rect 92528 115934 92580 115940
rect 92528 115876 92580 115882
rect 94000 115934 94052 115940
rect 94000 115876 94052 115882
rect 94012 108596 94040 115876
rect 94000 108590 94052 108596
rect 94000 108532 94052 108538
rect 97404 108522 97456 108528
rect 97404 108464 97456 108470
rect 97416 102544 97444 108464
rect 97404 102538 97456 102544
rect 97404 102480 97456 102486
rect 99704 102538 99756 102544
rect 99704 102480 99756 102486
rect 44872 100158 44924 100164
rect 44872 100100 44924 100106
rect 45792 100158 45844 100164
rect 45792 100100 45844 100106
rect 45804 99960 45832 100100
rect 45792 99954 45844 99960
rect 45792 99896 45844 99902
rect 45804 85612 45832 99896
rect 99716 99892 99744 102480
rect 540120 99960 540148 137960
rect 675164 137966 675216 137972
rect 675164 137908 675216 137914
rect 674888 132866 674940 132872
rect 674888 132808 674940 132814
rect 674900 130100 674928 132808
rect 675360 132804 675388 163748
rect 675440 157346 675492 157352
rect 675440 157288 675492 157294
rect 675452 132804 675480 157288
rect 675532 137966 675584 137972
rect 675532 137908 675584 137914
rect 675544 132872 675572 137908
rect 675532 132866 675584 132872
rect 675532 132808 675584 132814
rect 675348 132798 675400 132804
rect 675348 132740 675400 132746
rect 675440 132798 675492 132804
rect 675440 132740 675492 132746
rect 675072 132730 675124 132736
rect 675072 132672 675124 132678
rect 675084 130100 675112 132672
rect 675532 132594 675584 132600
rect 675532 132536 675584 132542
rect 675544 132276 675572 132536
rect 675176 132248 675572 132276
rect 675176 130294 675204 132248
rect 675254 130308 675310 130317
rect 675176 130266 675254 130294
rect 675254 130243 675310 130252
rect 674900 130072 675020 130100
rect 675084 130072 675296 130100
rect 674992 129964 675020 130072
rect 674992 129936 675204 129964
rect 674980 129126 675032 129132
rect 674980 129068 675032 129074
rect 674888 119946 674940 119952
rect 674888 119888 674940 119894
rect 674900 118728 674928 119888
rect 674888 118722 674940 118728
rect 674888 118664 674940 118670
rect 674900 117044 674928 118664
rect 674992 117180 675020 129068
rect 675176 124916 675204 129936
rect 675268 129132 675296 130072
rect 675256 129126 675308 129132
rect 675256 129068 675308 129074
rect 675164 124910 675216 124916
rect 675164 124852 675216 124858
rect 675268 124796 675296 125326
rect 675084 124768 675296 124796
rect 675084 119884 675112 124768
rect 675164 124706 675216 124712
rect 675164 124648 675216 124654
rect 675176 119952 675204 124648
rect 675164 119946 675216 119952
rect 675164 119888 675216 119894
rect 675072 119878 675124 119884
rect 675072 119820 675124 119826
rect 675070 119778 675126 119787
rect 675070 119713 675126 119722
rect 675084 117300 675112 119713
rect 675164 119674 675216 119680
rect 675164 119616 675216 119622
rect 675176 117316 675204 119616
rect 675268 118728 675296 119148
rect 675256 118722 675308 118728
rect 675256 118664 675308 118670
rect 675072 117294 675124 117300
rect 675176 117288 675282 117316
rect 675072 117236 675124 117242
rect 675532 117226 675584 117232
rect 674992 117152 675296 117180
rect 675532 117168 675584 117174
rect 674900 117016 675204 117044
rect 540108 99954 540160 99960
rect 540108 99896 540160 99902
rect 99704 99886 99756 99892
rect 99704 99828 99756 99834
rect 126844 99886 126896 99892
rect 126844 99828 126896 99834
rect 126856 95744 126884 99828
rect 126844 95738 126896 95744
rect 126844 95680 126896 95686
rect 130984 95670 131036 95676
rect 130984 95612 131036 95618
rect 130996 92004 131024 95612
rect 130984 91998 131036 92004
rect 130984 91940 131036 91946
rect 135032 91998 135084 92004
rect 135032 91940 135084 91946
rect 45148 85606 45200 85612
rect 45148 85548 45200 85554
rect 45792 85606 45844 85612
rect 45792 85548 45844 85554
rect 45160 84728 45188 85548
rect 45148 84722 45200 84728
rect 45148 84664 45200 84670
rect 135044 83640 135072 91940
rect 674796 86354 674848 86360
rect 674796 86296 674848 86302
rect 465496 85606 465548 85612
rect 465496 85548 465548 85554
rect 135032 83634 135084 83640
rect 135032 83576 135084 83582
rect 136044 83634 136096 83640
rect 136044 83576 136096 83582
rect 43950 76938 44006 76947
rect 43950 76873 44006 76882
rect 43964 76364 43992 76873
rect 43952 76358 44004 76364
rect 43952 76300 44004 76306
rect 136056 74664 136084 83576
rect 149752 76358 149804 76364
rect 149752 76300 149804 76306
rect 136044 74658 136096 74664
rect 136044 74600 136096 74606
rect 138804 74658 138856 74664
rect 138804 74600 138856 74606
rect 90872 72686 90924 72692
rect 90872 72628 90924 72634
rect 43032 45078 43084 45084
rect 43032 45020 43084 45026
rect 90884 44336 90912 72628
rect 138816 66232 138844 74600
rect 140552 67178 140604 67184
rect 140552 67120 140604 67126
rect 138804 66226 138856 66232
rect 138804 66168 138856 66174
rect 90872 44330 90924 44336
rect 90872 44272 90924 44278
rect 90884 40227 90912 44272
rect 90870 40218 90926 40227
rect 90870 40153 90926 40162
rect 134110 40218 134166 40227
rect 134110 40153 134112 40162
rect 134164 40153 134166 40162
rect 134112 40124 134164 40130
rect 140564 40068 140592 67120
rect 140644 66226 140696 66232
rect 140644 66168 140696 66174
rect 140656 62560 140684 66168
rect 140644 62554 140696 62560
rect 140644 62496 140696 62502
rect 142392 62554 142444 62560
rect 142392 62496 142444 62502
rect 142404 43384 142432 62496
rect 149764 44268 149792 76300
rect 183792 45146 183844 45152
rect 195844 45146 195896 45152
rect 183844 45094 183924 45100
rect 183792 45088 183924 45094
rect 195844 45088 195896 45094
rect 196672 45146 196724 45152
rect 196672 45088 196724 45094
rect 183804 45084 183924 45088
rect 183804 45078 183936 45084
rect 183804 45072 183884 45078
rect 183884 45020 183936 45026
rect 195200 44534 195252 44540
rect 195200 44476 195252 44482
rect 148924 44262 148976 44268
rect 148924 44204 148976 44210
rect 149752 44262 149804 44268
rect 149752 44204 149804 44210
rect 188392 44262 188444 44268
rect 188392 44204 188444 44210
rect 192716 44262 192768 44268
rect 192716 44204 192768 44210
rect 142392 43378 142444 43384
rect 142392 43320 142444 43326
rect 144968 43378 145020 43384
rect 144968 43320 145020 43326
rect 144980 42432 145008 43320
rect 144968 42426 145020 42432
rect 144968 42368 145020 42374
rect 144416 42358 144468 42364
rect 144416 42300 144468 42306
rect 142942 40218 142998 40227
rect 142942 40153 142998 40162
rect 143402 40218 143458 40227
rect 143402 40153 143404 40162
rect 140872 40120 140900 40151
rect 142948 40120 142976 40153
rect 143456 40153 143458 40162
rect 143404 40124 143456 40130
rect 144428 40120 144456 42300
rect 144980 40204 145008 42368
rect 148936 40363 148964 44204
rect 186552 44194 186604 44200
rect 186552 44136 186604 44142
rect 186564 41822 186592 44136
rect 188404 41822 188432 44204
rect 189128 41950 189180 41956
rect 189128 41892 189180 41898
rect 189140 41836 189168 41892
rect 189062 41808 189168 41836
rect 190902 41820 191008 41836
rect 192098 41820 192204 41836
rect 192728 41822 192756 44204
rect 194556 44194 194608 44200
rect 194556 44136 194608 44142
rect 193386 41820 193492 41836
rect 194568 41822 194596 44136
rect 195212 42432 195240 44476
rect 195200 42426 195252 42432
rect 195200 42368 195252 42374
rect 195212 41822 195240 42368
rect 195856 41822 195884 45088
rect 196684 44744 196712 45088
rect 218842 44842 218898 44851
rect 218842 44777 218844 44786
rect 218896 44777 218898 44786
rect 231630 44842 231686 44851
rect 231630 44777 231686 44786
rect 244602 44842 244658 44851
rect 244602 44777 244604 44786
rect 218844 44748 218896 44754
rect 231644 44744 231672 44777
rect 244656 44777 244658 44786
rect 257390 44842 257446 44851
rect 424922 44842 424978 44851
rect 273964 44812 274176 44828
rect 257390 44777 257446 44786
rect 273952 44806 274176 44812
rect 244604 44748 244656 44754
rect 257404 44744 257432 44777
rect 274004 44800 274176 44806
rect 273952 44748 274004 44754
rect 274148 44744 274176 44800
rect 417472 44806 417524 44812
rect 424922 44777 424924 44786
rect 417472 44748 417524 44754
rect 424976 44777 424978 44786
rect 437710 44842 437766 44851
rect 437710 44777 437766 44786
rect 424924 44748 424976 44754
rect 196672 44738 196724 44744
rect 196672 44680 196724 44686
rect 209552 44738 209604 44744
rect 209644 44738 209696 44744
rect 209604 44686 209644 44692
rect 209552 44680 209696 44686
rect 231632 44738 231684 44744
rect 231632 44680 231684 44686
rect 235312 44738 235364 44744
rect 235404 44738 235456 44744
rect 235364 44686 235404 44692
rect 235312 44680 235456 44686
rect 257392 44738 257444 44744
rect 257392 44680 257444 44686
rect 261072 44738 261124 44744
rect 261164 44738 261216 44744
rect 261124 44686 261164 44692
rect 261072 44680 261216 44686
rect 274136 44738 274188 44744
rect 307440 44738 307492 44744
rect 274136 44680 274188 44686
rect 209564 44664 209684 44680
rect 235324 44664 235444 44680
rect 261084 44664 261204 44680
rect 283164 44676 283376 44692
rect 307440 44680 307492 44686
rect 318112 44738 318164 44744
rect 318112 44680 318164 44686
rect 344792 44738 344844 44744
rect 344792 44680 344844 44686
rect 351784 44738 351836 44744
rect 351784 44680 351836 44686
rect 359236 44738 359288 44744
rect 359236 44680 359288 44686
rect 283152 44670 283376 44676
rect 283204 44664 283376 44670
rect 283152 44612 283204 44618
rect 283348 44608 283376 44664
rect 299620 44670 299672 44676
rect 299620 44612 299672 44618
rect 283336 44602 283388 44608
rect 283336 44544 283388 44550
rect 199524 44534 199576 44540
rect 199524 44476 199576 44482
rect 198880 44330 198932 44336
rect 198880 44272 198932 44278
rect 198328 41882 198380 41888
rect 196316 41830 198328 41836
rect 196316 41824 198380 41830
rect 196316 41820 198368 41824
rect 198892 41822 198920 44272
rect 199536 41822 199564 44476
rect 200720 44466 200772 44472
rect 200720 44408 200772 44414
rect 242764 44466 242816 44472
rect 242764 44408 242816 44414
rect 199984 41882 200036 41888
rect 200732 41836 200760 44408
rect 201364 44398 201416 44404
rect 201364 44340 201416 44346
rect 201376 44268 201404 44340
rect 201364 44262 201416 44268
rect 201364 44204 201416 44210
rect 200036 41830 200760 41836
rect 199984 41824 200760 41830
rect 199996 41822 200760 41824
rect 201376 41822 201404 44204
rect 242776 42432 242804 44408
rect 244512 44398 244564 44404
rect 244512 44340 244564 44346
rect 296952 44398 297004 44404
rect 296952 44340 297004 44346
rect 299436 44398 299488 44404
rect 299436 44340 299488 44346
rect 242764 42426 242816 42432
rect 242764 42368 242816 42374
rect 190902 41814 191020 41820
rect 190902 41808 190968 41814
rect 192098 41814 192216 41820
rect 192098 41808 192164 41814
rect 190968 41756 191020 41762
rect 193386 41814 193504 41820
rect 193386 41808 193452 41814
rect 192164 41756 192216 41762
rect 193452 41756 193504 41762
rect 196304 41814 198368 41820
rect 196356 41808 198368 41814
rect 199996 41808 200746 41822
rect 196304 41756 196356 41762
rect 148922 40354 148978 40363
rect 148922 40289 148978 40298
rect 144967 40176 145008 40204
rect 140860 40114 140912 40120
rect 140564 40062 140860 40068
rect 140564 40056 140912 40062
rect 142936 40114 142988 40120
rect 142936 40056 142988 40062
rect 144416 40114 144468 40120
rect 144416 40056 144468 40062
rect 140564 40040 140900 40056
rect 140872 39986 140900 40040
rect 142948 39918 142976 40056
rect 144428 39918 144456 40056
rect 144967 39986 144995 40176
rect 242776 39712 242804 42368
rect 244524 39955 244552 44340
rect 247088 44330 247140 44336
rect 247088 44272 247140 44278
rect 244510 39946 244566 39955
rect 244510 39881 244566 39890
rect 241108 39706 241160 39712
rect 88846 39674 88902 39683
rect 241108 39648 241160 39654
rect 242764 39706 242816 39712
rect 242764 39648 242816 39654
rect 247100 39660 247128 44272
rect 295112 44194 295164 44200
rect 295112 44136 295164 44142
rect 251320 43242 251372 43248
rect 251320 43184 251372 43190
rect 251332 42432 251360 43184
rect 251320 42426 251372 42432
rect 251320 42368 251372 42374
rect 251332 39955 251360 42368
rect 253804 42358 253856 42364
rect 253804 42300 253856 42306
rect 251964 41610 252016 41616
rect 251964 41552 252016 41558
rect 251976 40091 252004 41552
rect 251962 40082 252018 40091
rect 251962 40017 252018 40026
rect 251318 39946 251374 39955
rect 251318 39881 251374 39890
rect 253816 39712 253844 42300
rect 295124 41836 295152 44136
rect 296964 41836 296992 44340
rect 297596 43242 297648 43248
rect 297596 43184 297648 43190
rect 297608 42432 297636 43184
rect 297596 42426 297648 42432
rect 297596 42368 297648 42374
rect 297608 41836 297636 42368
rect 299448 41836 299476 44340
rect 299632 42500 299660 44612
rect 303760 44534 303812 44540
rect 303760 44476 303812 44482
rect 303116 44194 303168 44200
rect 303116 44136 303168 44142
rect 299620 42494 299672 42500
rect 299620 42436 299672 42442
rect 300632 42426 300684 42432
rect 300632 42368 300684 42374
rect 300644 41836 300672 42368
rect 303128 41836 303156 44136
rect 303772 42296 303800 44476
rect 306244 44466 306296 44472
rect 306244 44408 306296 44414
rect 305600 44398 305652 44404
rect 305600 44340 305652 44346
rect 304404 44262 304456 44268
rect 304404 44204 304456 44210
rect 304416 42500 304444 44204
rect 304404 42494 304456 42500
rect 304404 42436 304456 42442
rect 303760 42290 303812 42296
rect 303760 42232 303812 42238
rect 303772 41836 303800 42232
rect 304416 41836 304444 42436
rect 305612 41836 305640 44340
rect 306152 41950 306204 41956
rect 306256 41938 306284 44408
rect 307452 44336 307480 44680
rect 308084 44602 308136 44608
rect 308084 44544 308136 44550
rect 307440 44330 307492 44336
rect 307440 44272 307492 44278
rect 306204 41910 306284 41938
rect 306152 41892 306204 41898
rect 306256 41836 306284 41910
rect 307452 41836 307480 44272
rect 308096 42296 308124 44544
rect 318124 44540 318152 44680
rect 318112 44534 318164 44540
rect 318112 44476 318164 44482
rect 331084 44534 331136 44540
rect 331084 44476 331136 44482
rect 309280 44466 309332 44472
rect 309280 44408 309332 44414
rect 308084 42290 308136 42296
rect 308084 42232 308136 42238
rect 308096 41836 308124 42232
rect 309292 41836 309320 44408
rect 331096 44336 331124 44476
rect 344804 44404 344832 44680
rect 344792 44398 344844 44404
rect 344792 44340 344844 44346
rect 344884 44398 344936 44404
rect 344884 44340 344936 44346
rect 331084 44330 331136 44336
rect 334764 44330 334816 44336
rect 331084 44272 331136 44278
rect 334762 44298 334764 44307
rect 344896 44307 344924 44340
rect 351796 44336 351824 44680
rect 358592 44602 358644 44608
rect 358592 44544 358644 44550
rect 352428 44466 352480 44472
rect 352428 44408 352480 44414
rect 355464 44466 355516 44472
rect 355464 44408 355516 44414
rect 351784 44330 351836 44336
rect 334816 44298 334818 44307
rect 344882 44298 344938 44307
rect 338364 44268 338576 44284
rect 334762 44233 334818 44242
rect 338352 44262 338588 44268
rect 338404 44256 338536 44262
rect 338352 44204 338404 44210
rect 351784 44272 351836 44278
rect 344882 44233 344938 44242
rect 338536 44204 338588 44210
rect 349944 44194 349996 44200
rect 349944 44136 349996 44142
rect 295124 41808 295170 41836
rect 296964 41820 297176 41836
rect 296964 41814 297188 41820
rect 296964 41808 297136 41814
rect 297608 41808 297654 41836
rect 299448 41808 299494 41836
rect 300644 41820 302144 41836
rect 300644 41814 302156 41820
rect 300644 41808 302104 41814
rect 297136 41756 297188 41762
rect 303128 41808 303174 41836
rect 303772 41808 303818 41836
rect 304416 41808 304462 41836
rect 304876 41820 305014 41836
rect 304864 41814 305014 41820
rect 302104 41756 302156 41762
rect 304916 41808 305014 41814
rect 305612 41808 305658 41836
rect 306256 41808 306302 41836
rect 307452 41808 307498 41836
rect 308096 41808 308142 41836
rect 308694 41808 309338 41836
rect 349956 41822 349984 44136
rect 351796 41822 351824 44272
rect 352440 41822 352468 44408
rect 354268 44330 354320 44336
rect 354268 44272 354320 44278
rect 354280 41822 354308 44272
rect 355476 41836 355504 44408
rect 358604 44200 358632 44544
rect 359248 44268 359276 44680
rect 413884 44670 413936 44676
rect 413884 44612 413936 44618
rect 376992 44602 377044 44608
rect 377176 44602 377228 44608
rect 377044 44550 377176 44556
rect 376992 44544 377228 44550
rect 362824 44534 362876 44540
rect 377004 44528 377216 44544
rect 413896 44540 413924 44612
rect 413884 44534 413936 44540
rect 362824 44476 362876 44482
rect 413884 44476 413936 44482
rect 414068 44534 414120 44540
rect 414068 44476 414120 44482
rect 361076 44466 361128 44472
rect 361076 44408 361128 44414
rect 360432 44330 360484 44336
rect 360432 44272 360484 44278
rect 359236 44262 359288 44268
rect 359236 44204 359288 44210
rect 357948 44194 358000 44200
rect 357948 44136 358000 44142
rect 358592 44194 358644 44200
rect 358592 44136 358644 44142
rect 355476 41822 356778 41836
rect 357960 41822 357988 44136
rect 358604 41822 358632 44136
rect 359248 41822 359276 44204
rect 355490 41808 356778 41822
rect 359814 41820 359920 41836
rect 360444 41822 360472 44272
rect 361088 41836 361116 44408
rect 362836 44404 362864 44476
rect 364112 44466 364164 44472
rect 364112 44408 364164 44414
rect 407260 44466 407312 44472
rect 407260 44408 407312 44414
rect 410296 44466 410348 44472
rect 410296 44408 410348 44414
rect 412964 44466 413016 44472
rect 412964 44408 413016 44414
rect 362272 44398 362324 44404
rect 362272 44340 362324 44346
rect 362824 44398 362876 44404
rect 362824 44340 362876 44346
rect 362916 44398 362968 44404
rect 362916 44340 362968 44346
rect 360996 41822 361116 41836
rect 362284 41822 362312 44340
rect 362928 44200 362956 44340
rect 362916 44194 362968 44200
rect 362916 44136 362968 44142
rect 362928 41822 362956 44136
rect 364124 41836 364152 44408
rect 406616 44330 406668 44336
rect 406616 44272 406668 44278
rect 404776 44194 404828 44200
rect 404776 44136 404828 44142
rect 404788 41836 404816 44136
rect 406628 41836 406656 44272
rect 407272 41836 407300 44408
rect 409192 41882 409244 41888
rect 363494 41822 364152 41836
rect 360996 41820 361102 41822
rect 359814 41814 359932 41820
rect 359814 41808 359880 41814
rect 304864 41756 304916 41762
rect 359880 41756 359932 41762
rect 360984 41814 361102 41820
rect 361036 41808 361102 41814
rect 363494 41808 364138 41822
rect 404770 41808 404816 41836
rect 406610 41808 406656 41836
rect 407254 41808 407300 41836
rect 409094 41830 409192 41836
rect 410308 41836 410336 44408
rect 412976 44268 413004 44408
rect 413424 44398 413476 44404
rect 413424 44340 413476 44346
rect 410940 44262 410992 44268
rect 410940 44204 410992 44210
rect 412964 44262 413016 44268
rect 412964 44204 413016 44210
rect 410952 41836 410980 44204
rect 412780 44194 412832 44200
rect 412780 44136 412832 44142
rect 412228 41882 412280 41888
rect 409094 41824 409244 41830
rect 409094 41808 409232 41824
rect 410290 41820 410428 41836
rect 410290 41814 410440 41820
rect 410290 41808 410388 41814
rect 360984 41756 361036 41762
rect 410934 41808 410980 41836
rect 411412 41820 411578 41836
rect 411400 41814 411578 41820
rect 410388 41756 410440 41762
rect 411452 41808 411578 41814
rect 412130 41830 412228 41836
rect 412792 41836 412820 44136
rect 413436 41836 413464 44340
rect 414080 41836 414108 44476
rect 417484 44268 417512 44748
rect 437724 44744 437752 44777
rect 437712 44738 437764 44744
rect 437712 44680 437764 44686
rect 441392 44738 441444 44744
rect 450682 44706 450738 44715
rect 441444 44686 441616 44692
rect 441392 44680 441616 44686
rect 441404 44676 441616 44680
rect 441404 44670 441628 44676
rect 441404 44664 441576 44670
rect 463470 44706 463526 44715
rect 450682 44641 450684 44650
rect 441576 44612 441628 44618
rect 450736 44641 450738 44650
rect 459516 44670 459568 44676
rect 450684 44612 450736 44618
rect 463470 44641 463526 44650
rect 459516 44612 459568 44618
rect 419036 44466 419088 44472
rect 419036 44408 419088 44414
rect 417748 44398 417800 44404
rect 417748 44340 417800 44346
rect 417104 44262 417156 44268
rect 417104 44204 417156 44210
rect 417472 44262 417524 44268
rect 417472 44204 417524 44210
rect 415080 41882 415132 41888
rect 412130 41824 412280 41830
rect 412130 41808 412268 41824
rect 412774 41808 412820 41836
rect 413418 41808 413464 41836
rect 414062 41808 414108 41836
rect 414448 41820 414614 41836
rect 417116 41836 417144 44204
rect 417760 41836 417788 44340
rect 419048 41836 419076 44408
rect 419588 44194 419640 44200
rect 419588 44136 419640 44142
rect 419600 41836 419628 44136
rect 415132 41830 415258 41836
rect 415080 41824 415258 41830
rect 414436 41814 414614 41820
rect 411400 41756 411452 41762
rect 414488 41808 414614 41814
rect 415092 41808 415258 41824
rect 415736 41820 415902 41836
rect 415724 41814 415902 41820
rect 414436 41756 414488 41762
rect 415776 41808 415902 41814
rect 417098 41808 417144 41836
rect 417742 41808 417788 41836
rect 418128 41820 418294 41836
rect 418116 41814 418294 41820
rect 415724 41756 415776 41762
rect 418168 41808 418294 41814
rect 418938 41820 419076 41836
rect 418938 41814 419088 41820
rect 418938 41808 419036 41814
rect 418116 41756 418168 41762
rect 419582 41808 419628 41836
rect 459528 41822 459556 44612
rect 463484 44608 463512 44641
rect 463472 44602 463524 44608
rect 463472 44544 463524 44550
rect 465508 44472 465536 85548
rect 674808 83844 674836 86296
rect 675176 86292 675204 117016
rect 675164 86286 675216 86292
rect 675164 86228 675216 86234
rect 675268 86172 675296 117152
rect 675544 86360 675572 117168
rect 675532 86354 675584 86360
rect 675532 86296 675584 86302
rect 675084 86144 675296 86172
rect 674796 83838 674848 83844
rect 674796 83780 674848 83786
rect 674808 73712 674836 83780
rect 675084 83572 675112 86144
rect 675164 86082 675216 86088
rect 675164 86024 675216 86030
rect 675072 83566 675124 83572
rect 675072 83508 675124 83514
rect 675176 82636 675204 86024
rect 675256 83838 675308 83844
rect 675256 83780 675308 83786
rect 675268 83680 675296 83780
rect 675256 83566 675308 83572
rect 675256 83508 675308 83514
rect 675084 82608 675204 82636
rect 674888 82546 674940 82552
rect 674888 82488 674940 82494
rect 674900 74052 674928 82488
rect 675084 82364 675112 82608
rect 675268 82552 675296 83508
rect 675256 82546 675308 82552
rect 675256 82488 675308 82494
rect 675084 82336 675204 82364
rect 675176 78828 675204 82336
rect 675084 78800 675204 78828
rect 674888 74046 674940 74052
rect 674888 73988 674940 73994
rect 675084 73932 675112 78800
rect 674900 73904 675112 73932
rect 675176 78698 675282 78726
rect 674796 73706 674848 73712
rect 674796 73648 674848 73654
rect 674900 72148 674928 73904
rect 674980 73842 675032 73848
rect 675176 73796 675204 78698
rect 674980 73784 675032 73790
rect 674888 72142 674940 72148
rect 674888 72084 674940 72090
rect 674900 70260 674928 72084
rect 674992 70396 675020 73784
rect 675084 73768 675204 73796
rect 675084 73388 675112 73768
rect 675164 73706 675216 73712
rect 675164 73648 675216 73654
rect 675176 73576 675204 73648
rect 675164 73570 675216 73576
rect 675164 73512 675216 73518
rect 675084 73360 675204 73388
rect 675072 73298 675124 73304
rect 675072 73240 675124 73246
rect 675084 70532 675112 73240
rect 675176 70722 675204 73360
rect 675268 72148 675296 72558
rect 675256 72142 675308 72148
rect 675256 72084 675308 72090
rect 675176 70694 675282 70722
rect 675084 70504 675388 70532
rect 674992 70368 675296 70396
rect 674900 70232 675204 70260
rect 675176 45968 675204 70232
rect 670288 45962 670340 45968
rect 670288 45904 670340 45910
rect 675164 45962 675216 45968
rect 675164 45904 675216 45910
rect 515084 45146 515136 45152
rect 515084 45088 515136 45094
rect 516188 45146 516240 45152
rect 516188 45088 516240 45094
rect 527320 45146 527372 45152
rect 527320 45088 527372 45094
rect 540842 45114 540898 45123
rect 515096 44812 515124 45088
rect 515084 44806 515136 44812
rect 515084 44748 515136 44754
rect 467520 44670 467572 44676
rect 467520 44612 467572 44618
rect 471844 44670 471896 44676
rect 471844 44612 471896 44618
rect 473776 44670 473828 44676
rect 473776 44612 473828 44618
rect 473868 44670 473920 44676
rect 473868 44612 473920 44618
rect 480124 44670 480176 44676
rect 480124 44612 480176 44618
rect 489232 44670 489284 44676
rect 489232 44612 489284 44618
rect 462000 44466 462052 44472
rect 462000 44408 462052 44414
rect 465036 44466 465088 44472
rect 465036 44408 465088 44414
rect 465496 44466 465548 44472
rect 465496 44408 465548 44414
rect 461356 44330 461408 44336
rect 461356 44272 461408 44278
rect 461368 41822 461396 44272
rect 462012 41822 462040 44408
rect 464024 41882 464076 41888
rect 463866 41830 464024 41836
rect 465048 41859 465076 44408
rect 465680 44194 465732 44200
rect 465680 44136 465732 44142
rect 463866 41824 464076 41830
rect 465034 41850 465090 41859
rect 463866 41808 464064 41824
rect 465692 41822 465720 44136
rect 467060 41882 467112 41888
rect 466322 41850 466378 41859
rect 465034 41785 465090 41794
rect 466888 41842 467060 41870
rect 466888 41822 466916 41842
rect 467060 41824 467112 41830
rect 467532 41822 467560 44612
rect 468806 44570 468862 44579
rect 468806 44505 468808 44514
rect 468860 44505 468862 44514
rect 468808 44476 468860 44482
rect 468164 44398 468216 44404
rect 468164 44340 468216 44346
rect 468176 42296 468204 44340
rect 468164 42290 468216 42296
rect 468164 42232 468216 42238
rect 468176 41822 468204 42232
rect 468820 41822 468848 44476
rect 469266 41986 469322 41995
rect 469266 41921 469322 41930
rect 470554 41986 470610 41995
rect 470554 41921 470610 41930
rect 469280 41836 469308 41921
rect 469912 41882 469964 41888
rect 469280 41808 469386 41836
rect 469964 41842 470044 41870
rect 469912 41824 469964 41830
rect 470016 41822 470044 41842
rect 470568 41836 470596 41921
rect 470568 41808 470674 41836
rect 471856 41822 471884 44612
rect 473592 44466 473644 44472
rect 473592 44408 473644 44414
rect 472488 44398 472540 44404
rect 472488 44340 472540 44346
rect 472500 42296 472528 44340
rect 472488 42290 472540 42296
rect 472488 42232 472540 42238
rect 472500 41822 472528 42232
rect 473604 41995 473632 44408
rect 473788 44268 473816 44612
rect 473880 44336 473908 44612
rect 480136 44579 480164 44612
rect 489244 44579 489272 44612
rect 476350 44570 476406 44579
rect 476350 44505 476352 44514
rect 476404 44505 476406 44514
rect 480122 44570 480178 44579
rect 480122 44505 480178 44514
rect 489230 44570 489286 44579
rect 489230 44505 489286 44514
rect 515084 44534 515136 44540
rect 476352 44476 476404 44482
rect 515084 44476 515136 44482
rect 473868 44330 473920 44336
rect 473868 44272 473920 44278
rect 473776 44262 473828 44268
rect 473776 44204 473828 44210
rect 474328 44194 474380 44200
rect 474328 44136 474380 44142
rect 514348 44194 514400 44200
rect 514348 44136 514400 44142
rect 472946 41986 473002 41995
rect 472946 41921 473002 41930
rect 473590 41986 473646 41995
rect 473590 41921 473646 41930
rect 472960 41836 472988 41921
rect 473604 41836 473632 41921
rect 472960 41808 473066 41836
rect 473604 41808 473710 41836
rect 474340 41822 474368 44136
rect 514360 41822 514388 44136
rect 515096 43588 515124 44476
rect 515084 43582 515136 43588
rect 515084 43524 515136 43530
rect 516200 41822 516228 45088
rect 516832 44466 516884 44472
rect 516832 44408 516884 44414
rect 519868 44466 519920 44472
rect 519868 44408 519920 44414
rect 516844 41822 516872 44408
rect 518672 44330 518724 44336
rect 518672 44272 518724 44278
rect 518684 41822 518712 44272
rect 519880 41836 519908 44408
rect 522996 44398 523048 44404
rect 522996 44340 523048 44346
rect 523008 44200 523036 44340
rect 524836 44330 524888 44336
rect 524836 44272 524888 44278
rect 525940 44330 525992 44336
rect 525940 44272 525992 44278
rect 522352 44194 522404 44200
rect 522352 44136 522404 44142
rect 522996 44194 523048 44200
rect 522996 44136 523048 44142
rect 519960 41882 520012 41888
rect 519880 41830 519960 41836
rect 521248 41882 521300 41888
rect 519880 41824 520012 41830
rect 521182 41830 521248 41836
rect 521182 41824 521300 41830
rect 519880 41822 520000 41824
rect 519894 41808 520000 41822
rect 521182 41808 521288 41824
rect 522364 41822 522392 44136
rect 523008 41822 523036 44136
rect 523640 43582 523692 43588
rect 523640 43524 523692 43530
rect 523652 41822 523680 43524
rect 524284 41882 524336 41888
rect 524218 41830 524284 41836
rect 524218 41824 524336 41830
rect 524218 41808 524324 41824
rect 524848 41822 524876 44272
rect 525952 43588 525980 44272
rect 526676 44262 526728 44268
rect 526676 44204 526728 44210
rect 525940 43582 525992 43588
rect 525940 43524 525992 43530
rect 525572 41882 525624 41888
rect 525506 41830 525572 41836
rect 525506 41824 525624 41830
rect 525506 41808 525612 41824
rect 526688 41822 526716 44204
rect 527332 44200 527360 45088
rect 540842 45049 540844 45058
rect 540896 45049 540898 45058
rect 553630 45114 553686 45123
rect 553630 45049 553686 45058
rect 540844 45020 540896 45026
rect 553644 45016 553672 45049
rect 553632 45010 553684 45016
rect 553632 44952 553684 44958
rect 570204 44812 570324 44828
rect 595964 44812 596084 44828
rect 621724 44812 621844 44828
rect 647484 44812 647604 44828
rect 670300 44812 670328 45904
rect 570192 44806 570336 44812
rect 570244 44800 570284 44806
rect 570192 44748 570244 44754
rect 570284 44748 570336 44754
rect 592272 44806 592324 44812
rect 592272 44748 592324 44754
rect 595952 44806 596096 44812
rect 596004 44800 596044 44806
rect 595952 44748 596004 44754
rect 596044 44748 596096 44754
rect 618032 44806 618084 44812
rect 618032 44748 618084 44754
rect 621712 44806 621856 44812
rect 621764 44800 621804 44806
rect 621712 44748 621764 44754
rect 621804 44748 621856 44754
rect 643792 44806 643844 44812
rect 643792 44748 643844 44754
rect 647472 44806 647616 44812
rect 647524 44800 647564 44806
rect 647472 44748 647524 44754
rect 647564 44748 647616 44754
rect 669552 44806 669604 44812
rect 669552 44748 669604 44754
rect 670288 44806 670340 44812
rect 670288 44748 670340 44754
rect 579484 44738 579536 44744
rect 579482 44706 579484 44715
rect 592284 44715 592312 44748
rect 605244 44738 605296 44744
rect 579536 44706 579538 44715
rect 579482 44641 579538 44650
rect 592270 44706 592326 44715
rect 592270 44641 592326 44650
rect 605242 44706 605244 44715
rect 618044 44715 618072 44748
rect 631004 44738 631056 44744
rect 605296 44706 605298 44715
rect 605242 44641 605298 44650
rect 618030 44706 618086 44715
rect 618030 44641 618086 44650
rect 631002 44706 631004 44715
rect 643804 44715 643832 44748
rect 656764 44738 656816 44744
rect 631056 44706 631058 44715
rect 631002 44641 631058 44650
rect 643790 44706 643846 44715
rect 643790 44641 643846 44650
rect 656762 44706 656764 44715
rect 669564 44715 669592 44748
rect 656816 44706 656818 44715
rect 656762 44641 656818 44650
rect 669550 44706 669606 44715
rect 669550 44641 669606 44650
rect 568996 44330 569048 44336
rect 568996 44272 569048 44278
rect 527320 44194 527372 44200
rect 527320 44136 527372 44142
rect 527332 41822 527360 44136
rect 527780 41882 527832 41888
rect 527832 41830 528542 41836
rect 527780 41824 528542 41830
rect 527792 41808 528542 41824
rect 466322 41785 466378 41794
rect 419036 41756 419088 41762
rect 286924 41610 286976 41616
rect 286924 41552 286976 41558
rect 286936 41412 286964 41552
rect 286924 41406 286976 41412
rect 286924 41348 286976 41354
rect 251964 39706 252016 39712
rect 88846 39609 88902 39618
rect 241120 39374 241148 39648
rect 247100 39632 247220 39660
rect 251964 39648 252016 39654
rect 253804 39706 253856 39712
rect 253804 39648 253856 39654
rect 247192 39569 247220 39632
rect 251976 39374 252004 39648
rect 569008 39646 569036 44272
rect 630268 44262 630320 44268
rect 630268 44204 630320 44210
rect 579484 43242 579536 43248
rect 579484 43184 579536 43190
rect 579496 42364 579524 43184
rect 569088 42358 569140 42364
rect 569088 42300 569140 42306
rect 579484 42358 579536 42364
rect 579484 42300 579536 42306
rect 569100 40227 569128 42300
rect 569086 40218 569142 40227
rect 569086 40153 569142 40162
rect 579496 39660 579524 42300
rect 630280 40227 630308 44204
rect 675268 43248 675296 70368
rect 675360 45152 675388 70504
rect 675348 45146 675400 45152
rect 675348 45088 675400 45094
rect 675256 43242 675308 43248
rect 675256 43184 675308 43190
rect 630266 40218 630322 40227
rect 630266 40153 630322 40162
rect 622630 39810 622686 39819
rect 622630 39745 622686 39754
rect 579050 39632 579524 39660
rect 622644 39660 622672 39745
rect 622644 39632 622842 39660
<< via2 >>
rect 352150 997602 352206 997658
rect 353162 997466 353218 997522
rect 362178 997466 362234 997522
rect 364386 997466 364442 997522
rect 579390 997466 579446 997522
rect 581506 997466 581562 997522
rect 39718 917090 39774 917146
rect 39718 915186 39774 915242
rect 39350 903626 39406 903682
rect 39902 875746 39958 875802
rect 42294 914642 42350 914698
rect 42294 910834 42350 910890
rect 42202 875746 42258 875802
rect 39994 822706 40050 822762
rect 39994 822298 40050 822354
rect 41650 793602 41706 793658
rect 41926 789658 41982 789714
rect 42110 789522 42166 789578
rect 41650 785986 41706 786042
rect 41650 780682 41706 780738
rect 41558 780496 41614 780552
rect 41650 777962 41706 778018
rect 42110 743554 42166 743610
rect 41558 736540 41614 736596
rect 41558 735896 41614 735952
rect 42110 735896 42166 735952
rect 41650 733354 41706 733410
rect 41742 704794 41798 704850
rect 41650 704658 41706 704714
rect 41558 704468 41614 704524
rect 41558 696464 41614 696520
rect 42110 696362 42166 696418
rect 41650 692690 41706 692746
rect 42110 688882 42166 688938
rect 41926 682626 41982 682682
rect 41834 660050 41890 660106
rect 41558 659868 41614 659924
rect 41558 658010 41614 658066
rect 42018 653270 42074 653306
rect 42018 653250 42020 653270
rect 42020 653250 42072 653270
rect 42072 653250 42074 653270
rect 41650 652298 41706 652354
rect 42110 647946 42166 648002
rect 42110 646994 42166 647050
rect 41558 615714 41614 615770
rect 41742 644138 41798 644194
rect 41650 615442 41706 615498
rect 41558 615268 41614 615324
rect 41650 613810 41706 613866
rect 41558 607282 41614 607338
rect 41558 602930 41614 602986
rect 41558 602296 41614 602352
rect 41650 599802 41706 599858
rect 42110 599666 42166 599722
rect 41834 570970 41890 571026
rect 41650 570426 41706 570482
rect 41558 569028 41614 569084
rect 41650 563354 41706 563410
rect 41650 558050 41706 558106
rect 41558 557914 41614 557970
rect 42110 557914 42166 557970
rect 42110 557778 42166 557834
rect 41834 555330 41890 555386
rect 41926 555194 41982 555250
rect 42110 526498 42166 526554
rect 41558 526268 41614 526324
rect 42110 519018 42166 519074
rect 41558 518264 41614 518320
rect 41558 513940 41614 513996
rect 41558 513306 41614 513362
rect 41650 510722 41706 510778
rect 41926 510722 41982 510778
rect 39718 437826 39774 437882
rect 39534 423682 39590 423738
rect 39718 423682 39774 423738
rect 42110 381930 42166 381986
rect 41558 381696 41614 381752
rect 41742 379210 41798 379266
rect 41650 305770 41706 305826
rect 42110 297610 42166 297666
rect 41558 293340 41614 293396
rect 41558 292714 41614 292770
rect 41742 290130 41798 290186
rect 41650 287138 41706 287194
rect 102922 993542 102978 993578
rect 102922 993522 102924 993542
rect 102924 993522 102976 993542
rect 102976 993522 102978 993542
rect 115710 993522 115766 993578
rect 261162 993542 261218 993578
rect 261162 993522 261164 993542
rect 261164 993522 261216 993542
rect 261216 993522 261218 993542
rect 273950 993422 273952 993442
rect 273952 993422 274004 993442
rect 274004 993422 274006 993442
rect 273950 993386 274006 993422
rect 321882 993150 321884 993170
rect 321884 993150 321936 993170
rect 321936 993150 321938 993170
rect 321882 993114 321938 993150
rect 334670 993114 334726 993170
rect 347642 993150 347644 993170
rect 347644 993150 347696 993170
rect 347696 993150 347698 993170
rect 347642 993114 347698 993150
rect 360430 993114 360486 993170
rect 573962 997330 574018 997386
rect 406614 995426 406670 995482
rect 408822 995426 408878 995482
rect 413146 995426 413202 995482
rect 421150 995426 421206 995482
rect 373402 993150 373404 993170
rect 373404 993150 373456 993170
rect 373456 993150 373458 993170
rect 373402 993114 373458 993150
rect 386190 993114 386246 993170
rect 43030 879418 43086 879474
rect 42478 830050 42534 830106
rect 42386 822298 42442 822354
rect 42570 682626 42626 682682
rect 42662 658010 42718 658066
rect 42754 602930 42810 602986
rect 42478 476450 42534 476506
rect 42478 474818 42534 474874
rect 42386 472914 42442 472970
rect 675070 962786 675126 962842
rect 675254 962786 675310 962842
rect 675070 910970 675126 911026
rect 675070 905258 675126 905314
rect 677738 915594 677794 915650
rect 674978 822434 675034 822490
rect 674886 817674 674942 817730
rect 674886 813322 674942 813378
rect 674426 783810 674482 783866
rect 674886 783810 674942 783866
rect 674702 745186 674758 745242
rect 674886 745186 674942 745242
rect 674426 732266 674482 732322
rect 677278 822434 677334 822490
rect 675438 745186 675494 745242
rect 675714 745186 675770 745242
rect 675438 744370 675494 744426
rect 674886 732266 674942 732322
rect 675254 731994 675310 732050
rect 675254 721114 675310 721170
rect 675530 719482 675586 719538
rect 675438 719210 675494 719266
rect 674610 685346 674666 685402
rect 674426 592186 674482 592242
rect 674886 498638 674942 498674
rect 674886 498618 674888 498638
rect 674888 498618 674940 498638
rect 674940 498618 674942 498638
rect 674794 495218 674850 495274
rect 674610 493178 674666 493234
rect 42294 431298 42350 431354
rect 42294 292714 42350 292770
rect 41558 248106 41614 248162
rect 41742 245522 41798 245578
rect 41650 216690 41706 216746
rect 42110 215058 42166 215114
rect 41650 214106 41706 214162
rect 42110 209618 42166 209674
rect 41650 209210 41706 209266
rect 41558 204140 41614 204196
rect 41650 200914 41706 200970
rect 42110 172218 42166 172274
rect 41558 170228 41614 170284
rect 42294 248106 42350 248162
rect 42662 170178 42718 170234
rect 42202 120402 42258 120458
rect 42202 112922 42258 112978
rect 43030 112922 43086 112978
rect 42294 76882 42350 76938
rect 674978 493178 675034 493234
rect 675714 688882 675770 688938
rect 675254 685408 675310 685464
rect 675622 642098 675678 642154
rect 675346 641962 675402 642018
rect 675254 638834 675310 638890
rect 675254 628320 675310 628376
rect 675162 626322 675218 626378
rect 675530 626322 675586 626378
rect 675254 592186 675310 592242
rect 675162 583346 675218 583402
rect 675254 581714 675310 581770
rect 675346 579674 675402 579730
rect 677462 573146 677518 573202
rect 677738 550026 677794 550082
rect 675070 449658 675126 449714
rect 674978 428850 675034 428906
rect 674886 425062 674942 425098
rect 674886 425042 674888 425062
rect 674888 425042 674940 425062
rect 674940 425042 674942 425062
rect 674794 406546 674850 406602
rect 675070 401650 675126 401706
rect 677922 459858 677978 459914
rect 677738 452106 677794 452162
rect 677462 406546 677518 406602
rect 675162 356942 675164 356962
rect 675164 356942 675216 356962
rect 675216 356942 675218 356962
rect 675162 356906 675218 356942
rect 674978 356634 675034 356690
rect 674886 350106 674942 350162
rect 675254 350106 675310 350162
rect 675346 318962 675402 319018
rect 675254 316452 675310 316508
rect 675530 271090 675586 271146
rect 674886 212338 674942 212394
rect 675254 218458 675310 218514
rect 675254 218322 675310 218378
rect 675254 212338 675310 212394
rect 675254 189490 675310 189546
rect 675622 189354 675678 189410
rect 675254 130252 675310 130308
rect 675070 119722 675126 119778
rect 43950 76882 44006 76938
rect 90870 40162 90926 40218
rect 134110 40182 134166 40218
rect 134110 40162 134112 40182
rect 134112 40162 134164 40182
rect 134164 40162 134166 40182
rect 142942 40162 142998 40218
rect 143402 40182 143458 40218
rect 143402 40162 143404 40182
rect 143404 40162 143456 40182
rect 143456 40162 143458 40182
rect 218842 44806 218898 44842
rect 218842 44786 218844 44806
rect 218844 44786 218896 44806
rect 218896 44786 218898 44806
rect 231630 44786 231686 44842
rect 244602 44806 244658 44842
rect 244602 44786 244604 44806
rect 244604 44786 244656 44806
rect 244656 44786 244658 44806
rect 257390 44786 257446 44842
rect 424922 44806 424978 44842
rect 424922 44786 424924 44806
rect 424924 44786 424976 44806
rect 424976 44786 424978 44806
rect 437710 44786 437766 44842
rect 148922 40298 148978 40354
rect 244510 39890 244566 39946
rect 88846 39618 88902 39674
rect 251962 40026 252018 40082
rect 251318 39890 251374 39946
rect 334762 44278 334764 44298
rect 334764 44278 334816 44298
rect 334816 44278 334818 44298
rect 334762 44242 334818 44278
rect 344882 44242 344938 44298
rect 450682 44670 450738 44706
rect 450682 44650 450684 44670
rect 450684 44650 450736 44670
rect 450736 44650 450738 44670
rect 463470 44650 463526 44706
rect 465034 41794 465090 41850
rect 466322 41794 466378 41850
rect 468806 44534 468862 44570
rect 468806 44514 468808 44534
rect 468808 44514 468860 44534
rect 468860 44514 468862 44534
rect 469266 41930 469322 41986
rect 470554 41930 470610 41986
rect 476350 44534 476406 44570
rect 476350 44514 476352 44534
rect 476352 44514 476404 44534
rect 476404 44514 476406 44534
rect 480122 44514 480178 44570
rect 489230 44514 489286 44570
rect 472946 41930 473002 41986
rect 473590 41930 473646 41986
rect 540842 45078 540898 45114
rect 540842 45058 540844 45078
rect 540844 45058 540896 45078
rect 540896 45058 540898 45078
rect 553630 45058 553686 45114
rect 579482 44686 579484 44706
rect 579484 44686 579536 44706
rect 579536 44686 579538 44706
rect 579482 44650 579538 44686
rect 592270 44650 592326 44706
rect 605242 44686 605244 44706
rect 605244 44686 605296 44706
rect 605296 44686 605298 44706
rect 605242 44650 605298 44686
rect 618030 44650 618086 44706
rect 631002 44686 631004 44706
rect 631004 44686 631056 44706
rect 631056 44686 631058 44706
rect 631002 44650 631058 44686
rect 643790 44650 643846 44706
rect 656762 44686 656764 44706
rect 656764 44686 656816 44706
rect 656816 44686 656818 44706
rect 656762 44650 656818 44686
rect 669550 44650 669606 44706
rect 569086 40162 569142 40218
rect 630266 40162 630322 40218
rect 622630 39754 622686 39810
<< metal3 >>
rect 352145 997660 352211 997663
rect 352145 997658 352316 997660
rect 352145 997602 352150 997658
rect 352206 997630 352316 997658
rect 352206 997602 352346 997630
rect 352145 997600 352346 997602
rect 352145 997597 352211 997600
rect 352286 997524 352346 997600
rect 353157 997524 353223 997527
rect 352286 997522 353223 997524
rect 352286 997466 353162 997522
rect 353218 997466 353223 997522
rect 352286 997464 353223 997466
rect 353157 997461 353223 997464
rect 362173 997524 362239 997527
rect 364381 997524 364447 997527
rect 362173 997522 364447 997524
rect 362173 997466 362178 997522
rect 362234 997466 364386 997522
rect 364442 997466 364447 997522
rect 362173 997464 364447 997466
rect 362173 997461 362239 997464
rect 364381 997461 364447 997464
rect 569406 997388 569466 997630
rect 573957 997388 574023 997391
rect 574558 997388 574618 997630
rect 579385 997524 579451 997527
rect 581501 997524 581567 997527
rect 579385 997522 581567 997524
rect 579385 997466 579390 997522
rect 579446 997466 581506 997522
rect 581562 997466 581567 997522
rect 579385 997464 581567 997466
rect 579385 997461 579451 997464
rect 581501 997461 581567 997464
rect 569406 997386 574618 997388
rect 569406 997330 573962 997386
rect 574018 997330 574618 997386
rect 569406 997328 574618 997330
rect 573957 997325 574023 997328
rect 406609 995484 406675 995487
rect 408817 995484 408883 995487
rect 406609 995482 408883 995484
rect 406609 995426 406614 995482
rect 406670 995426 408822 995482
rect 408878 995426 408883 995482
rect 406609 995424 408883 995426
rect 406609 995421 406675 995424
rect 408817 995421 408883 995424
rect 413141 995484 413207 995487
rect 421145 995484 421211 995487
rect 413141 995482 421211 995484
rect 413141 995426 413146 995482
rect 413202 995426 421150 995482
rect 421206 995426 421211 995482
rect 413141 995424 421211 995426
rect 413141 995421 413207 995424
rect 421145 995421 421211 995424
rect 102917 993580 102983 993583
rect 115705 993580 115771 993583
rect 102917 993578 115771 993580
rect 102917 993522 102922 993578
rect 102978 993522 115710 993578
rect 115766 993522 115771 993578
rect 102917 993520 115771 993522
rect 102917 993517 102983 993520
rect 115705 993517 115771 993520
rect 261157 993580 261223 993583
rect 261157 993578 261266 993580
rect 261157 993522 261162 993578
rect 261218 993522 261266 993578
rect 261157 993517 261266 993522
rect 261206 993444 261266 993517
rect 273945 993444 274011 993447
rect 261206 993442 274011 993444
rect 261206 993386 273950 993442
rect 274006 993386 274011 993442
rect 261206 993384 274011 993386
rect 273945 993381 274011 993384
rect 321877 993172 321943 993175
rect 334665 993172 334731 993175
rect 321877 993170 334731 993172
rect 321877 993114 321882 993170
rect 321938 993114 334670 993170
rect 334726 993114 334731 993170
rect 321877 993112 334731 993114
rect 321877 993109 321943 993112
rect 334665 993109 334731 993112
rect 347637 993172 347703 993175
rect 360425 993172 360491 993175
rect 347637 993170 360491 993172
rect 347637 993114 347642 993170
rect 347698 993114 360430 993170
rect 360486 993114 360491 993170
rect 347637 993112 360491 993114
rect 347637 993109 347703 993112
rect 360425 993109 360491 993112
rect 373397 993172 373463 993175
rect 386185 993172 386251 993175
rect 373397 993170 386251 993172
rect 373397 993114 373402 993170
rect 373458 993114 386190 993170
rect 386246 993114 386251 993170
rect 373397 993112 386251 993114
rect 373397 993109 373463 993112
rect 386185 993109 386251 993112
rect 675065 962844 675131 962847
rect 675249 962844 675315 962847
rect 675065 962842 675315 962844
rect 675065 962786 675070 962842
rect 675126 962786 675254 962842
rect 675310 962786 675315 962842
rect 675065 962784 675315 962786
rect 675065 962781 675131 962784
rect 675249 962781 675315 962784
rect 39713 917148 39779 917151
rect 39332 917146 39779 917148
rect 39332 917090 39718 917146
rect 39774 917090 39779 917146
rect 39332 917088 39779 917090
rect 39713 917085 39779 917088
rect 677406 915590 677412 915654
rect 677476 915652 677482 915654
rect 677733 915652 677799 915655
rect 677476 915650 677799 915652
rect 677476 915594 677738 915650
rect 677794 915594 677799 915650
rect 677476 915592 677799 915594
rect 677476 915590 677482 915592
rect 677733 915589 677799 915592
rect 39713 915244 39779 915247
rect 39302 915242 39779 915244
rect 39302 915186 39718 915242
rect 39774 915186 39779 915242
rect 39302 915184 39779 915186
rect 39302 914700 39362 915184
rect 39713 915181 39779 915184
rect 42289 914700 42355 914703
rect 39302 914698 42355 914700
rect 39302 914670 42294 914698
rect 39332 914642 42294 914670
rect 42350 914642 42355 914698
rect 39332 914640 42355 914642
rect 42289 914637 42355 914640
rect 677598 912328 677996 912388
rect 677598 911844 677658 912328
rect 677598 911784 678026 911844
rect 675065 911028 675131 911031
rect 677966 911028 678026 911784
rect 675065 911026 678026 911028
rect 675065 910970 675070 911026
rect 675126 910970 678026 911026
rect 675065 910968 678026 910970
rect 675065 910965 675131 910968
rect 42289 910892 42355 910895
rect 39302 910890 42355 910892
rect 39302 910834 42294 910890
rect 42350 910834 42355 910890
rect 677966 910862 678026 910968
rect 39302 910832 42355 910834
rect 39302 909502 39362 910832
rect 42289 910829 42355 910832
rect 675065 905316 675131 905319
rect 675065 905314 678026 905316
rect 675065 905258 675070 905314
rect 675126 905258 678026 905314
rect 675065 905256 678026 905258
rect 675065 905253 675131 905256
rect 677966 904742 678026 905256
rect 39345 903684 39411 903687
rect 39846 903684 39852 903686
rect 39345 903682 39852 903684
rect 39345 903626 39350 903682
rect 39406 903626 39852 903682
rect 39345 903624 39852 903626
rect 39345 903621 39411 903624
rect 39846 903622 39852 903624
rect 39916 903622 39922 903686
rect 43025 879476 43091 879479
rect 39700 879474 43091 879476
rect 39700 879446 43030 879474
rect 39670 879418 43030 879446
rect 43086 879418 43091 879474
rect 39670 879416 43091 879418
rect 39670 875804 39730 879416
rect 43025 879413 43091 879416
rect 39897 875804 39963 875807
rect 42197 875804 42263 875807
rect 39670 875802 42263 875804
rect 39670 875746 39902 875802
rect 39958 875746 42202 875802
rect 42258 875746 42263 875802
rect 39670 875744 42263 875746
rect 39897 875741 39963 875744
rect 42197 875741 42263 875744
rect 42473 830108 42539 830111
rect 39516 830106 42539 830108
rect 39516 830050 42478 830106
rect 42534 830050 42539 830106
rect 39516 830048 42539 830050
rect 42473 830045 42539 830048
rect 39989 822764 40055 822767
rect 39486 822762 40055 822764
rect 39486 822706 39994 822762
rect 40050 822706 40055 822762
rect 39486 822704 40055 822706
rect 39486 822598 39546 822704
rect 39989 822701 40055 822704
rect 674973 822492 675039 822495
rect 677273 822492 677339 822495
rect 674973 822490 677339 822492
rect 674973 822434 674978 822490
rect 675034 822434 677278 822490
rect 677334 822434 677339 822490
rect 674973 822432 677339 822434
rect 674973 822429 675039 822432
rect 677273 822429 677339 822432
rect 39989 822356 40055 822359
rect 42381 822356 42447 822359
rect 39989 822354 42447 822356
rect 39989 822298 39994 822354
rect 40050 822298 42386 822354
rect 42442 822298 42447 822354
rect 39989 822296 42447 822298
rect 39989 822293 40055 822296
rect 42381 822293 42447 822296
rect 674881 817732 674947 817735
rect 674881 817730 677628 817732
rect 674881 817674 674886 817730
rect 674942 817674 677628 817730
rect 674881 817672 677628 817674
rect 674881 817669 674947 817672
rect 674881 813380 674947 813383
rect 674881 813378 677658 813380
rect 674881 813322 674886 813378
rect 674942 813322 677658 813378
rect 674881 813320 677658 813322
rect 674881 813317 674947 813320
rect 677598 812670 677658 813320
rect 41645 793660 41711 793663
rect 41870 793660 41876 793662
rect 41645 793658 41876 793660
rect 41645 793602 41650 793658
rect 41706 793602 41876 793658
rect 41645 793600 41876 793602
rect 41645 793597 41711 793600
rect 41870 793598 41876 793600
rect 41940 793598 41946 793662
rect 41921 789718 41987 789719
rect 41870 789716 41876 789718
rect 41830 789656 41876 789716
rect 41940 789714 41987 789718
rect 41982 789658 41987 789714
rect 41870 789654 41876 789656
rect 41940 789654 41987 789658
rect 41921 789653 41987 789654
rect 41686 789518 41692 789582
rect 41756 789580 41762 789582
rect 42105 789580 42171 789583
rect 41756 789578 42171 789580
rect 41756 789522 42110 789578
rect 42166 789522 42171 789578
rect 41756 789520 42171 789522
rect 41756 789518 41762 789520
rect 42105 789517 42171 789520
rect 41645 786046 41711 786047
rect 41645 786044 41692 786046
rect 41600 786042 41692 786044
rect 41600 785986 41650 786042
rect 41600 785984 41692 785986
rect 41645 785982 41692 785984
rect 41756 785982 41762 786046
rect 41645 785981 41711 785982
rect 674421 783868 674487 783871
rect 674881 783868 674947 783871
rect 674421 783866 674947 783868
rect 674421 783810 674426 783866
rect 674482 783810 674886 783866
rect 674942 783810 674947 783866
rect 674421 783808 674947 783810
rect 674421 783805 674487 783808
rect 674881 783805 674947 783808
rect 41645 780742 41711 780743
rect 41645 780740 41692 780742
rect 41600 780738 41692 780740
rect 41600 780682 41650 780738
rect 41600 780680 41692 780682
rect 41645 780678 41692 780680
rect 41756 780678 41762 780742
rect 41645 780677 41711 780678
rect 41134 780492 41140 780556
rect 41204 780554 41210 780556
rect 41553 780554 41619 780557
rect 41204 780552 41619 780554
rect 41204 780496 41558 780552
rect 41614 780496 41619 780552
rect 41204 780494 41619 780496
rect 41204 780492 41210 780494
rect 41553 780491 41619 780494
rect 41645 778022 41711 778023
rect 41645 778018 41692 778022
rect 41756 778020 41762 778022
rect 41645 777962 41650 778018
rect 41645 777958 41692 777962
rect 41756 777960 41802 778020
rect 41756 777958 41762 777960
rect 41645 777957 41711 777958
rect 674697 745244 674763 745247
rect 674881 745244 674947 745247
rect 674697 745242 674947 745244
rect 674697 745186 674702 745242
rect 674758 745186 674886 745242
rect 674942 745186 674947 745242
rect 674697 745184 674947 745186
rect 674697 745181 674763 745184
rect 674881 745181 674947 745184
rect 675433 745244 675499 745247
rect 675709 745244 675775 745247
rect 675433 745242 675775 745244
rect 675433 745186 675438 745242
rect 675494 745186 675714 745242
rect 675770 745186 675775 745242
rect 675433 745184 675775 745186
rect 675433 745181 675499 745184
rect 675709 745181 675775 745184
rect 675433 744428 675499 744431
rect 675566 744428 675572 744430
rect 675433 744426 675572 744428
rect 675433 744370 675438 744426
rect 675494 744370 675572 744426
rect 675433 744368 675572 744370
rect 675433 744365 675499 744368
rect 675566 744366 675572 744368
rect 675636 744366 675642 744430
rect 41870 743550 41876 743614
rect 41940 743612 41946 743614
rect 42105 743612 42171 743615
rect 41940 743610 42171 743612
rect 41940 743554 42110 743610
rect 42166 743554 42171 743610
rect 41940 743552 42171 743554
rect 41940 743550 41946 743552
rect 42105 743549 42171 743552
rect 41553 736598 41619 736601
rect 41870 736598 41876 736600
rect 41553 736596 41876 736598
rect 41553 736540 41558 736596
rect 41614 736540 41876 736596
rect 41553 736538 41876 736540
rect 41553 736535 41619 736538
rect 41870 736536 41876 736538
rect 41940 736536 41946 736600
rect 41134 735892 41140 735956
rect 41204 735954 41210 735956
rect 41553 735954 41619 735957
rect 42105 735954 42171 735957
rect 41204 735952 42171 735954
rect 41204 735896 41558 735952
rect 41614 735896 42110 735952
rect 42166 735896 42171 735952
rect 41204 735894 42171 735896
rect 41204 735892 41210 735894
rect 41553 735891 41619 735894
rect 42105 735891 42171 735894
rect 41645 733412 41711 733415
rect 41870 733412 41876 733414
rect 41645 733410 41876 733412
rect 41645 733354 41650 733410
rect 41706 733354 41876 733410
rect 41645 733352 41876 733354
rect 41645 733349 41711 733352
rect 41870 733350 41876 733352
rect 41940 733350 41946 733414
rect 674421 732324 674487 732327
rect 674881 732324 674947 732327
rect 674421 732322 674947 732324
rect 674421 732266 674426 732322
rect 674482 732266 674886 732322
rect 674942 732266 674947 732322
rect 674421 732264 674947 732266
rect 674421 732261 674487 732264
rect 674881 732261 674947 732264
rect 675249 732052 675315 732055
rect 675566 732052 675572 732054
rect 675249 732050 675572 732052
rect 675249 731994 675254 732050
rect 675310 731994 675572 732050
rect 675249 731992 675572 731994
rect 675249 731989 675315 731992
rect 675566 731990 675572 731992
rect 675636 731990 675642 732054
rect 675249 721172 675315 721175
rect 675382 721172 675388 721174
rect 675249 721170 675388 721172
rect 675249 721114 675254 721170
rect 675310 721114 675388 721170
rect 675249 721112 675388 721114
rect 675249 721109 675315 721112
rect 675382 721110 675388 721112
rect 675452 721110 675458 721174
rect 675525 719542 675591 719543
rect 675525 719540 675572 719542
rect 675480 719538 675572 719540
rect 675480 719482 675530 719538
rect 675480 719480 675572 719482
rect 675525 719478 675572 719480
rect 675636 719478 675642 719542
rect 675525 719477 675591 719478
rect 675433 719270 675499 719271
rect 675382 719268 675388 719270
rect 675342 719208 675388 719268
rect 675452 719266 675499 719270
rect 675494 719210 675499 719266
rect 675382 719206 675388 719208
rect 675452 719206 675499 719210
rect 675433 719205 675499 719206
rect 41737 704852 41803 704855
rect 41870 704852 41876 704854
rect 41737 704850 41876 704852
rect 41737 704794 41742 704850
rect 41798 704794 41876 704850
rect 41737 704792 41876 704794
rect 41737 704789 41803 704792
rect 41870 704790 41876 704792
rect 41940 704790 41946 704854
rect 41502 704654 41508 704718
rect 41572 704716 41578 704718
rect 41645 704716 41711 704719
rect 41572 704714 41711 704716
rect 41572 704658 41650 704714
rect 41706 704658 41711 704714
rect 41572 704656 41711 704658
rect 41572 704654 41578 704656
rect 41645 704653 41711 704656
rect 41553 704526 41619 704529
rect 41686 704526 41692 704528
rect 41553 704524 41692 704526
rect 41553 704468 41558 704524
rect 41614 704468 41692 704524
rect 41553 704466 41692 704468
rect 41553 704463 41619 704466
rect 41686 704464 41692 704466
rect 41756 704464 41762 704528
rect 41553 696522 41619 696525
rect 41686 696522 41692 696524
rect 41553 696520 41692 696522
rect 41553 696464 41558 696520
rect 41614 696464 41692 696520
rect 41553 696462 41692 696464
rect 41553 696459 41619 696462
rect 41686 696460 41692 696462
rect 41756 696460 41762 696524
rect 41870 696358 41876 696422
rect 41940 696420 41946 696422
rect 42105 696420 42171 696423
rect 41940 696418 42171 696420
rect 41940 696362 42110 696418
rect 42166 696362 42171 696418
rect 41940 696360 42171 696362
rect 41940 696358 41946 696360
rect 42105 696357 42171 696360
rect 41502 692686 41508 692750
rect 41572 692748 41578 692750
rect 41645 692748 41711 692751
rect 41572 692746 41711 692748
rect 41572 692690 41650 692746
rect 41706 692690 41711 692746
rect 41572 692688 41711 692690
rect 41572 692686 41578 692688
rect 41645 692685 41711 692688
rect 41502 688878 41508 688942
rect 41572 688940 41578 688942
rect 42105 688940 42171 688943
rect 41572 688938 42171 688940
rect 41572 688882 42110 688938
rect 42166 688882 42171 688938
rect 41572 688880 42171 688882
rect 41572 688878 41578 688880
rect 42105 688877 42171 688880
rect 675382 688878 675388 688942
rect 675452 688940 675458 688942
rect 675709 688940 675775 688943
rect 675452 688938 675775 688940
rect 675452 688882 675714 688938
rect 675770 688882 675775 688938
rect 675452 688880 675775 688882
rect 675452 688878 675458 688880
rect 675709 688877 675775 688880
rect 675249 685466 675315 685469
rect 675382 685466 675388 685468
rect 675249 685464 675388 685466
rect 675249 685408 675254 685464
rect 675310 685408 675388 685464
rect 674605 685404 674671 685407
rect 675249 685406 675388 685408
rect 675249 685404 675315 685406
rect 675382 685404 675388 685406
rect 675452 685404 675458 685468
rect 674605 685403 675315 685404
rect 674605 685402 675312 685403
rect 674605 685346 674610 685402
rect 674666 685346 675312 685402
rect 674605 685344 675312 685346
rect 674605 685341 674671 685344
rect 41921 682684 41987 682687
rect 42565 682684 42631 682687
rect 41921 682682 42631 682684
rect 41921 682626 41926 682682
rect 41982 682626 42570 682682
rect 42626 682626 42631 682682
rect 41921 682624 42631 682626
rect 41921 682621 41987 682624
rect 42565 682621 42631 682624
rect 41502 660046 41508 660110
rect 41572 660108 41578 660110
rect 41829 660108 41895 660111
rect 41572 660106 41895 660108
rect 41572 660050 41834 660106
rect 41890 660050 41895 660106
rect 41572 660048 41895 660050
rect 41572 660046 41578 660048
rect 41829 660045 41895 660048
rect 41553 659926 41619 659929
rect 41686 659926 41692 659928
rect 41553 659924 41692 659926
rect 41553 659868 41558 659924
rect 41614 659868 41692 659924
rect 41553 659866 41692 659868
rect 41553 659863 41619 659866
rect 41686 659864 41692 659866
rect 41756 659864 41762 659928
rect 41553 658070 41619 658071
rect 41502 658006 41508 658070
rect 41572 658068 41619 658070
rect 42657 658068 42723 658071
rect 41572 658066 42723 658068
rect 41614 658010 42662 658066
rect 42718 658010 42723 658066
rect 41572 658008 42723 658010
rect 41572 658006 41619 658008
rect 41553 658005 41619 658006
rect 42657 658005 42723 658008
rect 42013 653310 42079 653311
rect 42013 653306 42060 653310
rect 42124 653308 42130 653310
rect 42013 653250 42018 653306
rect 42013 653246 42060 653250
rect 42124 653248 42170 653308
rect 42124 653246 42130 653248
rect 42013 653245 42079 653246
rect 41645 652358 41711 652359
rect 41645 652356 41692 652358
rect 41600 652354 41692 652356
rect 41600 652298 41650 652354
rect 41600 652296 41692 652298
rect 41645 652294 41692 652296
rect 41756 652294 41762 652358
rect 41645 652293 41711 652294
rect 42105 648006 42171 648007
rect 42054 648004 42060 648006
rect 42014 647944 42060 648004
rect 42124 648002 42171 648006
rect 42166 647946 42171 648002
rect 42054 647942 42060 647944
rect 42124 647942 42171 647946
rect 42105 647941 42171 647942
rect 42105 647054 42171 647055
rect 42054 647052 42060 647054
rect 42014 646992 42060 647052
rect 42124 647050 42171 647054
rect 42166 646994 42171 647050
rect 42054 646990 42060 646992
rect 42124 646990 42171 646994
rect 42105 646989 42171 646990
rect 41737 644196 41803 644199
rect 42054 644196 42060 644198
rect 41737 644194 42060 644196
rect 41737 644138 41742 644194
rect 41798 644138 42060 644194
rect 41737 644136 42060 644138
rect 41737 644133 41803 644136
rect 42054 644134 42060 644136
rect 42124 644134 42130 644198
rect 675198 642094 675204 642158
rect 675268 642156 675274 642158
rect 675617 642156 675683 642159
rect 675268 642154 675683 642156
rect 675268 642098 675622 642154
rect 675678 642098 675683 642154
rect 675268 642096 675683 642098
rect 675268 642094 675274 642096
rect 675617 642093 675683 642096
rect 675014 641958 675020 642022
rect 675084 642020 675090 642022
rect 675341 642020 675407 642023
rect 675084 642018 675407 642020
rect 675084 641962 675346 642018
rect 675402 641962 675407 642018
rect 675084 641960 675407 641962
rect 675084 641958 675090 641960
rect 675341 641957 675407 641960
rect 675249 638894 675315 638895
rect 675198 638830 675204 638894
rect 675268 638892 675315 638894
rect 675268 638890 675360 638892
rect 675310 638834 675360 638890
rect 675268 638832 675360 638834
rect 675268 638830 675315 638832
rect 675249 638829 675315 638830
rect 675014 628316 675020 628380
rect 675084 628378 675090 628380
rect 675249 628378 675315 628381
rect 675382 628378 675388 628380
rect 675084 628376 675388 628378
rect 675084 628320 675254 628376
rect 675310 628320 675388 628376
rect 675084 628318 675388 628320
rect 675084 628316 675090 628318
rect 675249 628315 675315 628318
rect 675382 628316 675388 628318
rect 675452 628316 675458 628380
rect 675157 626382 675223 626383
rect 675157 626380 675204 626382
rect 675112 626378 675204 626380
rect 675112 626322 675162 626378
rect 675112 626320 675204 626322
rect 675157 626318 675204 626320
rect 675268 626318 675274 626382
rect 675382 626318 675388 626382
rect 675452 626380 675458 626382
rect 675525 626380 675591 626383
rect 675452 626378 675591 626380
rect 675452 626322 675530 626378
rect 675586 626322 675591 626378
rect 675452 626320 675591 626322
rect 675452 626318 675458 626320
rect 675157 626317 675223 626318
rect 675525 626317 675591 626320
rect 41553 615772 41619 615775
rect 41870 615772 41876 615774
rect 41553 615770 41876 615772
rect 41553 615714 41558 615770
rect 41614 615714 41876 615770
rect 41553 615712 41876 615714
rect 41553 615709 41619 615712
rect 41870 615710 41876 615712
rect 41940 615710 41946 615774
rect 41318 615438 41324 615502
rect 41388 615500 41394 615502
rect 41645 615500 41711 615503
rect 41388 615498 41711 615500
rect 41388 615442 41650 615498
rect 41706 615442 41711 615498
rect 41388 615440 41711 615442
rect 41388 615438 41394 615440
rect 41645 615437 41711 615440
rect 41553 615328 41619 615329
rect 41502 615326 41508 615328
rect 41462 615266 41508 615326
rect 41572 615324 41619 615328
rect 41614 615268 41619 615324
rect 41502 615264 41508 615266
rect 41572 615264 41619 615268
rect 41553 615263 41619 615264
rect 41645 613868 41711 613871
rect 41870 613868 41876 613870
rect 41645 613866 41876 613868
rect 41645 613810 41650 613866
rect 41706 613810 41876 613866
rect 41645 613808 41876 613810
rect 41645 613805 41711 613808
rect 41870 613806 41876 613808
rect 41940 613806 41946 613870
rect 41553 607342 41619 607343
rect 41502 607278 41508 607342
rect 41572 607340 41619 607342
rect 41572 607338 41664 607340
rect 41614 607282 41664 607338
rect 41572 607280 41664 607282
rect 41572 607278 41619 607280
rect 41553 607277 41619 607278
rect 41553 602988 41619 602991
rect 41686 602988 41692 602990
rect 41553 602986 41692 602988
rect 41553 602930 41558 602986
rect 41614 602930 41692 602986
rect 41553 602928 41692 602930
rect 41553 602925 41619 602928
rect 41686 602926 41692 602928
rect 41756 602988 41762 602990
rect 42749 602988 42815 602991
rect 41756 602986 42815 602988
rect 41756 602930 42754 602986
rect 42810 602930 42815 602986
rect 41756 602928 42815 602930
rect 41756 602926 41762 602928
rect 42749 602925 42815 602928
rect 41553 602356 41619 602357
rect 41502 602292 41508 602356
rect 41572 602354 41619 602356
rect 41572 602352 41664 602354
rect 41614 602296 41664 602352
rect 41572 602294 41664 602296
rect 41572 602292 41619 602294
rect 41553 602291 41619 602292
rect 41502 599798 41508 599862
rect 41572 599860 41578 599862
rect 41645 599860 41711 599863
rect 41572 599858 41711 599860
rect 41572 599802 41650 599858
rect 41706 599802 41711 599858
rect 41572 599800 41711 599802
rect 41572 599798 41578 599800
rect 41645 599797 41711 599800
rect 41686 599662 41692 599726
rect 41756 599724 41762 599726
rect 42105 599724 42171 599727
rect 41756 599722 42171 599724
rect 41756 599666 42110 599722
rect 42166 599666 42171 599722
rect 41756 599664 42171 599666
rect 41756 599662 41762 599664
rect 42105 599661 42171 599664
rect 674421 592244 674487 592247
rect 675249 592244 675315 592247
rect 674421 592242 675315 592244
rect 674421 592186 674426 592242
rect 674482 592186 675254 592242
rect 675310 592186 675315 592242
rect 674421 592184 675315 592186
rect 674421 592181 674487 592184
rect 675249 592181 675315 592184
rect 675157 583406 675223 583407
rect 675157 583402 675204 583406
rect 675268 583404 675274 583406
rect 675157 583346 675162 583402
rect 675157 583342 675204 583346
rect 675268 583344 675314 583404
rect 675268 583342 675274 583344
rect 675157 583341 675223 583342
rect 675249 581774 675315 581775
rect 675198 581710 675204 581774
rect 675268 581772 675315 581774
rect 675268 581770 675360 581772
rect 675310 581714 675360 581770
rect 675268 581712 675360 581714
rect 675268 581710 675315 581712
rect 675249 581709 675315 581710
rect 675198 579670 675204 579734
rect 675268 579732 675274 579734
rect 675341 579732 675407 579735
rect 675268 579730 675407 579732
rect 675268 579674 675346 579730
rect 675402 579674 675407 579730
rect 675268 579672 675407 579674
rect 675268 579670 675274 579672
rect 675341 579669 675407 579672
rect 677457 573206 677523 573207
rect 677406 573204 677412 573206
rect 677366 573144 677412 573204
rect 677476 573202 677523 573206
rect 677518 573146 677523 573202
rect 677406 573142 677412 573144
rect 677476 573142 677523 573146
rect 677457 573141 677523 573142
rect 41502 570966 41508 571030
rect 41572 571028 41578 571030
rect 41829 571028 41895 571031
rect 41572 571026 41895 571028
rect 41572 570970 41834 571026
rect 41890 570970 41895 571026
rect 41572 570968 41895 570970
rect 41572 570966 41578 570968
rect 41829 570965 41895 570968
rect 41645 570486 41711 570487
rect 41645 570482 41692 570486
rect 41756 570484 41762 570486
rect 41645 570426 41650 570482
rect 41645 570422 41692 570426
rect 41756 570424 41802 570484
rect 41756 570422 41762 570424
rect 41645 570421 41711 570422
rect 41553 569088 41619 569089
rect 41502 569024 41508 569088
rect 41572 569086 41619 569088
rect 42054 569086 42060 569088
rect 41572 569084 42060 569086
rect 41614 569028 42060 569084
rect 41572 569026 42060 569028
rect 41572 569024 41619 569026
rect 42054 569024 42060 569026
rect 42124 569024 42130 569088
rect 41553 569023 41619 569024
rect 41645 563414 41711 563415
rect 41645 563412 41692 563414
rect 41600 563410 41692 563412
rect 41600 563354 41650 563410
rect 41600 563352 41692 563354
rect 41645 563350 41692 563352
rect 41756 563350 41762 563414
rect 41645 563349 41711 563350
rect 41645 558110 41711 558111
rect 41645 558108 41692 558110
rect 41600 558106 41692 558108
rect 41600 558050 41650 558106
rect 41600 558048 41692 558050
rect 41645 558046 41692 558048
rect 41756 558046 41762 558110
rect 41645 558045 41711 558046
rect 41553 557972 41619 557975
rect 41870 557972 41876 557974
rect 41553 557970 41876 557972
rect 41553 557914 41558 557970
rect 41614 557914 41876 557970
rect 41553 557912 41876 557914
rect 41553 557909 41619 557912
rect 41870 557910 41876 557912
rect 41940 557972 41946 557974
rect 42105 557972 42171 557975
rect 41940 557970 42171 557972
rect 41940 557914 42110 557970
rect 42166 557914 42171 557970
rect 41940 557912 42171 557914
rect 41940 557910 41946 557912
rect 42105 557909 42171 557912
rect 42105 557838 42171 557839
rect 42054 557836 42060 557838
rect 42014 557776 42060 557836
rect 42124 557834 42171 557838
rect 42166 557778 42171 557834
rect 42054 557774 42060 557776
rect 42124 557774 42171 557778
rect 42105 557773 42171 557774
rect 41686 555326 41692 555390
rect 41756 555388 41762 555390
rect 41829 555388 41895 555391
rect 41756 555386 41895 555388
rect 41756 555330 41834 555386
rect 41890 555330 41895 555386
rect 41756 555328 41895 555330
rect 41756 555326 41762 555328
rect 41829 555325 41895 555328
rect 41921 555254 41987 555255
rect 41870 555190 41876 555254
rect 41940 555252 41987 555254
rect 41940 555250 42032 555252
rect 41982 555194 42032 555250
rect 41940 555192 42032 555194
rect 41940 555190 41987 555192
rect 41921 555189 41987 555190
rect 677406 550022 677412 550086
rect 677476 550084 677482 550086
rect 677733 550084 677799 550087
rect 677476 550082 677799 550084
rect 677476 550026 677738 550082
rect 677794 550026 677799 550082
rect 677476 550024 677799 550026
rect 677476 550022 677482 550024
rect 677733 550021 677799 550024
rect 42105 526558 42171 526559
rect 42054 526556 42060 526558
rect 42014 526496 42060 526556
rect 42124 526554 42171 526558
rect 42166 526498 42171 526554
rect 42054 526494 42060 526496
rect 42124 526494 42171 526498
rect 42105 526493 42171 526494
rect 41553 526328 41619 526329
rect 41502 526326 41508 526328
rect 41462 526266 41508 526326
rect 41572 526324 41619 526328
rect 41614 526268 41619 526324
rect 41502 526264 41508 526266
rect 41572 526264 41619 526268
rect 41553 526263 41619 526264
rect 41870 519014 41876 519078
rect 41940 519076 41946 519078
rect 42105 519076 42171 519079
rect 41940 519074 42171 519076
rect 41940 519018 42110 519074
rect 42166 519018 42171 519074
rect 41940 519016 42171 519018
rect 41940 519014 41946 519016
rect 42105 519013 42171 519016
rect 41553 518324 41619 518325
rect 41502 518260 41508 518324
rect 41572 518322 41619 518324
rect 41572 518320 41664 518322
rect 41614 518264 41664 518320
rect 41572 518262 41664 518264
rect 41572 518260 41619 518262
rect 41553 518259 41619 518260
rect 41553 513998 41619 514001
rect 41870 513998 41876 514000
rect 41553 513996 41876 513998
rect 41553 513940 41558 513996
rect 41614 513940 41876 513996
rect 41553 513938 41876 513940
rect 41553 513935 41619 513938
rect 41870 513936 41876 513938
rect 41940 513936 41946 514000
rect 41553 513366 41619 513367
rect 41502 513302 41508 513366
rect 41572 513364 41619 513366
rect 42054 513364 42060 513366
rect 41572 513362 42060 513364
rect 41614 513306 42060 513362
rect 41572 513304 42060 513306
rect 41572 513302 41619 513304
rect 42054 513302 42060 513304
rect 42124 513302 42130 513366
rect 41553 513301 41619 513302
rect 41502 510718 41508 510782
rect 41572 510780 41578 510782
rect 41645 510780 41711 510783
rect 41921 510782 41987 510783
rect 41870 510780 41876 510782
rect 41572 510778 41711 510780
rect 41572 510722 41650 510778
rect 41706 510722 41711 510778
rect 41572 510720 41711 510722
rect 41830 510720 41876 510780
rect 41940 510778 41987 510782
rect 41982 510722 41987 510778
rect 41572 510718 41578 510720
rect 41645 510717 41711 510720
rect 41870 510718 41876 510720
rect 41940 510718 41987 510722
rect 41921 510717 41987 510718
rect 674881 498676 674947 498679
rect 674881 498674 677628 498676
rect 674881 498618 674886 498674
rect 674942 498618 677628 498674
rect 674881 498616 677628 498618
rect 674881 498613 674947 498616
rect 674789 495276 674855 495279
rect 674789 495274 677628 495276
rect 674789 495218 674794 495274
rect 674850 495218 677628 495274
rect 674789 495216 677628 495218
rect 674789 495213 674855 495216
rect 674605 493236 674671 493239
rect 674973 493236 675039 493239
rect 674605 493234 677658 493236
rect 674605 493178 674610 493234
rect 674666 493178 674978 493234
rect 675034 493178 677658 493234
rect 674605 493176 677658 493178
rect 674605 493173 674671 493176
rect 674973 493173 675039 493176
rect 677598 492934 677658 493176
rect 39516 477128 39730 477188
rect 39670 476508 39730 477128
rect 42473 476508 42539 476511
rect 39670 476506 42539 476508
rect 39670 476450 42478 476506
rect 42534 476450 42539 476506
rect 39670 476448 42539 476450
rect 42473 476445 42539 476448
rect 42473 474876 42539 474879
rect 39670 474874 42539 474876
rect 39670 474818 42478 474874
rect 42534 474818 42539 474874
rect 39670 474816 42539 474818
rect 39670 474740 39730 474816
rect 42473 474813 42539 474816
rect 39516 474680 39730 474740
rect 42381 472972 42447 472975
rect 39670 472970 42447 472972
rect 39670 472914 42386 472970
rect 42442 472914 42447 472970
rect 39670 472912 42447 472914
rect 39670 472292 39730 472912
rect 42381 472909 42447 472912
rect 39516 472232 39730 472292
rect 677406 459854 677412 459918
rect 677476 459916 677482 459918
rect 677917 459916 677983 459919
rect 677476 459914 677983 459916
rect 677476 459858 677922 459914
rect 677978 459858 677983 459914
rect 677476 459856 677983 459858
rect 677476 459854 677482 459856
rect 677917 459853 677983 459856
rect 677733 452164 677799 452167
rect 677733 452162 677996 452164
rect 677733 452106 677738 452162
rect 677794 452106 677996 452162
rect 677733 452104 677996 452106
rect 677733 452101 677799 452104
rect 675065 449716 675131 449719
rect 675065 449714 677996 449716
rect 675065 449658 675070 449714
rect 675126 449686 677996 449714
rect 675126 449658 678026 449686
rect 675065 449656 678026 449658
rect 675065 449653 675131 449656
rect 677966 447238 678026 449656
rect 39713 437884 39779 437887
rect 39846 437884 39852 437886
rect 39713 437882 39852 437884
rect 39713 437826 39718 437882
rect 39774 437826 39852 437882
rect 39713 437824 39852 437826
rect 39713 437821 39779 437824
rect 39846 437822 39852 437824
rect 39916 437822 39922 437886
rect 42289 431356 42355 431359
rect 39332 431354 42355 431356
rect 39332 431326 42294 431354
rect 39302 431298 42294 431326
rect 42350 431298 42355 431354
rect 39302 431296 42355 431298
rect 39302 428878 39362 431296
rect 42289 431293 42355 431296
rect 674830 428846 674836 428910
rect 674900 428908 674906 428910
rect 674973 428908 675039 428911
rect 674900 428906 675039 428908
rect 674900 428850 674978 428906
rect 675034 428850 675039 428906
rect 674900 428848 675039 428850
rect 674900 428846 674906 428848
rect 674973 428845 675039 428848
rect 674881 425102 674947 425103
rect 674830 425038 674836 425102
rect 674900 425100 674947 425102
rect 674900 425098 674992 425100
rect 674942 425042 674992 425098
rect 674900 425040 674992 425042
rect 674900 425038 674947 425040
rect 674881 425037 674947 425038
rect 39529 423740 39595 423743
rect 39713 423740 39779 423743
rect 39332 423738 39779 423740
rect 39332 423682 39534 423738
rect 39590 423682 39718 423738
rect 39774 423682 39779 423738
rect 39332 423680 39779 423682
rect 39529 423677 39595 423680
rect 39713 423677 39779 423680
rect 674789 406604 674855 406607
rect 677457 406604 677523 406607
rect 674789 406602 677628 406604
rect 674789 406546 674794 406602
rect 674850 406546 677462 406602
rect 677518 406546 677628 406602
rect 674789 406544 677628 406546
rect 674789 406541 674855 406544
rect 677457 406541 677523 406544
rect 675065 401708 675131 401711
rect 675065 401706 677628 401708
rect 675065 401650 675070 401706
rect 675126 401650 677628 401706
rect 675065 401648 677628 401650
rect 675065 401645 675131 401648
rect 42105 381988 42171 381991
rect 41510 381986 42171 381988
rect 41510 381930 42110 381986
rect 42166 381930 42171 381986
rect 41510 381928 42171 381930
rect 41510 381757 41570 381928
rect 42105 381925 42171 381928
rect 41510 381756 41619 381757
rect 41502 381692 41508 381756
rect 41572 381754 41619 381756
rect 41572 381752 41664 381754
rect 41614 381696 41664 381752
rect 41572 381694 41664 381696
rect 41572 381692 41619 381694
rect 41553 381691 41619 381692
rect 41502 379206 41508 379270
rect 41572 379268 41578 379270
rect 41737 379268 41803 379271
rect 41572 379266 41803 379268
rect 41572 379210 41742 379266
rect 41798 379210 41803 379266
rect 41572 379208 41803 379210
rect 41572 379206 41578 379208
rect 41737 379205 41803 379208
rect 675157 356964 675223 356967
rect 675022 356962 675223 356964
rect 675022 356906 675162 356962
rect 675218 356906 675223 356962
rect 675022 356904 675223 356906
rect 675022 356695 675082 356904
rect 675157 356901 675223 356904
rect 674973 356690 675082 356695
rect 674973 356634 674978 356690
rect 675034 356634 675082 356690
rect 674973 356632 675082 356634
rect 674973 356629 675039 356632
rect 674881 350164 674947 350167
rect 675249 350164 675315 350167
rect 674881 350162 675315 350164
rect 674881 350106 674886 350162
rect 674942 350106 675254 350162
rect 675310 350106 675315 350162
rect 674881 350104 675315 350106
rect 674881 350101 674947 350104
rect 675249 350101 675315 350104
rect 675198 318958 675204 319022
rect 675268 319020 675274 319022
rect 675341 319020 675407 319023
rect 675268 319018 675407 319020
rect 675268 318962 675346 319018
rect 675402 318962 675407 319018
rect 675268 318960 675407 318962
rect 675268 318958 675274 318960
rect 675341 318957 675407 318960
rect 675249 316512 675315 316513
rect 675198 316448 675204 316512
rect 675268 316510 675315 316512
rect 675750 316510 675756 316512
rect 675268 316508 675756 316510
rect 675310 316452 675756 316508
rect 675268 316450 675756 316452
rect 675268 316448 675315 316450
rect 675750 316448 675756 316450
rect 675820 316448 675826 316512
rect 675249 316447 675315 316448
rect 41645 305830 41711 305831
rect 41645 305828 41692 305830
rect 41600 305826 41692 305828
rect 41600 305770 41650 305826
rect 41600 305768 41692 305770
rect 41645 305766 41692 305768
rect 41756 305766 41762 305830
rect 41645 305765 41711 305766
rect 41686 297606 41692 297670
rect 41756 297668 41762 297670
rect 42105 297668 42171 297671
rect 41756 297666 42171 297668
rect 41756 297610 42110 297666
rect 42166 297610 42171 297666
rect 41756 297608 42171 297610
rect 41756 297606 41762 297608
rect 42105 297605 42171 297608
rect 41553 293400 41619 293401
rect 41502 293336 41508 293400
rect 41572 293398 41619 293400
rect 41572 293396 41664 293398
rect 41614 293340 41664 293396
rect 41572 293338 41664 293340
rect 41572 293336 41619 293338
rect 41553 293335 41619 293336
rect 41553 292772 41619 292775
rect 41686 292772 41692 292774
rect 41553 292770 41692 292772
rect 41553 292714 41558 292770
rect 41614 292714 41692 292770
rect 41553 292712 41692 292714
rect 41553 292709 41619 292712
rect 41686 292710 41692 292712
rect 41756 292772 41762 292774
rect 42289 292772 42355 292775
rect 41756 292770 42355 292772
rect 41756 292714 42294 292770
rect 42350 292714 42355 292770
rect 41756 292712 42355 292714
rect 41756 292710 41762 292712
rect 42289 292709 42355 292712
rect 41737 290190 41803 290191
rect 41686 290188 41692 290190
rect 41646 290128 41692 290188
rect 41756 290186 41803 290190
rect 41798 290130 41803 290186
rect 41686 290126 41692 290128
rect 41756 290126 41803 290130
rect 41737 290125 41803 290126
rect 41502 287134 41508 287198
rect 41572 287196 41578 287198
rect 41645 287196 41711 287199
rect 41572 287194 41711 287196
rect 41572 287138 41650 287194
rect 41706 287138 41711 287194
rect 41572 287136 41711 287138
rect 41572 287134 41578 287136
rect 41645 287133 41711 287136
rect 675525 271148 675591 271151
rect 675934 271148 675940 271150
rect 675525 271146 675940 271148
rect 675525 271090 675530 271146
rect 675586 271090 675940 271146
rect 675525 271088 675940 271090
rect 675525 271085 675591 271088
rect 675934 271086 675940 271088
rect 676004 271086 676010 271150
rect 41553 248164 41619 248167
rect 41686 248164 41692 248166
rect 41553 248162 41692 248164
rect 41553 248106 41558 248162
rect 41614 248106 41692 248162
rect 41553 248104 41692 248106
rect 41553 248101 41619 248104
rect 41686 248102 41692 248104
rect 41756 248164 41762 248166
rect 42289 248164 42355 248167
rect 41756 248162 42355 248164
rect 41756 248106 42294 248162
rect 42350 248106 42355 248162
rect 41756 248104 42355 248106
rect 41756 248102 41762 248104
rect 42289 248101 42355 248104
rect 41737 245582 41803 245583
rect 41686 245580 41692 245582
rect 41646 245520 41692 245580
rect 41756 245578 41803 245582
rect 41798 245522 41803 245578
rect 41686 245518 41692 245520
rect 41756 245518 41803 245522
rect 41737 245517 41803 245518
rect 675249 218516 675315 218519
rect 675206 218514 675315 218516
rect 675206 218458 675254 218514
rect 675310 218458 675315 218514
rect 675206 218453 675315 218458
rect 675206 218383 675266 218453
rect 675206 218378 675315 218383
rect 675206 218322 675254 218378
rect 675310 218322 675315 218378
rect 675206 218320 675315 218322
rect 675249 218317 675315 218320
rect 41645 216750 41711 216751
rect 41645 216748 41692 216750
rect 41600 216746 41692 216748
rect 41600 216690 41650 216746
rect 41600 216688 41692 216690
rect 41645 216686 41692 216688
rect 41756 216686 41762 216750
rect 41645 216685 41711 216686
rect 41686 215054 41692 215118
rect 41756 215116 41762 215118
rect 42105 215116 42171 215119
rect 41756 215114 42171 215116
rect 41756 215058 42110 215114
rect 42166 215058 42171 215114
rect 41756 215056 42171 215058
rect 41756 215054 41762 215056
rect 42105 215053 42171 215056
rect 41645 214166 41711 214167
rect 41645 214164 41692 214166
rect 41600 214162 41692 214164
rect 41600 214106 41650 214162
rect 41600 214104 41692 214106
rect 41645 214102 41692 214104
rect 41756 214102 41762 214166
rect 41645 214101 41711 214102
rect 674881 212396 674947 212399
rect 675249 212396 675315 212399
rect 674881 212394 675315 212396
rect 674881 212338 674886 212394
rect 674942 212338 675254 212394
rect 675310 212338 675315 212394
rect 674881 212336 675315 212338
rect 674881 212333 674947 212336
rect 675249 212333 675315 212336
rect 41686 209614 41692 209678
rect 41756 209676 41762 209678
rect 42105 209676 42171 209679
rect 41756 209674 42171 209676
rect 41756 209618 42110 209674
rect 42166 209618 42171 209674
rect 41756 209616 42171 209618
rect 41756 209614 41762 209616
rect 42105 209613 42171 209616
rect 41502 209206 41508 209270
rect 41572 209268 41578 209270
rect 41645 209268 41711 209271
rect 41572 209266 41711 209268
rect 41572 209210 41650 209266
rect 41706 209210 41711 209266
rect 41572 209208 41711 209210
rect 41572 209206 41578 209208
rect 41645 209205 41711 209208
rect 41553 204200 41619 204201
rect 41502 204136 41508 204200
rect 41572 204198 41619 204200
rect 41572 204196 41664 204198
rect 41614 204140 41664 204196
rect 41572 204138 41664 204140
rect 41572 204136 41619 204138
rect 41553 204135 41619 204136
rect 41502 200910 41508 200974
rect 41572 200972 41578 200974
rect 41645 200972 41711 200975
rect 41572 200970 41711 200972
rect 41572 200914 41650 200970
rect 41706 200914 41711 200970
rect 41572 200912 41711 200914
rect 41572 200910 41578 200912
rect 41645 200909 41711 200912
rect 675249 189548 675315 189551
rect 675249 189546 675634 189548
rect 675249 189490 675254 189546
rect 675310 189490 675634 189546
rect 675249 189488 675634 189490
rect 675249 189485 675315 189488
rect 675574 189415 675634 189488
rect 675574 189410 675683 189415
rect 675574 189354 675622 189410
rect 675678 189354 675683 189410
rect 675574 189352 675683 189354
rect 675617 189349 675683 189352
rect 41686 172214 41692 172278
rect 41756 172276 41762 172278
rect 42105 172276 42171 172279
rect 41756 172274 42171 172276
rect 41756 172218 42110 172274
rect 42166 172218 42171 172274
rect 41756 172216 42171 172218
rect 41756 172214 41762 172216
rect 42105 172213 42171 172216
rect 41553 170286 41619 170289
rect 41686 170286 41692 170288
rect 41553 170284 41692 170286
rect 41553 170228 41558 170284
rect 41614 170228 41692 170284
rect 41553 170226 41692 170228
rect 41553 170223 41619 170226
rect 41686 170224 41692 170226
rect 41756 170236 41762 170288
rect 42657 170236 42723 170239
rect 41756 170234 42723 170236
rect 41756 170224 42662 170234
rect 41694 170178 42662 170224
rect 42718 170178 42723 170234
rect 41694 170176 42723 170178
rect 42657 170173 42723 170176
rect 675249 130312 675315 130313
rect 675198 130248 675204 130312
rect 675268 130310 675315 130312
rect 675268 130308 675360 130310
rect 675310 130252 675360 130308
rect 675268 130250 675360 130252
rect 675268 130248 675315 130250
rect 675249 130247 675315 130248
rect 42197 120460 42263 120463
rect 39516 120458 42263 120460
rect 39516 120402 42202 120458
rect 42258 120402 42263 120458
rect 39516 120400 42263 120402
rect 42197 120397 42263 120400
rect 675065 119780 675131 119783
rect 675198 119780 675204 119782
rect 675065 119778 675204 119780
rect 675065 119722 675070 119778
rect 675126 119722 675204 119778
rect 675065 119720 675204 119722
rect 675065 119717 675131 119720
rect 675198 119718 675204 119720
rect 675268 119718 675274 119782
rect 42197 112980 42263 112983
rect 43025 112980 43091 112983
rect 39700 112978 43091 112980
rect 39700 112922 42202 112978
rect 42258 112922 43030 112978
rect 43086 112922 43091 112978
rect 39700 112920 43091 112922
rect 42197 112917 42263 112920
rect 43025 112917 43091 112920
rect 42289 76940 42355 76943
rect 43945 76940 44011 76943
rect 39332 76938 44011 76940
rect 39332 76882 42294 76938
rect 42350 76882 43950 76938
rect 44006 76882 44011 76938
rect 39332 76880 44011 76882
rect 39670 76532 39730 76880
rect 42289 76877 42355 76880
rect 43945 76877 44011 76880
rect 39302 76472 39730 76532
rect 39302 74492 39362 76472
rect 39302 74462 39730 74492
rect 39332 74432 39730 74462
rect 39670 74084 39730 74432
rect 39302 74024 39730 74084
rect 39302 73646 39362 74024
rect 540837 45116 540903 45119
rect 553625 45116 553691 45119
rect 540837 45114 553691 45116
rect 540837 45058 540842 45114
rect 540898 45058 553630 45114
rect 553686 45058 553691 45114
rect 540837 45056 553691 45058
rect 540837 45053 540903 45056
rect 553625 45053 553691 45056
rect 218837 44844 218903 44847
rect 231625 44844 231691 44847
rect 218837 44842 231691 44844
rect 218837 44786 218842 44842
rect 218898 44786 231630 44842
rect 231686 44786 231691 44842
rect 218837 44784 231691 44786
rect 218837 44781 218903 44784
rect 231625 44781 231691 44784
rect 244597 44844 244663 44847
rect 257385 44844 257451 44847
rect 244597 44842 257451 44844
rect 244597 44786 244602 44842
rect 244658 44786 257390 44842
rect 257446 44786 257451 44842
rect 244597 44784 257451 44786
rect 244597 44781 244663 44784
rect 257385 44781 257451 44784
rect 424917 44844 424983 44847
rect 437705 44844 437771 44847
rect 424917 44842 437771 44844
rect 424917 44786 424922 44842
rect 424978 44786 437710 44842
rect 437766 44786 437771 44842
rect 424917 44784 437771 44786
rect 424917 44781 424983 44784
rect 437705 44781 437771 44784
rect 450677 44708 450743 44711
rect 463465 44708 463531 44711
rect 450677 44706 463531 44708
rect 450677 44650 450682 44706
rect 450738 44650 463470 44706
rect 463526 44650 463531 44706
rect 450677 44648 463531 44650
rect 450677 44645 450743 44648
rect 463465 44645 463531 44648
rect 579477 44708 579543 44711
rect 592265 44708 592331 44711
rect 579477 44706 592331 44708
rect 579477 44650 579482 44706
rect 579538 44650 592270 44706
rect 592326 44650 592331 44706
rect 579477 44648 592331 44650
rect 579477 44645 579543 44648
rect 592265 44645 592331 44648
rect 605237 44708 605303 44711
rect 618025 44708 618091 44711
rect 605237 44706 618091 44708
rect 605237 44650 605242 44706
rect 605298 44650 618030 44706
rect 618086 44650 618091 44706
rect 605237 44648 618091 44650
rect 605237 44645 605303 44648
rect 618025 44645 618091 44648
rect 630997 44708 631063 44711
rect 643785 44708 643851 44711
rect 630997 44706 643851 44708
rect 630997 44650 631002 44706
rect 631058 44650 643790 44706
rect 643846 44650 643851 44706
rect 630997 44648 643851 44650
rect 630997 44645 631063 44648
rect 643785 44645 643851 44648
rect 656757 44708 656823 44711
rect 669545 44708 669611 44711
rect 656757 44706 669611 44708
rect 656757 44650 656762 44706
rect 656818 44650 669550 44706
rect 669606 44650 669611 44706
rect 656757 44648 669611 44650
rect 656757 44645 656823 44648
rect 669545 44645 669611 44648
rect 468801 44572 468867 44575
rect 476345 44572 476411 44575
rect 468801 44570 476411 44572
rect 468801 44514 468806 44570
rect 468862 44514 476350 44570
rect 476406 44514 476411 44570
rect 468801 44512 476411 44514
rect 468801 44509 468867 44512
rect 476345 44509 476411 44512
rect 480117 44572 480183 44575
rect 489225 44572 489291 44575
rect 480117 44570 489291 44572
rect 480117 44514 480122 44570
rect 480178 44514 489230 44570
rect 489286 44514 489291 44570
rect 480117 44512 489291 44514
rect 480117 44509 480183 44512
rect 489225 44509 489291 44512
rect 334757 44300 334823 44303
rect 344877 44300 344943 44303
rect 334757 44298 344943 44300
rect 334757 44242 334762 44298
rect 334818 44242 344882 44298
rect 344938 44242 344943 44298
rect 334757 44240 344943 44242
rect 334757 44237 334823 44240
rect 344877 44237 344943 44240
rect 469261 41988 469327 41991
rect 470549 41988 470615 41991
rect 472941 41988 473007 41991
rect 473585 41988 473651 41991
rect 467470 41986 473651 41988
rect 467470 41930 469266 41986
rect 469322 41930 470554 41986
rect 470610 41930 472946 41986
rect 473002 41930 473590 41986
rect 473646 41930 473651 41986
rect 467470 41928 473651 41930
rect 465029 41852 465095 41855
rect 466317 41852 466383 41855
rect 467470 41852 467530 41928
rect 469261 41925 469327 41928
rect 470549 41925 470615 41928
rect 472941 41925 473007 41928
rect 473585 41925 473651 41928
rect 465029 41850 467530 41852
rect 465029 41794 465034 41850
rect 465090 41794 466322 41850
rect 466378 41794 467530 41850
rect 465029 41792 467530 41794
rect 465029 41789 465095 41792
rect 466317 41789 466383 41792
rect 84198 40432 623010 40492
rect 84198 40220 84258 40432
rect 148917 40356 148983 40359
rect 145702 40354 148983 40356
rect 145702 40298 148922 40354
rect 148978 40298 148983 40354
rect 145702 40296 148983 40298
rect 90865 40220 90931 40223
rect 134105 40220 134171 40223
rect 84014 40160 84258 40220
rect 88798 40218 90931 40220
rect 88798 40162 90870 40218
rect 90926 40162 90931 40218
rect 88798 40160 90931 40162
rect 84014 39646 84074 40160
rect 88798 39679 88858 40160
rect 90865 40157 90931 40160
rect 132958 40218 134171 40220
rect 132958 40162 134110 40218
rect 134166 40162 134171 40218
rect 132958 40160 134171 40162
rect 132958 39986 133018 40160
rect 134105 40157 134171 40160
rect 142937 40220 143003 40223
rect 143397 40220 143463 40223
rect 142937 40218 143322 40220
rect 142937 40162 142942 40218
rect 142998 40162 143322 40218
rect 142937 40160 143322 40162
rect 142937 40157 143003 40160
rect 143262 39986 143322 40160
rect 143397 40218 143874 40220
rect 143397 40162 143402 40218
rect 143458 40162 143874 40218
rect 143397 40160 143874 40162
rect 143397 40157 143463 40160
rect 143814 39986 143874 40160
rect 145702 40016 145762 40296
rect 148917 40293 148983 40296
rect 569081 40220 569147 40223
rect 569038 40218 569147 40220
rect 569038 40162 569086 40218
rect 569142 40162 569147 40218
rect 569038 40157 569147 40162
rect 251957 40084 252023 40087
rect 145684 39956 145762 40016
rect 248694 40082 252023 40084
rect 248694 40026 251962 40082
rect 252018 40026 252023 40082
rect 248694 40024 252023 40026
rect 244505 39948 244571 39951
rect 244505 39946 246362 39948
rect 244505 39890 244510 39946
rect 244566 39890 246362 39946
rect 244505 39888 246362 39890
rect 244505 39885 244571 39888
rect 88798 39674 88907 39679
rect 88798 39646 88846 39674
rect 88828 39618 88846 39646
rect 88902 39618 88907 39674
rect 88828 39616 88907 39618
rect 88841 39613 88907 39616
rect 246302 39540 246362 39888
rect 248694 39540 248754 40024
rect 251957 40021 252023 40024
rect 251313 39948 251379 39951
rect 246302 39480 248754 39540
rect 246302 39374 246362 39480
rect 248694 39374 248754 39480
rect 251270 39946 251379 39948
rect 251270 39890 251318 39946
rect 251374 39890 251379 39946
rect 251270 39885 251379 39890
rect 251270 39374 251330 39885
rect 569038 39646 569098 40157
rect 622625 39812 622691 39815
rect 622950 39812 623010 40432
rect 630261 40220 630327 40223
rect 630261 40218 630370 40220
rect 630261 40162 630266 40218
rect 630322 40162 630370 40218
rect 630261 40157 630370 40162
rect 622625 39810 623010 39812
rect 622625 39754 622630 39810
rect 622686 39754 623010 39810
rect 622625 39752 623010 39754
rect 622625 39749 622691 39752
rect 622950 39646 623010 39752
rect 630310 39646 630370 40157
<< via3 >>
rect 677412 915590 677476 915654
rect 39852 903622 39916 903686
rect 41876 793598 41940 793662
rect 41876 789714 41940 789718
rect 41876 789658 41926 789714
rect 41926 789658 41940 789714
rect 41876 789654 41940 789658
rect 41692 789518 41756 789582
rect 41692 786042 41756 786046
rect 41692 785986 41706 786042
rect 41706 785986 41756 786042
rect 41692 785982 41756 785986
rect 41692 780738 41756 780742
rect 41692 780682 41706 780738
rect 41706 780682 41756 780738
rect 41692 780678 41756 780682
rect 41140 780492 41204 780556
rect 41692 778018 41756 778022
rect 41692 777962 41706 778018
rect 41706 777962 41756 778018
rect 41692 777958 41756 777962
rect 675572 744366 675636 744430
rect 41876 743550 41940 743614
rect 41876 736536 41940 736600
rect 41140 735892 41204 735956
rect 41876 733350 41940 733414
rect 675572 731990 675636 732054
rect 675388 721110 675452 721174
rect 675572 719538 675636 719542
rect 675572 719482 675586 719538
rect 675586 719482 675636 719538
rect 675572 719478 675636 719482
rect 675388 719266 675452 719270
rect 675388 719210 675438 719266
rect 675438 719210 675452 719266
rect 675388 719206 675452 719210
rect 41876 704790 41940 704854
rect 41508 704654 41572 704718
rect 41692 704464 41756 704528
rect 41692 696460 41756 696524
rect 41876 696358 41940 696422
rect 41508 692686 41572 692750
rect 41508 688878 41572 688942
rect 675388 688878 675452 688942
rect 675388 685404 675452 685468
rect 41508 660046 41572 660110
rect 41692 659864 41756 659928
rect 41508 658066 41572 658070
rect 41508 658010 41558 658066
rect 41558 658010 41572 658066
rect 41508 658006 41572 658010
rect 42060 653306 42124 653310
rect 42060 653250 42074 653306
rect 42074 653250 42124 653306
rect 42060 653246 42124 653250
rect 41692 652354 41756 652358
rect 41692 652298 41706 652354
rect 41706 652298 41756 652354
rect 41692 652294 41756 652298
rect 42060 648002 42124 648006
rect 42060 647946 42110 648002
rect 42110 647946 42124 648002
rect 42060 647942 42124 647946
rect 42060 647050 42124 647054
rect 42060 646994 42110 647050
rect 42110 646994 42124 647050
rect 42060 646990 42124 646994
rect 42060 644134 42124 644198
rect 675204 642094 675268 642158
rect 675020 641958 675084 642022
rect 675204 638890 675268 638894
rect 675204 638834 675254 638890
rect 675254 638834 675268 638890
rect 675204 638830 675268 638834
rect 675020 628316 675084 628380
rect 675388 628316 675452 628380
rect 675204 626378 675268 626382
rect 675204 626322 675218 626378
rect 675218 626322 675268 626378
rect 675204 626318 675268 626322
rect 675388 626318 675452 626382
rect 41876 615710 41940 615774
rect 41324 615438 41388 615502
rect 41508 615324 41572 615328
rect 41508 615268 41558 615324
rect 41558 615268 41572 615324
rect 41508 615264 41572 615268
rect 41876 613806 41940 613870
rect 41508 607338 41572 607342
rect 41508 607282 41558 607338
rect 41558 607282 41572 607338
rect 41508 607278 41572 607282
rect 41692 602926 41756 602990
rect 41508 602352 41572 602356
rect 41508 602296 41558 602352
rect 41558 602296 41572 602352
rect 41508 602292 41572 602296
rect 41508 599798 41572 599862
rect 41692 599662 41756 599726
rect 675204 583402 675268 583406
rect 675204 583346 675218 583402
rect 675218 583346 675268 583402
rect 675204 583342 675268 583346
rect 675204 581770 675268 581774
rect 675204 581714 675254 581770
rect 675254 581714 675268 581770
rect 675204 581710 675268 581714
rect 675204 579670 675268 579734
rect 677412 573202 677476 573206
rect 677412 573146 677462 573202
rect 677462 573146 677476 573202
rect 677412 573142 677476 573146
rect 41508 570966 41572 571030
rect 41692 570482 41756 570486
rect 41692 570426 41706 570482
rect 41706 570426 41756 570482
rect 41692 570422 41756 570426
rect 41508 569084 41572 569088
rect 41508 569028 41558 569084
rect 41558 569028 41572 569084
rect 41508 569024 41572 569028
rect 42060 569024 42124 569088
rect 41692 563410 41756 563414
rect 41692 563354 41706 563410
rect 41706 563354 41756 563410
rect 41692 563350 41756 563354
rect 41692 558106 41756 558110
rect 41692 558050 41706 558106
rect 41706 558050 41756 558106
rect 41692 558046 41756 558050
rect 41876 557910 41940 557974
rect 42060 557834 42124 557838
rect 42060 557778 42110 557834
rect 42110 557778 42124 557834
rect 42060 557774 42124 557778
rect 41692 555326 41756 555390
rect 41876 555250 41940 555254
rect 41876 555194 41926 555250
rect 41926 555194 41940 555250
rect 41876 555190 41940 555194
rect 677412 550022 677476 550086
rect 42060 526554 42124 526558
rect 42060 526498 42110 526554
rect 42110 526498 42124 526554
rect 42060 526494 42124 526498
rect 41508 526324 41572 526328
rect 41508 526268 41558 526324
rect 41558 526268 41572 526324
rect 41508 526264 41572 526268
rect 41876 519014 41940 519078
rect 41508 518320 41572 518324
rect 41508 518264 41558 518320
rect 41558 518264 41572 518320
rect 41508 518260 41572 518264
rect 41876 513936 41940 514000
rect 41508 513362 41572 513366
rect 41508 513306 41558 513362
rect 41558 513306 41572 513362
rect 41508 513302 41572 513306
rect 42060 513302 42124 513366
rect 41508 510718 41572 510782
rect 41876 510778 41940 510782
rect 41876 510722 41926 510778
rect 41926 510722 41940 510778
rect 41876 510718 41940 510722
rect 677412 459854 677476 459918
rect 39852 437822 39916 437886
rect 674836 428846 674900 428910
rect 674836 425098 674900 425102
rect 674836 425042 674886 425098
rect 674886 425042 674900 425098
rect 674836 425038 674900 425042
rect 41508 381752 41572 381756
rect 41508 381696 41558 381752
rect 41558 381696 41572 381752
rect 41508 381692 41572 381696
rect 41508 379206 41572 379270
rect 675204 318958 675268 319022
rect 675204 316508 675268 316512
rect 675204 316452 675254 316508
rect 675254 316452 675268 316508
rect 675204 316448 675268 316452
rect 675756 316448 675820 316512
rect 41692 305826 41756 305830
rect 41692 305770 41706 305826
rect 41706 305770 41756 305826
rect 41692 305766 41756 305770
rect 41692 297606 41756 297670
rect 41508 293396 41572 293400
rect 41508 293340 41558 293396
rect 41558 293340 41572 293396
rect 41508 293336 41572 293340
rect 41692 292710 41756 292774
rect 41692 290186 41756 290190
rect 41692 290130 41742 290186
rect 41742 290130 41756 290186
rect 41692 290126 41756 290130
rect 41508 287134 41572 287198
rect 675940 271086 676004 271150
rect 41692 248102 41756 248166
rect 41692 245578 41756 245582
rect 41692 245522 41742 245578
rect 41742 245522 41756 245578
rect 41692 245518 41756 245522
rect 41692 216746 41756 216750
rect 41692 216690 41706 216746
rect 41706 216690 41756 216746
rect 41692 216686 41756 216690
rect 41692 215054 41756 215118
rect 41692 214162 41756 214166
rect 41692 214106 41706 214162
rect 41706 214106 41756 214162
rect 41692 214102 41756 214106
rect 41692 209614 41756 209678
rect 41508 209206 41572 209270
rect 41508 204196 41572 204200
rect 41508 204140 41558 204196
rect 41558 204140 41572 204196
rect 41508 204136 41572 204140
rect 41508 200910 41572 200974
rect 41692 172214 41756 172278
rect 41692 170224 41756 170288
rect 675204 130308 675268 130312
rect 675204 130252 675254 130308
rect 675254 130252 675268 130308
rect 675204 130248 675268 130252
rect 675204 119718 675268 119782
<< metal4 >>
rect 677411 915654 677477 915655
rect 677411 915590 677412 915654
rect 677476 915590 677477 915654
rect 677411 915589 677477 915590
rect 39851 903686 39917 903687
rect 39851 903622 39852 903686
rect 39916 903622 39917 903686
rect 39851 903621 39917 903622
rect 39854 437887 39914 903621
rect 41875 793662 41941 793663
rect 41875 793598 41876 793662
rect 41940 793598 41941 793662
rect 41875 793597 41941 793598
rect 41878 789719 41938 793597
rect 41875 789718 41941 789719
rect 41875 789654 41876 789718
rect 41940 789654 41941 789718
rect 41875 789653 41941 789654
rect 41691 789582 41757 789583
rect 41691 789518 41692 789582
rect 41756 789518 41757 789582
rect 41691 789517 41757 789518
rect 41694 786047 41754 789517
rect 41691 786046 41757 786047
rect 41691 785982 41692 786046
rect 41756 785982 41757 786046
rect 41691 785981 41757 785982
rect 41691 780742 41757 780743
rect 41691 780678 41692 780742
rect 41756 780678 41757 780742
rect 41691 780677 41757 780678
rect 41139 780556 41205 780557
rect 41139 780492 41140 780556
rect 41204 780492 41205 780556
rect 41139 780491 41205 780492
rect 41142 735957 41202 780491
rect 41694 778023 41754 780677
rect 41691 778022 41757 778023
rect 41691 777958 41692 778022
rect 41756 777958 41757 778022
rect 41691 777957 41757 777958
rect 675571 744430 675637 744431
rect 675571 744366 675572 744430
rect 675636 744366 675637 744430
rect 675571 744365 675637 744366
rect 41875 743614 41941 743615
rect 41875 743550 41876 743614
rect 41940 743550 41941 743614
rect 41875 743549 41941 743550
rect 41878 736601 41938 743549
rect 41875 736600 41941 736601
rect 41875 736536 41876 736600
rect 41940 736536 41941 736600
rect 41875 736535 41941 736536
rect 41139 735956 41205 735957
rect 41139 735892 41140 735956
rect 41204 735892 41205 735956
rect 41139 735891 41205 735892
rect 41878 733415 41938 736535
rect 41875 733414 41941 733415
rect 41875 733350 41876 733414
rect 41940 733350 41941 733414
rect 41875 733349 41941 733350
rect 675574 732055 675634 744365
rect 675571 732054 675637 732055
rect 675571 731990 675572 732054
rect 675636 731990 675637 732054
rect 675571 731989 675637 731990
rect 675387 721174 675453 721175
rect 675387 721110 675388 721174
rect 675452 721110 675453 721174
rect 675387 721109 675453 721110
rect 675390 719271 675450 721109
rect 675574 719543 675634 731989
rect 675571 719542 675637 719543
rect 675571 719478 675572 719542
rect 675636 719478 675637 719542
rect 675571 719477 675637 719478
rect 675387 719270 675453 719271
rect 675387 719206 675388 719270
rect 675452 719206 675453 719270
rect 675387 719205 675453 719206
rect 41875 704854 41941 704855
rect 41875 704790 41876 704854
rect 41940 704790 41941 704854
rect 41875 704789 41941 704790
rect 41507 704718 41573 704719
rect 41507 704654 41508 704718
rect 41572 704654 41573 704718
rect 41507 704653 41573 704654
rect 41510 692751 41570 704653
rect 41691 704528 41757 704529
rect 41691 704464 41692 704528
rect 41756 704464 41757 704528
rect 41691 704463 41757 704464
rect 41694 696525 41754 704463
rect 41691 696524 41757 696525
rect 41691 696460 41692 696524
rect 41756 696460 41757 696524
rect 41691 696459 41757 696460
rect 41878 696423 41938 704789
rect 41875 696422 41941 696423
rect 41875 696358 41876 696422
rect 41940 696358 41941 696422
rect 41875 696357 41941 696358
rect 41507 692750 41573 692751
rect 41507 692686 41508 692750
rect 41572 692686 41573 692750
rect 41507 692685 41573 692686
rect 41510 688943 41570 692685
rect 41507 688942 41573 688943
rect 41507 688878 41508 688942
rect 41572 688878 41573 688942
rect 41507 688877 41573 688878
rect 675387 688942 675453 688943
rect 675387 688878 675388 688942
rect 675452 688878 675453 688942
rect 675387 688877 675453 688878
rect 675390 685469 675450 688877
rect 675387 685468 675453 685469
rect 675387 685404 675388 685468
rect 675452 685404 675453 685468
rect 675387 685403 675453 685404
rect 41507 660110 41573 660111
rect 41507 660046 41508 660110
rect 41572 660046 41573 660110
rect 41507 660045 41573 660046
rect 41510 658071 41570 660045
rect 41691 659928 41757 659929
rect 41691 659864 41692 659928
rect 41756 659864 41757 659928
rect 41691 659863 41757 659864
rect 41507 658070 41573 658071
rect 41507 658006 41508 658070
rect 41572 658006 41573 658070
rect 41507 658005 41573 658006
rect 41694 652359 41754 659863
rect 42059 653310 42125 653311
rect 42059 653246 42060 653310
rect 42124 653246 42125 653310
rect 42059 653245 42125 653246
rect 41691 652358 41757 652359
rect 41691 652294 41692 652358
rect 41756 652294 41757 652358
rect 41691 652293 41757 652294
rect 42062 648007 42122 653245
rect 42059 648006 42125 648007
rect 42059 647942 42060 648006
rect 42124 647942 42125 648006
rect 42059 647941 42125 647942
rect 42059 647054 42125 647055
rect 42059 646990 42060 647054
rect 42124 646990 42125 647054
rect 42059 646989 42125 646990
rect 42062 644199 42122 646989
rect 42059 644198 42125 644199
rect 42059 644134 42060 644198
rect 42124 644134 42125 644198
rect 42059 644133 42125 644134
rect 675203 642158 675269 642159
rect 675203 642094 675204 642158
rect 675268 642094 675269 642158
rect 675203 642093 675269 642094
rect 675019 642022 675085 642023
rect 675019 641958 675020 642022
rect 675084 641958 675085 642022
rect 675019 641957 675085 641958
rect 675022 628381 675082 641957
rect 675206 638895 675266 642093
rect 675203 638894 675269 638895
rect 675203 638830 675204 638894
rect 675268 638830 675269 638894
rect 675203 638829 675269 638830
rect 675019 628380 675085 628381
rect 675019 628316 675020 628380
rect 675084 628316 675085 628380
rect 675019 628315 675085 628316
rect 675206 626383 675266 638829
rect 675387 628380 675453 628381
rect 675387 628316 675388 628380
rect 675452 628316 675453 628380
rect 675387 628315 675453 628316
rect 675390 626383 675450 628315
rect 675203 626382 675269 626383
rect 675203 626318 675204 626382
rect 675268 626318 675269 626382
rect 675203 626317 675269 626318
rect 675387 626382 675453 626383
rect 675387 626318 675388 626382
rect 675452 626318 675453 626382
rect 675387 626317 675453 626318
rect 41875 615774 41941 615775
rect 41875 615710 41876 615774
rect 41940 615710 41941 615774
rect 41875 615709 41941 615710
rect 41323 615502 41389 615503
rect 41323 615438 41324 615502
rect 41388 615438 41389 615502
rect 41323 615437 41389 615438
rect 41326 606932 41386 615437
rect 41507 615328 41573 615329
rect 41507 615264 41508 615328
rect 41572 615264 41573 615328
rect 41507 615263 41573 615264
rect 41510 607343 41570 615263
rect 41878 613871 41938 615709
rect 41875 613870 41941 613871
rect 41875 613806 41876 613870
rect 41940 613806 41941 613870
rect 41875 613805 41941 613806
rect 41507 607342 41573 607343
rect 41507 607278 41508 607342
rect 41572 607278 41573 607342
rect 41507 607277 41573 607278
rect 41326 606872 41570 606932
rect 41510 602357 41570 606872
rect 41691 602990 41757 602991
rect 41691 602926 41692 602990
rect 41756 602926 41757 602990
rect 41691 602925 41757 602926
rect 41507 602356 41573 602357
rect 41507 602292 41508 602356
rect 41572 602292 41573 602356
rect 41507 602291 41573 602292
rect 41510 599863 41570 602291
rect 41507 599862 41573 599863
rect 41507 599798 41508 599862
rect 41572 599798 41573 599862
rect 41507 599797 41573 599798
rect 41694 599727 41754 602925
rect 41691 599726 41757 599727
rect 41691 599662 41692 599726
rect 41756 599662 41757 599726
rect 41691 599661 41757 599662
rect 675203 583406 675269 583407
rect 675203 583342 675204 583406
rect 675268 583342 675269 583406
rect 675203 583341 675269 583342
rect 675206 581775 675266 583341
rect 675203 581774 675269 581775
rect 675203 581710 675204 581774
rect 675268 581710 675269 581774
rect 675203 581709 675269 581710
rect 675206 579735 675266 581709
rect 675203 579734 675269 579735
rect 675203 579670 675204 579734
rect 675268 579670 675269 579734
rect 675203 579669 675269 579670
rect 677414 573207 677474 915589
rect 677411 573206 677477 573207
rect 677411 573142 677412 573206
rect 677476 573142 677477 573206
rect 677411 573141 677477 573142
rect 41507 571030 41573 571031
rect 41507 570966 41508 571030
rect 41572 570966 41573 571030
rect 41507 570965 41573 570966
rect 41510 569089 41570 570965
rect 41691 570486 41757 570487
rect 41691 570422 41692 570486
rect 41756 570422 41757 570486
rect 41691 570421 41757 570422
rect 41507 569088 41573 569089
rect 41507 569024 41508 569088
rect 41572 569024 41573 569088
rect 41507 569023 41573 569024
rect 41694 563415 41754 570421
rect 42059 569088 42125 569089
rect 42059 569024 42060 569088
rect 42124 569024 42125 569088
rect 42059 569023 42125 569024
rect 41691 563414 41757 563415
rect 41691 563350 41692 563414
rect 41756 563350 41757 563414
rect 41691 563349 41757 563350
rect 41691 558110 41757 558111
rect 41691 558046 41692 558110
rect 41756 558046 41757 558110
rect 41691 558045 41757 558046
rect 41694 555391 41754 558045
rect 41875 557974 41941 557975
rect 41875 557910 41876 557974
rect 41940 557910 41941 557974
rect 41875 557909 41941 557910
rect 41691 555390 41757 555391
rect 41691 555326 41692 555390
rect 41756 555326 41757 555390
rect 41691 555325 41757 555326
rect 41878 555255 41938 557909
rect 42062 557839 42122 569023
rect 42059 557838 42125 557839
rect 42059 557774 42060 557838
rect 42124 557774 42125 557838
rect 42059 557773 42125 557774
rect 41875 555254 41941 555255
rect 41875 555190 41876 555254
rect 41940 555190 41941 555254
rect 41875 555189 41941 555190
rect 677411 550086 677477 550087
rect 677411 550022 677412 550086
rect 677476 550022 677477 550086
rect 677411 550021 677477 550022
rect 42059 526558 42125 526559
rect 42059 526494 42060 526558
rect 42124 526494 42125 526558
rect 42059 526493 42125 526494
rect 41507 526328 41573 526329
rect 41507 526264 41508 526328
rect 41572 526264 41573 526328
rect 41507 526263 41573 526264
rect 41510 518325 41570 526263
rect 41875 519078 41941 519079
rect 41875 519014 41876 519078
rect 41940 519014 41941 519078
rect 41875 519013 41941 519014
rect 41507 518324 41573 518325
rect 41507 518260 41508 518324
rect 41572 518260 41573 518324
rect 41507 518259 41573 518260
rect 41878 514001 41938 519013
rect 41875 514000 41941 514001
rect 41875 513936 41876 514000
rect 41940 513936 41941 514000
rect 41875 513935 41941 513936
rect 41507 513366 41573 513367
rect 41507 513302 41508 513366
rect 41572 513302 41573 513366
rect 41507 513301 41573 513302
rect 41510 510783 41570 513301
rect 41878 510783 41938 513935
rect 42062 513367 42122 526493
rect 42059 513366 42125 513367
rect 42059 513302 42060 513366
rect 42124 513302 42125 513366
rect 42059 513301 42125 513302
rect 41507 510782 41573 510783
rect 41507 510718 41508 510782
rect 41572 510718 41573 510782
rect 41507 510717 41573 510718
rect 41875 510782 41941 510783
rect 41875 510718 41876 510782
rect 41940 510718 41941 510782
rect 41875 510717 41941 510718
rect 677414 459919 677474 550021
rect 677411 459918 677477 459919
rect 677411 459854 677412 459918
rect 677476 459854 677477 459918
rect 677411 459853 677477 459854
rect 39851 437886 39917 437887
rect 39851 437822 39852 437886
rect 39916 437822 39917 437886
rect 39851 437821 39917 437822
rect 674835 428910 674901 428911
rect 674835 428846 674836 428910
rect 674900 428846 674901 428910
rect 674835 428845 674901 428846
rect 674838 425103 674898 428845
rect 674835 425102 674901 425103
rect 674835 425038 674836 425102
rect 674900 425038 674901 425102
rect 674835 425037 674901 425038
rect 41507 381756 41573 381757
rect 41507 381692 41508 381756
rect 41572 381692 41573 381756
rect 41507 381691 41573 381692
rect 41510 379271 41570 381691
rect 41507 379270 41573 379271
rect 41507 379206 41508 379270
rect 41572 379206 41573 379270
rect 41507 379205 41573 379206
rect 675203 319022 675269 319023
rect 675203 318958 675204 319022
rect 675268 318958 675269 319022
rect 675203 318957 675269 318958
rect 675206 316513 675266 318957
rect 675203 316512 675269 316513
rect 675203 316448 675204 316512
rect 675268 316448 675269 316512
rect 675203 316447 675269 316448
rect 675755 316512 675821 316513
rect 675755 316448 675756 316512
rect 675820 316448 675821 316512
rect 675755 316447 675821 316448
rect 675758 315892 675818 316447
rect 675758 315832 676002 315892
rect 41691 305830 41757 305831
rect 41691 305766 41692 305830
rect 41756 305766 41757 305830
rect 41691 305765 41757 305766
rect 41694 297671 41754 305765
rect 41691 297670 41757 297671
rect 41691 297606 41692 297670
rect 41756 297606 41757 297670
rect 41691 297605 41757 297606
rect 41507 293400 41573 293401
rect 41507 293336 41508 293400
rect 41572 293336 41573 293400
rect 41507 293335 41573 293336
rect 41510 287199 41570 293335
rect 41691 292774 41757 292775
rect 41691 292710 41692 292774
rect 41756 292710 41757 292774
rect 41691 292709 41757 292710
rect 41694 290191 41754 292709
rect 41691 290190 41757 290191
rect 41691 290126 41692 290190
rect 41756 290126 41757 290190
rect 41691 290125 41757 290126
rect 41507 287198 41573 287199
rect 41507 287134 41508 287198
rect 41572 287134 41573 287198
rect 41507 287133 41573 287134
rect 675942 271151 676002 315832
rect 675939 271150 676005 271151
rect 675939 271086 675940 271150
rect 676004 271086 676005 271150
rect 675939 271085 676005 271086
rect 41691 248166 41757 248167
rect 41691 248102 41692 248166
rect 41756 248102 41757 248166
rect 41691 248101 41757 248102
rect 41694 245583 41754 248101
rect 41691 245582 41757 245583
rect 41691 245518 41692 245582
rect 41756 245518 41757 245582
rect 41691 245517 41757 245518
rect 41691 216750 41757 216751
rect 41691 216686 41692 216750
rect 41756 216686 41757 216750
rect 41691 216685 41757 216686
rect 41694 215119 41754 216685
rect 41691 215118 41757 215119
rect 41691 215054 41692 215118
rect 41756 215054 41757 215118
rect 41691 215053 41757 215054
rect 41691 214166 41757 214167
rect 41691 214102 41692 214166
rect 41756 214102 41757 214166
rect 41691 214101 41757 214102
rect 41694 209679 41754 214101
rect 41691 209678 41757 209679
rect 41691 209614 41692 209678
rect 41756 209614 41757 209678
rect 41691 209613 41757 209614
rect 41507 209270 41573 209271
rect 41507 209206 41508 209270
rect 41572 209206 41573 209270
rect 41507 209205 41573 209206
rect 41510 204201 41570 209205
rect 41507 204200 41573 204201
rect 41507 204136 41508 204200
rect 41572 204136 41573 204200
rect 41507 204135 41573 204136
rect 41510 200975 41570 204135
rect 41507 200974 41573 200975
rect 41507 200910 41508 200974
rect 41572 200910 41573 200974
rect 41507 200909 41573 200910
rect 41691 172278 41757 172279
rect 41691 172214 41692 172278
rect 41756 172214 41757 172278
rect 41691 172213 41757 172214
rect 41694 170289 41754 172213
rect 41691 170288 41757 170289
rect 41691 170224 41692 170288
rect 41756 170224 41757 170288
rect 41691 170223 41757 170224
rect 675203 130312 675269 130313
rect 675203 130248 675204 130312
rect 675268 130248 675269 130312
rect 675203 130247 675269 130248
rect 675206 119783 675266 130247
rect 675203 119782 675269 119783
rect 675203 119718 675204 119782
rect 675268 119718 675269 119782
rect 675203 119717 675269 119718
use sky130_ef_io__corner_pad  mgmt_corner[0] /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform -1 0 39864 0 -1 40802
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_170 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform -1 0 43864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_346
timestamp 1605708945
transform 0 -1 39457 1 0 40802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_171
timestamp 1605708945
transform -1 0 47864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_172
timestamp 1605708945
transform -1 0 51864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_173
timestamp 1605708945
transform -1 0 55864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_174
timestamp 1605708945
transform -1 0 59864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_175
timestamp 1605708945
transform -1 0 63864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_176
timestamp 1605708945
transform -1 0 67864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_177
timestamp 1605708945
transform -1 0 71864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_178
timestamp 1605708945
transform -1 0 75864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  mgmt_vssa_hvclamp_pad /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform -1 0 93664 0 -1 39595
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_179 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform -1 0 77864 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_180 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform -1 0 78064 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_181
timestamp 1605708945
transform -1 0 78264 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_182
timestamp 1605708945
transform -1 0 78464 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_183
timestamp 1605708945
transform -1 0 78664 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_185
timestamp 1605708945
transform -1 0 97664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_186
timestamp 1605708945
transform -1 0 101664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_187
timestamp 1605708945
transform -1 0 105664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_188
timestamp 1605708945
transform -1 0 109664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_189
timestamp 1605708945
transform -1 0 113664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_190
timestamp 1605708945
transform -1 0 117664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_191
timestamp 1605708945
transform -1 0 121664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_192
timestamp 1605708945
transform -1 0 125664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_193
timestamp 1605708945
transform -1 0 129664 0 -1 39595
box 0 0 4000 39593
use sky130_fd_io__top_xres4v2  resetb_pad /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform -1 0 147464 0 -1 40002
box -103 0 15124 40000
use sky130_ef_io__com_bus_slice_10um  FILLER_194
timestamp 1605708945
transform -1 0 131664 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_195
timestamp 1605708945
transform -1 0 131864 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_196
timestamp 1605708945
transform -1 0 132064 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_197
timestamp 1605708945
transform -1 0 132264 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_198
timestamp 1605708945
transform -1 0 132464 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_200
timestamp 1605708945
transform -1 0 151464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_201
timestamp 1605708945
transform -1 0 155464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_202
timestamp 1605708945
transform -1 0 159464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_203
timestamp 1605708945
transform -1 0 163464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_204
timestamp 1605708945
transform -1 0 167464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_205
timestamp 1605708945
transform -1 0 171464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_206
timestamp 1605708945
transform -1 0 175464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_207
timestamp 1605708945
transform -1 0 179464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_208
timestamp 1605708945
transform -1 0 183464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_209
timestamp 1605708945
transform -1 0 185464 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad /home/xrex/usr/devel/pdks/sky130A/libs.tech/openlane/custom_cells/mag
timestamp 1605708945
transform -1 0 202265 0 -1 42194
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_210
timestamp 1605708945
transform -1 0 185664 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_211
timestamp 1605708945
transform -1 0 185864 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_212
timestamp 1605708945
transform -1 0 186064 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_213
timestamp 1605708945
transform -1 0 186264 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_215
timestamp 1605708945
transform -1 0 206264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_216
timestamp 1605708945
transform -1 0 210264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_217
timestamp 1605708945
transform -1 0 214264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_218
timestamp 1605708945
transform -1 0 218264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_219
timestamp 1605708945
transform -1 0 222264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_220
timestamp 1605708945
transform -1 0 226264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_221
timestamp 1605708945
transform -1 0 230264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_222
timestamp 1605708945
transform -1 0 234264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_223
timestamp 1605708945
transform -1 0 238264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_224
timestamp 1605708945
transform -1 0 240264 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_225
timestamp 1605708945
transform -1 0 240464 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_226
timestamp 1605708945
transform -1 0 240664 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_227
timestamp 1605708945
transform -1 0 240864 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__vssd_lvc_pad  mgmt_vssd_lvclmap_pad /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform -1 0 256064 0 -1 39595
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_228
timestamp 1605708945
transform -1 0 241064 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_230
timestamp 1605708945
transform -1 0 260064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_231
timestamp 1605708945
transform -1 0 264064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_232
timestamp 1605708945
transform -1 0 268064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_233
timestamp 1605708945
transform -1 0 272064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_234
timestamp 1605708945
transform -1 0 276064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_235
timestamp 1605708945
transform -1 0 280064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_236
timestamp 1605708945
transform -1 0 284064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_237
timestamp 1605708945
transform -1 0 288064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1605708945
transform -1 0 310865 0 -1 42194
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_238
timestamp 1605708945
transform -1 0 292064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_239
timestamp 1605708945
transform -1 0 294064 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_240
timestamp 1605708945
transform -1 0 294264 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_241
timestamp 1605708945
transform -1 0 294464 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_242
timestamp 1605708945
transform -1 0 294664 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_243
timestamp 1605708945
transform -1 0 294864 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_245
timestamp 1605708945
transform -1 0 314864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_246
timestamp 1605708945
transform -1 0 318864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_247
timestamp 1605708945
transform -1 0 322864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_248
timestamp 1605708945
transform -1 0 326864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_249
timestamp 1605708945
transform -1 0 330864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_250
timestamp 1605708945
transform -1 0 334864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_251
timestamp 1605708945
transform -1 0 338864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1605708945
transform -1 0 365665 0 -1 42194
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_252
timestamp 1605708945
transform -1 0 342864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_253
timestamp 1605708945
transform -1 0 346864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_254
timestamp 1605708945
transform -1 0 348864 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_255
timestamp 1605708945
transform -1 0 349064 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_256
timestamp 1605708945
transform -1 0 349264 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_257
timestamp 1605708945
transform -1 0 349464 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_258
timestamp 1605708945
transform -1 0 349664 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_260
timestamp 1605708945
transform -1 0 369664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_261
timestamp 1605708945
transform -1 0 373664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_262
timestamp 1605708945
transform -1 0 377664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_263
timestamp 1605708945
transform -1 0 381664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_264
timestamp 1605708945
transform -1 0 385664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_265
timestamp 1605708945
transform -1 0 389664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_266
timestamp 1605708945
transform -1 0 393664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_267
timestamp 1605708945
transform -1 0 397664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1605708945
transform -1 0 420465 0 -1 42194
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_268
timestamp 1605708945
transform -1 0 401664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_269
timestamp 1605708945
transform -1 0 403664 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_270
timestamp 1605708945
transform -1 0 403864 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_271
timestamp 1605708945
transform -1 0 404064 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_272
timestamp 1605708945
transform -1 0 404264 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_273
timestamp 1605708945
transform -1 0 404464 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_275
timestamp 1605708945
transform -1 0 424464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_276
timestamp 1605708945
transform -1 0 428464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_277
timestamp 1605708945
transform -1 0 432464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_278
timestamp 1605708945
transform -1 0 436464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_279
timestamp 1605708945
transform -1 0 440464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_280
timestamp 1605708945
transform -1 0 444464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_281
timestamp 1605708945
transform -1 0 448464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_282
timestamp 1605708945
transform -1 0 452464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_283
timestamp 1605708945
transform -1 0 456464 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1605708945
transform -1 0 475265 0 -1 42194
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_284
timestamp 1605708945
transform -1 0 458464 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_285
timestamp 1605708945
transform -1 0 458664 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_286
timestamp 1605708945
transform -1 0 458864 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_287
timestamp 1605708945
transform -1 0 459064 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_288
timestamp 1605708945
transform -1 0 459264 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_290
timestamp 1605708945
transform -1 0 479264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_291
timestamp 1605708945
transform -1 0 483264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_292
timestamp 1605708945
transform -1 0 487264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_293
timestamp 1605708945
transform -1 0 491264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_294
timestamp 1605708945
transform -1 0 495264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_295
timestamp 1605708945
transform -1 0 499264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_296
timestamp 1605708945
transform -1 0 503264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_297
timestamp 1605708945
transform -1 0 507264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1605708945
transform -1 0 530065 0 -1 42194
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_298
timestamp 1605708945
transform -1 0 511264 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_299
timestamp 1605708945
transform -1 0 513264 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_300
timestamp 1605708945
transform -1 0 513464 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_301
timestamp 1605708945
transform -1 0 513664 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_302
timestamp 1605708945
transform -1 0 513864 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_303
timestamp 1605708945
transform -1 0 514064 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_305
timestamp 1605708945
transform -1 0 534064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_306
timestamp 1605708945
transform -1 0 538064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_307
timestamp 1605708945
transform -1 0 542064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_308
timestamp 1605708945
transform -1 0 546064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_309
timestamp 1605708945
transform -1 0 550064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_310
timestamp 1605708945
transform -1 0 554064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_311
timestamp 1605708945
transform -1 0 558064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_312
timestamp 1605708945
transform -1 0 562064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_313
timestamp 1605708945
transform -1 0 566064 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__vssio_hvc_pad  mgmt_vssio_hvclamp_pad[1] /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform -1 0 583864 0 -1 39595
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_314
timestamp 1605708945
transform -1 0 568064 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_315
timestamp 1605708945
transform -1 0 568264 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_316
timestamp 1605708945
transform -1 0 568464 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_317
timestamp 1605708945
transform -1 0 568664 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_318
timestamp 1605708945
transform -1 0 568864 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_320
timestamp 1605708945
transform -1 0 587864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_321
timestamp 1605708945
transform -1 0 591864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_322
timestamp 1605708945
transform -1 0 595864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_323
timestamp 1605708945
transform -1 0 599864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_324
timestamp 1605708945
transform -1 0 603864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_325
timestamp 1605708945
transform -1 0 607864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_326
timestamp 1605708945
transform -1 0 611864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_327
timestamp 1605708945
transform -1 0 615864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_328
timestamp 1605708945
transform -1 0 619864 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_329
timestamp 1605708945
transform -1 0 621864 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__vdda_hvc_pad  mgmt_vdda_hvclamp_pad /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform -1 0 637664 0 -1 39595
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_330
timestamp 1605708945
transform -1 0 622064 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_331
timestamp 1605708945
transform -1 0 622264 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_332
timestamp 1605708945
transform -1 0 622464 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_333
timestamp 1605708945
transform -1 0 622664 0 -1 39595
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_335
timestamp 1605708945
transform -1 0 641664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_336
timestamp 1605708945
transform -1 0 645664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_337
timestamp 1605708945
transform -1 0 649664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_338
timestamp 1605708945
transform -1 0 653664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_339
timestamp 1605708945
transform -1 0 657664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_340
timestamp 1605708945
transform -1 0 661664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_341
timestamp 1605708945
transform -1 0 665664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_342
timestamp 1605708945
transform -1 0 669664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_343
timestamp 1605708945
transform -1 0 673664 0 -1 39595
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_344
timestamp 1605708945
transform -1 0 675664 0 -1 39595
box 0 0 2000 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1605708945
transform 0 1 676664 -1 0 40002
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_5um  FILLER_345 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform -1 0 676664 0 -1 39595
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_580
timestamp 1605708945
transform 0 1 677871 -1 0 44002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_347
timestamp 1605708945
transform 0 -1 39457 1 0 44802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_348
timestamp 1605708945
transform 0 -1 39457 1 0 48802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_349
timestamp 1605708945
transform 0 -1 39457 1 0 52802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_350
timestamp 1605708945
transform 0 -1 39457 1 0 56802
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  mgmt_vccd_lvclamp_pad /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform 0 -1 39457 1 0 69202
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_351
timestamp 1605708945
transform 0 -1 39457 1 0 60802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_352
timestamp 1605708945
transform 0 -1 39457 1 0 64802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_353
timestamp 1605708945
transform 0 -1 39457 1 0 68802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_354
timestamp 1605708945
transform 0 -1 39457 1 0 69002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_356
timestamp 1605708945
transform 0 -1 39457 1 0 84202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_581
timestamp 1605708945
transform 0 1 677871 -1 0 48002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_582
timestamp 1605708945
transform 0 1 677871 -1 0 52002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_583
timestamp 1605708945
transform 0 1 677871 -1 0 56002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_584
timestamp 1605708945
transform 0 1 677871 -1 0 60002
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[0]
timestamp 1605708945
transform 0 1 675272 -1 0 86403
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1605708945
transform 0 1 677871 -1 0 64002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1605708945
transform 0 1 677871 -1 0 68002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_587
timestamp 1605708945
transform 0 1 677871 -1 0 70002
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_588
timestamp 1605708945
transform 0 1 677871 -1 0 70202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_589
timestamp 1605708945
transform 0 1 677871 -1 0 70402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_357
timestamp 1605708945
transform 0 -1 39457 1 0 88202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_358
timestamp 1605708945
transform 0 -1 39457 1 0 92202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_359
timestamp 1605708945
transform 0 -1 39457 1 0 96202
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_pad  mgmt_vddio_hvclamp_pad[0] /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605708945
transform 0 -1 39457 1 0 112802
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_360
timestamp 1605708945
transform 0 -1 39457 1 0 100202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_361
timestamp 1605708945
transform 0 -1 39457 1 0 104202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_362
timestamp 1605708945
transform 0 -1 39457 1 0 108202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_363
timestamp 1605708945
transform 0 -1 39457 1 0 112202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_364
timestamp 1605708945
transform 0 -1 39457 1 0 112402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_365
timestamp 1605708945
transform 0 -1 39457 1 0 112602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_591
timestamp 1605708945
transform 0 1 677871 -1 0 90402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_592
timestamp 1605708945
transform 0 1 677871 -1 0 94402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_593
timestamp 1605708945
transform 0 1 677871 -1 0 98402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_594
timestamp 1605708945
transform 0 1 677871 -1 0 102402
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[1]
timestamp 1605708945
transform 0 1 675272 -1 0 133003
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1605708945
transform 0 1 677871 -1 0 106402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1605708945
transform 0 1 677871 -1 0 110402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_597
timestamp 1605708945
transform 0 1 677871 -1 0 114402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_598
timestamp 1605708945
transform 0 1 677871 -1 0 116402
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_599
timestamp 1605708945
transform 0 1 677871 -1 0 116602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_600
timestamp 1605708945
transform 0 1 677871 -1 0 116802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_601
timestamp 1605708945
transform 0 1 677871 -1 0 117002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_367
timestamp 1605708945
transform 0 -1 39457 1 0 127802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_368
timestamp 1605708945
transform 0 -1 39457 1 0 131802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_369
timestamp 1605708945
transform 0 -1 39457 1 0 135802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_370
timestamp 1605708945
transform 0 -1 39457 1 0 139802
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[19]
timestamp 1605708945
transform 0 -1 42056 1 0 156401
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_371
timestamp 1605708945
transform 0 -1 39457 1 0 143802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_372
timestamp 1605708945
transform 0 -1 39457 1 0 147802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_373
timestamp 1605708945
transform 0 -1 39457 1 0 151802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_374
timestamp 1605708945
transform 0 -1 39457 1 0 155802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_375
timestamp 1605708945
transform 0 -1 39457 1 0 156002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_376
timestamp 1605708945
transform 0 -1 39457 1 0 156202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_603
timestamp 1605708945
transform 0 1 677871 -1 0 137002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_604
timestamp 1605708945
transform 0 1 677871 -1 0 141002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1605708945
transform 0 1 677871 -1 0 145002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_606
timestamp 1605708945
transform 0 1 677871 -1 0 149002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_607
timestamp 1605708945
transform 0 1 677871 -1 0 153002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_608
timestamp 1605708945
transform 0 1 677871 -1 0 157002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_609
timestamp 1605708945
transform 0 1 677871 -1 0 161002
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[2]
timestamp 1605708945
transform 0 1 675272 -1 0 179603
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_610
timestamp 1605708945
transform 0 1 677871 -1 0 163002
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_611
timestamp 1605708945
transform 0 1 677871 -1 0 163202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_612
timestamp 1605708945
transform 0 1 677871 -1 0 163402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_613
timestamp 1605708945
transform 0 1 677871 -1 0 163602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_378
timestamp 1605708945
transform 0 -1 39457 1 0 172402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_379
timestamp 1605708945
transform 0 -1 39457 1 0 176402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_380
timestamp 1605708945
transform 0 -1 39457 1 0 180402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_381
timestamp 1605708945
transform 0 -1 39457 1 0 184402
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[18]
timestamp 1605708945
transform 0 -1 42056 1 0 200801
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_382
timestamp 1605708945
transform 0 -1 39457 1 0 188402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_383
timestamp 1605708945
transform 0 -1 39457 1 0 192402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1605708945
transform 0 -1 39457 1 0 196402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_385
timestamp 1605708945
transform 0 -1 39457 1 0 200402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_386
timestamp 1605708945
transform 0 -1 39457 1 0 200602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1605708945
transform 0 1 677871 -1 0 183602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_616
timestamp 1605708945
transform 0 1 677871 -1 0 187602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_617
timestamp 1605708945
transform 0 1 677871 -1 0 191602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1605708945
transform 0 1 677871 -1 0 195602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_619
timestamp 1605708945
transform 0 1 677871 -1 0 199602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_620
timestamp 1605708945
transform 0 1 677871 -1 0 203602
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[3]
timestamp 1605708945
transform 0 1 675272 -1 0 226203
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_621
timestamp 1605708945
transform 0 1 677871 -1 0 207602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_622
timestamp 1605708945
transform 0 1 677871 -1 0 209602
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_623
timestamp 1605708945
transform 0 1 677871 -1 0 209802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_624
timestamp 1605708945
transform 0 1 677871 -1 0 210002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_625
timestamp 1605708945
transform 0 1 677871 -1 0 210202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_388
timestamp 1605708945
transform 0 -1 39457 1 0 216802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_389
timestamp 1605708945
transform 0 -1 39457 1 0 220802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_390
timestamp 1605708945
transform 0 -1 39457 1 0 224802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_391
timestamp 1605708945
transform 0 -1 39457 1 0 228802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_392
timestamp 1605708945
transform 0 -1 39457 1 0 232802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_393
timestamp 1605708945
transform 0 -1 39457 1 0 236802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1605708945
transform 0 -1 39457 1 0 240802
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[17]
timestamp 1605708945
transform 0 -1 42056 1 0 245401
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_395
timestamp 1605708945
transform 0 -1 39457 1 0 244802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_396
timestamp 1605708945
transform 0 -1 39457 1 0 245002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_397
timestamp 1605708945
transform 0 -1 39457 1 0 245202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_627
timestamp 1605708945
transform 0 1 677871 -1 0 230202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1605708945
transform 0 1 677871 -1 0 234202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_629
timestamp 1605708945
transform 0 1 677871 -1 0 238202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_630
timestamp 1605708945
transform 0 1 677871 -1 0 242202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_631
timestamp 1605708945
transform 0 1 677871 -1 0 246202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_632
timestamp 1605708945
transform 0 1 677871 -1 0 250202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_633
timestamp 1605708945
transform 0 1 677871 -1 0 254202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_399
timestamp 1605708945
transform 0 -1 39457 1 0 261402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_400
timestamp 1605708945
transform 0 -1 39457 1 0 265402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_401
timestamp 1605708945
transform 0 -1 39457 1 0 269402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_402
timestamp 1605708945
transform 0 -1 39457 1 0 273402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_403
timestamp 1605708945
transform 0 -1 39457 1 0 277402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_404
timestamp 1605708945
transform 0 -1 39457 1 0 281402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1605708945
transform 0 -1 39457 1 0 285402
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[16]
timestamp 1605708945
transform 0 -1 42056 1 0 290001
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_406
timestamp 1605708945
transform 0 -1 39457 1 0 289402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_407
timestamp 1605708945
transform 0 -1 39457 1 0 289602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_408
timestamp 1605708945
transform 0 -1 39457 1 0 289802
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[4]
timestamp 1605708945
transform 0 1 675272 -1 0 272803
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_634
timestamp 1605708945
transform 0 1 677871 -1 0 256202
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_635
timestamp 1605708945
transform 0 1 677871 -1 0 256402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_636
timestamp 1605708945
transform 0 1 677871 -1 0 256602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_637
timestamp 1605708945
transform 0 1 677871 -1 0 256802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_639
timestamp 1605708945
transform 0 1 677871 -1 0 276802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_640
timestamp 1605708945
transform 0 1 677871 -1 0 280802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_641
timestamp 1605708945
transform 0 1 677871 -1 0 284802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_642
timestamp 1605708945
transform 0 1 677871 -1 0 288802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1605708945
transform 0 1 677871 -1 0 292802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_644
timestamp 1605708945
transform 0 1 677871 -1 0 296802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_410
timestamp 1605708945
transform 0 -1 39457 1 0 306002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_411
timestamp 1605708945
transform 0 -1 39457 1 0 310002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_412
timestamp 1605708945
transform 0 -1 39457 1 0 314002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_413
timestamp 1605708945
transform 0 -1 39457 1 0 318002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_414
timestamp 1605708945
transform 0 -1 39457 1 0 322002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1605708945
transform 0 -1 39457 1 0 326002
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[15]
timestamp 1605708945
transform 0 -1 42056 1 0 334401
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1605708945
transform 0 -1 39457 1 0 330002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_417
timestamp 1605708945
transform 0 -1 39457 1 0 334002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_418
timestamp 1605708945
transform 0 -1 39457 1 0 334202
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[5]
timestamp 1605708945
transform 0 1 675272 -1 0 319203
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_645
timestamp 1605708945
transform 0 1 677871 -1 0 300802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_646
timestamp 1605708945
transform 0 1 677871 -1 0 302802
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_647
timestamp 1605708945
transform 0 1 677871 -1 0 303002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_648
timestamp 1605708945
transform 0 1 677871 -1 0 303202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_650
timestamp 1605708945
transform 0 1 677871 -1 0 323202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_651
timestamp 1605708945
transform 0 1 677871 -1 0 327202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_652
timestamp 1605708945
transform 0 1 677871 -1 0 331202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_653
timestamp 1605708945
transform 0 1 677871 -1 0 335202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_654
timestamp 1605708945
transform 0 1 677871 -1 0 339202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_420
timestamp 1605708945
transform 0 -1 39457 1 0 350402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_421
timestamp 1605708945
transform 0 -1 39457 1 0 354402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_422
timestamp 1605708945
transform 0 -1 39457 1 0 358402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_423
timestamp 1605708945
transform 0 -1 39457 1 0 362402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_424
timestamp 1605708945
transform 0 -1 39457 1 0 366402
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[14]
timestamp 1605708945
transform 0 -1 42056 1 0 379001
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1605708945
transform 0 -1 39457 1 0 370402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1605708945
transform 0 -1 39457 1 0 374402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_427
timestamp 1605708945
transform 0 -1 39457 1 0 378402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_428
timestamp 1605708945
transform 0 -1 39457 1 0 378602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_429
timestamp 1605708945
transform 0 -1 39457 1 0 378802
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[6]
timestamp 1605708945
transform 0 1 675272 -1 0 365803
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_655
timestamp 1605708945
transform 0 1 677871 -1 0 343202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1605708945
transform 0 1 677871 -1 0 347202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_657
timestamp 1605708945
transform 0 1 677871 -1 0 349202
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_658
timestamp 1605708945
transform 0 1 677871 -1 0 349402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_659
timestamp 1605708945
transform 0 1 677871 -1 0 349602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_660
timestamp 1605708945
transform 0 1 677871 -1 0 349802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1605708945
transform 0 1 677871 -1 0 369802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_663
timestamp 1605708945
transform 0 1 677871 -1 0 373802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_664
timestamp 1605708945
transform 0 1 677871 -1 0 377802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1605708945
transform 0 1 677871 -1 0 381802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_431
timestamp 1605708945
transform 0 -1 39457 1 0 395002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_432
timestamp 1605708945
transform 0 -1 39457 1 0 399002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_433
timestamp 1605708945
transform 0 -1 39457 1 0 403002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_434
timestamp 1605708945
transform 0 -1 39457 1 0 407002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1605708945
transform 0 -1 39457 1 0 411002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1605708945
transform 0 -1 39457 1 0 415002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_437
timestamp 1605708945
transform 0 -1 39457 1 0 419002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1605708945
transform 0 1 677871 -1 0 385802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_667
timestamp 1605708945
transform 0 1 677871 -1 0 389802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_668
timestamp 1605708945
transform 0 1 677871 -1 0 393802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_669
timestamp 1605708945
transform 0 1 677871 -1 0 395802
box 0 0 2000 39593
use sky130_ef_io__vssa_hvc_pad  user1_vssa_hvclamp_pad[1]
timestamp 1605708945
transform 0 1 677871 -1 0 411402
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_670
timestamp 1605708945
transform 0 1 677871 -1 0 396002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_671
timestamp 1605708945
transform 0 1 677871 -1 0 396202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_672
timestamp 1605708945
transform 0 1 677871 -1 0 396402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_674
timestamp 1605708945
transform 0 1 677871 -1 0 415402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1605708945
transform 0 1 677871 -1 0 419402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_676
timestamp 1605708945
transform 0 1 677871 -1 0 423402
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_pad  user2_vssd_lvclmap_pad
timestamp 1605708945
transform 0 -1 39457 1 0 423602
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_438
timestamp 1605708945
transform 0 -1 39457 1 0 423002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_439
timestamp 1605708945
transform 0 -1 39457 1 0 423202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_440
timestamp 1605708945
transform 0 -1 39457 1 0 423402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_442
timestamp 1605708945
transform 0 -1 39457 1 0 438602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_443
timestamp 1605708945
transform 0 -1 39457 1 0 442602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_444
timestamp 1605708945
transform 0 -1 39457 1 0 446602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1605708945
transform 0 -1 39457 1 0 450602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1605708945
transform 0 -1 39457 1 0 454602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_447
timestamp 1605708945
transform 0 -1 39457 1 0 458602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_448
timestamp 1605708945
transform 0 -1 39457 1 0 462602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_677
timestamp 1605708945
transform 0 1 677871 -1 0 427402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_678
timestamp 1605708945
transform 0 1 677871 -1 0 431402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_679
timestamp 1605708945
transform 0 1 677871 -1 0 435402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_680
timestamp 1605708945
transform 0 1 677871 -1 0 439402
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_pad  user1_vssd_lvclmap_pad
timestamp 1605708945
transform 0 1 677871 -1 0 457002
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_681
timestamp 1605708945
transform 0 1 677871 -1 0 441402
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_682
timestamp 1605708945
transform 0 1 677871 -1 0 441602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_683
timestamp 1605708945
transform 0 1 677871 -1 0 441802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_684
timestamp 1605708945
transform 0 1 677871 -1 0 442002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_686
timestamp 1605708945
transform 0 1 677871 -1 0 461002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_687
timestamp 1605708945
transform 0 1 677871 -1 0 465002
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user2_vdda_hvclamp_pad
timestamp 1605708945
transform 0 -1 39457 1 0 467002
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_449
timestamp 1605708945
transform 0 -1 39457 1 0 466602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_450
timestamp 1605708945
transform 0 -1 39457 1 0 466802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_452
timestamp 1605708945
transform 0 -1 39457 1 0 482002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_453
timestamp 1605708945
transform 0 -1 39457 1 0 486002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_454
timestamp 1605708945
transform 0 -1 39457 1 0 490002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1605708945
transform 0 -1 39457 1 0 494002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1605708945
transform 0 -1 39457 1 0 498002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_457
timestamp 1605708945
transform 0 -1 39457 1 0 502002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_458
timestamp 1605708945
transform 0 -1 39457 1 0 506002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_688
timestamp 1605708945
transform 0 1 677871 -1 0 469002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_689
timestamp 1605708945
transform 0 1 677871 -1 0 473002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1605708945
transform 0 1 677871 -1 0 477002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_691
timestamp 1605708945
transform 0 1 677871 -1 0 481002
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user1_vdda_hvclamp_pad[1]
timestamp 1605708945
transform 0 1 677871 -1 0 502602
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_692
timestamp 1605708945
transform 0 1 677871 -1 0 485002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_693
timestamp 1605708945
transform 0 1 677871 -1 0 487002
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_694
timestamp 1605708945
transform 0 1 677871 -1 0 487202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_695
timestamp 1605708945
transform 0 1 677871 -1 0 487402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_696
timestamp 1605708945
transform 0 1 677871 -1 0 487602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_698
timestamp 1605708945
transform 0 1 677871 -1 0 506602
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[13]
timestamp 1605708945
transform 0 -1 42056 1 0 510601
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_459
timestamp 1605708945
transform 0 -1 39457 1 0 510002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_460
timestamp 1605708945
transform 0 -1 39457 1 0 510202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_461
timestamp 1605708945
transform 0 -1 39457 1 0 510402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_463
timestamp 1605708945
transform 0 -1 39457 1 0 526602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_464
timestamp 1605708945
transform 0 -1 39457 1 0 530602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1605708945
transform 0 -1 39457 1 0 534602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1605708945
transform 0 -1 39457 1 0 538602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_467
timestamp 1605708945
transform 0 -1 39457 1 0 542602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_468
timestamp 1605708945
transform 0 -1 39457 1 0 546602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_699
timestamp 1605708945
transform 0 1 677871 -1 0 510602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_700
timestamp 1605708945
transform 0 1 677871 -1 0 514602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_701
timestamp 1605708945
transform 0 1 677871 -1 0 518602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_702
timestamp 1605708945
transform 0 1 677871 -1 0 522602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1605708945
transform 0 1 677871 -1 0 526602
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[7]
timestamp 1605708945
transform 0 1 675272 -1 0 549003
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_704
timestamp 1605708945
transform 0 1 677871 -1 0 530602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_705
timestamp 1605708945
transform 0 1 677871 -1 0 532602
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_706
timestamp 1605708945
transform 0 1 677871 -1 0 532802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_707
timestamp 1605708945
transform 0 1 677871 -1 0 533002
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[12]
timestamp 1605708945
transform 0 -1 42056 1 0 555201
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_469
timestamp 1605708945
transform 0 -1 39457 1 0 550602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_470
timestamp 1605708945
transform 0 -1 39457 1 0 554602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_471
timestamp 1605708945
transform 0 -1 39457 1 0 554802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_472
timestamp 1605708945
transform 0 -1 39457 1 0 555002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_474
timestamp 1605708945
transform 0 -1 39457 1 0 571202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1605708945
transform 0 -1 39457 1 0 575202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1605708945
transform 0 -1 39457 1 0 579202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_477
timestamp 1605708945
transform 0 -1 39457 1 0 583202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_478
timestamp 1605708945
transform 0 -1 39457 1 0 587202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1605708945
transform 0 1 677871 -1 0 553002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_710
timestamp 1605708945
transform 0 1 677871 -1 0 557002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_711
timestamp 1605708945
transform 0 1 677871 -1 0 561002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1605708945
transform 0 1 677871 -1 0 565002
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[8]
timestamp 1605708945
transform 0 1 675272 -1 0 595603
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1605708945
transform 0 1 677871 -1 0 569002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_714
timestamp 1605708945
transform 0 1 677871 -1 0 573002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_715
timestamp 1605708945
transform 0 1 677871 -1 0 577002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_716
timestamp 1605708945
transform 0 1 677871 -1 0 579002
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_717
timestamp 1605708945
transform 0 1 677871 -1 0 579202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_718
timestamp 1605708945
transform 0 1 677871 -1 0 579402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_719
timestamp 1605708945
transform 0 1 677871 -1 0 579602
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[11]
timestamp 1605708945
transform 0 -1 42056 1 0 599601
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_479
timestamp 1605708945
transform 0 -1 39457 1 0 591202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_480
timestamp 1605708945
transform 0 -1 39457 1 0 595202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_481
timestamp 1605708945
transform 0 -1 39457 1 0 599202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_482
timestamp 1605708945
transform 0 -1 39457 1 0 599402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_484
timestamp 1605708945
transform 0 -1 39457 1 0 615602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1605708945
transform 0 -1 39457 1 0 619602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1605708945
transform 0 -1 39457 1 0 623602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_487
timestamp 1605708945
transform 0 -1 39457 1 0 627602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_488
timestamp 1605708945
transform 0 -1 39457 1 0 631602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_721
timestamp 1605708945
transform 0 1 677871 -1 0 599602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1605708945
transform 0 1 677871 -1 0 603602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_723
timestamp 1605708945
transform 0 1 677871 -1 0 607602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_724
timestamp 1605708945
transform 0 1 677871 -1 0 611602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_725
timestamp 1605708945
transform 0 1 677871 -1 0 615602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_726
timestamp 1605708945
transform 0 1 677871 -1 0 619602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_727
timestamp 1605708945
transform 0 1 677871 -1 0 623602
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[9]
timestamp 1605708945
transform 0 1 675272 -1 0 642203
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_728
timestamp 1605708945
transform 0 1 677871 -1 0 625602
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_729
timestamp 1605708945
transform 0 1 677871 -1 0 625802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_730
timestamp 1605708945
transform 0 1 677871 -1 0 626002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_731
timestamp 1605708945
transform 0 1 677871 -1 0 626202
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[10]
timestamp 1605708945
transform 0 -1 42056 1 0 644201
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_489
timestamp 1605708945
transform 0 -1 39457 1 0 635602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_490
timestamp 1605708945
transform 0 -1 39457 1 0 639602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_491
timestamp 1605708945
transform 0 -1 39457 1 0 643602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_492
timestamp 1605708945
transform 0 -1 39457 1 0 643802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_493
timestamp 1605708945
transform 0 -1 39457 1 0 644002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1605708945
transform 0 -1 39457 1 0 660202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1605708945
transform 0 -1 39457 1 0 664202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_497
timestamp 1605708945
transform 0 -1 39457 1 0 668202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_498
timestamp 1605708945
transform 0 -1 39457 1 0 672202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_733
timestamp 1605708945
transform 0 1 677871 -1 0 646202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_734
timestamp 1605708945
transform 0 1 677871 -1 0 650202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_735
timestamp 1605708945
transform 0 1 677871 -1 0 654202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_736
timestamp 1605708945
transform 0 1 677871 -1 0 658202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1605708945
transform 0 1 677871 -1 0 662202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_738
timestamp 1605708945
transform 0 1 677871 -1 0 666202
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[10]
timestamp 1605708945
transform 0 1 675272 -1 0 688803
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_739
timestamp 1605708945
transform 0 1 677871 -1 0 670202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_740
timestamp 1605708945
transform 0 1 677871 -1 0 672202
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_741
timestamp 1605708945
transform 0 1 677871 -1 0 672402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_742
timestamp 1605708945
transform 0 1 677871 -1 0 672602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_743
timestamp 1605708945
transform 0 1 677871 -1 0 672802
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[9]
timestamp 1605708945
transform 0 -1 42056 1 0 688801
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_499
timestamp 1605708945
transform 0 -1 39457 1 0 676202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_500
timestamp 1605708945
transform 0 -1 39457 1 0 680202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_501
timestamp 1605708945
transform 0 -1 39457 1 0 684202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_502
timestamp 1605708945
transform 0 -1 39457 1 0 688202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_503
timestamp 1605708945
transform 0 -1 39457 1 0 688402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_504
timestamp 1605708945
transform 0 -1 39457 1 0 688602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1605708945
transform 0 -1 39457 1 0 704802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_507
timestamp 1605708945
transform 0 -1 39457 1 0 708802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_508
timestamp 1605708945
transform 0 -1 39457 1 0 712802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_509
timestamp 1605708945
transform 0 -1 39457 1 0 716802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_745
timestamp 1605708945
transform 0 1 677871 -1 0 692802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_746
timestamp 1605708945
transform 0 1 677871 -1 0 696802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_747
timestamp 1605708945
transform 0 1 677871 -1 0 700802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_748
timestamp 1605708945
transform 0 1 677871 -1 0 704802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_749
timestamp 1605708945
transform 0 1 677871 -1 0 708802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1605708945
transform 0 1 677871 -1 0 712802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_751
timestamp 1605708945
transform 0 1 677871 -1 0 716802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_752
timestamp 1605708945
transform 0 1 677871 -1 0 718802
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[8]
timestamp 1605708945
transform 0 -1 42056 1 0 733201
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_510
timestamp 1605708945
transform 0 -1 39457 1 0 720802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_511
timestamp 1605708945
transform 0 -1 39457 1 0 724802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_512
timestamp 1605708945
transform 0 -1 39457 1 0 728802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_513
timestamp 1605708945
transform 0 -1 39457 1 0 732802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_514
timestamp 1605708945
transform 0 -1 39457 1 0 733002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1605708945
transform 0 -1 39457 1 0 749202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_517
timestamp 1605708945
transform 0 -1 39457 1 0 753202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_518
timestamp 1605708945
transform 0 -1 39457 1 0 757202
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[11]
timestamp 1605708945
transform 0 1 675272 -1 0 735403
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_753
timestamp 1605708945
transform 0 1 677871 -1 0 719002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_754
timestamp 1605708945
transform 0 1 677871 -1 0 719202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_755
timestamp 1605708945
transform 0 1 677871 -1 0 719402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_757
timestamp 1605708945
transform 0 1 677871 -1 0 739402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_758
timestamp 1605708945
transform 0 1 677871 -1 0 743402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1605708945
transform 0 1 677871 -1 0 747402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1605708945
transform 0 1 677871 -1 0 751402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_761
timestamp 1605708945
transform 0 1 677871 -1 0 755402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_762
timestamp 1605708945
transform 0 1 677871 -1 0 759402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_763
timestamp 1605708945
transform 0 1 677871 -1 0 763402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_519
timestamp 1605708945
transform 0 -1 39457 1 0 761202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_520
timestamp 1605708945
transform 0 -1 39457 1 0 765202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_521
timestamp 1605708945
transform 0 -1 39457 1 0 769202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_522
timestamp 1605708945
transform 0 -1 39457 1 0 773202
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[7]
timestamp 1605708945
transform 0 -1 42056 1 0 777801
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_523
timestamp 1605708945
transform 0 -1 39457 1 0 777202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_524
timestamp 1605708945
transform 0 -1 39457 1 0 777402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_525
timestamp 1605708945
transform 0 -1 39457 1 0 777602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_527
timestamp 1605708945
transform 0 -1 39457 1 0 793802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_528
timestamp 1605708945
transform 0 -1 39457 1 0 797802
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[12]
timestamp 1605708945
transform 0 1 675272 -1 0 781803
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_764
timestamp 1605708945
transform 0 1 677871 -1 0 765402
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_765
timestamp 1605708945
transform 0 1 677871 -1 0 765602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_766
timestamp 1605708945
transform 0 1 677871 -1 0 765802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_768
timestamp 1605708945
transform 0 1 677871 -1 0 785802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1605708945
transform 0 1 677871 -1 0 789802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_770
timestamp 1605708945
transform 0 1 677871 -1 0 793802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_771
timestamp 1605708945
transform 0 1 677871 -1 0 797802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_772
timestamp 1605708945
transform 0 1 677871 -1 0 801802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_529
timestamp 1605708945
transform 0 -1 39457 1 0 801802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_530
timestamp 1605708945
transform 0 -1 39457 1 0 805802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_531
timestamp 1605708945
transform 0 -1 39457 1 0 809802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_532
timestamp 1605708945
transform 0 -1 39457 1 0 813802
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user2_vssa_hvclamp_pad
timestamp 1605708945
transform 0 -1 39457 1 0 822402
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_533
timestamp 1605708945
transform 0 -1 39457 1 0 817802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_534
timestamp 1605708945
transform 0 -1 39457 1 0 821802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_535
timestamp 1605708945
transform 0 -1 39457 1 0 822002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_536
timestamp 1605708945
transform 0 -1 39457 1 0 822202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_538
timestamp 1605708945
transform 0 -1 39457 1 0 837402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_539
timestamp 1605708945
transform 0 -1 39457 1 0 841402
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user1_vdda_hvclamp_pad[0]
timestamp 1605708945
transform 0 1 677871 -1 0 827402
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_773
timestamp 1605708945
transform 0 1 677871 -1 0 805802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_774
timestamp 1605708945
transform 0 1 677871 -1 0 809802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_775
timestamp 1605708945
transform 0 1 677871 -1 0 811802
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_776
timestamp 1605708945
transform 0 1 677871 -1 0 812002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_777
timestamp 1605708945
transform 0 1 677871 -1 0 812202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_778
timestamp 1605708945
transform 0 1 677871 -1 0 812402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_780
timestamp 1605708945
transform 0 1 677871 -1 0 831402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_781
timestamp 1605708945
transform 0 1 677871 -1 0 835402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_782
timestamp 1605708945
transform 0 1 677871 -1 0 839402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_783
timestamp 1605708945
transform 0 1 677871 -1 0 843402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1605708945
transform 0 1 677871 -1 0 847402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_540
timestamp 1605708945
transform 0 -1 39457 1 0 845402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_541
timestamp 1605708945
transform 0 -1 39457 1 0 849402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_542
timestamp 1605708945
transform 0 -1 39457 1 0 853402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_543
timestamp 1605708945
transform 0 -1 39457 1 0 857402
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_pad  mgmt_vddio_hvclamp_pad[1]
timestamp 1605708945
transform 0 -1 39457 1 0 865802
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_544
timestamp 1605708945
transform 0 -1 39457 1 0 861402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_545
timestamp 1605708945
transform 0 -1 39457 1 0 865402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_546
timestamp 1605708945
transform 0 -1 39457 1 0 865602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_548
timestamp 1605708945
transform 0 -1 39457 1 0 880802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_549
timestamp 1605708945
transform 0 -1 39457 1 0 884802
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[13]
timestamp 1605708945
transform 0 1 675272 -1 0 874003
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1605708945
transform 0 1 677871 -1 0 851402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_786
timestamp 1605708945
transform 0 1 677871 -1 0 855402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_787
timestamp 1605708945
transform 0 1 677871 -1 0 857402
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_788
timestamp 1605708945
transform 0 1 677871 -1 0 857602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_789
timestamp 1605708945
transform 0 1 677871 -1 0 857802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_790
timestamp 1605708945
transform 0 1 677871 -1 0 858002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_792
timestamp 1605708945
transform 0 1 677871 -1 0 878002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_793
timestamp 1605708945
transform 0 1 677871 -1 0 882002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_794
timestamp 1605708945
transform 0 1 677871 -1 0 886002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_795
timestamp 1605708945
transform 0 1 677871 -1 0 890002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_550
timestamp 1605708945
transform 0 -1 39457 1 0 888802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_551
timestamp 1605708945
transform 0 -1 39457 1 0 892802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_552
timestamp 1605708945
transform 0 -1 39457 1 0 896802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_553
timestamp 1605708945
transform 0 -1 39457 1 0 900802
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  user2_vccd_lvclamp_pad
timestamp 1605708945
transform 0 -1 39457 1 0 909402
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_554
timestamp 1605708945
transform 0 -1 39457 1 0 904802
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_555
timestamp 1605708945
transform 0 -1 39457 1 0 908802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_556
timestamp 1605708945
transform 0 -1 39457 1 0 909002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_557
timestamp 1605708945
transform 0 -1 39457 1 0 909202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_559
timestamp 1605708945
transform 0 -1 39457 1 0 924402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_796
timestamp 1605708945
transform 0 1 677871 -1 0 894002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_797
timestamp 1605708945
transform 0 1 677871 -1 0 898002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_798
timestamp 1605708945
transform 0 1 677871 -1 0 902002
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  user1_vccd_lvclamp_pad
timestamp 1605708945
transform 0 1 677871 -1 0 919602
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_799
timestamp 1605708945
transform 0 1 677871 -1 0 904002
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_800
timestamp 1605708945
transform 0 1 677871 -1 0 904202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_801
timestamp 1605708945
transform 0 1 677871 -1 0 904402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_802
timestamp 1605708945
transform 0 1 677871 -1 0 904602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_804
timestamp 1605708945
transform 0 1 677871 -1 0 923602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_805
timestamp 1605708945
transform 0 1 677871 -1 0 927602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_806
timestamp 1605708945
transform 0 1 677871 -1 0 931602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_560
timestamp 1605708945
transform 0 -1 39457 1 0 928402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_561
timestamp 1605708945
transform 0 -1 39457 1 0 932402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_562
timestamp 1605708945
transform 0 -1 39457 1 0 936402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_563
timestamp 1605708945
transform 0 -1 39457 1 0 940402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_564
timestamp 1605708945
transform 0 -1 39457 1 0 944402
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[6]
timestamp 1605708945
transform 0 -1 42056 1 0 953001
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1605708945
transform 0 -1 39457 1 0 948402
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_566
timestamp 1605708945
transform 0 -1 39457 1 0 952402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_567
timestamp 1605708945
transform 0 -1 39457 1 0 952602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_568
timestamp 1605708945
transform 0 -1 39457 1 0 952802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_570
timestamp 1605708945
transform 0 -1 39457 1 0 969002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_807
timestamp 1605708945
transform 0 1 677871 -1 0 935602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_808
timestamp 1605708945
transform 0 1 677871 -1 0 939602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_809
timestamp 1605708945
transform 0 1 677871 -1 0 943602
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_810
timestamp 1605708945
transform 0 1 677871 -1 0 947602
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[14]
timestamp 1605708945
transform 0 1 675272 -1 0 966203
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_811
timestamp 1605708945
transform 0 1 677871 -1 0 949602
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_812
timestamp 1605708945
transform 0 1 677871 -1 0 949802
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_813
timestamp 1605708945
transform 0 1 677871 -1 0 950002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_814
timestamp 1605708945
transform 0 1 677871 -1 0 950202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_816
timestamp 1605708945
transform 0 1 677871 -1 0 970202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_817
timestamp 1605708945
transform 0 1 677871 -1 0 974202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_571
timestamp 1605708945
transform 0 -1 39457 1 0 973002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_572
timestamp 1605708945
transform 0 -1 39457 1 0 977002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_573
timestamp 1605708945
transform 0 -1 39457 1 0 981002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_574
timestamp 1605708945
transform 0 -1 39457 1 0 985002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1605708945
transform 0 -1 39457 1 0 989002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_576
timestamp 1605708945
transform 0 -1 39457 1 0 993002
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_577
timestamp 1605708945
transform 0 -1 39457 1 0 997002
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_578
timestamp 1605708945
transform 0 -1 39457 1 0 997202
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_579
timestamp 1605708945
transform 0 -1 39457 1 0 997402
box 0 0 200 39593
use sky130_ef_io__corner_pad  mgmt_corner[1]
timestamp 1605708945
transform 0 -1 40664 1 0 997602
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_5
timestamp 1605708945
transform 1 0 40664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1605708945
transform 1 0 44664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1605708945
transform 1 0 48664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1605708945
transform 1 0 52664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1605708945
transform 1 0 56664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1605708945
transform 1 0 60664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1605708945
transform 1 0 64664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1605708945
transform 1 0 68664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_13
timestamp 1605708945
transform 1 0 72664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[5]
timestamp 1605708945
transform 1 0 79063 0 1 995410
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_14
timestamp 1605708945
transform 1 0 76664 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15
timestamp 1605708945
transform 1 0 78664 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_16
timestamp 1605708945
transform 1 0 78864 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1605708945
transform 1 0 95064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1605708945
transform 1 0 99064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1605708945
transform 1 0 103064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1605708945
transform 1 0 107064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1605708945
transform 1 0 111064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1605708945
transform 1 0 115064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1605708945
transform 1 0 119064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1605708945
transform 1 0 123064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[4]
timestamp 1605708945
transform 1 0 133663 0 1 995410
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_26
timestamp 1605708945
transform 1 0 127064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_27
timestamp 1605708945
transform 1 0 131064 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_28
timestamp 1605708945
transform 1 0 133064 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_29
timestamp 1605708945
transform 1 0 133264 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_30
timestamp 1605708945
transform 1 0 133464 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1605708945
transform 1 0 149664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1605708945
transform 1 0 153664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1605708945
transform 1 0 157664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1605708945
transform 1 0 161664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1605708945
transform 1 0 165664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1605708945
transform 1 0 169664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_38
timestamp 1605708945
transform 1 0 173664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_39
timestamp 1605708945
transform 1 0 177664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_40
timestamp 1605708945
transform 1 0 181664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[3]
timestamp 1605708945
transform 1 0 188263 0 1 995410
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_41
timestamp 1605708945
transform 1 0 185664 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_42
timestamp 1605708945
transform 1 0 187664 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_43
timestamp 1605708945
transform 1 0 187864 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_44
timestamp 1605708945
transform 1 0 188064 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1605708945
transform 1 0 204264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_47
timestamp 1605708945
transform 1 0 208264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_48
timestamp 1605708945
transform 1 0 212264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1605708945
transform 1 0 216264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1605708945
transform 1 0 220264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1605708945
transform 1 0 224264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[2]
timestamp 1605708945
transform 1 0 242863 0 1 995410
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_52
timestamp 1605708945
transform 1 0 228264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_53
timestamp 1605708945
transform 1 0 232264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_54
timestamp 1605708945
transform 1 0 236264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_55
timestamp 1605708945
transform 1 0 240264 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_56
timestamp 1605708945
transform 1 0 242264 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_57
timestamp 1605708945
transform 1 0 242464 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_58
timestamp 1605708945
transform 1 0 242664 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1605708945
transform 1 0 258864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1605708945
transform 1 0 262864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1605708945
transform 1 0 266864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1605708945
transform 1 0 270864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1605708945
transform 1 0 274864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_65
timestamp 1605708945
transform 1 0 278864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_66
timestamp 1605708945
transform 1 0 282864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_67
timestamp 1605708945
transform 1 0 286864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_68
timestamp 1605708945
transform 1 0 290864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_69
timestamp 1605708945
transform 1 0 294864 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[1]
timestamp 1605708945
transform 1 0 297463 0 1 995410
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_70
timestamp 1605708945
transform 1 0 296864 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_71
timestamp 1605708945
transform 1 0 297064 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_72
timestamp 1605708945
transform 1 0 297264 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_74
timestamp 1605708945
transform 1 0 313464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_75
timestamp 1605708945
transform 1 0 317464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_76
timestamp 1605708945
transform 1 0 321464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_77
timestamp 1605708945
transform 1 0 325464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1605708945
transform 1 0 329464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_79
timestamp 1605708945
transform 1 0 333464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__vssio_hvc_pad  mgmt_vssio_hvclamp_pad[0]
timestamp 1605708945
transform 1 0 352064 0 1 998009
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_80
timestamp 1605708945
transform 1 0 337464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_81
timestamp 1605708945
transform 1 0 341464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_82
timestamp 1605708945
transform 1 0 345464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_83
timestamp 1605708945
transform 1 0 349464 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_84
timestamp 1605708945
transform 1 0 351464 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_85
timestamp 1605708945
transform 1 0 351664 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_86
timestamp 1605708945
transform 1 0 351864 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1605708945
transform 1 0 367064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1605708945
transform 1 0 371064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1605708945
transform 1 0 375064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1605708945
transform 1 0 379064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_92
timestamp 1605708945
transform 1 0 383064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_93
timestamp 1605708945
transform 1 0 387064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_94
timestamp 1605708945
transform 1 0 391064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_95
timestamp 1605708945
transform 1 0 395064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad[0]
timestamp 1605708945
transform 1 0 405463 0 1 995410
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_96
timestamp 1605708945
transform 1 0 399064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_97
timestamp 1605708945
transform 1 0 403064 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_98
timestamp 1605708945
transform 1 0 405064 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_99
timestamp 1605708945
transform 1 0 405264 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1605708945
transform 1 0 421464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1605708945
transform 1 0 425464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1605708945
transform 1 0 429464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1605708945
transform 1 0 433464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_105
timestamp 1605708945
transform 1 0 437464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_106
timestamp 1605708945
transform 1 0 441464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_107
timestamp 1605708945
transform 1 0 445464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_108
timestamp 1605708945
transform 1 0 449464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_109
timestamp 1605708945
transform 1 0 453464 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[17]
timestamp 1605708945
transform 1 0 460063 0 1 995410
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_110
timestamp 1605708945
transform 1 0 457464 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_111
timestamp 1605708945
transform 1 0 459464 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_112
timestamp 1605708945
transform 1 0 459664 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_113
timestamp 1605708945
transform 1 0 459864 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1605708945
transform 1 0 476064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_116
timestamp 1605708945
transform 1 0 480064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_117
timestamp 1605708945
transform 1 0 484064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_118
timestamp 1605708945
transform 1 0 488064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_119
timestamp 1605708945
transform 1 0 492064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_120
timestamp 1605708945
transform 1 0 496064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_121
timestamp 1605708945
transform 1 0 500064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_122
timestamp 1605708945
transform 1 0 504064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[16]
timestamp 1605708945
transform 1 0 514663 0 1 995410
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_123
timestamp 1605708945
transform 1 0 508064 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_124
timestamp 1605708945
transform 1 0 512064 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_125
timestamp 1605708945
transform 1 0 514064 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_126
timestamp 1605708945
transform 1 0 514264 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_127
timestamp 1605708945
transform 1 0 514464 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_129
timestamp 1605708945
transform 1 0 530664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_130
timestamp 1605708945
transform 1 0 534664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1605708945
transform 1 0 538664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_132
timestamp 1605708945
transform 1 0 542664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_133
timestamp 1605708945
transform 1 0 546664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_134
timestamp 1605708945
transform 1 0 550664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_135
timestamp 1605708945
transform 1 0 554664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_136
timestamp 1605708945
transform 1 0 558664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_137
timestamp 1605708945
transform 1 0 562664 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user1_vssa_hvclamp_pad[0]
timestamp 1605708945
transform 1 0 569264 0 1 998009
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_138
timestamp 1605708945
transform 1 0 566664 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_139
timestamp 1605708945
transform 1 0 568664 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_140
timestamp 1605708945
transform 1 0 568864 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_141
timestamp 1605708945
transform 1 0 569064 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_143
timestamp 1605708945
transform 1 0 584264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_144
timestamp 1605708945
transform 1 0 588264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_145
timestamp 1605708945
transform 1 0 592264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_146
timestamp 1605708945
transform 1 0 596264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_147
timestamp 1605708945
transform 1 0 600264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_148
timestamp 1605708945
transform 1 0 604264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad[15]
timestamp 1605708945
transform 1 0 622863 0 1 995410
box -137 0 16140 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_149
timestamp 1605708945
transform 1 0 608264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_150
timestamp 1605708945
transform 1 0 612264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_151
timestamp 1605708945
transform 1 0 616264 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_152
timestamp 1605708945
transform 1 0 620264 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_153
timestamp 1605708945
transform 1 0 622264 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_154
timestamp 1605708945
transform 1 0 622464 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_155
timestamp 1605708945
transform 1 0 622664 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_157
timestamp 1605708945
transform 1 0 638864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_158
timestamp 1605708945
transform 1 0 642864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_159
timestamp 1605708945
transform 1 0 646864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_160
timestamp 1605708945
transform 1 0 650864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_161
timestamp 1605708945
transform 1 0 654864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_162
timestamp 1605708945
transform 1 0 658864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_163
timestamp 1605708945
transform 1 0 662864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_164
timestamp 1605708945
transform 1 0 666864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_165
timestamp 1605708945
transform 1 0 670864 0 1 998009
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_166
timestamp 1605708945
transform 1 0 674864 0 1 998009
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_818
timestamp 1605708945
transform 0 1 677871 -1 0 978202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_819
timestamp 1605708945
transform 0 1 677871 -1 0 982202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_820
timestamp 1605708945
transform 0 1 677871 -1 0 986202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_821
timestamp 1605708945
transform 0 1 677871 -1 0 990202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_822
timestamp 1605708945
transform 0 1 677871 -1 0 994202
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_823
timestamp 1605708945
transform 0 1 677871 -1 0 996202
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_824
timestamp 1605708945
transform 0 1 677871 -1 0 996402
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_825
timestamp 1605708945
transform 0 1 677871 -1 0 996602
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_826
timestamp 1605708945
transform 0 1 677871 -1 0 996802
box 0 0 200 39593
use sky130_ef_io__corner_pad  user1_corner
timestamp 1605708945
transform 1 0 677464 0 1 996802
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_1um  FILLER_167
timestamp 1605708945
transform 1 0 676864 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_168
timestamp 1605708945
transform 1 0 677064 0 1 998009
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_169
timestamp 1605708945
transform 1 0 677264 0 1 998009
box 0 0 200 39593
<< properties >>
string FIXED_BBOX 1 1 16001 42193
string GDS_FILE ../gds/chip_io.gds
string GDS_END 35100088
string GDS_START 34501266
<< end >>
