magic
tech sky130A
magscale 1 2
timestamp 1624148281
<< checkpaint >>
rect -1260 -1260 718860 1038860
<< nwell >>
rect 0 969866 1211 970200
rect 0 967942 811 969866
rect 0 967284 775 967942
rect 0 967137 1082 967284
rect 0 966065 1205 967137
rect 0 962063 1241 965603
rect 0 960471 712 962063
rect 0 957279 1249 960471
rect 0 925714 34959 926068
rect 0 914174 354 925714
rect 0 913820 34959 914174
rect 0 883594 39863 883886
rect 0 883514 34377 883594
rect 0 871939 372 883514
rect 0 871567 13397 871939
rect 0 841394 39863 841686
rect 0 841314 34377 841394
rect 0 829739 372 841314
rect 0 829367 13397 829739
rect 0 800066 1211 800400
rect 0 798142 811 800066
rect 0 797484 775 798142
rect 0 797337 1082 797484
rect 0 796265 1205 797337
rect 0 792263 1241 795803
rect 0 790671 712 792263
rect 0 787479 1249 790671
rect 0 756866 1211 757200
rect 0 754942 811 756866
rect 0 754284 775 754942
rect 0 754137 1082 754284
rect 0 753065 1205 754137
rect 0 749063 1241 752603
rect 0 747471 712 749063
rect 0 744279 1249 747471
rect 0 713666 1211 714000
rect 0 711742 811 713666
rect 0 711084 775 711742
rect 0 710937 1082 711084
rect 0 709865 1205 710937
rect 0 705863 1241 709403
rect 0 704271 712 705863
rect 0 701079 1249 704271
rect 0 670466 1211 670800
rect 0 668542 811 670466
rect 0 667884 775 668542
rect 0 667737 1082 667884
rect 0 666665 1205 667737
rect 0 662663 1241 666203
rect 0 661071 712 662663
rect 0 657879 1249 661071
rect 0 627266 1211 627600
rect 0 625342 811 627266
rect 0 624684 775 625342
rect 0 624537 1082 624684
rect 0 623465 1205 624537
rect 0 619463 1241 623003
rect 0 617871 712 619463
rect 0 614679 1249 617871
rect 0 584066 1211 584400
rect 0 582142 811 584066
rect 0 581484 775 582142
rect 0 581337 1082 581484
rect 0 580265 1205 581337
rect 0 576263 1241 579803
rect 0 574671 712 576263
rect 0 571479 1249 574671
rect 0 540866 1211 541200
rect 0 538942 811 540866
rect 0 538284 775 538942
rect 0 538137 1082 538284
rect 0 537065 1205 538137
rect 0 533063 1241 536603
rect 0 531471 712 533063
rect 0 528279 1249 531471
rect 0 496794 39863 497086
rect 0 496714 34377 496794
rect 0 485139 372 496714
rect 0 484767 13397 485139
rect 0 454514 34959 454868
rect 0 442974 354 454514
rect 0 442620 34959 442974
rect 0 413266 1211 413600
rect 0 411342 811 413266
rect 0 410684 775 411342
rect 0 410537 1082 410684
rect 0 409465 1205 410537
rect 0 405463 1241 409003
rect 0 403871 712 405463
rect 0 400679 1249 403871
rect 0 370066 1211 370400
rect 0 368142 811 370066
rect 0 367484 775 368142
rect 0 367337 1082 367484
rect 0 366265 1205 367337
rect 0 362263 1241 365803
rect 0 360671 712 362263
rect 0 357479 1249 360671
rect 0 326866 1211 327200
rect 0 324942 811 326866
rect 0 324284 775 324942
rect 0 324137 1082 324284
rect 0 323065 1205 324137
rect 0 319063 1241 322603
rect 0 317471 712 319063
rect 0 314279 1249 317471
rect 0 283666 1211 284000
rect 0 281742 811 283666
rect 0 281084 775 281742
rect 0 280937 1082 281084
rect 0 279865 1205 280937
rect 0 275863 1241 279403
rect 0 274271 712 275863
rect 0 271079 1249 274271
rect 0 240466 1211 240800
rect 0 238542 811 240466
rect 0 237884 775 238542
rect 0 237737 1082 237884
rect 0 236665 1205 237737
rect 0 232663 1241 236203
rect 0 231071 712 232663
rect 0 227879 1249 231071
rect 0 197266 1211 197600
rect 0 195342 811 197266
rect 0 194684 775 195342
rect 0 194537 1082 194684
rect 0 193465 1205 194537
rect 0 189463 1241 193003
rect 0 187871 712 189463
rect 0 184679 1249 187871
rect 0 123994 39863 124286
rect 0 123914 34377 123994
rect 0 112339 372 123914
rect 0 111967 13397 112339
rect 0 81714 34959 82068
rect 0 70174 354 81714
rect 0 69820 34959 70174
<< obsli1 >>
rect 44 44 717556 1037541
<< metal1 >>
rect 145091 39934 145143 40000
<< obsm1 >>
rect 0 40056 717600 1037600
rect 0 39878 145035 40056
rect 145199 39878 717600 40056
rect 0 0 717600 39878
<< metal2 >>
rect 77049 995407 77105 995887
rect 77693 995407 77749 995887
rect 78337 995407 78393 995887
rect 80177 995407 80233 995887
rect 80729 995407 80785 995887
rect 81373 995407 81429 995887
rect 82017 995407 82073 995887
rect 82569 995407 82625 995887
rect 83213 995407 83269 995887
rect 84501 995407 84557 995887
rect 85053 995407 85109 995887
rect 85697 995407 85753 995887
rect 86341 995407 86397 995887
rect 87537 995407 87593 995887
rect 88733 995407 88789 995887
rect 89377 995407 89433 995887
rect 91217 995407 91273 995887
rect 128449 995407 128505 995887
rect 129093 995407 129149 995887
rect 129737 995407 129793 995887
rect 131577 995407 131633 995887
rect 132129 995407 132185 995887
rect 132773 995407 132829 995887
rect 133417 995407 133473 995887
rect 133969 995407 134025 995887
rect 134613 995407 134669 995887
rect 135901 995407 135957 995887
rect 136453 995407 136509 995887
rect 137097 995407 137153 995887
rect 137741 995407 137797 995887
rect 138937 995407 138993 995887
rect 140133 995407 140189 995887
rect 140777 995407 140833 995887
rect 142617 995407 142673 995887
rect 179849 995407 179905 995887
rect 180493 995407 180549 995887
rect 181137 995407 181193 995887
rect 182977 995407 183033 995887
rect 183529 995407 183585 995887
rect 184173 995407 184229 995887
rect 184817 995407 184873 995887
rect 185369 995407 185425 995887
rect 186013 995407 186069 995887
rect 187301 995407 187357 995887
rect 187853 995407 187909 995887
rect 188497 995407 188553 995887
rect 189141 995407 189197 995887
rect 190337 995407 190393 995887
rect 191533 995407 191589 995887
rect 192177 995407 192233 995887
rect 194017 995407 194073 995887
rect 231249 995407 231305 995887
rect 231893 995407 231949 995887
rect 232537 995407 232593 995887
rect 234377 995407 234433 995887
rect 234929 995407 234985 995887
rect 235573 995407 235629 995887
rect 236217 995407 236273 995887
rect 236769 995407 236825 995887
rect 237413 995407 237469 995887
rect 238701 995407 238757 995887
rect 239253 995407 239309 995887
rect 239897 995407 239953 995887
rect 240541 995407 240597 995887
rect 241737 995407 241793 995887
rect 242933 995407 242989 995887
rect 243577 995407 243633 995887
rect 245417 995407 245473 995887
rect 282849 995407 282905 995887
rect 283493 995407 283549 995887
rect 284137 995407 284193 995887
rect 285977 995407 286033 995887
rect 286529 995407 286585 995887
rect 287173 995407 287229 995887
rect 287817 995407 287873 995887
rect 288369 995407 288425 995887
rect 289013 995407 289069 995887
rect 290301 995407 290357 995887
rect 290853 995407 290909 995887
rect 291497 995407 291553 995887
rect 292141 995407 292197 995887
rect 293337 995407 293393 995887
rect 294533 995407 294589 995887
rect 295177 995407 295233 995887
rect 297017 995407 297073 995887
rect 384649 995407 384705 995887
rect 385293 995407 385349 995887
rect 385937 995407 385993 995887
rect 387777 995407 387833 995887
rect 388329 995407 388385 995887
rect 388973 995407 389029 995887
rect 389617 995407 389673 995887
rect 390169 995407 390225 995887
rect 390813 995407 390869 995887
rect 392101 995407 392157 995887
rect 392653 995407 392709 995887
rect 393297 995407 393353 995887
rect 393941 995407 393997 995887
rect 395137 995407 395193 995887
rect 396333 995407 396389 995887
rect 396977 995407 397033 995887
rect 398817 995407 398873 995887
rect 473649 995407 473705 995887
rect 474293 995407 474349 995887
rect 474937 995407 474993 995887
rect 476777 995407 476833 995887
rect 477329 995407 477385 995887
rect 477973 995407 478029 995887
rect 478617 995407 478673 995887
rect 479169 995407 479225 995887
rect 479813 995407 479869 995887
rect 481101 995407 481157 995887
rect 481653 995407 481709 995887
rect 482297 995407 482353 995887
rect 482941 995407 482997 995887
rect 484137 995407 484193 995887
rect 485333 995407 485389 995887
rect 485977 995407 486033 995887
rect 487817 995407 487873 995887
rect 525049 995407 525105 995887
rect 525693 995407 525749 995887
rect 526337 995407 526393 995887
rect 528177 995407 528233 995887
rect 528729 995407 528785 995887
rect 529373 995407 529429 995887
rect 530017 995407 530073 995887
rect 530569 995407 530625 995887
rect 531213 995407 531269 995887
rect 532501 995407 532557 995887
rect 533053 995407 533109 995887
rect 533697 995407 533753 995887
rect 534341 995407 534397 995887
rect 535537 995407 535593 995887
rect 536733 995407 536789 995887
rect 537377 995407 537433 995887
rect 539217 995407 539273 995887
rect 626849 995407 626905 995887
rect 627493 995407 627549 995887
rect 628137 995407 628193 995887
rect 629977 995407 630033 995887
rect 630529 995407 630585 995887
rect 631173 995407 631229 995887
rect 631817 995407 631873 995887
rect 632369 995407 632425 995887
rect 633013 995407 633069 995887
rect 634301 995407 634357 995887
rect 634853 995407 634909 995887
rect 635497 995407 635553 995887
rect 636141 995407 636197 995887
rect 637337 995407 637393 995887
rect 638533 995407 638589 995887
rect 639177 995407 639233 995887
rect 641017 995407 641073 995887
rect 41713 969217 42193 969273
rect 41713 967377 42193 967433
rect 41713 966733 42193 966789
rect 675407 966695 675887 966751
rect 675407 966051 675887 966107
rect 41713 965537 42193 965593
rect 675407 965407 675887 965463
rect 41713 964341 42193 964397
rect 41713 963697 42193 963753
rect 675407 963567 675887 963623
rect 41713 963053 42193 963109
rect 675407 963015 675887 963071
rect 41713 962501 42193 962557
rect 675407 962371 675887 962427
rect 675407 961727 675887 961783
rect 41713 961213 42193 961269
rect 675407 961175 675887 961231
rect 41713 960569 42193 960625
rect 675407 960531 675887 960587
rect 41713 960017 42193 960073
rect 41713 959373 42193 959429
rect 675407 959243 675887 959299
rect 41713 958729 42193 958785
rect 675407 958691 675887 958747
rect 41713 958177 42193 958233
rect 675407 958047 675887 958103
rect 675407 957403 675887 957459
rect 41713 956337 42193 956393
rect 675407 956207 675887 956263
rect 41713 955693 42193 955749
rect 41713 955049 42193 955105
rect 675407 955011 675887 955067
rect 675407 954367 675887 954423
rect 675407 952527 675887 952583
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 871975 675887 872031
rect 675407 871331 675887 871387
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675407 863327 675887 863383
rect 41713 799417 42193 799473
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 41713 791413 42193 791469
rect 41713 790769 42193 790825
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 782775 675887 782831
rect 675407 782131 675887 782187
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675407 774127 675887 774183
rect 41713 756217 42193 756273
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 41713 748213 42193 748269
rect 41713 747569 42193 747625
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 41713 743337 42193 743393
rect 675407 743295 675887 743351
rect 41713 742693 42193 742749
rect 675407 742651 675887 742707
rect 41713 742049 42193 742105
rect 675407 742007 675887 742063
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 737775 675887 737831
rect 675407 737131 675887 737187
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675407 729127 675887 729183
rect 41713 713017 42193 713073
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 41713 705013 42193 705069
rect 41713 704369 42193 704425
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 692775 675887 692831
rect 675407 692131 675887 692187
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675407 684127 675887 684183
rect 41713 669817 42193 669873
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 41713 661813 42193 661869
rect 41713 661169 42193 661225
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 647575 675887 647631
rect 675407 646931 675887 646987
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675407 638927 675887 638983
rect 41713 626617 42193 626673
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 41713 618613 42193 618669
rect 41713 617969 42193 618025
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 602575 675887 602631
rect 675407 601931 675887 601987
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675407 593927 675887 593983
rect 41713 583417 42193 583473
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 41713 575413 42193 575469
rect 41713 574769 42193 574825
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675407 557375 675887 557431
rect 675407 556731 675887 556787
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675407 548727 675887 548783
rect 41713 540217 42193 540273
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 41713 532213 42193 532269
rect 41713 531569 42193 531625
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 41713 412617 42193 412673
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 41713 404613 42193 404669
rect 41713 403969 42193 404025
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675407 380175 675887 380231
rect 675407 379531 675887 379587
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675407 371527 675887 371583
rect 41713 369417 42193 369473
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 41713 361413 42193 361469
rect 41713 360769 42193 360825
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 334975 675887 335031
rect 675407 334331 675887 334387
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 41713 326217 42193 326273
rect 675407 326327 675887 326383
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 41713 318213 42193 318269
rect 41713 317569 42193 317625
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 289975 675887 290031
rect 675407 289331 675887 289387
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 41713 283017 42193 283073
rect 675407 281327 675887 281383
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 41713 275013 42193 275069
rect 41713 274369 42193 274425
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 244975 675887 245031
rect 675407 244331 675887 244387
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 41713 239817 42193 239873
rect 675407 238167 675887 238223
rect 41713 237977 42193 238033
rect 41713 237333 42193 237389
rect 675407 236327 675887 236383
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 41713 231813 42193 231869
rect 41713 231169 42193 231225
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 199775 675887 199831
rect 675407 199131 675887 199187
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 41713 196617 42193 196673
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 41713 194777 42193 194833
rect 675407 194807 675887 194863
rect 41713 194133 42193 194189
rect 41713 192937 42193 192993
rect 675407 192967 675887 193023
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 675407 191127 675887 191183
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 41713 188613 42193 188669
rect 41713 187969 42193 188025
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 154775 675887 154831
rect 675407 154131 675887 154187
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675407 146127 675887 146183
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675407 109575 675887 109631
rect 675407 108931 675887 108987
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675407 100927 675887 100983
rect 187327 41713 187383 42193
rect 194043 41713 194099 42193
rect 302643 41713 302699 42193
rect 306967 41713 307023 42193
rect 310095 41713 310151 42193
rect 357443 41713 357499 42193
rect 361767 41713 361823 42193
rect 364895 41713 364951 42193
rect 405527 41713 405583 42193
rect 412243 41713 412299 42193
rect 416567 41713 416623 42193
rect 419695 41713 419751 42193
rect 460327 41713 460383 42193
rect 467043 41713 467099 42193
rect 471367 41713 471423 42193
rect 474495 41713 474551 42193
rect 515127 41713 515183 42193
rect 520647 41713 520703 42193
rect 521843 41713 521899 42193
rect 524971 41713 525027 42193
rect 526167 41713 526223 42193
rect 529295 41713 529351 42193
rect 141667 39934 141813 40000
rect 145091 39706 145143 40000
<< obsm2 >>
rect 0 995943 717600 1037600
rect 0 995351 76993 995943
rect 77161 995351 77637 995943
rect 77805 995351 78281 995943
rect 78449 995351 80121 995943
rect 80289 995351 80673 995943
rect 80841 995351 81317 995943
rect 81485 995351 81961 995943
rect 82129 995351 82513 995943
rect 82681 995351 83157 995943
rect 83325 995351 84445 995943
rect 84613 995351 84997 995943
rect 85165 995351 85641 995943
rect 85809 995351 86285 995943
rect 86453 995351 87481 995943
rect 87649 995351 88677 995943
rect 88845 995351 89321 995943
rect 89489 995351 91161 995943
rect 91329 995351 128393 995943
rect 128561 995351 129037 995943
rect 129205 995351 129681 995943
rect 129849 995351 131521 995943
rect 131689 995351 132073 995943
rect 132241 995351 132717 995943
rect 132885 995351 133361 995943
rect 133529 995351 133913 995943
rect 134081 995351 134557 995943
rect 134725 995351 135845 995943
rect 136013 995351 136397 995943
rect 136565 995351 137041 995943
rect 137209 995351 137685 995943
rect 137853 995351 138881 995943
rect 139049 995351 140077 995943
rect 140245 995351 140721 995943
rect 140889 995351 142561 995943
rect 142729 995351 179793 995943
rect 179961 995351 180437 995943
rect 180605 995351 181081 995943
rect 181249 995351 182921 995943
rect 183089 995351 183473 995943
rect 183641 995351 184117 995943
rect 184285 995351 184761 995943
rect 184929 995351 185313 995943
rect 185481 995351 185957 995943
rect 186125 995351 187245 995943
rect 187413 995351 187797 995943
rect 187965 995351 188441 995943
rect 188609 995351 189085 995943
rect 189253 995351 190281 995943
rect 190449 995351 191477 995943
rect 191645 995351 192121 995943
rect 192289 995351 193961 995943
rect 194129 995351 231193 995943
rect 231361 995351 231837 995943
rect 232005 995351 232481 995943
rect 232649 995351 234321 995943
rect 234489 995351 234873 995943
rect 235041 995351 235517 995943
rect 235685 995351 236161 995943
rect 236329 995351 236713 995943
rect 236881 995351 237357 995943
rect 237525 995351 238645 995943
rect 238813 995351 239197 995943
rect 239365 995351 239841 995943
rect 240009 995351 240485 995943
rect 240653 995351 241681 995943
rect 241849 995351 242877 995943
rect 243045 995351 243521 995943
rect 243689 995351 245361 995943
rect 245529 995351 282793 995943
rect 282961 995351 283437 995943
rect 283605 995351 284081 995943
rect 284249 995351 285921 995943
rect 286089 995351 286473 995943
rect 286641 995351 287117 995943
rect 287285 995351 287761 995943
rect 287929 995351 288313 995943
rect 288481 995351 288957 995943
rect 289125 995351 290245 995943
rect 290413 995351 290797 995943
rect 290965 995351 291441 995943
rect 291609 995351 292085 995943
rect 292253 995351 293281 995943
rect 293449 995351 294477 995943
rect 294645 995351 295121 995943
rect 295289 995351 296961 995943
rect 297129 995351 384593 995943
rect 384761 995351 385237 995943
rect 385405 995351 385881 995943
rect 386049 995351 387721 995943
rect 387889 995351 388273 995943
rect 388441 995351 388917 995943
rect 389085 995351 389561 995943
rect 389729 995351 390113 995943
rect 390281 995351 390757 995943
rect 390925 995351 392045 995943
rect 392213 995351 392597 995943
rect 392765 995351 393241 995943
rect 393409 995351 393885 995943
rect 394053 995351 395081 995943
rect 395249 995351 396277 995943
rect 396445 995351 396921 995943
rect 397089 995351 398761 995943
rect 398929 995351 473593 995943
rect 473761 995351 474237 995943
rect 474405 995351 474881 995943
rect 475049 995351 476721 995943
rect 476889 995351 477273 995943
rect 477441 995351 477917 995943
rect 478085 995351 478561 995943
rect 478729 995351 479113 995943
rect 479281 995351 479757 995943
rect 479925 995351 481045 995943
rect 481213 995351 481597 995943
rect 481765 995351 482241 995943
rect 482409 995351 482885 995943
rect 483053 995351 484081 995943
rect 484249 995351 485277 995943
rect 485445 995351 485921 995943
rect 486089 995351 487761 995943
rect 487929 995351 524993 995943
rect 525161 995351 525637 995943
rect 525805 995351 526281 995943
rect 526449 995351 528121 995943
rect 528289 995351 528673 995943
rect 528841 995351 529317 995943
rect 529485 995351 529961 995943
rect 530129 995351 530513 995943
rect 530681 995351 531157 995943
rect 531325 995351 532445 995943
rect 532613 995351 532997 995943
rect 533165 995351 533641 995943
rect 533809 995351 534285 995943
rect 534453 995351 535481 995943
rect 535649 995351 536677 995943
rect 536845 995351 537321 995943
rect 537489 995351 539161 995943
rect 539329 995351 626793 995943
rect 626961 995351 627437 995943
rect 627605 995351 628081 995943
rect 628249 995351 629921 995943
rect 630089 995351 630473 995943
rect 630641 995351 631117 995943
rect 631285 995351 631761 995943
rect 631929 995351 632313 995943
rect 632481 995351 632957 995943
rect 633125 995351 634245 995943
rect 634413 995351 634797 995943
rect 634965 995351 635441 995943
rect 635609 995351 636085 995943
rect 636253 995351 637281 995943
rect 637449 995351 638477 995943
rect 638645 995351 639121 995943
rect 639289 995351 640961 995943
rect 641129 995351 717600 995943
rect 0 969329 717600 995351
rect 0 969161 41657 969329
rect 42249 969161 717600 969329
rect 0 967489 717600 969161
rect 0 967321 41657 967489
rect 42249 967321 717600 967489
rect 0 966845 717600 967321
rect 0 966677 41657 966845
rect 42249 966807 717600 966845
rect 42249 966677 675351 966807
rect 0 966639 675351 966677
rect 675943 966639 717600 966807
rect 0 966163 717600 966639
rect 0 965995 675351 966163
rect 675943 965995 717600 966163
rect 0 965649 717600 965995
rect 0 965481 41657 965649
rect 42249 965519 717600 965649
rect 42249 965481 675351 965519
rect 0 965351 675351 965481
rect 675943 965351 717600 965519
rect 0 964453 717600 965351
rect 0 964285 41657 964453
rect 42249 964285 717600 964453
rect 0 963809 717600 964285
rect 0 963641 41657 963809
rect 42249 963679 717600 963809
rect 42249 963641 675351 963679
rect 0 963511 675351 963641
rect 675943 963511 717600 963679
rect 0 963165 717600 963511
rect 0 962997 41657 963165
rect 42249 963127 717600 963165
rect 42249 962997 675351 963127
rect 0 962959 675351 962997
rect 675943 962959 717600 963127
rect 0 962613 717600 962959
rect 0 962445 41657 962613
rect 42249 962483 717600 962613
rect 42249 962445 675351 962483
rect 0 962315 675351 962445
rect 675943 962315 717600 962483
rect 0 961839 717600 962315
rect 0 961671 675351 961839
rect 675943 961671 717600 961839
rect 0 961325 717600 961671
rect 0 961157 41657 961325
rect 42249 961287 717600 961325
rect 42249 961157 675351 961287
rect 0 961119 675351 961157
rect 675943 961119 717600 961287
rect 0 960681 717600 961119
rect 0 960513 41657 960681
rect 42249 960643 717600 960681
rect 42249 960513 675351 960643
rect 0 960475 675351 960513
rect 675943 960475 717600 960643
rect 0 960129 717600 960475
rect 0 959961 41657 960129
rect 42249 959961 717600 960129
rect 0 959485 717600 959961
rect 0 959317 41657 959485
rect 42249 959355 717600 959485
rect 42249 959317 675351 959355
rect 0 959187 675351 959317
rect 675943 959187 717600 959355
rect 0 958841 717600 959187
rect 0 958673 41657 958841
rect 42249 958803 717600 958841
rect 42249 958673 675351 958803
rect 0 958635 675351 958673
rect 675943 958635 717600 958803
rect 0 958289 717600 958635
rect 0 958121 41657 958289
rect 42249 958159 717600 958289
rect 42249 958121 675351 958159
rect 0 957991 675351 958121
rect 675943 957991 717600 958159
rect 0 957515 717600 957991
rect 0 957347 675351 957515
rect 675943 957347 717600 957515
rect 0 956449 717600 957347
rect 0 956281 41657 956449
rect 42249 956319 717600 956449
rect 42249 956281 675351 956319
rect 0 956151 675351 956281
rect 675943 956151 717600 956319
rect 0 955805 717600 956151
rect 0 955637 41657 955805
rect 42249 955637 717600 955805
rect 0 955161 717600 955637
rect 0 954993 41657 955161
rect 42249 955123 717600 955161
rect 42249 954993 675351 955123
rect 0 954955 675351 954993
rect 675943 954955 717600 955123
rect 0 954479 717600 954955
rect 0 954311 675351 954479
rect 675943 954311 717600 954479
rect 0 952639 717600 954311
rect 0 952471 675351 952639
rect 675943 952471 717600 952639
rect 0 877607 717600 952471
rect 0 877439 675351 877607
rect 675943 877439 717600 877607
rect 0 876963 717600 877439
rect 0 876795 675351 876963
rect 675943 876795 717600 876963
rect 0 876319 717600 876795
rect 0 876151 675351 876319
rect 675943 876151 717600 876319
rect 0 874479 717600 876151
rect 0 874311 675351 874479
rect 675943 874311 717600 874479
rect 0 873927 717600 874311
rect 0 873759 675351 873927
rect 675943 873759 717600 873927
rect 0 873283 717600 873759
rect 0 873115 675351 873283
rect 675943 873115 717600 873283
rect 0 872639 717600 873115
rect 0 872471 675351 872639
rect 675943 872471 717600 872639
rect 0 872087 717600 872471
rect 0 871919 675351 872087
rect 675943 871919 717600 872087
rect 0 871443 717600 871919
rect 0 871275 675351 871443
rect 675943 871275 717600 871443
rect 0 870155 717600 871275
rect 0 869987 675351 870155
rect 675943 869987 717600 870155
rect 0 869603 717600 869987
rect 0 869435 675351 869603
rect 675943 869435 717600 869603
rect 0 868959 717600 869435
rect 0 868791 675351 868959
rect 675943 868791 717600 868959
rect 0 868315 717600 868791
rect 0 868147 675351 868315
rect 675943 868147 717600 868315
rect 0 867119 717600 868147
rect 0 866951 675351 867119
rect 675943 866951 717600 867119
rect 0 865923 717600 866951
rect 0 865755 675351 865923
rect 675943 865755 717600 865923
rect 0 865279 717600 865755
rect 0 865111 675351 865279
rect 675943 865111 717600 865279
rect 0 863439 717600 865111
rect 0 863271 675351 863439
rect 675943 863271 717600 863439
rect 0 799529 717600 863271
rect 0 799361 41657 799529
rect 42249 799361 717600 799529
rect 0 797689 717600 799361
rect 0 797521 41657 797689
rect 42249 797521 717600 797689
rect 0 797045 717600 797521
rect 0 796877 41657 797045
rect 42249 796877 717600 797045
rect 0 795849 717600 796877
rect 0 795681 41657 795849
rect 42249 795681 717600 795849
rect 0 794653 717600 795681
rect 0 794485 41657 794653
rect 42249 794485 717600 794653
rect 0 794009 717600 794485
rect 0 793841 41657 794009
rect 42249 793841 717600 794009
rect 0 793365 717600 793841
rect 0 793197 41657 793365
rect 42249 793197 717600 793365
rect 0 792813 717600 793197
rect 0 792645 41657 792813
rect 42249 792645 717600 792813
rect 0 791525 717600 792645
rect 0 791357 41657 791525
rect 42249 791357 717600 791525
rect 0 790881 717600 791357
rect 0 790713 41657 790881
rect 42249 790713 717600 790881
rect 0 790329 717600 790713
rect 0 790161 41657 790329
rect 42249 790161 717600 790329
rect 0 789685 717600 790161
rect 0 789517 41657 789685
rect 42249 789517 717600 789685
rect 0 789041 717600 789517
rect 0 788873 41657 789041
rect 42249 788873 717600 789041
rect 0 788489 717600 788873
rect 0 788321 41657 788489
rect 42249 788407 717600 788489
rect 42249 788321 675351 788407
rect 0 788239 675351 788321
rect 675943 788239 717600 788407
rect 0 787763 717600 788239
rect 0 787595 675351 787763
rect 675943 787595 717600 787763
rect 0 787119 717600 787595
rect 0 786951 675351 787119
rect 675943 786951 717600 787119
rect 0 786649 717600 786951
rect 0 786481 41657 786649
rect 42249 786481 717600 786649
rect 0 786005 717600 786481
rect 0 785837 41657 786005
rect 42249 785837 717600 786005
rect 0 785361 717600 785837
rect 0 785193 41657 785361
rect 42249 785279 717600 785361
rect 42249 785193 675351 785279
rect 0 785111 675351 785193
rect 675943 785111 717600 785279
rect 0 784727 717600 785111
rect 0 784559 675351 784727
rect 675943 784559 717600 784727
rect 0 784083 717600 784559
rect 0 783915 675351 784083
rect 675943 783915 717600 784083
rect 0 783439 717600 783915
rect 0 783271 675351 783439
rect 675943 783271 717600 783439
rect 0 782887 717600 783271
rect 0 782719 675351 782887
rect 675943 782719 717600 782887
rect 0 782243 717600 782719
rect 0 782075 675351 782243
rect 675943 782075 717600 782243
rect 0 780955 717600 782075
rect 0 780787 675351 780955
rect 675943 780787 717600 780955
rect 0 780403 717600 780787
rect 0 780235 675351 780403
rect 675943 780235 717600 780403
rect 0 779759 717600 780235
rect 0 779591 675351 779759
rect 675943 779591 717600 779759
rect 0 779115 717600 779591
rect 0 778947 675351 779115
rect 675943 778947 717600 779115
rect 0 777919 717600 778947
rect 0 777751 675351 777919
rect 675943 777751 717600 777919
rect 0 776723 717600 777751
rect 0 776555 675351 776723
rect 675943 776555 717600 776723
rect 0 776079 717600 776555
rect 0 775911 675351 776079
rect 675943 775911 717600 776079
rect 0 774239 717600 775911
rect 0 774071 675351 774239
rect 675943 774071 717600 774239
rect 0 756329 717600 774071
rect 0 756161 41657 756329
rect 42249 756161 717600 756329
rect 0 754489 717600 756161
rect 0 754321 41657 754489
rect 42249 754321 717600 754489
rect 0 753845 717600 754321
rect 0 753677 41657 753845
rect 42249 753677 717600 753845
rect 0 752649 717600 753677
rect 0 752481 41657 752649
rect 42249 752481 717600 752649
rect 0 751453 717600 752481
rect 0 751285 41657 751453
rect 42249 751285 717600 751453
rect 0 750809 717600 751285
rect 0 750641 41657 750809
rect 42249 750641 717600 750809
rect 0 750165 717600 750641
rect 0 749997 41657 750165
rect 42249 749997 717600 750165
rect 0 749613 717600 749997
rect 0 749445 41657 749613
rect 42249 749445 717600 749613
rect 0 748325 717600 749445
rect 0 748157 41657 748325
rect 42249 748157 717600 748325
rect 0 747681 717600 748157
rect 0 747513 41657 747681
rect 42249 747513 717600 747681
rect 0 747129 717600 747513
rect 0 746961 41657 747129
rect 42249 746961 717600 747129
rect 0 746485 717600 746961
rect 0 746317 41657 746485
rect 42249 746317 717600 746485
rect 0 745841 717600 746317
rect 0 745673 41657 745841
rect 42249 745673 717600 745841
rect 0 745289 717600 745673
rect 0 745121 41657 745289
rect 42249 745121 717600 745289
rect 0 743449 717600 745121
rect 0 743281 41657 743449
rect 42249 743407 717600 743449
rect 42249 743281 675351 743407
rect 0 743239 675351 743281
rect 675943 743239 717600 743407
rect 0 742805 717600 743239
rect 0 742637 41657 742805
rect 42249 742763 717600 742805
rect 42249 742637 675351 742763
rect 0 742595 675351 742637
rect 675943 742595 717600 742763
rect 0 742161 717600 742595
rect 0 741993 41657 742161
rect 42249 742119 717600 742161
rect 42249 741993 675351 742119
rect 0 741951 675351 741993
rect 675943 741951 717600 742119
rect 0 740279 717600 741951
rect 0 740111 675351 740279
rect 675943 740111 717600 740279
rect 0 739727 717600 740111
rect 0 739559 675351 739727
rect 675943 739559 717600 739727
rect 0 739083 717600 739559
rect 0 738915 675351 739083
rect 675943 738915 717600 739083
rect 0 738439 717600 738915
rect 0 738271 675351 738439
rect 675943 738271 717600 738439
rect 0 737887 717600 738271
rect 0 737719 675351 737887
rect 675943 737719 717600 737887
rect 0 737243 717600 737719
rect 0 737075 675351 737243
rect 675943 737075 717600 737243
rect 0 735955 717600 737075
rect 0 735787 675351 735955
rect 675943 735787 717600 735955
rect 0 735403 717600 735787
rect 0 735235 675351 735403
rect 675943 735235 717600 735403
rect 0 734759 717600 735235
rect 0 734591 675351 734759
rect 675943 734591 717600 734759
rect 0 734115 717600 734591
rect 0 733947 675351 734115
rect 675943 733947 717600 734115
rect 0 732919 717600 733947
rect 0 732751 675351 732919
rect 675943 732751 717600 732919
rect 0 731723 717600 732751
rect 0 731555 675351 731723
rect 675943 731555 717600 731723
rect 0 731079 717600 731555
rect 0 730911 675351 731079
rect 675943 730911 717600 731079
rect 0 729239 717600 730911
rect 0 729071 675351 729239
rect 675943 729071 717600 729239
rect 0 713129 717600 729071
rect 0 712961 41657 713129
rect 42249 712961 717600 713129
rect 0 711289 717600 712961
rect 0 711121 41657 711289
rect 42249 711121 717600 711289
rect 0 710645 717600 711121
rect 0 710477 41657 710645
rect 42249 710477 717600 710645
rect 0 709449 717600 710477
rect 0 709281 41657 709449
rect 42249 709281 717600 709449
rect 0 708253 717600 709281
rect 0 708085 41657 708253
rect 42249 708085 717600 708253
rect 0 707609 717600 708085
rect 0 707441 41657 707609
rect 42249 707441 717600 707609
rect 0 706965 717600 707441
rect 0 706797 41657 706965
rect 42249 706797 717600 706965
rect 0 706413 717600 706797
rect 0 706245 41657 706413
rect 42249 706245 717600 706413
rect 0 705125 717600 706245
rect 0 704957 41657 705125
rect 42249 704957 717600 705125
rect 0 704481 717600 704957
rect 0 704313 41657 704481
rect 42249 704313 717600 704481
rect 0 703929 717600 704313
rect 0 703761 41657 703929
rect 42249 703761 717600 703929
rect 0 703285 717600 703761
rect 0 703117 41657 703285
rect 42249 703117 717600 703285
rect 0 702641 717600 703117
rect 0 702473 41657 702641
rect 42249 702473 717600 702641
rect 0 702089 717600 702473
rect 0 701921 41657 702089
rect 42249 701921 717600 702089
rect 0 700249 717600 701921
rect 0 700081 41657 700249
rect 42249 700081 717600 700249
rect 0 699605 717600 700081
rect 0 699437 41657 699605
rect 42249 699437 717600 699605
rect 0 698961 717600 699437
rect 0 698793 41657 698961
rect 42249 698793 717600 698961
rect 0 698407 717600 698793
rect 0 698239 675351 698407
rect 675943 698239 717600 698407
rect 0 697763 717600 698239
rect 0 697595 675351 697763
rect 675943 697595 717600 697763
rect 0 697119 717600 697595
rect 0 696951 675351 697119
rect 675943 696951 717600 697119
rect 0 695279 717600 696951
rect 0 695111 675351 695279
rect 675943 695111 717600 695279
rect 0 694727 717600 695111
rect 0 694559 675351 694727
rect 675943 694559 717600 694727
rect 0 694083 717600 694559
rect 0 693915 675351 694083
rect 675943 693915 717600 694083
rect 0 693439 717600 693915
rect 0 693271 675351 693439
rect 675943 693271 717600 693439
rect 0 692887 717600 693271
rect 0 692719 675351 692887
rect 675943 692719 717600 692887
rect 0 692243 717600 692719
rect 0 692075 675351 692243
rect 675943 692075 717600 692243
rect 0 690955 717600 692075
rect 0 690787 675351 690955
rect 675943 690787 717600 690955
rect 0 690403 717600 690787
rect 0 690235 675351 690403
rect 675943 690235 717600 690403
rect 0 689759 717600 690235
rect 0 689591 675351 689759
rect 675943 689591 717600 689759
rect 0 689115 717600 689591
rect 0 688947 675351 689115
rect 675943 688947 717600 689115
rect 0 687919 717600 688947
rect 0 687751 675351 687919
rect 675943 687751 717600 687919
rect 0 686723 717600 687751
rect 0 686555 675351 686723
rect 675943 686555 717600 686723
rect 0 686079 717600 686555
rect 0 685911 675351 686079
rect 675943 685911 717600 686079
rect 0 684239 717600 685911
rect 0 684071 675351 684239
rect 675943 684071 717600 684239
rect 0 669929 717600 684071
rect 0 669761 41657 669929
rect 42249 669761 717600 669929
rect 0 668089 717600 669761
rect 0 667921 41657 668089
rect 42249 667921 717600 668089
rect 0 667445 717600 667921
rect 0 667277 41657 667445
rect 42249 667277 717600 667445
rect 0 666249 717600 667277
rect 0 666081 41657 666249
rect 42249 666081 717600 666249
rect 0 665053 717600 666081
rect 0 664885 41657 665053
rect 42249 664885 717600 665053
rect 0 664409 717600 664885
rect 0 664241 41657 664409
rect 42249 664241 717600 664409
rect 0 663765 717600 664241
rect 0 663597 41657 663765
rect 42249 663597 717600 663765
rect 0 663213 717600 663597
rect 0 663045 41657 663213
rect 42249 663045 717600 663213
rect 0 661925 717600 663045
rect 0 661757 41657 661925
rect 42249 661757 717600 661925
rect 0 661281 717600 661757
rect 0 661113 41657 661281
rect 42249 661113 717600 661281
rect 0 660729 717600 661113
rect 0 660561 41657 660729
rect 42249 660561 717600 660729
rect 0 660085 717600 660561
rect 0 659917 41657 660085
rect 42249 659917 717600 660085
rect 0 659441 717600 659917
rect 0 659273 41657 659441
rect 42249 659273 717600 659441
rect 0 658889 717600 659273
rect 0 658721 41657 658889
rect 42249 658721 717600 658889
rect 0 657049 717600 658721
rect 0 656881 41657 657049
rect 42249 656881 717600 657049
rect 0 656405 717600 656881
rect 0 656237 41657 656405
rect 42249 656237 717600 656405
rect 0 655761 717600 656237
rect 0 655593 41657 655761
rect 42249 655593 717600 655761
rect 0 653207 717600 655593
rect 0 653039 675351 653207
rect 675943 653039 717600 653207
rect 0 652563 717600 653039
rect 0 652395 675351 652563
rect 675943 652395 717600 652563
rect 0 651919 717600 652395
rect 0 651751 675351 651919
rect 675943 651751 717600 651919
rect 0 650079 717600 651751
rect 0 649911 675351 650079
rect 675943 649911 717600 650079
rect 0 649527 717600 649911
rect 0 649359 675351 649527
rect 675943 649359 717600 649527
rect 0 648883 717600 649359
rect 0 648715 675351 648883
rect 675943 648715 717600 648883
rect 0 648239 717600 648715
rect 0 648071 675351 648239
rect 675943 648071 717600 648239
rect 0 647687 717600 648071
rect 0 647519 675351 647687
rect 675943 647519 717600 647687
rect 0 647043 717600 647519
rect 0 646875 675351 647043
rect 675943 646875 717600 647043
rect 0 645755 717600 646875
rect 0 645587 675351 645755
rect 675943 645587 717600 645755
rect 0 645203 717600 645587
rect 0 645035 675351 645203
rect 675943 645035 717600 645203
rect 0 644559 717600 645035
rect 0 644391 675351 644559
rect 675943 644391 717600 644559
rect 0 643915 717600 644391
rect 0 643747 675351 643915
rect 675943 643747 717600 643915
rect 0 642719 717600 643747
rect 0 642551 675351 642719
rect 675943 642551 717600 642719
rect 0 641523 717600 642551
rect 0 641355 675351 641523
rect 675943 641355 717600 641523
rect 0 640879 717600 641355
rect 0 640711 675351 640879
rect 675943 640711 717600 640879
rect 0 639039 717600 640711
rect 0 638871 675351 639039
rect 675943 638871 717600 639039
rect 0 626729 717600 638871
rect 0 626561 41657 626729
rect 42249 626561 717600 626729
rect 0 624889 717600 626561
rect 0 624721 41657 624889
rect 42249 624721 717600 624889
rect 0 624245 717600 624721
rect 0 624077 41657 624245
rect 42249 624077 717600 624245
rect 0 623049 717600 624077
rect 0 622881 41657 623049
rect 42249 622881 717600 623049
rect 0 621853 717600 622881
rect 0 621685 41657 621853
rect 42249 621685 717600 621853
rect 0 621209 717600 621685
rect 0 621041 41657 621209
rect 42249 621041 717600 621209
rect 0 620565 717600 621041
rect 0 620397 41657 620565
rect 42249 620397 717600 620565
rect 0 620013 717600 620397
rect 0 619845 41657 620013
rect 42249 619845 717600 620013
rect 0 618725 717600 619845
rect 0 618557 41657 618725
rect 42249 618557 717600 618725
rect 0 618081 717600 618557
rect 0 617913 41657 618081
rect 42249 617913 717600 618081
rect 0 617529 717600 617913
rect 0 617361 41657 617529
rect 42249 617361 717600 617529
rect 0 616885 717600 617361
rect 0 616717 41657 616885
rect 42249 616717 717600 616885
rect 0 616241 717600 616717
rect 0 616073 41657 616241
rect 42249 616073 717600 616241
rect 0 615689 717600 616073
rect 0 615521 41657 615689
rect 42249 615521 717600 615689
rect 0 613849 717600 615521
rect 0 613681 41657 613849
rect 42249 613681 717600 613849
rect 0 613205 717600 613681
rect 0 613037 41657 613205
rect 42249 613037 717600 613205
rect 0 612561 717600 613037
rect 0 612393 41657 612561
rect 42249 612393 717600 612561
rect 0 608207 717600 612393
rect 0 608039 675351 608207
rect 675943 608039 717600 608207
rect 0 607563 717600 608039
rect 0 607395 675351 607563
rect 675943 607395 717600 607563
rect 0 606919 717600 607395
rect 0 606751 675351 606919
rect 675943 606751 717600 606919
rect 0 605079 717600 606751
rect 0 604911 675351 605079
rect 675943 604911 717600 605079
rect 0 604527 717600 604911
rect 0 604359 675351 604527
rect 675943 604359 717600 604527
rect 0 603883 717600 604359
rect 0 603715 675351 603883
rect 675943 603715 717600 603883
rect 0 603239 717600 603715
rect 0 603071 675351 603239
rect 675943 603071 717600 603239
rect 0 602687 717600 603071
rect 0 602519 675351 602687
rect 675943 602519 717600 602687
rect 0 602043 717600 602519
rect 0 601875 675351 602043
rect 675943 601875 717600 602043
rect 0 600755 717600 601875
rect 0 600587 675351 600755
rect 675943 600587 717600 600755
rect 0 600203 717600 600587
rect 0 600035 675351 600203
rect 675943 600035 717600 600203
rect 0 599559 717600 600035
rect 0 599391 675351 599559
rect 675943 599391 717600 599559
rect 0 598915 717600 599391
rect 0 598747 675351 598915
rect 675943 598747 717600 598915
rect 0 597719 717600 598747
rect 0 597551 675351 597719
rect 675943 597551 717600 597719
rect 0 596523 717600 597551
rect 0 596355 675351 596523
rect 675943 596355 717600 596523
rect 0 595879 717600 596355
rect 0 595711 675351 595879
rect 675943 595711 717600 595879
rect 0 594039 717600 595711
rect 0 593871 675351 594039
rect 675943 593871 717600 594039
rect 0 583529 717600 593871
rect 0 583361 41657 583529
rect 42249 583361 717600 583529
rect 0 581689 717600 583361
rect 0 581521 41657 581689
rect 42249 581521 717600 581689
rect 0 581045 717600 581521
rect 0 580877 41657 581045
rect 42249 580877 717600 581045
rect 0 579849 717600 580877
rect 0 579681 41657 579849
rect 42249 579681 717600 579849
rect 0 578653 717600 579681
rect 0 578485 41657 578653
rect 42249 578485 717600 578653
rect 0 578009 717600 578485
rect 0 577841 41657 578009
rect 42249 577841 717600 578009
rect 0 577365 717600 577841
rect 0 577197 41657 577365
rect 42249 577197 717600 577365
rect 0 576813 717600 577197
rect 0 576645 41657 576813
rect 42249 576645 717600 576813
rect 0 575525 717600 576645
rect 0 575357 41657 575525
rect 42249 575357 717600 575525
rect 0 574881 717600 575357
rect 0 574713 41657 574881
rect 42249 574713 717600 574881
rect 0 574329 717600 574713
rect 0 574161 41657 574329
rect 42249 574161 717600 574329
rect 0 573685 717600 574161
rect 0 573517 41657 573685
rect 42249 573517 717600 573685
rect 0 573041 717600 573517
rect 0 572873 41657 573041
rect 42249 572873 717600 573041
rect 0 572489 717600 572873
rect 0 572321 41657 572489
rect 42249 572321 717600 572489
rect 0 570649 717600 572321
rect 0 570481 41657 570649
rect 42249 570481 717600 570649
rect 0 570005 717600 570481
rect 0 569837 41657 570005
rect 42249 569837 717600 570005
rect 0 569361 717600 569837
rect 0 569193 41657 569361
rect 42249 569193 717600 569361
rect 0 563007 717600 569193
rect 0 562839 675351 563007
rect 675943 562839 717600 563007
rect 0 562363 717600 562839
rect 0 562195 675351 562363
rect 675943 562195 717600 562363
rect 0 561719 717600 562195
rect 0 561551 675351 561719
rect 675943 561551 717600 561719
rect 0 559879 717600 561551
rect 0 559711 675351 559879
rect 675943 559711 717600 559879
rect 0 559327 717600 559711
rect 0 559159 675351 559327
rect 675943 559159 717600 559327
rect 0 558683 717600 559159
rect 0 558515 675351 558683
rect 675943 558515 717600 558683
rect 0 558039 717600 558515
rect 0 557871 675351 558039
rect 675943 557871 717600 558039
rect 0 557487 717600 557871
rect 0 557319 675351 557487
rect 675943 557319 717600 557487
rect 0 556843 717600 557319
rect 0 556675 675351 556843
rect 675943 556675 717600 556843
rect 0 555555 717600 556675
rect 0 555387 675351 555555
rect 675943 555387 717600 555555
rect 0 555003 717600 555387
rect 0 554835 675351 555003
rect 675943 554835 717600 555003
rect 0 554359 717600 554835
rect 0 554191 675351 554359
rect 675943 554191 717600 554359
rect 0 553715 717600 554191
rect 0 553547 675351 553715
rect 675943 553547 717600 553715
rect 0 552519 717600 553547
rect 0 552351 675351 552519
rect 675943 552351 717600 552519
rect 0 551323 717600 552351
rect 0 551155 675351 551323
rect 675943 551155 717600 551323
rect 0 550679 717600 551155
rect 0 550511 675351 550679
rect 675943 550511 717600 550679
rect 0 548839 717600 550511
rect 0 548671 675351 548839
rect 675943 548671 717600 548839
rect 0 540329 717600 548671
rect 0 540161 41657 540329
rect 42249 540161 717600 540329
rect 0 538489 717600 540161
rect 0 538321 41657 538489
rect 42249 538321 717600 538489
rect 0 537845 717600 538321
rect 0 537677 41657 537845
rect 42249 537677 717600 537845
rect 0 536649 717600 537677
rect 0 536481 41657 536649
rect 42249 536481 717600 536649
rect 0 535453 717600 536481
rect 0 535285 41657 535453
rect 42249 535285 717600 535453
rect 0 534809 717600 535285
rect 0 534641 41657 534809
rect 42249 534641 717600 534809
rect 0 534165 717600 534641
rect 0 533997 41657 534165
rect 42249 533997 717600 534165
rect 0 533613 717600 533997
rect 0 533445 41657 533613
rect 42249 533445 717600 533613
rect 0 532325 717600 533445
rect 0 532157 41657 532325
rect 42249 532157 717600 532325
rect 0 531681 717600 532157
rect 0 531513 41657 531681
rect 42249 531513 717600 531681
rect 0 531129 717600 531513
rect 0 530961 41657 531129
rect 42249 530961 717600 531129
rect 0 530485 717600 530961
rect 0 530317 41657 530485
rect 42249 530317 717600 530485
rect 0 529841 717600 530317
rect 0 529673 41657 529841
rect 42249 529673 717600 529841
rect 0 529289 717600 529673
rect 0 529121 41657 529289
rect 42249 529121 717600 529289
rect 0 527449 717600 529121
rect 0 527281 41657 527449
rect 42249 527281 717600 527449
rect 0 526805 717600 527281
rect 0 526637 41657 526805
rect 42249 526637 717600 526805
rect 0 526161 717600 526637
rect 0 525993 41657 526161
rect 42249 525993 717600 526161
rect 0 412729 717600 525993
rect 0 412561 41657 412729
rect 42249 412561 717600 412729
rect 0 410889 717600 412561
rect 0 410721 41657 410889
rect 42249 410721 717600 410889
rect 0 410245 717600 410721
rect 0 410077 41657 410245
rect 42249 410077 717600 410245
rect 0 409049 717600 410077
rect 0 408881 41657 409049
rect 42249 408881 717600 409049
rect 0 407853 717600 408881
rect 0 407685 41657 407853
rect 42249 407685 717600 407853
rect 0 407209 717600 407685
rect 0 407041 41657 407209
rect 42249 407041 717600 407209
rect 0 406565 717600 407041
rect 0 406397 41657 406565
rect 42249 406397 717600 406565
rect 0 406013 717600 406397
rect 0 405845 41657 406013
rect 42249 405845 717600 406013
rect 0 404725 717600 405845
rect 0 404557 41657 404725
rect 42249 404557 717600 404725
rect 0 404081 717600 404557
rect 0 403913 41657 404081
rect 42249 403913 717600 404081
rect 0 403529 717600 403913
rect 0 403361 41657 403529
rect 42249 403361 717600 403529
rect 0 402885 717600 403361
rect 0 402717 41657 402885
rect 42249 402717 717600 402885
rect 0 402241 717600 402717
rect 0 402073 41657 402241
rect 42249 402073 717600 402241
rect 0 401689 717600 402073
rect 0 401521 41657 401689
rect 42249 401521 717600 401689
rect 0 399849 717600 401521
rect 0 399681 41657 399849
rect 42249 399681 717600 399849
rect 0 399205 717600 399681
rect 0 399037 41657 399205
rect 42249 399037 717600 399205
rect 0 398561 717600 399037
rect 0 398393 41657 398561
rect 42249 398393 717600 398561
rect 0 385807 717600 398393
rect 0 385639 675351 385807
rect 675943 385639 717600 385807
rect 0 385163 717600 385639
rect 0 384995 675351 385163
rect 675943 384995 717600 385163
rect 0 384519 717600 384995
rect 0 384351 675351 384519
rect 675943 384351 717600 384519
rect 0 382679 717600 384351
rect 0 382511 675351 382679
rect 675943 382511 717600 382679
rect 0 382127 717600 382511
rect 0 381959 675351 382127
rect 675943 381959 717600 382127
rect 0 381483 717600 381959
rect 0 381315 675351 381483
rect 675943 381315 717600 381483
rect 0 380839 717600 381315
rect 0 380671 675351 380839
rect 675943 380671 717600 380839
rect 0 380287 717600 380671
rect 0 380119 675351 380287
rect 675943 380119 717600 380287
rect 0 379643 717600 380119
rect 0 379475 675351 379643
rect 675943 379475 717600 379643
rect 0 378355 717600 379475
rect 0 378187 675351 378355
rect 675943 378187 717600 378355
rect 0 377803 717600 378187
rect 0 377635 675351 377803
rect 675943 377635 717600 377803
rect 0 377159 717600 377635
rect 0 376991 675351 377159
rect 675943 376991 717600 377159
rect 0 376515 717600 376991
rect 0 376347 675351 376515
rect 675943 376347 717600 376515
rect 0 375319 717600 376347
rect 0 375151 675351 375319
rect 675943 375151 717600 375319
rect 0 373479 717600 375151
rect 0 373311 675351 373479
rect 675943 373311 717600 373479
rect 0 371639 717600 373311
rect 0 371471 675351 371639
rect 675943 371471 717600 371639
rect 0 369529 717600 371471
rect 0 369361 41657 369529
rect 42249 369361 717600 369529
rect 0 367689 717600 369361
rect 0 367521 41657 367689
rect 42249 367521 717600 367689
rect 0 367045 717600 367521
rect 0 366877 41657 367045
rect 42249 366877 717600 367045
rect 0 365849 717600 366877
rect 0 365681 41657 365849
rect 42249 365681 717600 365849
rect 0 364653 717600 365681
rect 0 364485 41657 364653
rect 42249 364485 717600 364653
rect 0 364009 717600 364485
rect 0 363841 41657 364009
rect 42249 363841 717600 364009
rect 0 363365 717600 363841
rect 0 363197 41657 363365
rect 42249 363197 717600 363365
rect 0 362813 717600 363197
rect 0 362645 41657 362813
rect 42249 362645 717600 362813
rect 0 361525 717600 362645
rect 0 361357 41657 361525
rect 42249 361357 717600 361525
rect 0 360881 717600 361357
rect 0 360713 41657 360881
rect 42249 360713 717600 360881
rect 0 360329 717600 360713
rect 0 360161 41657 360329
rect 42249 360161 717600 360329
rect 0 359685 717600 360161
rect 0 359517 41657 359685
rect 42249 359517 717600 359685
rect 0 359041 717600 359517
rect 0 358873 41657 359041
rect 42249 358873 717600 359041
rect 0 358489 717600 358873
rect 0 358321 41657 358489
rect 42249 358321 717600 358489
rect 0 356649 717600 358321
rect 0 356481 41657 356649
rect 42249 356481 717600 356649
rect 0 356005 717600 356481
rect 0 355837 41657 356005
rect 42249 355837 717600 356005
rect 0 355361 717600 355837
rect 0 355193 41657 355361
rect 42249 355193 717600 355361
rect 0 340607 717600 355193
rect 0 340439 675351 340607
rect 675943 340439 717600 340607
rect 0 339963 717600 340439
rect 0 339795 675351 339963
rect 675943 339795 717600 339963
rect 0 339319 717600 339795
rect 0 339151 675351 339319
rect 675943 339151 717600 339319
rect 0 337479 717600 339151
rect 0 337311 675351 337479
rect 675943 337311 717600 337479
rect 0 336927 717600 337311
rect 0 336759 675351 336927
rect 675943 336759 717600 336927
rect 0 336283 717600 336759
rect 0 336115 675351 336283
rect 675943 336115 717600 336283
rect 0 335639 717600 336115
rect 0 335471 675351 335639
rect 675943 335471 717600 335639
rect 0 335087 717600 335471
rect 0 334919 675351 335087
rect 675943 334919 717600 335087
rect 0 334443 717600 334919
rect 0 334275 675351 334443
rect 675943 334275 717600 334443
rect 0 333155 717600 334275
rect 0 332987 675351 333155
rect 675943 332987 717600 333155
rect 0 332603 717600 332987
rect 0 332435 675351 332603
rect 675943 332435 717600 332603
rect 0 331959 717600 332435
rect 0 331791 675351 331959
rect 675943 331791 717600 331959
rect 0 331315 717600 331791
rect 0 331147 675351 331315
rect 675943 331147 717600 331315
rect 0 330119 717600 331147
rect 0 329951 675351 330119
rect 675943 329951 717600 330119
rect 0 328279 717600 329951
rect 0 328111 675351 328279
rect 675943 328111 717600 328279
rect 0 326439 717600 328111
rect 0 326329 675351 326439
rect 0 326161 41657 326329
rect 42249 326271 675351 326329
rect 675943 326271 717600 326439
rect 42249 326161 717600 326271
rect 0 324489 717600 326161
rect 0 324321 41657 324489
rect 42249 324321 717600 324489
rect 0 323845 717600 324321
rect 0 323677 41657 323845
rect 42249 323677 717600 323845
rect 0 322649 717600 323677
rect 0 322481 41657 322649
rect 42249 322481 717600 322649
rect 0 321453 717600 322481
rect 0 321285 41657 321453
rect 42249 321285 717600 321453
rect 0 320809 717600 321285
rect 0 320641 41657 320809
rect 42249 320641 717600 320809
rect 0 320165 717600 320641
rect 0 319997 41657 320165
rect 42249 319997 717600 320165
rect 0 319613 717600 319997
rect 0 319445 41657 319613
rect 42249 319445 717600 319613
rect 0 318325 717600 319445
rect 0 318157 41657 318325
rect 42249 318157 717600 318325
rect 0 317681 717600 318157
rect 0 317513 41657 317681
rect 42249 317513 717600 317681
rect 0 317129 717600 317513
rect 0 316961 41657 317129
rect 42249 316961 717600 317129
rect 0 316485 717600 316961
rect 0 316317 41657 316485
rect 42249 316317 717600 316485
rect 0 315841 717600 316317
rect 0 315673 41657 315841
rect 42249 315673 717600 315841
rect 0 315289 717600 315673
rect 0 315121 41657 315289
rect 42249 315121 717600 315289
rect 0 313449 717600 315121
rect 0 313281 41657 313449
rect 42249 313281 717600 313449
rect 0 312805 717600 313281
rect 0 312637 41657 312805
rect 42249 312637 717600 312805
rect 0 312161 717600 312637
rect 0 311993 41657 312161
rect 42249 311993 717600 312161
rect 0 295607 717600 311993
rect 0 295439 675351 295607
rect 675943 295439 717600 295607
rect 0 294963 717600 295439
rect 0 294795 675351 294963
rect 675943 294795 717600 294963
rect 0 294319 717600 294795
rect 0 294151 675351 294319
rect 675943 294151 717600 294319
rect 0 292479 717600 294151
rect 0 292311 675351 292479
rect 675943 292311 717600 292479
rect 0 291927 717600 292311
rect 0 291759 675351 291927
rect 675943 291759 717600 291927
rect 0 291283 717600 291759
rect 0 291115 675351 291283
rect 675943 291115 717600 291283
rect 0 290639 717600 291115
rect 0 290471 675351 290639
rect 675943 290471 717600 290639
rect 0 290087 717600 290471
rect 0 289919 675351 290087
rect 675943 289919 717600 290087
rect 0 289443 717600 289919
rect 0 289275 675351 289443
rect 675943 289275 717600 289443
rect 0 288155 717600 289275
rect 0 287987 675351 288155
rect 675943 287987 717600 288155
rect 0 287603 717600 287987
rect 0 287435 675351 287603
rect 675943 287435 717600 287603
rect 0 286959 717600 287435
rect 0 286791 675351 286959
rect 675943 286791 717600 286959
rect 0 286315 717600 286791
rect 0 286147 675351 286315
rect 675943 286147 717600 286315
rect 0 285119 717600 286147
rect 0 284951 675351 285119
rect 675943 284951 717600 285119
rect 0 283279 717600 284951
rect 0 283129 675351 283279
rect 0 282961 41657 283129
rect 42249 283111 675351 283129
rect 675943 283111 717600 283279
rect 42249 282961 717600 283111
rect 0 281439 717600 282961
rect 0 281289 675351 281439
rect 0 281121 41657 281289
rect 42249 281271 675351 281289
rect 675943 281271 717600 281439
rect 42249 281121 717600 281271
rect 0 280645 717600 281121
rect 0 280477 41657 280645
rect 42249 280477 717600 280645
rect 0 279449 717600 280477
rect 0 279281 41657 279449
rect 42249 279281 717600 279449
rect 0 278253 717600 279281
rect 0 278085 41657 278253
rect 42249 278085 717600 278253
rect 0 277609 717600 278085
rect 0 277441 41657 277609
rect 42249 277441 717600 277609
rect 0 276965 717600 277441
rect 0 276797 41657 276965
rect 42249 276797 717600 276965
rect 0 276413 717600 276797
rect 0 276245 41657 276413
rect 42249 276245 717600 276413
rect 0 275125 717600 276245
rect 0 274957 41657 275125
rect 42249 274957 717600 275125
rect 0 274481 717600 274957
rect 0 274313 41657 274481
rect 42249 274313 717600 274481
rect 0 273929 717600 274313
rect 0 273761 41657 273929
rect 42249 273761 717600 273929
rect 0 273285 717600 273761
rect 0 273117 41657 273285
rect 42249 273117 717600 273285
rect 0 272641 717600 273117
rect 0 272473 41657 272641
rect 42249 272473 717600 272641
rect 0 272089 717600 272473
rect 0 271921 41657 272089
rect 42249 271921 717600 272089
rect 0 270249 717600 271921
rect 0 270081 41657 270249
rect 42249 270081 717600 270249
rect 0 269605 717600 270081
rect 0 269437 41657 269605
rect 42249 269437 717600 269605
rect 0 268961 717600 269437
rect 0 268793 41657 268961
rect 42249 268793 717600 268961
rect 0 250607 717600 268793
rect 0 250439 675351 250607
rect 675943 250439 717600 250607
rect 0 249963 717600 250439
rect 0 249795 675351 249963
rect 675943 249795 717600 249963
rect 0 249319 717600 249795
rect 0 249151 675351 249319
rect 675943 249151 717600 249319
rect 0 247479 717600 249151
rect 0 247311 675351 247479
rect 675943 247311 717600 247479
rect 0 246927 717600 247311
rect 0 246759 675351 246927
rect 675943 246759 717600 246927
rect 0 246283 717600 246759
rect 0 246115 675351 246283
rect 675943 246115 717600 246283
rect 0 245639 717600 246115
rect 0 245471 675351 245639
rect 675943 245471 717600 245639
rect 0 245087 717600 245471
rect 0 244919 675351 245087
rect 675943 244919 717600 245087
rect 0 244443 717600 244919
rect 0 244275 675351 244443
rect 675943 244275 717600 244443
rect 0 243155 717600 244275
rect 0 242987 675351 243155
rect 675943 242987 717600 243155
rect 0 242603 717600 242987
rect 0 242435 675351 242603
rect 675943 242435 717600 242603
rect 0 241959 717600 242435
rect 0 241791 675351 241959
rect 675943 241791 717600 241959
rect 0 241315 717600 241791
rect 0 241147 675351 241315
rect 675943 241147 717600 241315
rect 0 240119 717600 241147
rect 0 239951 675351 240119
rect 675943 239951 717600 240119
rect 0 239929 717600 239951
rect 0 239761 41657 239929
rect 42249 239761 717600 239929
rect 0 238279 717600 239761
rect 0 238111 675351 238279
rect 675943 238111 717600 238279
rect 0 238089 717600 238111
rect 0 237921 41657 238089
rect 42249 237921 717600 238089
rect 0 237445 717600 237921
rect 0 237277 41657 237445
rect 42249 237277 717600 237445
rect 0 236439 717600 237277
rect 0 236271 675351 236439
rect 675943 236271 717600 236439
rect 0 236249 717600 236271
rect 0 236081 41657 236249
rect 42249 236081 717600 236249
rect 0 235053 717600 236081
rect 0 234885 41657 235053
rect 42249 234885 717600 235053
rect 0 234409 717600 234885
rect 0 234241 41657 234409
rect 42249 234241 717600 234409
rect 0 233765 717600 234241
rect 0 233597 41657 233765
rect 42249 233597 717600 233765
rect 0 233213 717600 233597
rect 0 233045 41657 233213
rect 42249 233045 717600 233213
rect 0 231925 717600 233045
rect 0 231757 41657 231925
rect 42249 231757 717600 231925
rect 0 231281 717600 231757
rect 0 231113 41657 231281
rect 42249 231113 717600 231281
rect 0 230729 717600 231113
rect 0 230561 41657 230729
rect 42249 230561 717600 230729
rect 0 230085 717600 230561
rect 0 229917 41657 230085
rect 42249 229917 717600 230085
rect 0 229441 717600 229917
rect 0 229273 41657 229441
rect 42249 229273 717600 229441
rect 0 228889 717600 229273
rect 0 228721 41657 228889
rect 42249 228721 717600 228889
rect 0 227049 717600 228721
rect 0 226881 41657 227049
rect 42249 226881 717600 227049
rect 0 226405 717600 226881
rect 0 226237 41657 226405
rect 42249 226237 717600 226405
rect 0 225761 717600 226237
rect 0 225593 41657 225761
rect 42249 225593 717600 225761
rect 0 205407 717600 225593
rect 0 205239 675351 205407
rect 675943 205239 717600 205407
rect 0 204763 717600 205239
rect 0 204595 675351 204763
rect 675943 204595 717600 204763
rect 0 204119 717600 204595
rect 0 203951 675351 204119
rect 675943 203951 717600 204119
rect 0 202279 717600 203951
rect 0 202111 675351 202279
rect 675943 202111 717600 202279
rect 0 201727 717600 202111
rect 0 201559 675351 201727
rect 675943 201559 717600 201727
rect 0 201083 717600 201559
rect 0 200915 675351 201083
rect 675943 200915 717600 201083
rect 0 200439 717600 200915
rect 0 200271 675351 200439
rect 675943 200271 717600 200439
rect 0 199887 717600 200271
rect 0 199719 675351 199887
rect 675943 199719 717600 199887
rect 0 199243 717600 199719
rect 0 199075 675351 199243
rect 675943 199075 717600 199243
rect 0 197955 717600 199075
rect 0 197787 675351 197955
rect 675943 197787 717600 197955
rect 0 197403 717600 197787
rect 0 197235 675351 197403
rect 675943 197235 717600 197403
rect 0 196759 717600 197235
rect 0 196729 675351 196759
rect 0 196561 41657 196729
rect 42249 196591 675351 196729
rect 675943 196591 717600 196759
rect 42249 196561 717600 196591
rect 0 196115 717600 196561
rect 0 195947 675351 196115
rect 675943 195947 717600 196115
rect 0 194919 717600 195947
rect 0 194889 675351 194919
rect 0 194721 41657 194889
rect 42249 194751 675351 194889
rect 675943 194751 717600 194919
rect 42249 194721 717600 194751
rect 0 194245 717600 194721
rect 0 194077 41657 194245
rect 42249 194077 717600 194245
rect 0 193079 717600 194077
rect 0 193049 675351 193079
rect 0 192881 41657 193049
rect 42249 192911 675351 193049
rect 675943 192911 717600 193079
rect 42249 192881 717600 192911
rect 0 191853 717600 192881
rect 0 191685 41657 191853
rect 42249 191685 717600 191853
rect 0 191239 717600 191685
rect 0 191209 675351 191239
rect 0 191041 41657 191209
rect 42249 191071 675351 191209
rect 675943 191071 717600 191239
rect 42249 191041 717600 191071
rect 0 190565 717600 191041
rect 0 190397 41657 190565
rect 42249 190397 717600 190565
rect 0 190013 717600 190397
rect 0 189845 41657 190013
rect 42249 189845 717600 190013
rect 0 188725 717600 189845
rect 0 188557 41657 188725
rect 42249 188557 717600 188725
rect 0 188081 717600 188557
rect 0 187913 41657 188081
rect 42249 187913 717600 188081
rect 0 187529 717600 187913
rect 0 187361 41657 187529
rect 42249 187361 717600 187529
rect 0 186885 717600 187361
rect 0 186717 41657 186885
rect 42249 186717 717600 186885
rect 0 186241 717600 186717
rect 0 186073 41657 186241
rect 42249 186073 717600 186241
rect 0 185689 717600 186073
rect 0 185521 41657 185689
rect 42249 185521 717600 185689
rect 0 183849 717600 185521
rect 0 183681 41657 183849
rect 42249 183681 717600 183849
rect 0 183205 717600 183681
rect 0 183037 41657 183205
rect 42249 183037 717600 183205
rect 0 182561 717600 183037
rect 0 182393 41657 182561
rect 42249 182393 717600 182561
rect 0 160407 717600 182393
rect 0 160239 675351 160407
rect 675943 160239 717600 160407
rect 0 159763 717600 160239
rect 0 159595 675351 159763
rect 675943 159595 717600 159763
rect 0 159119 717600 159595
rect 0 158951 675351 159119
rect 675943 158951 717600 159119
rect 0 157279 717600 158951
rect 0 157111 675351 157279
rect 675943 157111 717600 157279
rect 0 156727 717600 157111
rect 0 156559 675351 156727
rect 675943 156559 717600 156727
rect 0 156083 717600 156559
rect 0 155915 675351 156083
rect 675943 155915 717600 156083
rect 0 155439 717600 155915
rect 0 155271 675351 155439
rect 675943 155271 717600 155439
rect 0 154887 717600 155271
rect 0 154719 675351 154887
rect 675943 154719 717600 154887
rect 0 154243 717600 154719
rect 0 154075 675351 154243
rect 675943 154075 717600 154243
rect 0 152955 717600 154075
rect 0 152787 675351 152955
rect 675943 152787 717600 152955
rect 0 152403 717600 152787
rect 0 152235 675351 152403
rect 675943 152235 717600 152403
rect 0 151759 717600 152235
rect 0 151591 675351 151759
rect 675943 151591 717600 151759
rect 0 151115 717600 151591
rect 0 150947 675351 151115
rect 675943 150947 717600 151115
rect 0 149919 717600 150947
rect 0 149751 675351 149919
rect 675943 149751 717600 149919
rect 0 148079 717600 149751
rect 0 147911 675351 148079
rect 675943 147911 717600 148079
rect 0 146239 717600 147911
rect 0 146071 675351 146239
rect 675943 146071 717600 146239
rect 0 115207 717600 146071
rect 0 115039 675351 115207
rect 675943 115039 717600 115207
rect 0 114563 717600 115039
rect 0 114395 675351 114563
rect 675943 114395 717600 114563
rect 0 113919 717600 114395
rect 0 113751 675351 113919
rect 675943 113751 717600 113919
rect 0 112079 717600 113751
rect 0 111911 675351 112079
rect 675943 111911 717600 112079
rect 0 111527 717600 111911
rect 0 111359 675351 111527
rect 675943 111359 717600 111527
rect 0 110883 717600 111359
rect 0 110715 675351 110883
rect 675943 110715 717600 110883
rect 0 110239 717600 110715
rect 0 110071 675351 110239
rect 675943 110071 717600 110239
rect 0 109687 717600 110071
rect 0 109519 675351 109687
rect 675943 109519 717600 109687
rect 0 109043 717600 109519
rect 0 108875 675351 109043
rect 675943 108875 717600 109043
rect 0 107755 717600 108875
rect 0 107587 675351 107755
rect 675943 107587 717600 107755
rect 0 107203 717600 107587
rect 0 107035 675351 107203
rect 675943 107035 717600 107203
rect 0 106559 717600 107035
rect 0 106391 675351 106559
rect 675943 106391 717600 106559
rect 0 105915 717600 106391
rect 0 105747 675351 105915
rect 675943 105747 717600 105915
rect 0 104719 717600 105747
rect 0 104551 675351 104719
rect 675943 104551 717600 104719
rect 0 102879 717600 104551
rect 0 102711 675351 102879
rect 675943 102711 717600 102879
rect 0 101039 717600 102711
rect 0 100871 675351 101039
rect 675943 100871 717600 101039
rect 0 42249 717600 100871
rect 0 41657 187271 42249
rect 187439 41657 193987 42249
rect 194155 41657 302587 42249
rect 302755 41657 306911 42249
rect 307079 41657 310039 42249
rect 310207 41657 357387 42249
rect 357555 41657 361711 42249
rect 361879 41657 364839 42249
rect 365007 41657 405471 42249
rect 405639 41657 412187 42249
rect 412355 41657 416511 42249
rect 416679 41657 419639 42249
rect 419807 41657 460271 42249
rect 460439 41657 466987 42249
rect 467155 41657 471311 42249
rect 471479 41657 474439 42249
rect 474607 41657 515071 42249
rect 515239 41657 520591 42249
rect 520759 41657 521787 42249
rect 521955 41657 524915 42249
rect 525083 41657 526111 42249
rect 526279 41657 529239 42249
rect 529407 41657 717600 42249
rect 0 40056 717600 41657
rect 0 39878 141611 40056
rect 141869 39878 145035 40056
rect 0 39650 145035 39878
rect 145199 39650 717600 40056
rect 0 0 717600 39650
<< metal3 >>
rect 333499 997600 338279 1002770
rect 343478 997600 348258 1002770
rect 575699 997600 580479 1004112
rect 585678 997600 590458 1004952
rect 38220 922151 39600 926940
rect 678000 917700 679380 922500
rect 38220 912100 39600 916900
rect 678000 907660 679380 912449
rect 32648 837678 40000 842458
rect 32698 827699 40000 832479
rect 677600 828521 680592 833301
rect 677600 818542 680592 823322
rect 37008 493078 40000 497858
rect 37008 483099 40000 487879
rect 678000 469900 685920 474700
rect 678000 459860 685920 464649
rect 31680 450951 39600 455740
rect 31680 440900 39600 445700
rect 36040 120278 40000 125058
rect 36040 110299 40000 115079
rect 38220 78151 39600 82940
rect 38220 68100 39600 72900
rect 78942 32648 83722 40000
rect 88921 32698 93701 40000
rect 141667 37818 141813 40000
rect 241260 31680 246049 39600
rect 251300 31680 256100 39600
rect 569142 34830 573922 40000
rect 579121 34830 583901 40000
rect 622942 37008 627722 40000
rect 632921 37008 637701 40000
<< obsm3 >>
rect 0 1005032 717600 1037600
rect 0 1004192 585598 1005032
rect 0 1002850 575619 1004192
rect 0 997520 333419 1002850
rect 338359 997520 343398 1002850
rect 348338 997520 575619 1002850
rect 580559 997520 585598 1004192
rect 590538 997520 717600 1005032
rect 0 927020 717600 997520
rect 0 922071 38140 927020
rect 39680 922580 717600 927020
rect 39680 922071 677920 922580
rect 0 917620 677920 922071
rect 679460 917620 717600 922580
rect 0 916980 717600 917620
rect 0 912020 38140 916980
rect 39680 912529 717600 916980
rect 39680 912020 677920 912529
rect 0 907580 677920 912020
rect 679460 907580 717600 912529
rect 0 842538 717600 907580
rect 0 837598 32568 842538
rect 40080 837598 717600 842538
rect 0 833381 717600 837598
rect 0 832559 677520 833381
rect 0 827619 32618 832559
rect 40080 828441 677520 832559
rect 680672 828441 717600 833381
rect 40080 827619 717600 828441
rect 0 823402 717600 827619
rect 0 818462 677520 823402
rect 680672 818462 717600 823402
rect 0 497938 717600 818462
rect 0 492998 36928 497938
rect 40080 492998 717600 497938
rect 0 487959 717600 492998
rect 0 483019 36928 487959
rect 40080 483019 717600 487959
rect 0 474780 717600 483019
rect 0 469820 677920 474780
rect 686000 469820 717600 474780
rect 0 464729 717600 469820
rect 0 459780 677920 464729
rect 686000 459780 717600 464729
rect 0 455820 717600 459780
rect 0 450871 31600 455820
rect 39680 450871 717600 455820
rect 0 445780 717600 450871
rect 0 440820 31600 445780
rect 39680 440820 717600 445780
rect 0 125138 717600 440820
rect 0 120198 35960 125138
rect 40080 120198 717600 125138
rect 0 115159 717600 120198
rect 0 110219 35960 115159
rect 40080 110219 717600 115159
rect 0 83020 717600 110219
rect 0 78071 38140 83020
rect 39680 78071 717600 83020
rect 0 72980 717600 78071
rect 0 68020 38140 72980
rect 39680 68020 717600 72980
rect 0 40080 717600 68020
rect 0 32568 78862 40080
rect 83802 32618 88841 40080
rect 93781 37738 141587 40080
rect 141893 39680 569062 40080
rect 141893 37738 241180 39680
rect 93781 32618 241180 37738
rect 83802 32568 241180 32618
rect 0 31600 241180 32568
rect 246129 31600 251220 39680
rect 256180 34750 569062 39680
rect 574002 34750 579041 40080
rect 583981 36928 622862 40080
rect 627802 36928 632841 40080
rect 637781 36928 717600 40080
rect 583981 34750 717600 36928
rect 256180 31600 717600 34750
rect 0 0 717600 31600
<< metal4 >>
rect 333400 1032757 333654 1037599
rect 348146 1032757 348400 1037599
rect 575600 1008881 575854 1008947
rect 590346 1008881 590600 1008947
rect 575600 1007929 575854 1008165
rect 590346 1007929 590600 1008165
rect 575600 1007147 575854 1007213
rect 590346 1007147 590600 1007213
rect 575600 1004947 575854 1005637
rect 590346 1004947 590600 1005637
rect 333400 1002767 333654 1003697
rect 348146 1002767 348400 1003697
rect 37293 926746 38223 927000
rect 679377 922346 680307 922600
rect 37293 912000 38223 912254
rect 679377 907600 680307 907854
rect 28653 842346 28719 842600
rect 29435 842346 29671 842600
rect 30387 842346 30453 842600
rect 31963 842346 32653 842600
rect 680587 833207 681277 833399
rect 28653 827600 28719 827854
rect 29435 827600 29671 827854
rect 30387 827600 30453 827854
rect 31963 827600 32653 827854
rect 680587 818400 681277 818592
rect 36323 497807 37013 497999
rect 36323 483000 37013 483192
rect 685917 474546 686847 474800
rect 685917 459800 686847 460054
rect 30753 455546 31683 455800
rect 30753 440800 31683 441054
rect 21000 124946 25992 125200
rect 35113 124946 36043 125200
rect 21000 110200 25992 110454
rect 35113 110200 36043 110454
rect 37293 82746 38223 83000
rect 37293 68000 38223 68254
rect 622800 36323 622992 37013
rect 637607 36323 637799 37013
rect 78800 31963 79054 32653
rect 93546 31963 93800 32653
rect 241200 30753 241454 31683
rect 255946 30753 256200 31683
rect 78800 30387 79054 30453
rect 93546 30387 93800 30453
rect 78800 29435 79054 29671
rect 93546 29435 93800 29671
rect 78800 28653 79054 28719
rect 93546 28653 93800 28719
<< obsm4 >>
rect 0 1032677 333320 1037600
rect 333734 1032677 348066 1037600
rect 348480 1032677 717600 1037600
rect 0 1009027 717600 1032677
rect 0 1008801 575520 1009027
rect 575934 1008801 590266 1009027
rect 590680 1008801 717600 1009027
rect 0 1008245 717600 1008801
rect 0 1007849 575520 1008245
rect 575934 1007849 590266 1008245
rect 590680 1007849 717600 1008245
rect 0 1007293 717600 1007849
rect 0 1007067 575520 1007293
rect 575934 1007067 590266 1007293
rect 590680 1007067 717600 1007293
rect 0 1005717 717600 1007067
rect 0 1004867 575520 1005717
rect 575934 1004867 590266 1005717
rect 590680 1004867 717600 1005717
rect 0 1003777 717600 1004867
rect 0 1002687 333320 1003777
rect 333734 1002687 348066 1003777
rect 348480 1002687 717600 1003777
rect 0 927080 717600 1002687
rect 0 926666 37213 927080
rect 38303 926666 717600 927080
rect 0 922680 717600 926666
rect 0 922266 679297 922680
rect 680387 922266 717600 922680
rect 0 912334 717600 922266
rect 0 911920 37213 912334
rect 38303 911920 717600 912334
rect 0 907934 717600 911920
rect 0 907520 679297 907934
rect 680387 907520 717600 907934
rect 0 842680 717600 907520
rect 0 842266 28573 842680
rect 28799 842266 29355 842680
rect 29751 842266 30307 842680
rect 30533 842266 31883 842680
rect 32733 842266 717600 842680
rect 0 833479 717600 842266
rect 0 833127 680507 833479
rect 681357 833127 717600 833479
rect 0 827934 717600 833127
rect 0 827520 28573 827934
rect 28799 827520 29355 827934
rect 29751 827520 30307 827934
rect 30533 827520 31883 827934
rect 32733 827520 717600 827934
rect 0 818672 717600 827520
rect 0 818320 680507 818672
rect 681357 818320 717600 818672
rect 0 498079 717600 818320
rect 0 497727 36243 498079
rect 37093 497727 717600 498079
rect 0 483272 717600 497727
rect 0 482920 36243 483272
rect 37093 482920 717600 483272
rect 0 474880 717600 482920
rect 0 474466 685837 474880
rect 686927 474466 717600 474880
rect 0 460134 717600 474466
rect 0 459720 685837 460134
rect 686927 459720 717600 460134
rect 0 455880 717600 459720
rect 0 455466 30673 455880
rect 31763 455466 717600 455880
rect 0 441134 717600 455466
rect 0 440720 30673 441134
rect 31763 440720 717600 441134
rect 0 125280 717600 440720
rect 0 124866 20920 125280
rect 26072 124866 35033 125280
rect 36123 124866 717600 125280
rect 0 110534 717600 124866
rect 0 110120 20920 110534
rect 26072 110120 35033 110534
rect 36123 110120 717600 110534
rect 0 83080 717600 110120
rect 0 82666 37213 83080
rect 38303 82666 717600 83080
rect 0 68334 717600 82666
rect 0 67920 37213 68334
rect 38303 67920 717600 68334
rect 0 37093 717600 67920
rect 0 36243 622720 37093
rect 623072 36243 637527 37093
rect 637879 36243 717600 37093
rect 0 32733 717600 36243
rect 0 31883 78720 32733
rect 79134 31883 93466 32733
rect 93880 31883 717600 32733
rect 0 31763 717600 31883
rect 0 30673 241120 31763
rect 241534 30673 255866 31763
rect 256280 30673 717600 31763
rect 0 30533 717600 30673
rect 0 30307 78720 30533
rect 79134 30307 93466 30533
rect 93880 30307 717600 30533
rect 0 29751 717600 30307
rect 0 29355 78720 29751
rect 79134 29355 93466 29751
rect 93880 29355 717600 29751
rect 0 28799 717600 29355
rect 0 28573 78720 28799
rect 79134 28573 93466 28799
rect 93880 28573 717600 28799
rect 0 0 717600 28573
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030789
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 575600 1007147 575854 1008947
rect 590346 1007147 590600 1008947
rect 575600 1004968 575854 1005616
rect 590346 1004968 590600 1005616
rect 333400 1002787 333654 1003677
rect 348146 1002787 348400 1003677
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 37313 926746 38203 927000
rect 6167 914054 19620 924934
rect 679397 922346 680287 922600
rect 37313 912000 38203 912254
rect 697980 909666 711433 920546
rect 679397 907600 680287 907854
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 28653 842346 30453 842600
rect 31983 842346 32631 842600
rect 6811 829010 18976 841178
rect 680607 833207 681257 833399
rect 28653 827600 30453 827854
rect 31983 827600 32631 827854
rect 698624 819822 710789 831990
rect 680607 818400 681257 818592
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 36343 497807 36993 497999
rect 6811 484410 18976 496578
rect 36343 483000 36993 483192
rect 685937 474546 686827 474800
rect 697980 461866 711433 472746
rect 685937 459800 686827 460054
rect 30773 455546 31663 455800
rect 6167 442854 19620 453734
rect 30773 440800 31663 441054
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 21003 124946 25993 125200
rect 35133 124946 36023 125200
rect 6811 111610 18976 123778
rect 21003 110200 25993 110454
rect 35133 110200 36023 110454
rect 698512 101240 711002 113760
rect 37313 82746 38203 83000
rect 6167 70054 19620 80934
rect 37313 68000 38203 68254
rect 622800 36343 622992 36993
rect 637607 36343 637799 36993
rect 78800 31983 79054 32631
rect 93546 31983 93800 32631
rect 241200 30773 241454 31663
rect 78800 28653 79054 30453
rect 255946 30773 256200 31663
rect 93546 28653 93800 30453
rect 80222 6811 92390 18976
rect 136703 7133 144159 18319
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
<< obsm5 >>
rect 0 1031322 717600 1037600
rect 0 1018192 78120 1031322
rect 91280 1018192 129520 1031322
rect 142680 1018192 180920 1031322
rect 194080 1018192 232320 1031322
rect 245480 1018192 283920 1031322
rect 297080 1031109 385720 1031322
rect 297080 1018304 334490 1031109
rect 347298 1018304 385720 1031109
rect 297080 1018192 385720 1018304
rect 398880 1018192 474720 1031322
rect 487880 1018192 526120 1031322
rect 539280 1031109 627920 1031322
rect 539280 1018304 576690 1031109
rect 589498 1018304 627920 1031109
rect 539280 1018192 627920 1018304
rect 641080 1018192 717600 1031322
rect 0 1009267 717600 1018192
rect 0 1006827 575280 1009267
rect 576174 1006827 590026 1009267
rect 590920 1006827 717600 1009267
rect 0 1005936 717600 1006827
rect 0 1004648 575280 1005936
rect 576174 1004648 590026 1005936
rect 590920 1004648 717600 1005936
rect 0 1003997 717600 1004648
rect 0 1002467 333080 1003997
rect 333974 1002467 347826 1003997
rect 348720 1002467 717600 1003997
rect 0 969280 717600 1002467
rect 0 956120 6278 969280
rect 19408 965680 717600 969280
rect 19408 956120 698192 965680
rect 0 952520 698192 956120
rect 711322 952520 717600 965680
rect 0 927320 717600 952520
rect 0 926426 36993 927320
rect 38523 926426 717600 927320
rect 0 925254 717600 926426
rect 0 913734 5847 925254
rect 19940 922920 717600 925254
rect 19940 922026 679077 922920
rect 680607 922026 717600 922920
rect 19940 920866 717600 922026
rect 19940 913734 697660 920866
rect 0 912574 697660 913734
rect 0 911680 36993 912574
rect 38523 911680 697660 912574
rect 0 909346 697660 911680
rect 711753 909346 717600 920866
rect 0 908174 717600 909346
rect 0 907280 679077 908174
rect 680607 907280 717600 908174
rect 0 883698 717600 907280
rect 0 870890 6491 883698
rect 19296 876480 717600 883698
rect 19296 870890 698192 876480
rect 0 863320 698192 870890
rect 711322 863320 717600 876480
rect 0 842920 717600 863320
rect 0 842026 28333 842920
rect 30773 842026 31663 842920
rect 32951 842026 717600 842920
rect 0 841498 717600 842026
rect 0 828690 6491 841498
rect 19296 833719 717600 841498
rect 19296 832887 680287 833719
rect 681577 832887 717600 833719
rect 19296 832310 717600 832887
rect 19296 828690 698304 832310
rect 0 828174 698304 828690
rect 0 827280 28333 828174
rect 30773 827280 31663 828174
rect 32951 827280 698304 828174
rect 0 819502 698304 827280
rect 711109 819502 717600 832310
rect 0 818912 717600 819502
rect 0 818080 680287 818912
rect 681577 818080 717600 818912
rect 0 799480 717600 818080
rect 0 786320 6278 799480
rect 19408 787280 717600 799480
rect 19408 786320 698192 787280
rect 0 774120 698192 786320
rect 711322 774120 717600 787280
rect 0 756280 717600 774120
rect 0 743120 6278 756280
rect 19408 743120 717600 756280
rect 0 742280 717600 743120
rect 0 729120 698192 742280
rect 711322 729120 717600 742280
rect 0 713080 717600 729120
rect 0 699920 6278 713080
rect 19408 699920 717600 713080
rect 0 697280 717600 699920
rect 0 684120 698192 697280
rect 711322 684120 717600 697280
rect 0 669880 717600 684120
rect 0 656720 6278 669880
rect 19408 656720 717600 669880
rect 0 652080 717600 656720
rect 0 638920 698192 652080
rect 711322 638920 717600 652080
rect 0 626680 717600 638920
rect 0 613520 6278 626680
rect 19408 613520 717600 626680
rect 0 607080 717600 613520
rect 0 593920 698192 607080
rect 711322 593920 717600 607080
rect 0 583480 717600 593920
rect 0 570320 6278 583480
rect 19408 570320 717600 583480
rect 0 561880 717600 570320
rect 0 548720 698192 561880
rect 711322 548720 717600 561880
rect 0 540280 717600 548720
rect 0 527120 6278 540280
rect 19408 527120 717600 540280
rect 0 517710 717600 527120
rect 0 504902 698304 517710
rect 711109 504902 717600 517710
rect 0 498319 717600 504902
rect 0 497487 36023 498319
rect 37313 497487 717600 498319
rect 0 496898 717600 497487
rect 0 484090 6491 496898
rect 19296 484090 717600 496898
rect 0 483512 717600 484090
rect 0 482680 36023 483512
rect 37313 482680 717600 483512
rect 0 475120 717600 482680
rect 0 474226 685617 475120
rect 687147 474226 717600 475120
rect 0 473066 717600 474226
rect 0 461546 697660 473066
rect 711753 461546 717600 473066
rect 0 460374 717600 461546
rect 0 459480 685617 460374
rect 687147 459480 717600 460374
rect 0 456120 717600 459480
rect 0 455226 30453 456120
rect 31983 455226 717600 456120
rect 0 454054 717600 455226
rect 0 442534 5847 454054
rect 19940 442534 717600 454054
rect 0 441374 717600 442534
rect 0 440480 30453 441374
rect 31983 440480 717600 441374
rect 0 429510 717600 440480
rect 0 416702 698304 429510
rect 711109 416702 717600 429510
rect 0 412680 717600 416702
rect 0 399520 6278 412680
rect 19408 399520 717600 412680
rect 0 384680 717600 399520
rect 0 371520 698192 384680
rect 711322 371520 717600 384680
rect 0 369480 717600 371520
rect 0 356320 6278 369480
rect 19408 356320 717600 369480
rect 0 339480 717600 356320
rect 0 326320 698192 339480
rect 711322 326320 717600 339480
rect 0 326280 717600 326320
rect 0 313120 6278 326280
rect 19408 313120 717600 326280
rect 0 294480 717600 313120
rect 0 283080 698192 294480
rect 0 269920 6278 283080
rect 19408 281320 698192 283080
rect 711322 281320 717600 294480
rect 19408 269920 717600 281320
rect 0 249480 717600 269920
rect 0 239880 698192 249480
rect 0 226720 6278 239880
rect 19408 236320 698192 239880
rect 711322 236320 717600 249480
rect 19408 226720 717600 236320
rect 0 204280 717600 226720
rect 0 196680 698192 204280
rect 0 183520 6278 196680
rect 19408 191120 698192 196680
rect 711322 191120 717600 204280
rect 19408 183520 717600 191120
rect 0 159280 717600 183520
rect 0 146120 698192 159280
rect 711322 146120 717600 159280
rect 0 125520 717600 146120
rect 0 124626 20683 125520
rect 26313 124626 34813 125520
rect 36343 124626 717600 125520
rect 0 124098 717600 124626
rect 0 111290 6491 124098
rect 19296 114080 717600 124098
rect 19296 111290 698192 114080
rect 0 110774 698192 111290
rect 0 109880 20683 110774
rect 26313 109880 34813 110774
rect 36343 109880 698192 110774
rect 0 100920 698192 109880
rect 711322 100920 717600 114080
rect 0 83320 717600 100920
rect 0 82426 36993 83320
rect 38523 82426 717600 83320
rect 0 81254 717600 82426
rect 0 69734 5847 81254
rect 19940 69734 717600 81254
rect 0 68574 717600 69734
rect 0 67680 36993 68574
rect 38523 67680 717600 68574
rect 0 37313 717600 67680
rect 0 36023 622480 37313
rect 623312 36023 637287 37313
rect 638119 36023 717600 37313
rect 0 32951 717600 36023
rect 0 31663 78480 32951
rect 79374 31663 93226 32951
rect 94120 31983 717600 32951
rect 94120 31663 240880 31983
rect 0 30773 240880 31663
rect 0 28333 78480 30773
rect 79374 28333 93226 30773
rect 94120 30453 240880 30773
rect 241774 30453 255626 31983
rect 256520 30453 717600 31983
rect 94120 28333 717600 30453
rect 0 19940 717600 28333
rect 0 19408 242946 19940
rect 0 19296 187320 19408
rect 0 6491 79902 19296
rect 92710 18639 187320 19296
rect 92710 6813 136383 18639
rect 144479 6813 187320 18639
rect 92710 6491 187320 6813
rect 0 6278 187320 6491
rect 200480 6278 242946 19408
rect 0 5847 242946 6278
rect 254466 19408 717600 19940
rect 254466 6278 295920 19408
rect 309080 6278 350720 19408
rect 363880 6278 405520 19408
rect 418680 6278 460320 19408
rect 473480 6278 515120 19408
rect 528280 19296 717600 19408
rect 528280 6491 570102 19296
rect 582910 6491 623902 19296
rect 636710 6491 717600 19296
rect 528280 6278 717600 6491
rect 254466 5847 717600 6278
rect 0 0 717600 5847
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 1 nsew signal input
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 2 nsew signal output
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 4 nsew signal output
rlabel metal2 s 361767 41713 361823 42193 6 flash_clk_core
port 5 nsew signal input
rlabel metal2 s 357443 41713 357499 42193 6 flash_clk_ieb_core
port 6 nsew signal input
rlabel metal2 s 364895 41713 364951 42193 6 flash_clk_oeb_core
port 7 nsew signal input
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 8 nsew signal output
rlabel metal2 s 306967 41713 307023 42193 6 flash_csb_core
port 9 nsew signal input
rlabel metal2 s 302643 41713 302699 42193 6 flash_csb_ieb_core
port 10 nsew signal input
rlabel metal2 s 310095 41713 310151 42193 6 flash_csb_oeb_core
port 11 nsew signal input
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 12 nsew signal bidirectional
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 13 nsew signal output
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 14 nsew signal input
rlabel metal2 s 412243 41713 412299 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 419695 41713 419751 42193 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 17 nsew signal bidirectional
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 18 nsew signal output
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 19 nsew signal input
rlabel metal2 s 467043 41713 467099 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 474495 41713 474551 42193 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 22 nsew signal bidirectional
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 23 nsew signal output
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 24 nsew signal input
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 25 nsew signal input
rlabel metal2 s 524971 41713 525027 42193 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 27 nsew signal input
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 28 nsew signal input
rlabel metal2 s 675407 551211 675887 551267 6 mprj_analog_io[0]
port 292 nsew signal bidirectional
rlabel metal2 s 485333 995407 485389 995887 6 mprj_analog_io[10]
port 172 nsew signal bidirectional
rlabel metal2 s 396333 995407 396389 995887 6 mprj_analog_io[11]
port 346 nsew signal bidirectional
rlabel metal2 s 294533 995407 294589 995887 6 mprj_analog_io[12]
port 544 nsew signal bidirectional
rlabel metal2 s 242933 995407 242989 995887 6 mprj_analog_io[13]
port 562 nsew signal bidirectional
rlabel metal2 s 191533 995407 191589 995887 6 mprj_analog_io[14]
port 580 nsew signal bidirectional
rlabel metal2 s 140133 995407 140189 995887 6 mprj_analog_io[15]
port 598 nsew signal bidirectional
rlabel metal2 s 88733 995407 88789 995887 6 mprj_analog_io[16]
port 616 nsew signal bidirectional
rlabel metal2 s 41713 966733 42193 966789 6 mprj_analog_io[17]
port 634 nsew signal bidirectional
rlabel metal2 s 41713 796933 42193 796989 6 mprj_analog_io[18]
port 652 nsew signal bidirectional
rlabel metal2 s 41713 753733 42193 753789 6 mprj_analog_io[19]
port 670 nsew signal bidirectional
rlabel metal2 s 675407 596411 675887 596467 6 mprj_analog_io[1]
port 310 nsew signal bidirectional
rlabel metal2 s 41713 710533 42193 710589 6 mprj_analog_io[20]
port 688 nsew signal bidirectional
rlabel metal2 s 41713 667333 42193 667389 6 mprj_analog_io[21]
port 364 nsew signal bidirectional
rlabel metal2 s 41713 624133 42193 624189 6 mprj_analog_io[22]
port 382 nsew signal bidirectional
rlabel metal2 s 41713 580933 42193 580989 6 mprj_analog_io[23]
port 400 nsew signal bidirectional
rlabel metal2 s 41713 537733 42193 537789 6 mprj_analog_io[24]
port 418 nsew signal bidirectional
rlabel metal2 s 41713 410133 42193 410189 6 mprj_analog_io[25]
port 436 nsew signal bidirectional
rlabel metal2 s 41713 366933 42193 366989 6 mprj_analog_io[26]
port 454 nsew signal bidirectional
rlabel metal2 s 41713 323733 42193 323789 6 mprj_analog_io[27]
port 472 nsew signal bidirectional
rlabel metal2 s 41713 280533 42193 280589 6 mprj_analog_io[28]
port 490 nsew signal bidirectional
rlabel metal2 s 41713 237333 42193 237389 6 mprj_analog_io[29]
port 508 nsew signal bidirectional
rlabel metal2 s 675407 641411 675887 641467 6 mprj_analog_io[2]
port 328 nsew signal bidirectional
rlabel metal2 s 41713 194133 42193 194189 6 mprj_analog_io[30]
port 526 nsew signal bidirectional
rlabel metal2 s 675407 686611 675887 686667 6 mprj_analog_io[3]
port 46 nsew signal bidirectional
rlabel metal2 s 675407 731611 675887 731667 6 mprj_analog_io[4]
port 64 nsew signal bidirectional
rlabel metal2 s 675407 776611 675887 776667 6 mprj_analog_io[5]
port 82 nsew signal bidirectional
rlabel metal2 s 675407 865811 675887 865867 6 mprj_analog_io[6]
port 100 nsew signal bidirectional
rlabel metal2 s 675407 955011 675887 955067 6 mprj_analog_io[7]
port 118 nsew signal bidirectional
rlabel metal2 s 638533 995407 638589 995887 6 mprj_analog_io[8]
port 136 nsew signal bidirectional
rlabel metal2 s 536733 995407 536789 995887 6 mprj_analog_io[9]
port 154 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 29 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 47 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 65 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 83 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 101 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 119 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 137 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 155 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 173 nsew signal bidirectional
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 347 nsew signal bidirectional
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 545 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 190 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 563 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 581 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 599 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 617 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 635 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 653 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 671 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 689 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 365 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 383 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 207 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 401 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 419 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 437 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 455 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 473 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 491 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 509 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 527 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 224 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 241 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 258 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 275 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 293 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 311 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 329 nsew signal bidirectional
rlabel metal2 s 675407 105803 675887 105859 6 mprj_io_analog_en[0]
port 30 nsew signal input
rlabel metal2 s 675407 689003 675887 689059 6 mprj_io_analog_en[10]
port 48 nsew signal input
rlabel metal2 s 675407 734003 675887 734059 6 mprj_io_analog_en[11]
port 66 nsew signal input
rlabel metal2 s 675407 779003 675887 779059 6 mprj_io_analog_en[12]
port 84 nsew signal input
rlabel metal2 s 675407 868203 675887 868259 6 mprj_io_analog_en[13]
port 102 nsew signal input
rlabel metal2 s 675407 957403 675887 957459 6 mprj_io_analog_en[14]
port 120 nsew signal input
rlabel metal2 s 636141 995407 636197 995887 6 mprj_io_analog_en[15]
port 138 nsew signal input
rlabel metal2 s 534341 995407 534397 995887 6 mprj_io_analog_en[16]
port 156 nsew signal input
rlabel metal2 s 482941 995407 482997 995887 6 mprj_io_analog_en[17]
port 174 nsew signal input
rlabel metal2 s 393941 995407 393997 995887 6 mprj_io_analog_en[18]
port 348 nsew signal input
rlabel metal2 s 292141 995407 292197 995887 6 mprj_io_analog_en[19]
port 546 nsew signal input
rlabel metal2 s 675407 151003 675887 151059 6 mprj_io_analog_en[1]
port 191 nsew signal input
rlabel metal2 s 240541 995407 240597 995887 6 mprj_io_analog_en[20]
port 564 nsew signal input
rlabel metal2 s 189141 995407 189197 995887 6 mprj_io_analog_en[21]
port 582 nsew signal input
rlabel metal2 s 137741 995407 137797 995887 6 mprj_io_analog_en[22]
port 600 nsew signal input
rlabel metal2 s 86341 995407 86397 995887 6 mprj_io_analog_en[23]
port 618 nsew signal input
rlabel metal2 s 41713 964341 42193 964397 6 mprj_io_analog_en[24]
port 636 nsew signal input
rlabel metal2 s 41713 794541 42193 794597 6 mprj_io_analog_en[25]
port 654 nsew signal input
rlabel metal2 s 41713 751341 42193 751397 6 mprj_io_analog_en[26]
port 672 nsew signal input
rlabel metal2 s 41713 708141 42193 708197 6 mprj_io_analog_en[27]
port 690 nsew signal input
rlabel metal2 s 41713 664941 42193 664997 6 mprj_io_analog_en[28]
port 366 nsew signal input
rlabel metal2 s 41713 621741 42193 621797 6 mprj_io_analog_en[29]
port 384 nsew signal input
rlabel metal2 s 675407 196003 675887 196059 6 mprj_io_analog_en[2]
port 208 nsew signal input
rlabel metal2 s 41713 578541 42193 578597 6 mprj_io_analog_en[30]
port 402 nsew signal input
rlabel metal2 s 41713 535341 42193 535397 6 mprj_io_analog_en[31]
port 420 nsew signal input
rlabel metal2 s 41713 407741 42193 407797 6 mprj_io_analog_en[32]
port 438 nsew signal input
rlabel metal2 s 41713 364541 42193 364597 6 mprj_io_analog_en[33]
port 456 nsew signal input
rlabel metal2 s 41713 321341 42193 321397 6 mprj_io_analog_en[34]
port 474 nsew signal input
rlabel metal2 s 41713 278141 42193 278197 6 mprj_io_analog_en[35]
port 492 nsew signal input
rlabel metal2 s 41713 234941 42193 234997 6 mprj_io_analog_en[36]
port 510 nsew signal input
rlabel metal2 s 41713 191741 42193 191797 6 mprj_io_analog_en[37]
port 528 nsew signal input
rlabel metal2 s 675407 241203 675887 241259 6 mprj_io_analog_en[3]
port 225 nsew signal input
rlabel metal2 s 675407 286203 675887 286259 6 mprj_io_analog_en[4]
port 242 nsew signal input
rlabel metal2 s 675407 331203 675887 331259 6 mprj_io_analog_en[5]
port 259 nsew signal input
rlabel metal2 s 675407 376403 675887 376459 6 mprj_io_analog_en[6]
port 276 nsew signal input
rlabel metal2 s 675407 553603 675887 553659 6 mprj_io_analog_en[7]
port 294 nsew signal input
rlabel metal2 s 675407 598803 675887 598859 6 mprj_io_analog_en[8]
port 312 nsew signal input
rlabel metal2 s 675407 643803 675887 643859 6 mprj_io_analog_en[9]
port 330 nsew signal input
rlabel metal2 s 675407 107091 675887 107147 6 mprj_io_analog_pol[0]
port 31 nsew signal input
rlabel metal2 s 675407 690291 675887 690347 6 mprj_io_analog_pol[10]
port 49 nsew signal input
rlabel metal2 s 675407 735291 675887 735347 6 mprj_io_analog_pol[11]
port 67 nsew signal input
rlabel metal2 s 675407 780291 675887 780347 6 mprj_io_analog_pol[12]
port 85 nsew signal input
rlabel metal2 s 675407 869491 675887 869547 6 mprj_io_analog_pol[13]
port 103 nsew signal input
rlabel metal2 s 675407 958691 675887 958747 6 mprj_io_analog_pol[14]
port 121 nsew signal input
rlabel metal2 s 634853 995407 634909 995887 6 mprj_io_analog_pol[15]
port 139 nsew signal input
rlabel metal2 s 533053 995407 533109 995887 6 mprj_io_analog_pol[16]
port 157 nsew signal input
rlabel metal2 s 481653 995407 481709 995887 6 mprj_io_analog_pol[17]
port 175 nsew signal input
rlabel metal2 s 392653 995407 392709 995887 6 mprj_io_analog_pol[18]
port 349 nsew signal input
rlabel metal2 s 290853 995407 290909 995887 6 mprj_io_analog_pol[19]
port 547 nsew signal input
rlabel metal2 s 675407 152291 675887 152347 6 mprj_io_analog_pol[1]
port 192 nsew signal input
rlabel metal2 s 239253 995407 239309 995887 6 mprj_io_analog_pol[20]
port 565 nsew signal input
rlabel metal2 s 187853 995407 187909 995887 6 mprj_io_analog_pol[21]
port 583 nsew signal input
rlabel metal2 s 136453 995407 136509 995887 6 mprj_io_analog_pol[22]
port 601 nsew signal input
rlabel metal2 s 85053 995407 85109 995887 6 mprj_io_analog_pol[23]
port 619 nsew signal input
rlabel metal2 s 41713 963053 42193 963109 6 mprj_io_analog_pol[24]
port 637 nsew signal input
rlabel metal2 s 41713 793253 42193 793309 6 mprj_io_analog_pol[25]
port 655 nsew signal input
rlabel metal2 s 41713 750053 42193 750109 6 mprj_io_analog_pol[26]
port 673 nsew signal input
rlabel metal2 s 41713 706853 42193 706909 6 mprj_io_analog_pol[27]
port 691 nsew signal input
rlabel metal2 s 41713 663653 42193 663709 6 mprj_io_analog_pol[28]
port 367 nsew signal input
rlabel metal2 s 41713 620453 42193 620509 6 mprj_io_analog_pol[29]
port 385 nsew signal input
rlabel metal2 s 675407 197291 675887 197347 6 mprj_io_analog_pol[2]
port 209 nsew signal input
rlabel metal2 s 41713 577253 42193 577309 6 mprj_io_analog_pol[30]
port 403 nsew signal input
rlabel metal2 s 41713 534053 42193 534109 6 mprj_io_analog_pol[31]
port 421 nsew signal input
rlabel metal2 s 41713 406453 42193 406509 6 mprj_io_analog_pol[32]
port 439 nsew signal input
rlabel metal2 s 41713 363253 42193 363309 6 mprj_io_analog_pol[33]
port 457 nsew signal input
rlabel metal2 s 41713 320053 42193 320109 6 mprj_io_analog_pol[34]
port 475 nsew signal input
rlabel metal2 s 41713 276853 42193 276909 6 mprj_io_analog_pol[35]
port 493 nsew signal input
rlabel metal2 s 41713 233653 42193 233709 6 mprj_io_analog_pol[36]
port 511 nsew signal input
rlabel metal2 s 41713 190453 42193 190509 6 mprj_io_analog_pol[37]
port 529 nsew signal input
rlabel metal2 s 675407 242491 675887 242547 6 mprj_io_analog_pol[3]
port 226 nsew signal input
rlabel metal2 s 675407 287491 675887 287547 6 mprj_io_analog_pol[4]
port 243 nsew signal input
rlabel metal2 s 675407 332491 675887 332547 6 mprj_io_analog_pol[5]
port 260 nsew signal input
rlabel metal2 s 675407 377691 675887 377747 6 mprj_io_analog_pol[6]
port 277 nsew signal input
rlabel metal2 s 675407 554891 675887 554947 6 mprj_io_analog_pol[7]
port 295 nsew signal input
rlabel metal2 s 675407 600091 675887 600147 6 mprj_io_analog_pol[8]
port 313 nsew signal input
rlabel metal2 s 675407 645091 675887 645147 6 mprj_io_analog_pol[9]
port 331 nsew signal input
rlabel metal2 s 675407 110127 675887 110183 6 mprj_io_analog_sel[0]
port 32 nsew signal input
rlabel metal2 s 675407 693327 675887 693383 6 mprj_io_analog_sel[10]
port 50 nsew signal input
rlabel metal2 s 675407 738327 675887 738383 6 mprj_io_analog_sel[11]
port 68 nsew signal input
rlabel metal2 s 675407 783327 675887 783383 6 mprj_io_analog_sel[12]
port 86 nsew signal input
rlabel metal2 s 675407 872527 675887 872583 6 mprj_io_analog_sel[13]
port 104 nsew signal input
rlabel metal2 s 675407 961727 675887 961783 6 mprj_io_analog_sel[14]
port 122 nsew signal input
rlabel metal2 s 631817 995407 631873 995887 6 mprj_io_analog_sel[15]
port 140 nsew signal input
rlabel metal2 s 530017 995407 530073 995887 6 mprj_io_analog_sel[16]
port 158 nsew signal input
rlabel metal2 s 478617 995407 478673 995887 6 mprj_io_analog_sel[17]
port 176 nsew signal input
rlabel metal2 s 389617 995407 389673 995887 6 mprj_io_analog_sel[18]
port 350 nsew signal input
rlabel metal2 s 287817 995407 287873 995887 6 mprj_io_analog_sel[19]
port 548 nsew signal input
rlabel metal2 s 675407 155327 675887 155383 6 mprj_io_analog_sel[1]
port 193 nsew signal input
rlabel metal2 s 236217 995407 236273 995887 6 mprj_io_analog_sel[20]
port 566 nsew signal input
rlabel metal2 s 184817 995407 184873 995887 6 mprj_io_analog_sel[21]
port 584 nsew signal input
rlabel metal2 s 133417 995407 133473 995887 6 mprj_io_analog_sel[22]
port 602 nsew signal input
rlabel metal2 s 82017 995407 82073 995887 6 mprj_io_analog_sel[23]
port 620 nsew signal input
rlabel metal2 s 41713 960017 42193 960073 6 mprj_io_analog_sel[24]
port 638 nsew signal input
rlabel metal2 s 41713 790217 42193 790273 6 mprj_io_analog_sel[25]
port 656 nsew signal input
rlabel metal2 s 41713 747017 42193 747073 6 mprj_io_analog_sel[26]
port 674 nsew signal input
rlabel metal2 s 41713 703817 42193 703873 6 mprj_io_analog_sel[27]
port 692 nsew signal input
rlabel metal2 s 41713 660617 42193 660673 6 mprj_io_analog_sel[28]
port 368 nsew signal input
rlabel metal2 s 41713 617417 42193 617473 6 mprj_io_analog_sel[29]
port 386 nsew signal input
rlabel metal2 s 675407 200327 675887 200383 6 mprj_io_analog_sel[2]
port 210 nsew signal input
rlabel metal2 s 41713 574217 42193 574273 6 mprj_io_analog_sel[30]
port 404 nsew signal input
rlabel metal2 s 41713 531017 42193 531073 6 mprj_io_analog_sel[31]
port 422 nsew signal input
rlabel metal2 s 41713 403417 42193 403473 6 mprj_io_analog_sel[32]
port 440 nsew signal input
rlabel metal2 s 41713 360217 42193 360273 6 mprj_io_analog_sel[33]
port 458 nsew signal input
rlabel metal2 s 41713 317017 42193 317073 6 mprj_io_analog_sel[34]
port 476 nsew signal input
rlabel metal2 s 41713 273817 42193 273873 6 mprj_io_analog_sel[35]
port 494 nsew signal input
rlabel metal2 s 41713 230617 42193 230673 6 mprj_io_analog_sel[36]
port 512 nsew signal input
rlabel metal2 s 41713 187417 42193 187473 6 mprj_io_analog_sel[37]
port 530 nsew signal input
rlabel metal2 s 675407 245527 675887 245583 6 mprj_io_analog_sel[3]
port 227 nsew signal input
rlabel metal2 s 675407 290527 675887 290583 6 mprj_io_analog_sel[4]
port 244 nsew signal input
rlabel metal2 s 675407 335527 675887 335583 6 mprj_io_analog_sel[5]
port 261 nsew signal input
rlabel metal2 s 675407 380727 675887 380783 6 mprj_io_analog_sel[6]
port 278 nsew signal input
rlabel metal2 s 675407 557927 675887 557983 6 mprj_io_analog_sel[7]
port 296 nsew signal input
rlabel metal2 s 675407 603127 675887 603183 6 mprj_io_analog_sel[8]
port 314 nsew signal input
rlabel metal2 s 675407 648127 675887 648183 6 mprj_io_analog_sel[9]
port 332 nsew signal input
rlabel metal2 s 675407 106447 675887 106503 6 mprj_io_dm[0]
port 33 nsew signal input
rlabel metal2 s 41713 365737 42193 365793 6 mprj_io_dm[100]
port 459 nsew signal input
rlabel metal2 s 41713 359573 42193 359629 6 mprj_io_dm[101]
port 460 nsew signal input
rlabel metal2 s 41713 320697 42193 320753 6 mprj_io_dm[102]
port 477 nsew signal input
rlabel metal2 s 41713 322537 42193 322593 6 mprj_io_dm[103]
port 478 nsew signal input
rlabel metal2 s 41713 316373 42193 316429 6 mprj_io_dm[104]
port 479 nsew signal input
rlabel metal2 s 41713 277497 42193 277553 6 mprj_io_dm[105]
port 495 nsew signal input
rlabel metal2 s 41713 279337 42193 279393 6 mprj_io_dm[106]
port 496 nsew signal input
rlabel metal2 s 41713 273173 42193 273229 6 mprj_io_dm[107]
port 497 nsew signal input
rlabel metal2 s 41713 234297 42193 234353 6 mprj_io_dm[108]
port 513 nsew signal input
rlabel metal2 s 41713 236137 42193 236193 6 mprj_io_dm[109]
port 514 nsew signal input
rlabel metal2 s 675407 240007 675887 240063 6 mprj_io_dm[10]
port 228 nsew signal input
rlabel metal2 s 41713 229973 42193 230029 6 mprj_io_dm[110]
port 515 nsew signal input
rlabel metal2 s 41713 191097 42193 191153 6 mprj_io_dm[111]
port 531 nsew signal input
rlabel metal2 s 41713 192937 42193 192993 6 mprj_io_dm[112]
port 532 nsew signal input
rlabel metal2 s 41713 186773 42193 186829 6 mprj_io_dm[113]
port 533 nsew signal input
rlabel metal2 s 675407 246171 675887 246227 6 mprj_io_dm[11]
port 229 nsew signal input
rlabel metal2 s 675407 286847 675887 286903 6 mprj_io_dm[12]
port 245 nsew signal input
rlabel metal2 s 675407 285007 675887 285063 6 mprj_io_dm[13]
port 246 nsew signal input
rlabel metal2 s 675407 291171 675887 291227 6 mprj_io_dm[14]
port 247 nsew signal input
rlabel metal2 s 675407 331847 675887 331903 6 mprj_io_dm[15]
port 262 nsew signal input
rlabel metal2 s 675407 330007 675887 330063 6 mprj_io_dm[16]
port 263 nsew signal input
rlabel metal2 s 675407 336171 675887 336227 6 mprj_io_dm[17]
port 264 nsew signal input
rlabel metal2 s 675407 377047 675887 377103 6 mprj_io_dm[18]
port 279 nsew signal input
rlabel metal2 s 675407 375207 675887 375263 6 mprj_io_dm[19]
port 280 nsew signal input
rlabel metal2 s 675407 104607 675887 104663 6 mprj_io_dm[1]
port 34 nsew signal input
rlabel metal2 s 675407 381371 675887 381427 6 mprj_io_dm[20]
port 281 nsew signal input
rlabel metal2 s 675407 554247 675887 554303 6 mprj_io_dm[21]
port 297 nsew signal input
rlabel metal2 s 675407 552407 675887 552463 6 mprj_io_dm[22]
port 298 nsew signal input
rlabel metal2 s 675407 558571 675887 558627 6 mprj_io_dm[23]
port 299 nsew signal input
rlabel metal2 s 675407 599447 675887 599503 6 mprj_io_dm[24]
port 315 nsew signal input
rlabel metal2 s 675407 597607 675887 597663 6 mprj_io_dm[25]
port 316 nsew signal input
rlabel metal2 s 675407 603771 675887 603827 6 mprj_io_dm[26]
port 317 nsew signal input
rlabel metal2 s 675407 644447 675887 644503 6 mprj_io_dm[27]
port 333 nsew signal input
rlabel metal2 s 675407 642607 675887 642663 6 mprj_io_dm[28]
port 334 nsew signal input
rlabel metal2 s 675407 648771 675887 648827 6 mprj_io_dm[29]
port 335 nsew signal input
rlabel metal2 s 675407 110771 675887 110827 6 mprj_io_dm[2]
port 35 nsew signal input
rlabel metal2 s 675407 689647 675887 689703 6 mprj_io_dm[30]
port 51 nsew signal input
rlabel metal2 s 675407 687807 675887 687863 6 mprj_io_dm[31]
port 52 nsew signal input
rlabel metal2 s 675407 693971 675887 694027 6 mprj_io_dm[32]
port 53 nsew signal input
rlabel metal2 s 675407 734647 675887 734703 6 mprj_io_dm[33]
port 69 nsew signal input
rlabel metal2 s 675407 732807 675887 732863 6 mprj_io_dm[34]
port 70 nsew signal input
rlabel metal2 s 675407 738971 675887 739027 6 mprj_io_dm[35]
port 71 nsew signal input
rlabel metal2 s 675407 779647 675887 779703 6 mprj_io_dm[36]
port 87 nsew signal input
rlabel metal2 s 675407 777807 675887 777863 6 mprj_io_dm[37]
port 88 nsew signal input
rlabel metal2 s 675407 783971 675887 784027 6 mprj_io_dm[38]
port 89 nsew signal input
rlabel metal2 s 675407 868847 675887 868903 6 mprj_io_dm[39]
port 105 nsew signal input
rlabel metal2 s 675407 151647 675887 151703 6 mprj_io_dm[3]
port 194 nsew signal input
rlabel metal2 s 675407 867007 675887 867063 6 mprj_io_dm[40]
port 106 nsew signal input
rlabel metal2 s 675407 873171 675887 873227 6 mprj_io_dm[41]
port 107 nsew signal input
rlabel metal2 s 675407 958047 675887 958103 6 mprj_io_dm[42]
port 123 nsew signal input
rlabel metal2 s 675407 956207 675887 956263 6 mprj_io_dm[43]
port 124 nsew signal input
rlabel metal2 s 675407 962371 675887 962427 6 mprj_io_dm[44]
port 125 nsew signal input
rlabel metal2 s 635497 995407 635553 995887 6 mprj_io_dm[45]
port 141 nsew signal input
rlabel metal2 s 637337 995407 637393 995887 6 mprj_io_dm[46]
port 142 nsew signal input
rlabel metal2 s 631173 995407 631229 995887 6 mprj_io_dm[47]
port 143 nsew signal input
rlabel metal2 s 533697 995407 533753 995887 6 mprj_io_dm[48]
port 159 nsew signal input
rlabel metal2 s 535537 995407 535593 995887 6 mprj_io_dm[49]
port 160 nsew signal input
rlabel metal2 s 675407 149807 675887 149863 6 mprj_io_dm[4]
port 195 nsew signal input
rlabel metal2 s 529373 995407 529429 995887 6 mprj_io_dm[50]
port 161 nsew signal input
rlabel metal2 s 482297 995407 482353 995887 6 mprj_io_dm[51]
port 177 nsew signal input
rlabel metal2 s 484137 995407 484193 995887 6 mprj_io_dm[52]
port 178 nsew signal input
rlabel metal2 s 477973 995407 478029 995887 6 mprj_io_dm[53]
port 179 nsew signal input
rlabel metal2 s 393297 995407 393353 995887 6 mprj_io_dm[54]
port 351 nsew signal input
rlabel metal2 s 395137 995407 395193 995887 6 mprj_io_dm[55]
port 352 nsew signal input
rlabel metal2 s 388973 995407 389029 995887 6 mprj_io_dm[56]
port 353 nsew signal input
rlabel metal2 s 291497 995407 291553 995887 6 mprj_io_dm[57]
port 549 nsew signal input
rlabel metal2 s 293337 995407 293393 995887 6 mprj_io_dm[58]
port 550 nsew signal input
rlabel metal2 s 287173 995407 287229 995887 6 mprj_io_dm[59]
port 551 nsew signal input
rlabel metal2 s 675407 155971 675887 156027 6 mprj_io_dm[5]
port 196 nsew signal input
rlabel metal2 s 239897 995407 239953 995887 6 mprj_io_dm[60]
port 567 nsew signal input
rlabel metal2 s 241737 995407 241793 995887 6 mprj_io_dm[61]
port 568 nsew signal input
rlabel metal2 s 235573 995407 235629 995887 6 mprj_io_dm[62]
port 569 nsew signal input
rlabel metal2 s 188497 995407 188553 995887 6 mprj_io_dm[63]
port 585 nsew signal input
rlabel metal2 s 190337 995407 190393 995887 6 mprj_io_dm[64]
port 586 nsew signal input
rlabel metal2 s 184173 995407 184229 995887 6 mprj_io_dm[65]
port 587 nsew signal input
rlabel metal2 s 137097 995407 137153 995887 6 mprj_io_dm[66]
port 603 nsew signal input
rlabel metal2 s 138937 995407 138993 995887 6 mprj_io_dm[67]
port 604 nsew signal input
rlabel metal2 s 132773 995407 132829 995887 6 mprj_io_dm[68]
port 605 nsew signal input
rlabel metal2 s 85697 995407 85753 995887 6 mprj_io_dm[69]
port 621 nsew signal input
rlabel metal2 s 675407 196647 675887 196703 6 mprj_io_dm[6]
port 211 nsew signal input
rlabel metal2 s 87537 995407 87593 995887 6 mprj_io_dm[70]
port 622 nsew signal input
rlabel metal2 s 81373 995407 81429 995887 6 mprj_io_dm[71]
port 623 nsew signal input
rlabel metal2 s 41713 963697 42193 963753 6 mprj_io_dm[72]
port 639 nsew signal input
rlabel metal2 s 41713 965537 42193 965593 6 mprj_io_dm[73]
port 640 nsew signal input
rlabel metal2 s 41713 959373 42193 959429 6 mprj_io_dm[74]
port 641 nsew signal input
rlabel metal2 s 41713 793897 42193 793953 6 mprj_io_dm[75]
port 657 nsew signal input
rlabel metal2 s 41713 795737 42193 795793 6 mprj_io_dm[76]
port 658 nsew signal input
rlabel metal2 s 41713 789573 42193 789629 6 mprj_io_dm[77]
port 659 nsew signal input
rlabel metal2 s 41713 750697 42193 750753 6 mprj_io_dm[78]
port 675 nsew signal input
rlabel metal2 s 41713 752537 42193 752593 6 mprj_io_dm[79]
port 676 nsew signal input
rlabel metal2 s 675407 194807 675887 194863 6 mprj_io_dm[7]
port 212 nsew signal input
rlabel metal2 s 41713 746373 42193 746429 6 mprj_io_dm[80]
port 677 nsew signal input
rlabel metal2 s 41713 707497 42193 707553 6 mprj_io_dm[81]
port 693 nsew signal input
rlabel metal2 s 41713 709337 42193 709393 6 mprj_io_dm[82]
port 694 nsew signal input
rlabel metal2 s 41713 703173 42193 703229 6 mprj_io_dm[83]
port 695 nsew signal input
rlabel metal2 s 41713 664297 42193 664353 6 mprj_io_dm[84]
port 369 nsew signal input
rlabel metal2 s 41713 666137 42193 666193 6 mprj_io_dm[85]
port 370 nsew signal input
rlabel metal2 s 41713 659973 42193 660029 6 mprj_io_dm[86]
port 371 nsew signal input
rlabel metal2 s 41713 621097 42193 621153 6 mprj_io_dm[87]
port 387 nsew signal input
rlabel metal2 s 41713 622937 42193 622993 6 mprj_io_dm[88]
port 388 nsew signal input
rlabel metal2 s 41713 616773 42193 616829 6 mprj_io_dm[89]
port 389 nsew signal input
rlabel metal2 s 675407 200971 675887 201027 6 mprj_io_dm[8]
port 213 nsew signal input
rlabel metal2 s 41713 577897 42193 577953 6 mprj_io_dm[90]
port 405 nsew signal input
rlabel metal2 s 41713 579737 42193 579793 6 mprj_io_dm[91]
port 406 nsew signal input
rlabel metal2 s 41713 573573 42193 573629 6 mprj_io_dm[92]
port 407 nsew signal input
rlabel metal2 s 41713 534697 42193 534753 6 mprj_io_dm[93]
port 423 nsew signal input
rlabel metal2 s 41713 536537 42193 536593 6 mprj_io_dm[94]
port 424 nsew signal input
rlabel metal2 s 41713 530373 42193 530429 6 mprj_io_dm[95]
port 425 nsew signal input
rlabel metal2 s 41713 407097 42193 407153 6 mprj_io_dm[96]
port 441 nsew signal input
rlabel metal2 s 41713 408937 42193 408993 6 mprj_io_dm[97]
port 442 nsew signal input
rlabel metal2 s 41713 402773 42193 402829 6 mprj_io_dm[98]
port 443 nsew signal input
rlabel metal2 s 41713 363897 42193 363953 6 mprj_io_dm[99]
port 461 nsew signal input
rlabel metal2 s 675407 241847 675887 241903 6 mprj_io_dm[9]
port 230 nsew signal input
rlabel metal2 s 675407 108931 675887 108987 6 mprj_io_enh[0]
port 36 nsew signal input
rlabel metal2 s 675407 692131 675887 692187 6 mprj_io_enh[10]
port 54 nsew signal input
rlabel metal2 s 675407 737131 675887 737187 6 mprj_io_enh[11]
port 72 nsew signal input
rlabel metal2 s 675407 782131 675887 782187 6 mprj_io_enh[12]
port 90 nsew signal input
rlabel metal2 s 675407 871331 675887 871387 6 mprj_io_enh[13]
port 108 nsew signal input
rlabel metal2 s 675407 960531 675887 960587 6 mprj_io_enh[14]
port 126 nsew signal input
rlabel metal2 s 633013 995407 633069 995887 6 mprj_io_enh[15]
port 144 nsew signal input
rlabel metal2 s 531213 995407 531269 995887 6 mprj_io_enh[16]
port 162 nsew signal input
rlabel metal2 s 479813 995407 479869 995887 6 mprj_io_enh[17]
port 180 nsew signal input
rlabel metal2 s 390813 995407 390869 995887 6 mprj_io_enh[18]
port 354 nsew signal input
rlabel metal2 s 289013 995407 289069 995887 6 mprj_io_enh[19]
port 552 nsew signal input
rlabel metal2 s 675407 154131 675887 154187 6 mprj_io_enh[1]
port 197 nsew signal input
rlabel metal2 s 237413 995407 237469 995887 6 mprj_io_enh[20]
port 570 nsew signal input
rlabel metal2 s 186013 995407 186069 995887 6 mprj_io_enh[21]
port 588 nsew signal input
rlabel metal2 s 134613 995407 134669 995887 6 mprj_io_enh[22]
port 606 nsew signal input
rlabel metal2 s 83213 995407 83269 995887 6 mprj_io_enh[23]
port 624 nsew signal input
rlabel metal2 s 41713 961213 42193 961269 6 mprj_io_enh[24]
port 642 nsew signal input
rlabel metal2 s 41713 791413 42193 791469 6 mprj_io_enh[25]
port 660 nsew signal input
rlabel metal2 s 41713 748213 42193 748269 6 mprj_io_enh[26]
port 678 nsew signal input
rlabel metal2 s 41713 705013 42193 705069 6 mprj_io_enh[27]
port 696 nsew signal input
rlabel metal2 s 41713 661813 42193 661869 6 mprj_io_enh[28]
port 372 nsew signal input
rlabel metal2 s 41713 618613 42193 618669 6 mprj_io_enh[29]
port 390 nsew signal input
rlabel metal2 s 675407 199131 675887 199187 6 mprj_io_enh[2]
port 214 nsew signal input
rlabel metal2 s 41713 575413 42193 575469 6 mprj_io_enh[30]
port 408 nsew signal input
rlabel metal2 s 41713 532213 42193 532269 6 mprj_io_enh[31]
port 426 nsew signal input
rlabel metal2 s 41713 404613 42193 404669 6 mprj_io_enh[32]
port 444 nsew signal input
rlabel metal2 s 41713 361413 42193 361469 6 mprj_io_enh[33]
port 462 nsew signal input
rlabel metal2 s 41713 318213 42193 318269 6 mprj_io_enh[34]
port 480 nsew signal input
rlabel metal2 s 41713 275013 42193 275069 6 mprj_io_enh[35]
port 498 nsew signal input
rlabel metal2 s 41713 231813 42193 231869 6 mprj_io_enh[36]
port 516 nsew signal input
rlabel metal2 s 41713 188613 42193 188669 6 mprj_io_enh[37]
port 534 nsew signal input
rlabel metal2 s 675407 244331 675887 244387 6 mprj_io_enh[3]
port 231 nsew signal input
rlabel metal2 s 675407 289331 675887 289387 6 mprj_io_enh[4]
port 248 nsew signal input
rlabel metal2 s 675407 334331 675887 334387 6 mprj_io_enh[5]
port 265 nsew signal input
rlabel metal2 s 675407 379531 675887 379587 6 mprj_io_enh[6]
port 282 nsew signal input
rlabel metal2 s 675407 556731 675887 556787 6 mprj_io_enh[7]
port 300 nsew signal input
rlabel metal2 s 675407 601931 675887 601987 6 mprj_io_enh[8]
port 318 nsew signal input
rlabel metal2 s 675407 646931 675887 646987 6 mprj_io_enh[9]
port 336 nsew signal input
rlabel metal2 s 675407 109575 675887 109631 6 mprj_io_hldh_n[0]
port 37 nsew signal input
rlabel metal2 s 675407 692775 675887 692831 6 mprj_io_hldh_n[10]
port 55 nsew signal input
rlabel metal2 s 675407 737775 675887 737831 6 mprj_io_hldh_n[11]
port 73 nsew signal input
rlabel metal2 s 675407 782775 675887 782831 6 mprj_io_hldh_n[12]
port 91 nsew signal input
rlabel metal2 s 675407 871975 675887 872031 6 mprj_io_hldh_n[13]
port 109 nsew signal input
rlabel metal2 s 675407 961175 675887 961231 6 mprj_io_hldh_n[14]
port 127 nsew signal input
rlabel metal2 s 632369 995407 632425 995887 6 mprj_io_hldh_n[15]
port 145 nsew signal input
rlabel metal2 s 530569 995407 530625 995887 6 mprj_io_hldh_n[16]
port 163 nsew signal input
rlabel metal2 s 479169 995407 479225 995887 6 mprj_io_hldh_n[17]
port 181 nsew signal input
rlabel metal2 s 390169 995407 390225 995887 6 mprj_io_hldh_n[18]
port 355 nsew signal input
rlabel metal2 s 288369 995407 288425 995887 6 mprj_io_hldh_n[19]
port 553 nsew signal input
rlabel metal2 s 675407 154775 675887 154831 6 mprj_io_hldh_n[1]
port 198 nsew signal input
rlabel metal2 s 236769 995407 236825 995887 6 mprj_io_hldh_n[20]
port 571 nsew signal input
rlabel metal2 s 185369 995407 185425 995887 6 mprj_io_hldh_n[21]
port 589 nsew signal input
rlabel metal2 s 133969 995407 134025 995887 6 mprj_io_hldh_n[22]
port 607 nsew signal input
rlabel metal2 s 82569 995407 82625 995887 6 mprj_io_hldh_n[23]
port 625 nsew signal input
rlabel metal2 s 41713 960569 42193 960625 6 mprj_io_hldh_n[24]
port 643 nsew signal input
rlabel metal2 s 41713 790769 42193 790825 6 mprj_io_hldh_n[25]
port 661 nsew signal input
rlabel metal2 s 41713 747569 42193 747625 6 mprj_io_hldh_n[26]
port 679 nsew signal input
rlabel metal2 s 41713 704369 42193 704425 6 mprj_io_hldh_n[27]
port 697 nsew signal input
rlabel metal2 s 41713 661169 42193 661225 6 mprj_io_hldh_n[28]
port 373 nsew signal input
rlabel metal2 s 41713 617969 42193 618025 6 mprj_io_hldh_n[29]
port 391 nsew signal input
rlabel metal2 s 675407 199775 675887 199831 6 mprj_io_hldh_n[2]
port 215 nsew signal input
rlabel metal2 s 41713 574769 42193 574825 6 mprj_io_hldh_n[30]
port 409 nsew signal input
rlabel metal2 s 41713 531569 42193 531625 6 mprj_io_hldh_n[31]
port 427 nsew signal input
rlabel metal2 s 41713 403969 42193 404025 6 mprj_io_hldh_n[32]
port 445 nsew signal input
rlabel metal2 s 41713 360769 42193 360825 6 mprj_io_hldh_n[33]
port 463 nsew signal input
rlabel metal2 s 41713 317569 42193 317625 6 mprj_io_hldh_n[34]
port 481 nsew signal input
rlabel metal2 s 41713 274369 42193 274425 6 mprj_io_hldh_n[35]
port 499 nsew signal input
rlabel metal2 s 41713 231169 42193 231225 6 mprj_io_hldh_n[36]
port 517 nsew signal input
rlabel metal2 s 41713 187969 42193 188025 6 mprj_io_hldh_n[37]
port 535 nsew signal input
rlabel metal2 s 675407 244975 675887 245031 6 mprj_io_hldh_n[3]
port 232 nsew signal input
rlabel metal2 s 675407 289975 675887 290031 6 mprj_io_hldh_n[4]
port 249 nsew signal input
rlabel metal2 s 675407 334975 675887 335031 6 mprj_io_hldh_n[5]
port 266 nsew signal input
rlabel metal2 s 675407 380175 675887 380231 6 mprj_io_hldh_n[6]
port 283 nsew signal input
rlabel metal2 s 675407 557375 675887 557431 6 mprj_io_hldh_n[7]
port 301 nsew signal input
rlabel metal2 s 675407 602575 675887 602631 6 mprj_io_hldh_n[8]
port 319 nsew signal input
rlabel metal2 s 675407 647575 675887 647631 6 mprj_io_hldh_n[9]
port 337 nsew signal input
rlabel metal2 s 675407 111415 675887 111471 6 mprj_io_holdover[0]
port 38 nsew signal input
rlabel metal2 s 675407 694615 675887 694671 6 mprj_io_holdover[10]
port 56 nsew signal input
rlabel metal2 s 675407 739615 675887 739671 6 mprj_io_holdover[11]
port 74 nsew signal input
rlabel metal2 s 675407 784615 675887 784671 6 mprj_io_holdover[12]
port 92 nsew signal input
rlabel metal2 s 675407 873815 675887 873871 6 mprj_io_holdover[13]
port 110 nsew signal input
rlabel metal2 s 675407 963015 675887 963071 6 mprj_io_holdover[14]
port 128 nsew signal input
rlabel metal2 s 630529 995407 630585 995887 6 mprj_io_holdover[15]
port 146 nsew signal input
rlabel metal2 s 528729 995407 528785 995887 6 mprj_io_holdover[16]
port 164 nsew signal input
rlabel metal2 s 477329 995407 477385 995887 6 mprj_io_holdover[17]
port 182 nsew signal input
rlabel metal2 s 388329 995407 388385 995887 6 mprj_io_holdover[18]
port 356 nsew signal input
rlabel metal2 s 286529 995407 286585 995887 6 mprj_io_holdover[19]
port 554 nsew signal input
rlabel metal2 s 675407 156615 675887 156671 6 mprj_io_holdover[1]
port 199 nsew signal input
rlabel metal2 s 234929 995407 234985 995887 6 mprj_io_holdover[20]
port 572 nsew signal input
rlabel metal2 s 183529 995407 183585 995887 6 mprj_io_holdover[21]
port 590 nsew signal input
rlabel metal2 s 132129 995407 132185 995887 6 mprj_io_holdover[22]
port 608 nsew signal input
rlabel metal2 s 80729 995407 80785 995887 6 mprj_io_holdover[23]
port 626 nsew signal input
rlabel metal2 s 41713 958729 42193 958785 6 mprj_io_holdover[24]
port 644 nsew signal input
rlabel metal2 s 41713 788929 42193 788985 6 mprj_io_holdover[25]
port 662 nsew signal input
rlabel metal2 s 41713 745729 42193 745785 6 mprj_io_holdover[26]
port 680 nsew signal input
rlabel metal2 s 41713 702529 42193 702585 6 mprj_io_holdover[27]
port 698 nsew signal input
rlabel metal2 s 41713 659329 42193 659385 6 mprj_io_holdover[28]
port 374 nsew signal input
rlabel metal2 s 41713 616129 42193 616185 6 mprj_io_holdover[29]
port 392 nsew signal input
rlabel metal2 s 675407 201615 675887 201671 6 mprj_io_holdover[2]
port 216 nsew signal input
rlabel metal2 s 41713 572929 42193 572985 6 mprj_io_holdover[30]
port 410 nsew signal input
rlabel metal2 s 41713 529729 42193 529785 6 mprj_io_holdover[31]
port 428 nsew signal input
rlabel metal2 s 41713 402129 42193 402185 6 mprj_io_holdover[32]
port 446 nsew signal input
rlabel metal2 s 41713 358929 42193 358985 6 mprj_io_holdover[33]
port 464 nsew signal input
rlabel metal2 s 41713 315729 42193 315785 6 mprj_io_holdover[34]
port 482 nsew signal input
rlabel metal2 s 41713 272529 42193 272585 6 mprj_io_holdover[35]
port 500 nsew signal input
rlabel metal2 s 41713 229329 42193 229385 6 mprj_io_holdover[36]
port 518 nsew signal input
rlabel metal2 s 41713 186129 42193 186185 6 mprj_io_holdover[37]
port 536 nsew signal input
rlabel metal2 s 675407 246815 675887 246871 6 mprj_io_holdover[3]
port 233 nsew signal input
rlabel metal2 s 675407 291815 675887 291871 6 mprj_io_holdover[4]
port 250 nsew signal input
rlabel metal2 s 675407 336815 675887 336871 6 mprj_io_holdover[5]
port 267 nsew signal input
rlabel metal2 s 675407 382015 675887 382071 6 mprj_io_holdover[6]
port 284 nsew signal input
rlabel metal2 s 675407 559215 675887 559271 6 mprj_io_holdover[7]
port 302 nsew signal input
rlabel metal2 s 675407 604415 675887 604471 6 mprj_io_holdover[8]
port 320 nsew signal input
rlabel metal2 s 675407 649415 675887 649471 6 mprj_io_holdover[9]
port 338 nsew signal input
rlabel metal2 s 675407 114451 675887 114507 6 mprj_io_ib_mode_sel[0]
port 39 nsew signal input
rlabel metal2 s 675407 697651 675887 697707 6 mprj_io_ib_mode_sel[10]
port 57 nsew signal input
rlabel metal2 s 675407 742651 675887 742707 6 mprj_io_ib_mode_sel[11]
port 75 nsew signal input
rlabel metal2 s 675407 787651 675887 787707 6 mprj_io_ib_mode_sel[12]
port 93 nsew signal input
rlabel metal2 s 675407 876851 675887 876907 6 mprj_io_ib_mode_sel[13]
port 111 nsew signal input
rlabel metal2 s 675407 966051 675887 966107 6 mprj_io_ib_mode_sel[14]
port 129 nsew signal input
rlabel metal2 s 627493 995407 627549 995887 6 mprj_io_ib_mode_sel[15]
port 147 nsew signal input
rlabel metal2 s 525693 995407 525749 995887 6 mprj_io_ib_mode_sel[16]
port 165 nsew signal input
rlabel metal2 s 474293 995407 474349 995887 6 mprj_io_ib_mode_sel[17]
port 183 nsew signal input
rlabel metal2 s 385293 995407 385349 995887 6 mprj_io_ib_mode_sel[18]
port 357 nsew signal input
rlabel metal2 s 283493 995407 283549 995887 6 mprj_io_ib_mode_sel[19]
port 555 nsew signal input
rlabel metal2 s 675407 159651 675887 159707 6 mprj_io_ib_mode_sel[1]
port 200 nsew signal input
rlabel metal2 s 231893 995407 231949 995887 6 mprj_io_ib_mode_sel[20]
port 573 nsew signal input
rlabel metal2 s 180493 995407 180549 995887 6 mprj_io_ib_mode_sel[21]
port 591 nsew signal input
rlabel metal2 s 129093 995407 129149 995887 6 mprj_io_ib_mode_sel[22]
port 609 nsew signal input
rlabel metal2 s 77693 995407 77749 995887 6 mprj_io_ib_mode_sel[23]
port 627 nsew signal input
rlabel metal2 s 41713 955693 42193 955749 6 mprj_io_ib_mode_sel[24]
port 645 nsew signal input
rlabel metal2 s 41713 785893 42193 785949 6 mprj_io_ib_mode_sel[25]
port 663 nsew signal input
rlabel metal2 s 41713 742693 42193 742749 6 mprj_io_ib_mode_sel[26]
port 681 nsew signal input
rlabel metal2 s 41713 699493 42193 699549 6 mprj_io_ib_mode_sel[27]
port 699 nsew signal input
rlabel metal2 s 41713 656293 42193 656349 6 mprj_io_ib_mode_sel[28]
port 375 nsew signal input
rlabel metal2 s 41713 613093 42193 613149 6 mprj_io_ib_mode_sel[29]
port 393 nsew signal input
rlabel metal2 s 675407 204651 675887 204707 6 mprj_io_ib_mode_sel[2]
port 217 nsew signal input
rlabel metal2 s 41713 569893 42193 569949 6 mprj_io_ib_mode_sel[30]
port 411 nsew signal input
rlabel metal2 s 41713 526693 42193 526749 6 mprj_io_ib_mode_sel[31]
port 429 nsew signal input
rlabel metal2 s 41713 399093 42193 399149 6 mprj_io_ib_mode_sel[32]
port 447 nsew signal input
rlabel metal2 s 41713 355893 42193 355949 6 mprj_io_ib_mode_sel[33]
port 465 nsew signal input
rlabel metal2 s 41713 312693 42193 312749 6 mprj_io_ib_mode_sel[34]
port 483 nsew signal input
rlabel metal2 s 41713 269493 42193 269549 6 mprj_io_ib_mode_sel[35]
port 501 nsew signal input
rlabel metal2 s 41713 226293 42193 226349 6 mprj_io_ib_mode_sel[36]
port 519 nsew signal input
rlabel metal2 s 41713 183093 42193 183149 6 mprj_io_ib_mode_sel[37]
port 537 nsew signal input
rlabel metal2 s 675407 249851 675887 249907 6 mprj_io_ib_mode_sel[3]
port 234 nsew signal input
rlabel metal2 s 675407 294851 675887 294907 6 mprj_io_ib_mode_sel[4]
port 251 nsew signal input
rlabel metal2 s 675407 339851 675887 339907 6 mprj_io_ib_mode_sel[5]
port 268 nsew signal input
rlabel metal2 s 675407 385051 675887 385107 6 mprj_io_ib_mode_sel[6]
port 285 nsew signal input
rlabel metal2 s 675407 562251 675887 562307 6 mprj_io_ib_mode_sel[7]
port 303 nsew signal input
rlabel metal2 s 675407 607451 675887 607507 6 mprj_io_ib_mode_sel[8]
port 321 nsew signal input
rlabel metal2 s 675407 652451 675887 652507 6 mprj_io_ib_mode_sel[9]
port 339 nsew signal input
rlabel metal2 s 675407 100927 675887 100983 6 mprj_io_in[0]
port 45 nsew signal output
rlabel metal2 s 675407 684127 675887 684183 6 mprj_io_in[10]
port 63 nsew signal output
rlabel metal2 s 675407 729127 675887 729183 6 mprj_io_in[11]
port 81 nsew signal output
rlabel metal2 s 675407 774127 675887 774183 6 mprj_io_in[12]
port 99 nsew signal output
rlabel metal2 s 675407 863327 675887 863383 6 mprj_io_in[13]
port 117 nsew signal output
rlabel metal2 s 675407 952527 675887 952583 6 mprj_io_in[14]
port 135 nsew signal output
rlabel metal2 s 641017 995407 641073 995887 6 mprj_io_in[15]
port 153 nsew signal output
rlabel metal2 s 539217 995407 539273 995887 6 mprj_io_in[16]
port 171 nsew signal output
rlabel metal2 s 487817 995407 487873 995887 6 mprj_io_in[17]
port 189 nsew signal output
rlabel metal2 s 398817 995407 398873 995887 6 mprj_io_in[18]
port 363 nsew signal output
rlabel metal2 s 297017 995407 297073 995887 6 mprj_io_in[19]
port 561 nsew signal output
rlabel metal2 s 675407 146127 675887 146183 6 mprj_io_in[1]
port 206 nsew signal output
rlabel metal2 s 245417 995407 245473 995887 6 mprj_io_in[20]
port 579 nsew signal output
rlabel metal2 s 194017 995407 194073 995887 6 mprj_io_in[21]
port 597 nsew signal output
rlabel metal2 s 142617 995407 142673 995887 6 mprj_io_in[22]
port 615 nsew signal output
rlabel metal2 s 91217 995407 91273 995887 6 mprj_io_in[23]
port 633 nsew signal output
rlabel metal2 s 41713 969217 42193 969273 6 mprj_io_in[24]
port 651 nsew signal output
rlabel metal2 s 41713 799417 42193 799473 6 mprj_io_in[25]
port 669 nsew signal output
rlabel metal2 s 41713 756217 42193 756273 6 mprj_io_in[26]
port 687 nsew signal output
rlabel metal2 s 41713 713017 42193 713073 6 mprj_io_in[27]
port 705 nsew signal output
rlabel metal2 s 41713 669817 42193 669873 6 mprj_io_in[28]
port 381 nsew signal output
rlabel metal2 s 41713 626617 42193 626673 6 mprj_io_in[29]
port 399 nsew signal output
rlabel metal2 s 675407 191127 675887 191183 6 mprj_io_in[2]
port 223 nsew signal output
rlabel metal2 s 41713 583417 42193 583473 6 mprj_io_in[30]
port 417 nsew signal output
rlabel metal2 s 41713 540217 42193 540273 6 mprj_io_in[31]
port 435 nsew signal output
rlabel metal2 s 41713 412617 42193 412673 6 mprj_io_in[32]
port 453 nsew signal output
rlabel metal2 s 41713 369417 42193 369473 6 mprj_io_in[33]
port 471 nsew signal output
rlabel metal2 s 41713 326217 42193 326273 6 mprj_io_in[34]
port 489 nsew signal output
rlabel metal2 s 41713 283017 42193 283073 6 mprj_io_in[35]
port 507 nsew signal output
rlabel metal2 s 41713 239817 42193 239873 6 mprj_io_in[36]
port 525 nsew signal output
rlabel metal2 s 41713 196617 42193 196673 6 mprj_io_in[37]
port 543 nsew signal output
rlabel metal2 s 675407 236327 675887 236383 6 mprj_io_in[3]
port 240 nsew signal output
rlabel metal2 s 675407 281327 675887 281383 6 mprj_io_in[4]
port 257 nsew signal output
rlabel metal2 s 675407 326327 675887 326383 6 mprj_io_in[5]
port 274 nsew signal output
rlabel metal2 s 675407 371527 675887 371583 6 mprj_io_in[6]
port 291 nsew signal output
rlabel metal2 s 675407 548727 675887 548783 6 mprj_io_in[7]
port 309 nsew signal output
rlabel metal2 s 675407 593927 675887 593983 6 mprj_io_in[8]
port 327 nsew signal output
rlabel metal2 s 675407 638927 675887 638983 6 mprj_io_in[9]
port 345 nsew signal output
rlabel metal2 s 675407 107643 675887 107699 6 mprj_io_inp_dis[0]
port 40 nsew signal input
rlabel metal2 s 675407 690843 675887 690899 6 mprj_io_inp_dis[10]
port 58 nsew signal input
rlabel metal2 s 675407 735843 675887 735899 6 mprj_io_inp_dis[11]
port 76 nsew signal input
rlabel metal2 s 675407 780843 675887 780899 6 mprj_io_inp_dis[12]
port 94 nsew signal input
rlabel metal2 s 675407 870043 675887 870099 6 mprj_io_inp_dis[13]
port 112 nsew signal input
rlabel metal2 s 675407 959243 675887 959299 6 mprj_io_inp_dis[14]
port 130 nsew signal input
rlabel metal2 s 634301 995407 634357 995887 6 mprj_io_inp_dis[15]
port 148 nsew signal input
rlabel metal2 s 532501 995407 532557 995887 6 mprj_io_inp_dis[16]
port 166 nsew signal input
rlabel metal2 s 481101 995407 481157 995887 6 mprj_io_inp_dis[17]
port 184 nsew signal input
rlabel metal2 s 392101 995407 392157 995887 6 mprj_io_inp_dis[18]
port 358 nsew signal input
rlabel metal2 s 290301 995407 290357 995887 6 mprj_io_inp_dis[19]
port 556 nsew signal input
rlabel metal2 s 675407 152843 675887 152899 6 mprj_io_inp_dis[1]
port 201 nsew signal input
rlabel metal2 s 238701 995407 238757 995887 6 mprj_io_inp_dis[20]
port 574 nsew signal input
rlabel metal2 s 187301 995407 187357 995887 6 mprj_io_inp_dis[21]
port 592 nsew signal input
rlabel metal2 s 135901 995407 135957 995887 6 mprj_io_inp_dis[22]
port 610 nsew signal input
rlabel metal2 s 84501 995407 84557 995887 6 mprj_io_inp_dis[23]
port 628 nsew signal input
rlabel metal2 s 41713 962501 42193 962557 6 mprj_io_inp_dis[24]
port 646 nsew signal input
rlabel metal2 s 41713 792701 42193 792757 6 mprj_io_inp_dis[25]
port 664 nsew signal input
rlabel metal2 s 41713 749501 42193 749557 6 mprj_io_inp_dis[26]
port 682 nsew signal input
rlabel metal2 s 41713 706301 42193 706357 6 mprj_io_inp_dis[27]
port 700 nsew signal input
rlabel metal2 s 41713 663101 42193 663157 6 mprj_io_inp_dis[28]
port 376 nsew signal input
rlabel metal2 s 41713 619901 42193 619957 6 mprj_io_inp_dis[29]
port 394 nsew signal input
rlabel metal2 s 675407 197843 675887 197899 6 mprj_io_inp_dis[2]
port 218 nsew signal input
rlabel metal2 s 41713 576701 42193 576757 6 mprj_io_inp_dis[30]
port 412 nsew signal input
rlabel metal2 s 41713 533501 42193 533557 6 mprj_io_inp_dis[31]
port 430 nsew signal input
rlabel metal2 s 41713 405901 42193 405957 6 mprj_io_inp_dis[32]
port 448 nsew signal input
rlabel metal2 s 41713 362701 42193 362757 6 mprj_io_inp_dis[33]
port 466 nsew signal input
rlabel metal2 s 41713 319501 42193 319557 6 mprj_io_inp_dis[34]
port 484 nsew signal input
rlabel metal2 s 41713 276301 42193 276357 6 mprj_io_inp_dis[35]
port 502 nsew signal input
rlabel metal2 s 41713 233101 42193 233157 6 mprj_io_inp_dis[36]
port 520 nsew signal input
rlabel metal2 s 41713 189901 42193 189957 6 mprj_io_inp_dis[37]
port 538 nsew signal input
rlabel metal2 s 675407 243043 675887 243099 6 mprj_io_inp_dis[3]
port 235 nsew signal input
rlabel metal2 s 675407 288043 675887 288099 6 mprj_io_inp_dis[4]
port 252 nsew signal input
rlabel metal2 s 675407 333043 675887 333099 6 mprj_io_inp_dis[5]
port 269 nsew signal input
rlabel metal2 s 675407 378243 675887 378299 6 mprj_io_inp_dis[6]
port 286 nsew signal input
rlabel metal2 s 675407 555443 675887 555499 6 mprj_io_inp_dis[7]
port 304 nsew signal input
rlabel metal2 s 675407 600643 675887 600699 6 mprj_io_inp_dis[8]
port 322 nsew signal input
rlabel metal2 s 675407 645643 675887 645699 6 mprj_io_inp_dis[9]
port 340 nsew signal input
rlabel metal2 s 675407 115095 675887 115151 6 mprj_io_oeb[0]
port 41 nsew signal input
rlabel metal2 s 675407 698295 675887 698351 6 mprj_io_oeb[10]
port 59 nsew signal input
rlabel metal2 s 675407 743295 675887 743351 6 mprj_io_oeb[11]
port 77 nsew signal input
rlabel metal2 s 675407 788295 675887 788351 6 mprj_io_oeb[12]
port 95 nsew signal input
rlabel metal2 s 675407 877495 675887 877551 6 mprj_io_oeb[13]
port 113 nsew signal input
rlabel metal2 s 675407 966695 675887 966751 6 mprj_io_oeb[14]
port 131 nsew signal input
rlabel metal2 s 626849 995407 626905 995887 6 mprj_io_oeb[15]
port 149 nsew signal input
rlabel metal2 s 525049 995407 525105 995887 6 mprj_io_oeb[16]
port 167 nsew signal input
rlabel metal2 s 473649 995407 473705 995887 6 mprj_io_oeb[17]
port 185 nsew signal input
rlabel metal2 s 384649 995407 384705 995887 6 mprj_io_oeb[18]
port 359 nsew signal input
rlabel metal2 s 282849 995407 282905 995887 6 mprj_io_oeb[19]
port 557 nsew signal input
rlabel metal2 s 675407 160295 675887 160351 6 mprj_io_oeb[1]
port 202 nsew signal input
rlabel metal2 s 231249 995407 231305 995887 6 mprj_io_oeb[20]
port 575 nsew signal input
rlabel metal2 s 179849 995407 179905 995887 6 mprj_io_oeb[21]
port 593 nsew signal input
rlabel metal2 s 128449 995407 128505 995887 6 mprj_io_oeb[22]
port 611 nsew signal input
rlabel metal2 s 77049 995407 77105 995887 6 mprj_io_oeb[23]
port 629 nsew signal input
rlabel metal2 s 41713 955049 42193 955105 6 mprj_io_oeb[24]
port 647 nsew signal input
rlabel metal2 s 41713 785249 42193 785305 6 mprj_io_oeb[25]
port 665 nsew signal input
rlabel metal2 s 41713 742049 42193 742105 6 mprj_io_oeb[26]
port 683 nsew signal input
rlabel metal2 s 41713 698849 42193 698905 6 mprj_io_oeb[27]
port 701 nsew signal input
rlabel metal2 s 41713 655649 42193 655705 6 mprj_io_oeb[28]
port 377 nsew signal input
rlabel metal2 s 41713 612449 42193 612505 6 mprj_io_oeb[29]
port 395 nsew signal input
rlabel metal2 s 675407 205295 675887 205351 6 mprj_io_oeb[2]
port 219 nsew signal input
rlabel metal2 s 41713 569249 42193 569305 6 mprj_io_oeb[30]
port 413 nsew signal input
rlabel metal2 s 41713 526049 42193 526105 6 mprj_io_oeb[31]
port 431 nsew signal input
rlabel metal2 s 41713 398449 42193 398505 6 mprj_io_oeb[32]
port 449 nsew signal input
rlabel metal2 s 41713 355249 42193 355305 6 mprj_io_oeb[33]
port 467 nsew signal input
rlabel metal2 s 41713 312049 42193 312105 6 mprj_io_oeb[34]
port 485 nsew signal input
rlabel metal2 s 41713 268849 42193 268905 6 mprj_io_oeb[35]
port 503 nsew signal input
rlabel metal2 s 41713 225649 42193 225705 6 mprj_io_oeb[36]
port 521 nsew signal input
rlabel metal2 s 41713 182449 42193 182505 6 mprj_io_oeb[37]
port 539 nsew signal input
rlabel metal2 s 675407 250495 675887 250551 6 mprj_io_oeb[3]
port 236 nsew signal input
rlabel metal2 s 675407 295495 675887 295551 6 mprj_io_oeb[4]
port 253 nsew signal input
rlabel metal2 s 675407 340495 675887 340551 6 mprj_io_oeb[5]
port 270 nsew signal input
rlabel metal2 s 675407 385695 675887 385751 6 mprj_io_oeb[6]
port 287 nsew signal input
rlabel metal2 s 675407 562895 675887 562951 6 mprj_io_oeb[7]
port 305 nsew signal input
rlabel metal2 s 675407 608095 675887 608151 6 mprj_io_oeb[8]
port 323 nsew signal input
rlabel metal2 s 675407 653095 675887 653151 6 mprj_io_oeb[9]
port 341 nsew signal input
rlabel metal2 s 675407 111967 675887 112023 6 mprj_io_out[0]
port 42 nsew signal input
rlabel metal2 s 675407 695167 675887 695223 6 mprj_io_out[10]
port 60 nsew signal input
rlabel metal2 s 675407 740167 675887 740223 6 mprj_io_out[11]
port 78 nsew signal input
rlabel metal2 s 675407 785167 675887 785223 6 mprj_io_out[12]
port 96 nsew signal input
rlabel metal2 s 675407 874367 675887 874423 6 mprj_io_out[13]
port 114 nsew signal input
rlabel metal2 s 675407 963567 675887 963623 6 mprj_io_out[14]
port 132 nsew signal input
rlabel metal2 s 629977 995407 630033 995887 6 mprj_io_out[15]
port 150 nsew signal input
rlabel metal2 s 528177 995407 528233 995887 6 mprj_io_out[16]
port 168 nsew signal input
rlabel metal2 s 476777 995407 476833 995887 6 mprj_io_out[17]
port 186 nsew signal input
rlabel metal2 s 387777 995407 387833 995887 6 mprj_io_out[18]
port 360 nsew signal input
rlabel metal2 s 285977 995407 286033 995887 6 mprj_io_out[19]
port 558 nsew signal input
rlabel metal2 s 675407 157167 675887 157223 6 mprj_io_out[1]
port 203 nsew signal input
rlabel metal2 s 234377 995407 234433 995887 6 mprj_io_out[20]
port 576 nsew signal input
rlabel metal2 s 182977 995407 183033 995887 6 mprj_io_out[21]
port 594 nsew signal input
rlabel metal2 s 131577 995407 131633 995887 6 mprj_io_out[22]
port 612 nsew signal input
rlabel metal2 s 80177 995407 80233 995887 6 mprj_io_out[23]
port 630 nsew signal input
rlabel metal2 s 41713 958177 42193 958233 6 mprj_io_out[24]
port 648 nsew signal input
rlabel metal2 s 41713 788377 42193 788433 6 mprj_io_out[25]
port 666 nsew signal input
rlabel metal2 s 41713 745177 42193 745233 6 mprj_io_out[26]
port 684 nsew signal input
rlabel metal2 s 41713 701977 42193 702033 6 mprj_io_out[27]
port 702 nsew signal input
rlabel metal2 s 41713 658777 42193 658833 6 mprj_io_out[28]
port 378 nsew signal input
rlabel metal2 s 41713 615577 42193 615633 6 mprj_io_out[29]
port 396 nsew signal input
rlabel metal2 s 675407 202167 675887 202223 6 mprj_io_out[2]
port 220 nsew signal input
rlabel metal2 s 41713 572377 42193 572433 6 mprj_io_out[30]
port 414 nsew signal input
rlabel metal2 s 41713 529177 42193 529233 6 mprj_io_out[31]
port 432 nsew signal input
rlabel metal2 s 41713 401577 42193 401633 6 mprj_io_out[32]
port 450 nsew signal input
rlabel metal2 s 41713 358377 42193 358433 6 mprj_io_out[33]
port 468 nsew signal input
rlabel metal2 s 41713 315177 42193 315233 6 mprj_io_out[34]
port 486 nsew signal input
rlabel metal2 s 41713 271977 42193 272033 6 mprj_io_out[35]
port 504 nsew signal input
rlabel metal2 s 41713 228777 42193 228833 6 mprj_io_out[36]
port 522 nsew signal input
rlabel metal2 s 41713 185577 42193 185633 6 mprj_io_out[37]
port 540 nsew signal input
rlabel metal2 s 675407 247367 675887 247423 6 mprj_io_out[3]
port 237 nsew signal input
rlabel metal2 s 675407 292367 675887 292423 6 mprj_io_out[4]
port 254 nsew signal input
rlabel metal2 s 675407 337367 675887 337423 6 mprj_io_out[5]
port 271 nsew signal input
rlabel metal2 s 675407 382567 675887 382623 6 mprj_io_out[6]
port 288 nsew signal input
rlabel metal2 s 675407 559767 675887 559823 6 mprj_io_out[7]
port 306 nsew signal input
rlabel metal2 s 675407 604967 675887 605023 6 mprj_io_out[8]
port 324 nsew signal input
rlabel metal2 s 675407 649967 675887 650023 6 mprj_io_out[9]
port 342 nsew signal input
rlabel metal2 s 675407 102767 675887 102823 6 mprj_io_slow_sel[0]
port 43 nsew signal input
rlabel metal2 s 675407 685967 675887 686023 6 mprj_io_slow_sel[10]
port 61 nsew signal input
rlabel metal2 s 675407 730967 675887 731023 6 mprj_io_slow_sel[11]
port 79 nsew signal input
rlabel metal2 s 675407 775967 675887 776023 6 mprj_io_slow_sel[12]
port 97 nsew signal input
rlabel metal2 s 675407 865167 675887 865223 6 mprj_io_slow_sel[13]
port 115 nsew signal input
rlabel metal2 s 675407 954367 675887 954423 6 mprj_io_slow_sel[14]
port 133 nsew signal input
rlabel metal2 s 639177 995407 639233 995887 6 mprj_io_slow_sel[15]
port 151 nsew signal input
rlabel metal2 s 537377 995407 537433 995887 6 mprj_io_slow_sel[16]
port 169 nsew signal input
rlabel metal2 s 485977 995407 486033 995887 6 mprj_io_slow_sel[17]
port 187 nsew signal input
rlabel metal2 s 396977 995407 397033 995887 6 mprj_io_slow_sel[18]
port 361 nsew signal input
rlabel metal2 s 295177 995407 295233 995887 6 mprj_io_slow_sel[19]
port 559 nsew signal input
rlabel metal2 s 675407 147967 675887 148023 6 mprj_io_slow_sel[1]
port 204 nsew signal input
rlabel metal2 s 243577 995407 243633 995887 6 mprj_io_slow_sel[20]
port 577 nsew signal input
rlabel metal2 s 192177 995407 192233 995887 6 mprj_io_slow_sel[21]
port 595 nsew signal input
rlabel metal2 s 140777 995407 140833 995887 6 mprj_io_slow_sel[22]
port 613 nsew signal input
rlabel metal2 s 89377 995407 89433 995887 6 mprj_io_slow_sel[23]
port 631 nsew signal input
rlabel metal2 s 41713 967377 42193 967433 6 mprj_io_slow_sel[24]
port 649 nsew signal input
rlabel metal2 s 41713 797577 42193 797633 6 mprj_io_slow_sel[25]
port 667 nsew signal input
rlabel metal2 s 41713 754377 42193 754433 6 mprj_io_slow_sel[26]
port 685 nsew signal input
rlabel metal2 s 41713 711177 42193 711233 6 mprj_io_slow_sel[27]
port 703 nsew signal input
rlabel metal2 s 41713 667977 42193 668033 6 mprj_io_slow_sel[28]
port 379 nsew signal input
rlabel metal2 s 41713 624777 42193 624833 6 mprj_io_slow_sel[29]
port 397 nsew signal input
rlabel metal2 s 675407 192967 675887 193023 6 mprj_io_slow_sel[2]
port 221 nsew signal input
rlabel metal2 s 41713 581577 42193 581633 6 mprj_io_slow_sel[30]
port 415 nsew signal input
rlabel metal2 s 41713 538377 42193 538433 6 mprj_io_slow_sel[31]
port 433 nsew signal input
rlabel metal2 s 41713 410777 42193 410833 6 mprj_io_slow_sel[32]
port 451 nsew signal input
rlabel metal2 s 41713 367577 42193 367633 6 mprj_io_slow_sel[33]
port 469 nsew signal input
rlabel metal2 s 41713 324377 42193 324433 6 mprj_io_slow_sel[34]
port 487 nsew signal input
rlabel metal2 s 41713 281177 42193 281233 6 mprj_io_slow_sel[35]
port 505 nsew signal input
rlabel metal2 s 41713 237977 42193 238033 6 mprj_io_slow_sel[36]
port 523 nsew signal input
rlabel metal2 s 41713 194777 42193 194833 6 mprj_io_slow_sel[37]
port 541 nsew signal input
rlabel metal2 s 675407 238167 675887 238223 6 mprj_io_slow_sel[3]
port 238 nsew signal input
rlabel metal2 s 675407 283167 675887 283223 6 mprj_io_slow_sel[4]
port 255 nsew signal input
rlabel metal2 s 675407 328167 675887 328223 6 mprj_io_slow_sel[5]
port 272 nsew signal input
rlabel metal2 s 675407 373367 675887 373423 6 mprj_io_slow_sel[6]
port 289 nsew signal input
rlabel metal2 s 675407 550567 675887 550623 6 mprj_io_slow_sel[7]
port 307 nsew signal input
rlabel metal2 s 675407 595767 675887 595823 6 mprj_io_slow_sel[8]
port 325 nsew signal input
rlabel metal2 s 675407 640767 675887 640823 6 mprj_io_slow_sel[9]
port 343 nsew signal input
rlabel metal2 s 675407 113807 675887 113863 6 mprj_io_vtrip_sel[0]
port 44 nsew signal input
rlabel metal2 s 675407 697007 675887 697063 6 mprj_io_vtrip_sel[10]
port 62 nsew signal input
rlabel metal2 s 675407 742007 675887 742063 6 mprj_io_vtrip_sel[11]
port 80 nsew signal input
rlabel metal2 s 675407 787007 675887 787063 6 mprj_io_vtrip_sel[12]
port 98 nsew signal input
rlabel metal2 s 675407 876207 675887 876263 6 mprj_io_vtrip_sel[13]
port 116 nsew signal input
rlabel metal2 s 675407 965407 675887 965463 6 mprj_io_vtrip_sel[14]
port 134 nsew signal input
rlabel metal2 s 628137 995407 628193 995887 6 mprj_io_vtrip_sel[15]
port 152 nsew signal input
rlabel metal2 s 526337 995407 526393 995887 6 mprj_io_vtrip_sel[16]
port 170 nsew signal input
rlabel metal2 s 474937 995407 474993 995887 6 mprj_io_vtrip_sel[17]
port 188 nsew signal input
rlabel metal2 s 385937 995407 385993 995887 6 mprj_io_vtrip_sel[18]
port 362 nsew signal input
rlabel metal2 s 284137 995407 284193 995887 6 mprj_io_vtrip_sel[19]
port 560 nsew signal input
rlabel metal2 s 675407 159007 675887 159063 6 mprj_io_vtrip_sel[1]
port 205 nsew signal input
rlabel metal2 s 232537 995407 232593 995887 6 mprj_io_vtrip_sel[20]
port 578 nsew signal input
rlabel metal2 s 181137 995407 181193 995887 6 mprj_io_vtrip_sel[21]
port 596 nsew signal input
rlabel metal2 s 129737 995407 129793 995887 6 mprj_io_vtrip_sel[22]
port 614 nsew signal input
rlabel metal2 s 78337 995407 78393 995887 6 mprj_io_vtrip_sel[23]
port 632 nsew signal input
rlabel metal2 s 41713 956337 42193 956393 6 mprj_io_vtrip_sel[24]
port 650 nsew signal input
rlabel metal2 s 41713 786537 42193 786593 6 mprj_io_vtrip_sel[25]
port 668 nsew signal input
rlabel metal2 s 41713 743337 42193 743393 6 mprj_io_vtrip_sel[26]
port 686 nsew signal input
rlabel metal2 s 41713 700137 42193 700193 6 mprj_io_vtrip_sel[27]
port 704 nsew signal input
rlabel metal2 s 41713 656937 42193 656993 6 mprj_io_vtrip_sel[28]
port 380 nsew signal input
rlabel metal2 s 41713 613737 42193 613793 6 mprj_io_vtrip_sel[29]
port 398 nsew signal input
rlabel metal2 s 675407 204007 675887 204063 6 mprj_io_vtrip_sel[2]
port 222 nsew signal input
rlabel metal2 s 41713 570537 42193 570593 6 mprj_io_vtrip_sel[30]
port 416 nsew signal input
rlabel metal2 s 41713 527337 42193 527393 6 mprj_io_vtrip_sel[31]
port 434 nsew signal input
rlabel metal2 s 41713 399737 42193 399793 6 mprj_io_vtrip_sel[32]
port 452 nsew signal input
rlabel metal2 s 41713 356537 42193 356593 6 mprj_io_vtrip_sel[33]
port 470 nsew signal input
rlabel metal2 s 41713 313337 42193 313393 6 mprj_io_vtrip_sel[34]
port 488 nsew signal input
rlabel metal2 s 41713 270137 42193 270193 6 mprj_io_vtrip_sel[35]
port 506 nsew signal input
rlabel metal2 s 41713 226937 42193 226993 6 mprj_io_vtrip_sel[36]
port 524 nsew signal input
rlabel metal2 s 41713 183737 42193 183793 6 mprj_io_vtrip_sel[37]
port 542 nsew signal input
rlabel metal2 s 675407 249207 675887 249263 6 mprj_io_vtrip_sel[3]
port 239 nsew signal input
rlabel metal2 s 675407 294207 675887 294263 6 mprj_io_vtrip_sel[4]
port 256 nsew signal input
rlabel metal2 s 675407 339207 675887 339263 6 mprj_io_vtrip_sel[5]
port 273 nsew signal input
rlabel metal2 s 675407 384407 675887 384463 6 mprj_io_vtrip_sel[6]
port 290 nsew signal input
rlabel metal2 s 675407 561607 675887 561663 6 mprj_io_vtrip_sel[7]
port 308 nsew signal input
rlabel metal2 s 675407 606807 675887 606863 6 mprj_io_vtrip_sel[8]
port 326 nsew signal input
rlabel metal2 s 675407 651807 675887 651863 6 mprj_io_vtrip_sel[9]
port 344 nsew signal input
rlabel metal2 s 194043 41713 194099 42193 6 por
port 3 nsew signal input
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 1580 nsew signal input
rlabel metal2 s 145091 39934 145143 40000 6 porb_h
port 1580 nsew signal input
rlabel metal1 s 145091 39934 145143 40000 6 porb_h
port 1580 nsew signal input
rlabel metal5 s 136703 7133 144159 18319 6 resetb
port 706 nsew signal input
rlabel metal3 s 141667 37818 141813 39199 6 resetb_core_h
port 1582 nsew signal output
rlabel metal3 s 141667 38031 141813 39999 6 resetb_core_h
port 1582 nsew signal output
rlabel metal3 s 141667 39934 141813 40000 6 resetb_core_h
port 1582 nsew signal output
rlabel metal2 s 141667 39934 141813 40000 6 resetb_core_h
port 1582 nsew signal output
rlabel metal4 s 37293 68000 38223 68254 6 vccd
port 1583 nsew signal bidirectional
rlabel metal4 s 37293 82746 38223 83000 6 vccd
port 1583 nsew signal bidirectional
rlabel metal5 s 37313 68000 38203 68254 6 vccd
port 1583 nsew signal bidirectional
rlabel metal5 s 37313 82746 38203 83000 6 vccd
port 1583 nsew signal bidirectional
rlabel metal3 s 38220 68100 39600 72900 6 vccd
port 1583 nsew signal bidirectional
rlabel metal3 s 38220 78151 39600 82940 6 vccd
port 1583 nsew signal bidirectional
rlabel metal4 s 679377 922346 680307 922600 6 vccd1
port 1584 nsew signal bidirectional
rlabel metal4 s 679377 907600 680307 907854 6 vccd1
port 1584 nsew signal bidirectional
rlabel metal5 s 679397 922346 680287 922600 6 vccd1
port 1584 nsew signal bidirectional
rlabel metal5 s 679397 907600 680287 907854 6 vccd1
port 1584 nsew signal bidirectional
rlabel metal3 s 678000 917700 679380 922500 6 vccd1
port 1584 nsew signal bidirectional
rlabel metal3 s 678000 907660 679380 912449 6 vccd1
port 1584 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1_pad
port 1585 nsew
rlabel metal4 s 37293 912000 38223 912254 6 vccd2
port 1586 nsew signal bidirectional
rlabel metal4 s 37293 926746 38223 927000 6 vccd2
port 1586 nsew signal bidirectional
rlabel metal5 s 37313 912000 38203 912254 6 vccd2
port 1586 nsew signal bidirectional
rlabel metal5 s 37313 926746 38203 927000 6 vccd2
port 1586 nsew signal bidirectional
rlabel metal3 s 38220 912100 39600 916900 6 vccd2
port 1586 nsew signal bidirectional
rlabel metal3 s 38220 922151 39600 926940 6 vccd2
port 1586 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2_pad
port 1587 nsew
rlabel metal5 s 6167 70054 19620 80934 6 vccd_pad
port 1588 nsew
rlabel metal4 s 637607 36323 637799 37013 6 vdda
port 1589 nsew signal bidirectional
rlabel metal4 s 622800 36323 622992 37013 6 vdda
port 1589 nsew signal bidirectional
rlabel metal5 s 637607 36343 637799 36993 6 vdda
port 1589 nsew signal bidirectional
rlabel metal5 s 622800 36343 622992 36993 6 vdda
port 1589 nsew signal bidirectional
rlabel metal3 s 632921 37008 637701 40000 6 vdda
port 1589 nsew signal bidirectional
rlabel metal3 s 622942 37008 627722 40000 6 vdda
port 1589 nsew signal bidirectional
rlabel metal4 s 680587 833207 681277 833399 6 vdda1
port 1590 nsew signal bidirectional
rlabel metal4 s 680587 818400 681277 818592 6 vdda1
port 1590 nsew signal bidirectional
rlabel metal5 s 680607 833207 681257 833399 6 vdda1
port 1590 nsew signal bidirectional
rlabel metal5 s 680607 818400 681257 818592 6 vdda1
port 1590 nsew signal bidirectional
rlabel metal3 s 677600 828521 680592 833301 6 vdda1
port 1590 nsew signal bidirectional
rlabel metal3 s 677600 818542 680592 823322 6 vdda1
port 1590 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1_pad
port 1591 nsew
rlabel metal4 s 36323 483000 37013 483192 6 vdda2
port 1592 nsew signal bidirectional
rlabel metal4 s 36323 497807 37013 497999 6 vdda2
port 1592 nsew signal bidirectional
rlabel metal5 s 36343 483000 36993 483192 6 vdda2
port 1592 nsew signal bidirectional
rlabel metal5 s 36343 497807 36993 497999 6 vdda2
port 1592 nsew signal bidirectional
rlabel metal3 s 37008 483099 40000 487879 6 vdda2
port 1592 nsew signal bidirectional
rlabel metal3 s 37008 493078 40000 497858 6 vdda2
port 1592 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2_pad
port 1593 nsew
rlabel metal5 s 624222 6811 636390 18976 6 vdda_pad
port 1594 nsew
rlabel metal4 s 21000 110200 25992 110454 6 vddio
port 1595 nsew signal bidirectional
rlabel metal4 s 35113 110200 36043 110454 6 vddio
port 1595 nsew signal bidirectional
rlabel metal4 s 21000 124946 25992 125200 6 vddio
port 1595 nsew signal bidirectional
rlabel metal4 s 35113 124946 36043 125200 6 vddio
port 1595 nsew signal bidirectional
rlabel metal5 s 35133 110200 36023 110454 6 vddio
port 1595 nsew signal bidirectional
rlabel metal5 s 21003 110200 25993 110454 6 vddio
port 1595 nsew signal bidirectional
rlabel metal5 s 35133 124946 36023 125200 6 vddio
port 1595 nsew signal bidirectional
rlabel metal5 s 21003 124946 25993 125200 6 vddio
port 1595 nsew signal bidirectional
rlabel metal3 s 36040 110299 40000 115079 6 vddio
port 1595 nsew signal bidirectional
rlabel metal3 s 36040 120278 40000 125058 6 vddio
port 1595 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio_pad
port 1596 nsew
rlabel metal4 s 93546 31963 93800 32653 6 vssa
port 1597 nsew signal bidirectional
rlabel metal4 s 93546 28653 93800 28719 6 vssa
port 1597 nsew signal bidirectional
rlabel metal4 s 93546 29435 93800 29671 6 vssa
port 1597 nsew signal bidirectional
rlabel metal4 s 93546 30387 93800 30453 6 vssa
port 1597 nsew signal bidirectional
rlabel metal4 s 78800 31963 79054 32653 6 vssa
port 1597 nsew signal bidirectional
rlabel metal4 s 78800 30387 79054 30453 6 vssa
port 1597 nsew signal bidirectional
rlabel metal4 s 78800 28653 79054 28719 6 vssa
port 1597 nsew signal bidirectional
rlabel metal4 s 78800 29435 79054 29671 6 vssa
port 1597 nsew signal bidirectional
rlabel metal5 s 93546 31983 93800 32631 6 vssa
port 1597 nsew signal bidirectional
rlabel metal5 s 93546 28653 93800 30453 6 vssa
port 1597 nsew signal bidirectional
rlabel metal5 s 78800 31983 79054 32631 6 vssa
port 1597 nsew signal bidirectional
rlabel metal5 s 78800 28653 79054 30453 6 vssa
port 1597 nsew signal bidirectional
rlabel metal3 s 78942 32648 83722 40000 6 vssa
port 1597 nsew signal bidirectional
rlabel metal3 s 88921 32698 93701 40000 6 vssa
port 1597 nsew signal bidirectional
rlabel metal4 s 575600 1004947 575854 1005637 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal4 s 575600 1008881 575854 1008947 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal4 s 575600 1007929 575854 1008165 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal4 s 575600 1007147 575854 1007213 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal4 s 590346 1004947 590600 1005637 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal4 s 590346 1007147 590600 1007213 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal4 s 590346 1008881 590600 1008947 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal4 s 590346 1007929 590600 1008165 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal5 s 575600 1004968 575854 1005616 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal5 s 575600 1007147 575854 1008947 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal5 s 590346 1004968 590600 1005616 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal5 s 590346 1007147 590600 1008947 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal3 s 585678 997600 590458 1004952 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal3 s 575699 997600 580479 1004112 6 vssa1
port 1598 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1_pad
port 1599 nsew
rlabel metal4 s 31963 827600 32653 827854 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal4 s 28653 827600 28719 827854 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal4 s 29435 827600 29671 827854 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal4 s 30387 827600 30453 827854 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal4 s 31963 842346 32653 842600 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal4 s 30387 842346 30453 842600 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal4 s 28653 842346 28719 842600 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal4 s 29435 842346 29671 842600 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal5 s 31983 827600 32631 827854 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal5 s 28653 827600 30453 827854 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal5 s 31983 842346 32631 842600 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal5 s 28653 842346 30453 842600 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal3 s 32648 837678 40000 842458 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal3 s 32698 827699 40000 832479 6 vssa2
port 1600 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2_pad
port 1601 nsew
rlabel metal5 s 80222 6811 92390 18976 6 vssa_pad
port 1602 nsew
rlabel metal4 s 255946 30753 256200 31683 6 vssd
port 1603 nsew signal bidirectional
rlabel metal4 s 241200 30753 241454 31683 6 vssd
port 1603 nsew signal bidirectional
rlabel metal5 s 255946 30773 256200 31663 6 vssd
port 1603 nsew signal bidirectional
rlabel metal5 s 241200 30773 241454 31663 6 vssd
port 1603 nsew signal bidirectional
rlabel metal3 s 251300 31680 256100 39600 6 vssd
port 1603 nsew signal bidirectional
rlabel metal3 s 241260 31680 246049 39600 6 vssd
port 1603 nsew signal bidirectional
rlabel metal4 s 685917 474546 686847 474800 6 vssd1
port 1604 nsew signal bidirectional
rlabel metal4 s 685917 459800 686847 460054 6 vssd1
port 1604 nsew signal bidirectional
rlabel metal5 s 685937 474546 686827 474800 6 vssd1
port 1604 nsew signal bidirectional
rlabel metal5 s 685937 459800 686827 460054 6 vssd1
port 1604 nsew signal bidirectional
rlabel metal3 s 678000 469900 685920 474700 6 vssd1
port 1604 nsew signal bidirectional
rlabel metal3 s 678000 459860 685920 464649 6 vssd1
port 1604 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1_pad
port 1605 nsew
rlabel metal4 s 30753 440800 31683 441054 6 vssd2
port 1606 nsew signal bidirectional
rlabel metal4 s 30753 455546 31683 455800 6 vssd2
port 1606 nsew signal bidirectional
rlabel metal5 s 30773 440800 31663 441054 6 vssd2
port 1606 nsew signal bidirectional
rlabel metal5 s 30773 455546 31663 455800 6 vssd2
port 1606 nsew signal bidirectional
rlabel metal3 s 31680 440900 39600 445700 6 vssd2
port 1606 nsew signal bidirectional
rlabel metal3 s 31680 450951 39600 455740 6 vssd2
port 1606 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2_pad
port 1607 nsew
rlabel metal5 s 243266 6167 254146 19620 6 vssd_pad
port 1608 nsew
rlabel metal4 s 333400 1002767 333654 1003697 6 vssio
port 1609 nsew signal bidirectional
rlabel metal4 s 333400 1032757 333654 1037599 6 vssio
port 1609 nsew signal bidirectional
rlabel metal4 s 348146 1032757 348400 1037599 6 vssio
port 1609 nsew signal bidirectional
rlabel metal4 s 348146 1002767 348400 1003697 6 vssio
port 1609 nsew signal bidirectional
rlabel metal5 s 333400 1002787 333654 1003677 6 vssio
port 1609 nsew signal bidirectional
rlabel metal5 s 348146 1002787 348400 1003677 6 vssio
port 1609 nsew signal bidirectional
rlabel metal3 s 343478 997600 348258 1002770 6 vssio
port 1609 nsew signal bidirectional
rlabel metal3 s 333499 997600 338279 1002770 6 vssio
port 1609 nsew signal bidirectional
rlabel metal4 s 348250 1032757 348400 1037599 6 vssio
port 1609 nsew signal bidirectional
rlabel metal4 s 333526 1035920 333528 1035922 6 vssio
port 1609 nsew signal bidirectional
rlabel metal3 s 579121 34830 583901 40000 6 vssio
port 1609 nsew signal bidirectional
rlabel metal3 s 569142 34830 573922 40000 6 vssio
port 1609 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio_pad
port 1610 nsew
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_pad2
port 1611 nsew
rlabel metal5 s 6811 871210 18976 883378 6 vddio_pad2
port 1612 nsew
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_pad2
port 1613 nsew
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_pad2
port 1614 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 717600 1037600
string GDS_FILE ../gds/chip_io.gds
string GDS_END 36571438
string GDS_START 36076930
string LEFview TRUE
<< end >>
