.subckt sky130_fd_io__condiode A C 
.ends
