magic
tech sky130A
magscale 1 2
timestamp 1623348513
<< obsli1 >>
rect 26 669 770 770
rect 26 127 127 669
rect 189 535 607 607
rect 189 261 261 535
rect 319 319 477 477
rect 535 261 607 535
rect 189 189 607 261
rect 669 127 770 669
rect 26 26 770 127
<< obsm1 >>
rect 315 315 481 481
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 26 26 770 795
string LEFview TRUE
<< end >>
