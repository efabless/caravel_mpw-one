magic
tech sky130A
magscale 12 1
timestamp 1598785768
<< metal5 >>
rect 0 45 15 105
rect 30 45 45 105
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
