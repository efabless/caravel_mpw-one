* NGSPICE file created from storage.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sram_1rw1r_32_256_8_sky130 abstract view
.subckt sram_1rw1r_32_256_8_sky130 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5]
+ din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24]
+ din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0] addr0[1]
+ addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr1[0] addr1[1] addr1[2]
+ addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] csb0 csb1 web0 clk0 clk1 wmask0[0]
+ wmask0[1] wmask0[2] wmask0[3] dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5]
+ dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14]
+ dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22]
+ dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30]
+ dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4] dout1[5] dout1[6] dout1[7]
+ dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16]
+ dout1[17] dout1[18] dout1[19] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24]
+ dout1[25] dout1[26] dout1[27] dout1[28] dout1[29] dout1[30] dout1[31] vdd gnd
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

.subckt storage mgmt_addr[0] mgmt_addr[1] mgmt_addr[2] mgmt_addr[3] mgmt_addr[4] mgmt_addr[5]
+ mgmt_addr[6] mgmt_addr[7] mgmt_addr_ro[0] mgmt_addr_ro[1] mgmt_addr_ro[2] mgmt_addr_ro[3]
+ mgmt_addr_ro[4] mgmt_addr_ro[5] mgmt_addr_ro[6] mgmt_addr_ro[7] mgmt_clk mgmt_ena[0]
+ mgmt_ena[1] mgmt_ena_ro mgmt_rdata[0] mgmt_rdata[10] mgmt_rdata[11] mgmt_rdata[12]
+ mgmt_rdata[13] mgmt_rdata[14] mgmt_rdata[15] mgmt_rdata[16] mgmt_rdata[17] mgmt_rdata[18]
+ mgmt_rdata[19] mgmt_rdata[1] mgmt_rdata[20] mgmt_rdata[21] mgmt_rdata[22] mgmt_rdata[23]
+ mgmt_rdata[24] mgmt_rdata[25] mgmt_rdata[26] mgmt_rdata[27] mgmt_rdata[28] mgmt_rdata[29]
+ mgmt_rdata[2] mgmt_rdata[30] mgmt_rdata[31] mgmt_rdata[32] mgmt_rdata[33] mgmt_rdata[34]
+ mgmt_rdata[35] mgmt_rdata[36] mgmt_rdata[37] mgmt_rdata[38] mgmt_rdata[39] mgmt_rdata[3]
+ mgmt_rdata[40] mgmt_rdata[41] mgmt_rdata[42] mgmt_rdata[43] mgmt_rdata[44] mgmt_rdata[45]
+ mgmt_rdata[46] mgmt_rdata[47] mgmt_rdata[48] mgmt_rdata[49] mgmt_rdata[4] mgmt_rdata[50]
+ mgmt_rdata[51] mgmt_rdata[52] mgmt_rdata[53] mgmt_rdata[54] mgmt_rdata[55] mgmt_rdata[56]
+ mgmt_rdata[57] mgmt_rdata[58] mgmt_rdata[59] mgmt_rdata[5] mgmt_rdata[60] mgmt_rdata[61]
+ mgmt_rdata[62] mgmt_rdata[63] mgmt_rdata[6] mgmt_rdata[7] mgmt_rdata[8] mgmt_rdata[9]
+ mgmt_rdata_ro[0] mgmt_rdata_ro[10] mgmt_rdata_ro[11] mgmt_rdata_ro[12] mgmt_rdata_ro[13]
+ mgmt_rdata_ro[14] mgmt_rdata_ro[15] mgmt_rdata_ro[16] mgmt_rdata_ro[17] mgmt_rdata_ro[18]
+ mgmt_rdata_ro[19] mgmt_rdata_ro[1] mgmt_rdata_ro[20] mgmt_rdata_ro[21] mgmt_rdata_ro[22]
+ mgmt_rdata_ro[23] mgmt_rdata_ro[24] mgmt_rdata_ro[25] mgmt_rdata_ro[26] mgmt_rdata_ro[27]
+ mgmt_rdata_ro[28] mgmt_rdata_ro[29] mgmt_rdata_ro[2] mgmt_rdata_ro[30] mgmt_rdata_ro[31]
+ mgmt_rdata_ro[3] mgmt_rdata_ro[4] mgmt_rdata_ro[5] mgmt_rdata_ro[6] mgmt_rdata_ro[7]
+ mgmt_rdata_ro[8] mgmt_rdata_ro[9] mgmt_wdata[0] mgmt_wdata[10] mgmt_wdata[11] mgmt_wdata[12]
+ mgmt_wdata[13] mgmt_wdata[14] mgmt_wdata[15] mgmt_wdata[16] mgmt_wdata[17] mgmt_wdata[18]
+ mgmt_wdata[19] mgmt_wdata[1] mgmt_wdata[20] mgmt_wdata[21] mgmt_wdata[22] mgmt_wdata[23]
+ mgmt_wdata[24] mgmt_wdata[25] mgmt_wdata[26] mgmt_wdata[27] mgmt_wdata[28] mgmt_wdata[29]
+ mgmt_wdata[2] mgmt_wdata[30] mgmt_wdata[31] mgmt_wdata[3] mgmt_wdata[4] mgmt_wdata[5]
+ mgmt_wdata[6] mgmt_wdata[7] mgmt_wdata[8] mgmt_wdata[9] mgmt_wen[0] mgmt_wen[1]
+ mgmt_wen_mask[0] mgmt_wen_mask[1] mgmt_wen_mask[2] mgmt_wen_mask[3] mgmt_wen_mask[4]
+ mgmt_wen_mask[5] mgmt_wen_mask[6] mgmt_wen_mask[7] VPWR VGND
XFILLER_283_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_329_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[23] mgmt_wdata[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_340_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_280_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_250_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_326_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_308_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_302_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_250_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_252_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_302_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_277_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_293_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_296_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_343_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_287_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_288_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_SRAM_1_din0[22] mgmt_wdata[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_280_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_296_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_310_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_283_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_299_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_1_din0[21] mgmt_wdata[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_265_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_280_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_314_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_286_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_299_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_274_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[20] mgmt_wdata[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_280_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_332_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_314_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_250_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[7] mgmt_addr_ro[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSRAM_0 mgmt_wdata[0] mgmt_wdata[1] mgmt_wdata[2] mgmt_wdata[3] mgmt_wdata[4] mgmt_wdata[5]
+ mgmt_wdata[6] mgmt_wdata[7] mgmt_wdata[8] mgmt_wdata[9] mgmt_wdata[10] mgmt_wdata[11]
+ mgmt_wdata[12] mgmt_wdata[13] mgmt_wdata[14] mgmt_wdata[15] mgmt_wdata[16] mgmt_wdata[17]
+ mgmt_wdata[18] mgmt_wdata[19] mgmt_wdata[20] mgmt_wdata[21] mgmt_wdata[22] mgmt_wdata[23]
+ mgmt_wdata[24] mgmt_wdata[25] mgmt_wdata[26] mgmt_wdata[27] mgmt_wdata[28] mgmt_wdata[29]
+ mgmt_wdata[30] mgmt_wdata[31] mgmt_addr[0] mgmt_addr[1] mgmt_addr[2] mgmt_addr[3]
+ mgmt_addr[4] mgmt_addr[5] mgmt_addr[6] mgmt_addr[7] mgmt_addr_ro[0] mgmt_addr_ro[1]
+ mgmt_addr_ro[2] mgmt_addr_ro[3] mgmt_addr_ro[4] mgmt_addr_ro[5] mgmt_addr_ro[6]
+ mgmt_addr_ro[7] mgmt_ena[0] mgmt_ena_ro mgmt_wen[0] mgmt_clk mgmt_clk mgmt_wen_mask[0]
+ mgmt_wen_mask[1] mgmt_wen_mask[2] mgmt_wen_mask[3] mgmt_rdata[0] mgmt_rdata[1] mgmt_rdata[2]
+ mgmt_rdata[3] mgmt_rdata[4] mgmt_rdata[5] mgmt_rdata[6] mgmt_rdata[7] mgmt_rdata[8]
+ mgmt_rdata[9] mgmt_rdata[10] mgmt_rdata[11] mgmt_rdata[12] mgmt_rdata[13] mgmt_rdata[14]
+ mgmt_rdata[15] mgmt_rdata[16] mgmt_rdata[17] mgmt_rdata[18] mgmt_rdata[19] mgmt_rdata[20]
+ mgmt_rdata[21] mgmt_rdata[22] mgmt_rdata[23] mgmt_rdata[24] mgmt_rdata[25] mgmt_rdata[26]
+ mgmt_rdata[27] mgmt_rdata[28] mgmt_rdata[29] mgmt_rdata[30] mgmt_rdata[31] mgmt_rdata_ro[0]
+ mgmt_rdata_ro[1] mgmt_rdata_ro[2] mgmt_rdata_ro[3] mgmt_rdata_ro[4] mgmt_rdata_ro[5]
+ mgmt_rdata_ro[6] mgmt_rdata_ro[7] mgmt_rdata_ro[8] mgmt_rdata_ro[9] mgmt_rdata_ro[10]
+ mgmt_rdata_ro[11] mgmt_rdata_ro[12] mgmt_rdata_ro[13] mgmt_rdata_ro[14] mgmt_rdata_ro[15]
+ mgmt_rdata_ro[16] mgmt_rdata_ro[17] mgmt_rdata_ro[18] mgmt_rdata_ro[19] mgmt_rdata_ro[20]
+ mgmt_rdata_ro[21] mgmt_rdata_ro[22] mgmt_rdata_ro[23] mgmt_rdata_ro[24] mgmt_rdata_ro[25]
+ mgmt_rdata_ro[26] mgmt_rdata_ro[27] mgmt_rdata_ro[28] mgmt_rdata_ro[29] mgmt_rdata_ro[30]
+ mgmt_rdata_ro[31] VPWR VGND sram_1rw1r_32_256_8_sky130
XFILLER_7_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_299_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_338_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_clk0 mgmt_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_256_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_286_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_322_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_305_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_addr1[6] mgmt_addr_ro[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSRAM_1 mgmt_wdata[0] mgmt_wdata[1] mgmt_wdata[2] mgmt_wdata[3] mgmt_wdata[4] mgmt_wdata[5]
+ mgmt_wdata[6] mgmt_wdata[7] mgmt_wdata[8] mgmt_wdata[9] mgmt_wdata[10] mgmt_wdata[11]
+ mgmt_wdata[12] mgmt_wdata[13] mgmt_wdata[14] mgmt_wdata[15] mgmt_wdata[16] mgmt_wdata[17]
+ mgmt_wdata[18] mgmt_wdata[19] mgmt_wdata[20] mgmt_wdata[21] mgmt_wdata[22] mgmt_wdata[23]
+ mgmt_wdata[24] mgmt_wdata[25] mgmt_wdata[26] mgmt_wdata[27] mgmt_wdata[28] mgmt_wdata[29]
+ mgmt_wdata[30] mgmt_wdata[31] mgmt_addr[0] mgmt_addr[1] mgmt_addr[2] mgmt_addr[3]
+ mgmt_addr[4] mgmt_addr[5] mgmt_addr[6] mgmt_addr[7] SRAM_1/addr1[0] SRAM_1/addr1[1]
+ SRAM_1/addr1[2] SRAM_1/addr1[3] SRAM_1/addr1[4] SRAM_1/addr1[5] SRAM_1/addr1[6]
+ SRAM_1/addr1[7] mgmt_ena[1] SRAM_1/csb1 mgmt_wen[1] mgmt_clk SRAM_1/clk1 mgmt_wen_mask[4]
+ mgmt_wen_mask[5] mgmt_wen_mask[6] mgmt_wen_mask[7] mgmt_rdata[32] mgmt_rdata[33]
+ mgmt_rdata[34] mgmt_rdata[35] mgmt_rdata[36] mgmt_rdata[37] mgmt_rdata[38] mgmt_rdata[39]
+ mgmt_rdata[40] mgmt_rdata[41] mgmt_rdata[42] mgmt_rdata[43] mgmt_rdata[44] mgmt_rdata[45]
+ mgmt_rdata[46] mgmt_rdata[47] mgmt_rdata[48] mgmt_rdata[49] mgmt_rdata[50] mgmt_rdata[51]
+ mgmt_rdata[52] mgmt_rdata[53] mgmt_rdata[54] mgmt_rdata[55] mgmt_rdata[56] mgmt_rdata[57]
+ mgmt_rdata[58] mgmt_rdata[59] mgmt_rdata[60] mgmt_rdata[61] mgmt_rdata[62] mgmt_rdata[63]
+ SRAM_1/dout1[0] SRAM_1/dout1[1] SRAM_1/dout1[2] SRAM_1/dout1[3] SRAM_1/dout1[4]
+ SRAM_1/dout1[5] SRAM_1/dout1[6] SRAM_1/dout1[7] SRAM_1/dout1[8] SRAM_1/dout1[9]
+ SRAM_1/dout1[10] SRAM_1/dout1[11] SRAM_1/dout1[12] SRAM_1/dout1[13] SRAM_1/dout1[14]
+ SRAM_1/dout1[15] SRAM_1/dout1[16] SRAM_1/dout1[17] SRAM_1/dout1[18] SRAM_1/dout1[19]
+ SRAM_1/dout1[20] SRAM_1/dout1[21] SRAM_1/dout1[22] SRAM_1/dout1[23] SRAM_1/dout1[24]
+ SRAM_1/dout1[25] SRAM_1/dout1[26] SRAM_1/dout1[27] SRAM_1/dout1[28] SRAM_1/dout1[29]
+ SRAM_1/dout1[30] SRAM_1/dout1[31] VPWR VGND sram_1rw1r_32_256_8_sky130
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_299_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_302_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_295_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[29] mgmt_wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_294_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_313_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_clk1 mgmt_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_256_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_310_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_308_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_307_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[5] mgmt_addr_ro[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_310_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_289_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[28] mgmt_wdata[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_308_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_324_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_280_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_271_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_326_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_319_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_261_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[4] mgmt_addr_ro[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_313_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_316_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_332_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_327_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[27] mgmt_wdata[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_324_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_324_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_296_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_340_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_271_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_wmask0[3] mgmt_wen_mask[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_316_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_SRAM_0_addr1[3] mgmt_addr_ro[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_310_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_332_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_327_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_253_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[26] mgmt_wdata[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_340_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_289_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_250_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_SRAM_1_wmask0[2] mgmt_wen_mask[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_261_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_252_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_307_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_322_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[2] mgmt_addr_ro[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_321_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_256_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_343_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_286_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_253_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_1_csb0 mgmt_ena[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_SRAM_0_din0[25] mgmt_wdata[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_292_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_291_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_264_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_274_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_329_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_273_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_340_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_wmask0[1] mgmt_wen_mask[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_261_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr1[1] mgmt_addr_ro[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_256_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_298_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_253_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_din0[24] mgmt_wdata[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_292_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_283_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_264_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_264_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_280_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_256_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_294_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_261_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_1_wmask0[0] mgmt_wen_mask[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_316_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_261_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_0_addr1[0] mgmt_addr_ro[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_272_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_272_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_257_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[23] mgmt_wdata[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_282_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_280_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_280_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_337_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_343_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_330_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_259_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_334_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_316_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_267_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_283_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_286_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_278_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[22] mgmt_wdata[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_294_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_291_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_259_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_343_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_249_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_275_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_252_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_286_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_283_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_286_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[21] mgmt_wdata[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_294_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_294_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_259_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_273_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_291_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_255_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_304_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[9] mgmt_wdata[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[19] mgmt_wdata[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_255_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[20] mgmt_wdata[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_276_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_282_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_270_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_335_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_304_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_297_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_1_din0[8] mgmt_wdata[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[18] mgmt_wdata[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_279_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_268_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_282_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_300_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_312_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[7] mgmt_wdata[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[17] mgmt_wdata[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_310_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_285_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_284_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_260_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_wmask0[3] mgmt_wen_mask[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_334_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_300_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_316_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_307_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_1_addr0[7] mgmt_addr[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_1_din0[6] mgmt_wdata[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[16] mgmt_wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_300_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_303_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_253_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_wmask0[2] mgmt_wen_mask[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_334_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_261_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_316_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_252_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_307_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_addr0[6] mgmt_addr[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_311_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[5] mgmt_wdata[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_306_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_322_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_1_din0[15] mgmt_wdata[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_300_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_317_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_303_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_276_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_wmask0[1] mgmt_wen_mask[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_258_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_314_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_342_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_270_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_261_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_309_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_330_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_addr0[5] mgmt_addr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_306_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[31] mgmt_wdata[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[4] mgmt_wdata[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_276_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_300_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_297_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_1_din0[14] mgmt_wdata[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_317_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_wmask0[0] mgmt_wen_mask[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_258_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_330_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_325_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_315_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_330_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_1_addr0[4] mgmt_addr[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_336_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_312_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[30] mgmt_wdata[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_1_din0[3] mgmt_wdata[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[13] mgmt_wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_288_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_317_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_291_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_csb0 mgmt_ena[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_301_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_337_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_258_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_254_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_339_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_319_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_263_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_addr0[3] mgmt_addr[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_336_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_262_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[2] mgmt_wdata[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_331_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[12] mgmt_wdata[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_281_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_SRAM_0_csb1 mgmt_ena_ro VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_282_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_254_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_264_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_304_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_255_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_249_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_251_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_1_addr0[2] mgmt_addr[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_306_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_262_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_1_din0[1] mgmt_wdata[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[11] mgmt_wdata[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_312_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_270_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_320_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_263_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_281_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_324_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_260_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_1_addr0[1] mgmt_addr[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_306_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[0] mgmt_wdata[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_300_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[10] mgmt_wdata[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_0_din0[9] mgmt_wdata[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_267_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_293_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_268_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_276_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_258_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_249_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_263_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_265_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_276_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_1_addr0[0] mgmt_addr[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_297_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_SRAM_1_web0 mgmt_wen[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_294_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_din0[8] mgmt_wdata[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_284_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_276_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_334_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_258_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_281_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_263_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_318_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_330_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_292_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_292_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[19] mgmt_wdata[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_311_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_SRAM_0_din0[7] mgmt_wdata[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_339_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_336_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_257_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_318_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_260_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_321_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_312_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_SRAM_0_din0[18] mgmt_wdata[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_303_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_297_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_288_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_298_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_279_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[6] mgmt_wdata[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_287_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_293_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_258_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_272_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[17] mgmt_wdata[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_266_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_320_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_311_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[5] mgmt_wdata[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_293_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_290_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_258_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_342_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_addr0[7] mgmt_addr[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_315_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_323_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_306_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[16] mgmt_wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_305_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_288_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[4] mgmt_wdata[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_342_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr0[6] mgmt_addr[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_324_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_315_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_306_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[15] mgmt_wdata[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_301_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_312_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_din0[3] mgmt_wdata[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_288_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_307_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_clk0 mgmt_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_266_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_320_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_304_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_263_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_SRAM_0_addr0[5] mgmt_addr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[31] mgmt_wdata[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_332_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_260_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_314_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[14] mgmt_wdata[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_320_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_302_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_312_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_343_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_0_din0[2] mgmt_wdata[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_287_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_307_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_318_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[29] mgmt_wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_335_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_320_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_256_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr0[4] mgmt_addr[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_318_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_din0[30] mgmt_wdata[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_din0[13] mgmt_wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_305_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_320_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_326_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_299_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[1] mgmt_wdata[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_278_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_318_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_318_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_336_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[28] mgmt_wdata[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_327_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_263_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr0[3] mgmt_addr[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_254_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_309_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_315_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_331_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[12] mgmt_wdata[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_305_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_320_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_326_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_299_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_302_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_din0[0] mgmt_wdata[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_278_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_279_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_290_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_334_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_1_din0[27] mgmt_wdata[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_272_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_263_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_SRAM_0_addr0[2] mgmt_addr[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_308_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_261_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_314_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_SRAM_0_din0[11] mgmt_wdata[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_342_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_252_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_252_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_263_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_341_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[26] mgmt_wdata[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_280_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_260_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_260_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_SRAM_0_addr0[1] mgmt_addr[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_262_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_254_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_314_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_250_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_SRAM_0_din0[10] mgmt_wdata[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_266_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_293_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_334_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_339_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_258_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_266_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_308_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_265_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[25] mgmt_wdata[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_269_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_0_addr0[0] mgmt_addr[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_314_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_250_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_266_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_SRAM_0_web0 mgmt_wen[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_263_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_284_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_274_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_266_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_SRAM_1_din0[24] mgmt_wdata[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_324_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_257_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_271_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_326_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_271_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_314_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_250_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_282_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_302_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_332_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_290_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

