magic
tech sky130A
magscale 1 2
timestamp 1607712712
<< obsli1 >>
rect 0 0 4992 4087
<< obsm1 >>
rect 0 0 4992 4935
<< metal2 >>
rect 4244 4200 4300 5000
rect 596 0 652 800
<< obsm2 >>
rect 598 4144 4188 4935
rect 4356 4144 4396 4935
rect 598 856 4396 4144
rect 708 0 4396 856
<< obsm3 >>
rect 673 0 4401 4917
<< metal4 >>
rect 673 -51 993 4935
rect 1507 -51 1827 4935
rect 2340 -51 2660 4935
rect 3173 -51 3493 4935
rect 4007 -51 4327 4935
<< obsm4 >>
rect 1907 0 2260 4935
rect 2740 0 3093 4935
rect 3573 0 3927 4935
<< metal5 >>
rect 0 3956 4992 4276
rect 0 3122 4992 3442
rect 0 2289 4992 2609
rect 0 1456 4992 1776
rect 0 622 4992 942
<< labels >>
rlabel metal2 s 4244 4200 4300 5000 6 A
port 1 nsew signal input
rlabel metal2 s 596 0 652 800 6 X
port 2 nsew signal output
rlabel metal4 s 4007 -51 4327 4935 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 2340 -51 2660 4935 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 673 -51 993 4935 6 VPWR
port 5 nsew power bidirectional
rlabel metal5 s 0 3956 4992 4276 6 VPWR
port 6 nsew power bidirectional
rlabel metal5 s 0 2289 4992 2609 6 VPWR
port 7 nsew power bidirectional
rlabel metal5 s 0 622 4992 942 6 VPWR
port 8 nsew power bidirectional
rlabel metal4 s 3173 -51 3493 4935 6 VGND
port 9 nsew ground bidirectional
rlabel metal4 s 1507 -51 1827 4935 6 VGND
port 10 nsew ground bidirectional
rlabel metal5 s 0 3122 4992 3442 6 VGND
port 11 nsew ground bidirectional
rlabel metal5 s 0 1456 4992 1776 6 VGND
port 12 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 5000 5000
string LEFview TRUE
<< end >>
