magic
tech sky130A
magscale 1 2
timestamp 1607630556
<< metal1 >>
rect 84010 995596 84016 995648
rect 84068 995636 84074 995648
rect 91738 995636 91744 995648
rect 84068 995608 91744 995636
rect 84068 995596 84074 995608
rect 91738 995596 91744 995608
rect 91796 995596 91802 995648
rect 531958 995596 531964 995648
rect 532016 995636 532022 995648
rect 539686 995636 539692 995648
rect 532016 995608 539692 995636
rect 532016 995596 532022 995608
rect 539686 995596 539692 995608
rect 539744 995596 539750 995648
rect 135346 995460 135352 995512
rect 135404 995500 135410 995512
rect 143166 995500 143172 995512
rect 135404 995472 143172 995500
rect 135404 995460 135410 995472
rect 143166 995460 143172 995472
rect 143224 995460 143230 995512
rect 633802 995460 633808 995512
rect 633860 995500 633866 995512
rect 641530 995500 641536 995512
rect 633860 995472 641536 995500
rect 633860 995460 633866 995472
rect 641530 995460 641536 995472
rect 641588 995460 641594 995512
rect 238202 995392 238208 995444
rect 238260 995432 238266 995444
rect 245930 995432 245936 995444
rect 238260 995404 245936 995432
rect 238260 995392 238266 995404
rect 245930 995392 245936 995404
rect 245988 995392 245994 995444
rect 289630 995256 289636 995308
rect 289688 995296 289694 995308
rect 297634 995296 297640 995308
rect 289688 995268 297640 995296
rect 289688 995256 289694 995268
rect 297634 995256 297640 995268
rect 297692 995256 297698 995308
rect 391474 995256 391480 995308
rect 391532 995296 391538 995308
rect 399478 995296 399484 995308
rect 391532 995268 399484 995296
rect 391532 995256 391538 995268
rect 399478 995256 399484 995268
rect 399536 995256 399542 995308
rect 480438 995256 480444 995308
rect 480496 995296 480502 995308
rect 488442 995296 488448 995308
rect 480496 995268 488448 995296
rect 480496 995256 480502 995268
rect 488442 995256 488448 995268
rect 488500 995256 488506 995308
rect 589550 992264 589556 992316
rect 589608 992304 589614 992316
rect 674742 992304 674748 992316
rect 589608 992276 674748 992304
rect 589608 992264 589614 992276
rect 674742 992264 674748 992276
rect 674800 992264 674806 992316
rect 44082 992196 44088 992248
rect 44140 992236 44146 992248
rect 329558 992236 329564 992248
rect 44140 992208 329564 992236
rect 44140 992196 44146 992208
rect 329558 992196 329564 992208
rect 329616 992196 329622 992248
rect 585042 992196 585048 992248
rect 585100 992236 585106 992248
rect 675202 992236 675208 992248
rect 585100 992208 675208 992236
rect 585100 992196 585106 992208
rect 675202 992196 675208 992208
rect 675260 992196 675266 992248
rect 78858 990768 78864 990820
rect 78916 990808 78922 990820
rect 130286 990808 130292 990820
rect 78916 990780 130292 990808
rect 78916 990768 78922 990780
rect 130286 990768 130292 990780
rect 130344 990808 130350 990820
rect 132402 990808 132408 990820
rect 130344 990780 132408 990808
rect 130344 990768 130350 990780
rect 132402 990768 132408 990780
rect 132460 990768 132466 990820
rect 181714 990768 181720 990820
rect 181772 990808 181778 990820
rect 233050 990808 233056 990820
rect 181772 990780 233056 990808
rect 181772 990768 181778 990780
rect 233050 990768 233056 990780
rect 233108 990768 233114 990820
rect 285306 990808 285312 990820
rect 275940 990780 285312 990808
rect 79502 990700 79508 990752
rect 79560 990740 79566 990752
rect 130930 990740 130936 990752
rect 79560 990712 130936 990740
rect 79560 990700 79566 990712
rect 130930 990700 130936 990712
rect 130988 990740 130994 990752
rect 182358 990740 182364 990752
rect 130988 990712 182364 990740
rect 130988 990700 130994 990712
rect 182358 990700 182364 990712
rect 182416 990740 182422 990752
rect 187694 990740 187700 990752
rect 182416 990712 187700 990740
rect 182416 990700 182422 990712
rect 187694 990700 187700 990712
rect 187752 990700 187758 990752
rect 206922 990700 206928 990752
rect 206980 990740 206986 990752
rect 226334 990740 226340 990752
rect 206980 990712 226340 990740
rect 206980 990700 206986 990712
rect 226334 990700 226340 990712
rect 226392 990700 226398 990752
rect 256602 990740 256608 990752
rect 237392 990712 256608 990740
rect 88334 990632 88340 990684
rect 88392 990672 88398 990684
rect 89990 990672 89996 990684
rect 88392 990644 89996 990672
rect 88392 990632 88398 990644
rect 89990 990632 89996 990644
rect 90048 990672 90054 990684
rect 141418 990672 141424 990684
rect 90048 990644 141424 990672
rect 90048 990632 90054 990644
rect 141418 990632 141424 990644
rect 141476 990672 141482 990684
rect 192846 990672 192852 990684
rect 141476 990644 192852 990672
rect 141476 990632 141482 990644
rect 192846 990632 192852 990644
rect 192904 990672 192910 990684
rect 192904 990644 226380 990672
rect 192904 990632 192910 990644
rect 132402 990564 132408 990616
rect 132460 990604 132466 990616
rect 181714 990604 181720 990616
rect 132460 990576 181720 990604
rect 132460 990564 132466 990576
rect 181714 990564 181720 990576
rect 181772 990564 181778 990616
rect 186682 990564 186688 990616
rect 186740 990604 186746 990616
rect 194686 990604 194692 990616
rect 186740 990576 194692 990604
rect 186740 990564 186746 990576
rect 194686 990564 194692 990576
rect 194744 990564 194750 990616
rect 226352 990604 226380 990644
rect 233602 990604 233608 990616
rect 226352 990576 233608 990604
rect 233602 990564 233608 990576
rect 233660 990564 233666 990616
rect 237392 990604 237420 990712
rect 256602 990700 256608 990712
rect 256660 990700 256666 990752
rect 275940 990740 275968 990780
rect 285306 990768 285312 990780
rect 285364 990768 285370 990820
rect 295702 990768 295708 990820
rect 295760 990808 295766 990820
rect 295760 990780 324176 990808
rect 295760 990768 295766 990780
rect 256712 990712 275968 990740
rect 246942 990632 246948 990684
rect 247000 990672 247006 990684
rect 256712 990672 256740 990712
rect 295518 990700 295524 990752
rect 295576 990740 295582 990752
rect 314654 990740 314660 990752
rect 295576 990712 314660 990740
rect 295576 990700 295582 990712
rect 314654 990700 314660 990712
rect 314712 990700 314718 990752
rect 324148 990740 324176 990780
rect 324222 990768 324228 990820
rect 324280 990808 324286 990820
rect 333882 990808 333888 990820
rect 324280 990780 333888 990808
rect 324280 990768 324286 990780
rect 333882 990768 333888 990780
rect 333940 990768 333946 990820
rect 343634 990768 343640 990820
rect 343692 990808 343698 990820
rect 353294 990808 353300 990820
rect 343692 990780 353300 990808
rect 343692 990768 343698 990780
rect 353294 990768 353300 990780
rect 353352 990768 353358 990820
rect 387150 990808 387156 990820
rect 386524 990780 387156 990808
rect 324314 990740 324320 990752
rect 324148 990712 324320 990740
rect 324314 990700 324320 990712
rect 324372 990700 324378 990752
rect 333974 990700 333980 990752
rect 334032 990740 334038 990752
rect 357802 990740 357808 990752
rect 334032 990712 357808 990740
rect 334032 990700 334038 990712
rect 357802 990700 357808 990712
rect 357860 990700 357866 990752
rect 372338 990700 372344 990752
rect 372396 990740 372402 990752
rect 386524 990740 386552 990780
rect 387150 990768 387156 990780
rect 387208 990808 387214 990820
rect 475378 990808 475384 990820
rect 387208 990780 475384 990808
rect 387208 990768 387214 990780
rect 475378 990768 475384 990780
rect 475436 990768 475442 990820
rect 475470 990768 475476 990820
rect 475528 990808 475534 990820
rect 526898 990808 526904 990820
rect 475528 990780 526904 990808
rect 475528 990768 475534 990780
rect 526898 990768 526904 990780
rect 526956 990808 526962 990820
rect 545942 990808 545948 990820
rect 526956 990780 545948 990808
rect 526956 990768 526962 990780
rect 545942 990768 545948 990780
rect 546000 990768 546006 990820
rect 546402 990768 546408 990820
rect 546460 990808 546466 990820
rect 628650 990808 628656 990820
rect 546460 990780 628656 990808
rect 546460 990768 546466 990780
rect 628650 990768 628656 990780
rect 628708 990768 628714 990820
rect 372396 990712 375880 990740
rect 372396 990700 372402 990712
rect 247000 990644 256740 990672
rect 247000 990632 247006 990644
rect 353294 990632 353300 990684
rect 353352 990672 353358 990684
rect 353352 990644 353432 990672
rect 353352 990632 353358 990644
rect 233804 990576 237420 990604
rect 233050 990496 233056 990548
rect 233108 990536 233114 990548
rect 233804 990536 233832 990576
rect 244366 990564 244372 990616
rect 244424 990604 244430 990616
rect 256694 990604 256700 990616
rect 244424 990576 256700 990604
rect 244424 990564 244430 990576
rect 256694 990564 256700 990576
rect 256752 990564 256758 990616
rect 284570 990604 284576 990616
rect 270512 990576 284576 990604
rect 233108 990508 233832 990536
rect 233108 990496 233114 990508
rect 256602 990496 256608 990548
rect 256660 990536 256666 990548
rect 270512 990536 270540 990576
rect 284570 990564 284576 990576
rect 284628 990564 284634 990616
rect 284662 990564 284668 990616
rect 284720 990604 284726 990616
rect 289814 990604 289820 990616
rect 284720 990576 289820 990604
rect 284720 990564 284726 990576
rect 289814 990564 289820 990576
rect 289872 990564 289878 990616
rect 309042 990564 309048 990616
rect 309100 990604 309106 990616
rect 315942 990604 315948 990616
rect 309100 990576 315948 990604
rect 309100 990564 309106 990576
rect 315942 990564 315948 990576
rect 316000 990564 316006 990616
rect 343634 990604 343640 990616
rect 328472 990576 343640 990604
rect 256660 990508 270540 990536
rect 256660 990496 256666 990508
rect 187694 990428 187700 990480
rect 187752 990468 187758 990480
rect 206922 990468 206928 990480
rect 187752 990440 206928 990468
rect 187752 990428 187758 990440
rect 206922 990428 206928 990440
rect 206980 990428 206986 990480
rect 295794 990428 295800 990480
rect 295852 990468 295858 990480
rect 309042 990468 309048 990480
rect 295852 990440 309048 990468
rect 295852 990428 295858 990440
rect 309042 990428 309048 990440
rect 309100 990428 309106 990480
rect 314654 990428 314660 990480
rect 314712 990468 314718 990480
rect 324222 990468 324228 990480
rect 314712 990440 324228 990468
rect 314712 990428 314718 990440
rect 324222 990428 324228 990440
rect 324280 990428 324286 990480
rect 324314 990428 324320 990480
rect 324372 990468 324378 990480
rect 328472 990468 328500 990576
rect 343634 990564 343640 990576
rect 343692 990564 343698 990616
rect 343726 990564 343732 990616
rect 343784 990604 343790 990616
rect 353404 990604 353432 990644
rect 357986 990632 357992 990684
rect 358044 990672 358050 990684
rect 372246 990672 372252 990684
rect 358044 990644 372252 990672
rect 358044 990632 358050 990644
rect 372246 990632 372252 990644
rect 372304 990632 372310 990684
rect 375852 990672 375880 990712
rect 386432 990712 386552 990740
rect 386432 990672 386460 990712
rect 488442 990700 488448 990752
rect 488500 990740 488506 990752
rect 527542 990740 527548 990752
rect 488500 990712 527548 990740
rect 488500 990700 488506 990712
rect 527542 990700 527548 990712
rect 527600 990740 527606 990752
rect 629294 990740 629300 990752
rect 527600 990712 629300 990740
rect 527600 990700 527606 990712
rect 629294 990700 629300 990712
rect 629352 990700 629358 990752
rect 475470 990672 475476 990684
rect 375852 990644 386460 990672
rect 390848 990644 475476 990672
rect 372338 990604 372344 990616
rect 343784 990576 347636 990604
rect 353404 990576 372344 990604
rect 343784 990564 343790 990576
rect 324372 990440 328500 990468
rect 347608 990468 347636 990576
rect 372338 990564 372344 990576
rect 372396 990564 372402 990616
rect 386506 990604 386512 990616
rect 372632 990576 386512 990604
rect 372246 990496 372252 990548
rect 372304 990536 372310 990548
rect 372632 990536 372660 990576
rect 386506 990564 386512 990576
rect 386564 990604 386570 990616
rect 390848 990604 390876 990644
rect 475470 990632 475476 990644
rect 475528 990632 475534 990684
rect 546310 990632 546316 990684
rect 546368 990672 546374 990684
rect 563054 990672 563060 990684
rect 546368 990644 563060 990672
rect 546368 990632 546374 990644
rect 563054 990632 563060 990644
rect 563112 990632 563118 990684
rect 386564 990576 390876 990604
rect 386564 990564 386570 990576
rect 486694 990564 486700 990616
rect 486752 990604 486758 990616
rect 486752 990576 537616 990604
rect 486752 990564 486758 990576
rect 372304 990508 372660 990536
rect 372304 990496 372310 990508
rect 475378 990496 475384 990548
rect 475436 990536 475442 990548
rect 476114 990536 476120 990548
rect 475436 990508 476120 990536
rect 475436 990496 475442 990508
rect 476114 990496 476120 990508
rect 476172 990536 476178 990548
rect 488350 990536 488356 990548
rect 476172 990508 488356 990536
rect 476172 990496 476178 990508
rect 488350 990496 488356 990508
rect 488408 990496 488414 990548
rect 537588 990536 537616 990576
rect 582282 990564 582288 990616
rect 582340 990604 582346 990616
rect 582340 990576 585180 990604
rect 582340 990564 582346 990576
rect 585152 990548 585180 990576
rect 587986 990564 587992 990616
rect 588044 990604 588050 990616
rect 623682 990604 623688 990616
rect 588044 990576 623688 990604
rect 588044 990564 588050 990576
rect 623682 990564 623688 990576
rect 623740 990564 623746 990616
rect 537846 990536 537852 990548
rect 537588 990508 537852 990536
rect 537846 990496 537852 990508
rect 537904 990496 537910 990548
rect 585134 990496 585140 990548
rect 585192 990496 585198 990548
rect 623866 990496 623872 990548
rect 623924 990536 623930 990548
rect 639782 990536 639788 990548
rect 623924 990508 639788 990536
rect 623924 990496 623930 990508
rect 639782 990496 639788 990508
rect 639840 990496 639846 990548
rect 353202 990468 353208 990480
rect 347608 990440 353208 990468
rect 324372 990428 324378 990440
rect 353202 990428 353208 990440
rect 353260 990428 353266 990480
rect 353386 990428 353392 990480
rect 353444 990468 353450 990480
rect 364334 990468 364340 990480
rect 353444 990440 364340 990468
rect 353444 990428 353450 990440
rect 364334 990428 364340 990440
rect 364392 990428 364398 990480
rect 397638 990428 397644 990480
rect 397696 990468 397702 990480
rect 405642 990468 405648 990480
rect 397696 990440 405648 990468
rect 397696 990428 397702 990440
rect 405642 990428 405648 990440
rect 405700 990428 405706 990480
rect 537864 990468 537892 990496
rect 546310 990468 546316 990480
rect 537864 990440 546316 990468
rect 546310 990428 546316 990440
rect 546368 990428 546374 990480
rect 226334 990360 226340 990412
rect 226392 990400 226398 990412
rect 233694 990400 233700 990412
rect 226392 990372 233700 990400
rect 226392 990360 226398 990372
rect 233694 990360 233700 990372
rect 233752 990400 233758 990412
rect 246942 990400 246948 990412
rect 233752 990372 246948 990400
rect 233752 990360 233758 990372
rect 246942 990360 246948 990372
rect 247000 990360 247006 990412
rect 285306 990360 285312 990412
rect 285364 990400 285370 990412
rect 295702 990400 295708 990412
rect 285364 990372 295708 990400
rect 285364 990360 285370 990372
rect 295702 990360 295708 990372
rect 295760 990360 295766 990412
rect 233602 990292 233608 990344
rect 233660 990332 233666 990344
rect 244366 990332 244372 990344
rect 233660 990304 244372 990332
rect 233660 990292 233666 990304
rect 244366 990292 244372 990304
rect 244424 990292 244430 990344
rect 256694 990292 256700 990344
rect 256752 990332 256758 990344
rect 295812 990332 295840 990428
rect 424962 990360 424968 990412
rect 425020 990400 425026 990412
rect 430482 990400 430488 990412
rect 425020 990372 430488 990400
rect 425020 990360 425026 990372
rect 430482 990360 430488 990372
rect 430540 990360 430546 990412
rect 430574 990360 430580 990412
rect 430632 990400 430638 990412
rect 430632 990372 434668 990400
rect 430632 990360 430638 990372
rect 256752 990304 295840 990332
rect 256752 990292 256758 990304
rect 383562 990292 383568 990344
rect 383620 990332 383626 990344
rect 397638 990332 397644 990344
rect 383620 990304 397644 990332
rect 383620 990292 383626 990304
rect 397638 990292 397644 990304
rect 397696 990292 397702 990344
rect 405642 990292 405648 990344
rect 405700 990332 405706 990344
rect 434640 990332 434668 990372
rect 463602 990360 463608 990412
rect 463660 990400 463666 990412
rect 469122 990400 469128 990412
rect 463660 990372 469128 990400
rect 463660 990360 463666 990372
rect 469122 990360 469128 990372
rect 469180 990360 469186 990412
rect 469214 990360 469220 990412
rect 469272 990400 469278 990412
rect 471974 990400 471980 990412
rect 469272 990372 471980 990400
rect 469272 990360 469278 990372
rect 471974 990360 471980 990372
rect 472032 990360 472038 990412
rect 444374 990332 444380 990344
rect 405700 990304 405780 990332
rect 434640 990304 444380 990332
rect 405700 990292 405706 990304
rect 405752 990276 405780 990304
rect 444374 990292 444380 990304
rect 444432 990292 444438 990344
rect 315942 990224 315948 990276
rect 316000 990264 316006 990276
rect 325694 990264 325700 990276
rect 316000 990236 325700 990264
rect 316000 990224 316006 990236
rect 325694 990224 325700 990236
rect 325752 990224 325758 990276
rect 405734 990224 405740 990276
rect 405792 990224 405798 990276
rect 471974 990224 471980 990276
rect 472032 990264 472038 990276
rect 486694 990264 486700 990276
rect 472032 990236 486700 990264
rect 472032 990224 472038 990236
rect 486694 990224 486700 990236
rect 486752 990224 486758 990276
rect 42334 990156 42340 990208
rect 42392 990196 42398 990208
rect 79502 990196 79508 990208
rect 42392 990168 79508 990196
rect 42392 990156 42398 990168
rect 79502 990156 79508 990168
rect 79560 990156 79566 990208
rect 639782 990156 639788 990208
rect 639840 990196 639846 990208
rect 673638 990196 673644 990208
rect 639840 990168 673644 990196
rect 639840 990156 639846 990168
rect 673638 990156 673644 990168
rect 673696 990156 673702 990208
rect 42242 990088 42248 990140
rect 42300 990128 42306 990140
rect 78858 990128 78864 990140
rect 42300 990100 78864 990128
rect 42300 990088 42306 990100
rect 78858 990088 78864 990100
rect 78916 990088 78922 990140
rect 88334 990088 88340 990140
rect 88392 990088 88398 990140
rect 325694 990088 325700 990140
rect 325752 990128 325758 990140
rect 343726 990128 343732 990140
rect 325752 990100 343732 990128
rect 325752 990088 325758 990100
rect 343726 990088 343732 990100
rect 343784 990088 343790 990140
rect 628650 990088 628656 990140
rect 628708 990088 628714 990140
rect 629294 990088 629300 990140
rect 629352 990128 629358 990140
rect 673546 990128 673552 990140
rect 629352 990100 673552 990128
rect 629352 990088 629358 990100
rect 673546 990088 673552 990100
rect 673604 990088 673610 990140
rect 42518 990020 42524 990072
rect 42576 990060 42582 990072
rect 88352 990060 88380 990088
rect 42576 990032 88380 990060
rect 628668 990060 628696 990088
rect 673454 990060 673460 990072
rect 628668 990032 673460 990060
rect 42576 990020 42582 990032
rect 673454 990020 673460 990032
rect 673512 990020 673518 990072
rect 674834 985260 674840 985312
rect 674892 985300 674898 985312
rect 675110 985300 675116 985312
rect 674892 985272 675116 985300
rect 674892 985260 674898 985272
rect 675110 985260 675116 985272
rect 675168 985260 675174 985312
rect 41782 969348 41788 969400
rect 41840 969388 41846 969400
rect 42426 969388 42432 969400
rect 41840 969360 42432 969388
rect 41840 969348 41846 969360
rect 42426 969348 42432 969360
rect 42484 969348 42490 969400
rect 42518 968532 42524 968584
rect 42576 968532 42582 968584
rect 41782 968464 41788 968516
rect 41840 968504 41846 968516
rect 42536 968504 42564 968532
rect 42702 968504 42708 968516
rect 41840 968476 42708 968504
rect 41840 968464 41846 968476
rect 42702 968464 42708 968476
rect 42760 968464 42766 968516
rect 42518 966016 42524 966068
rect 42576 966056 42582 966068
rect 42702 966056 42708 966068
rect 42576 966028 42708 966056
rect 42576 966016 42582 966028
rect 42702 966016 42708 966028
rect 42760 966016 42766 966068
rect 674650 966016 674656 966068
rect 674708 966056 674714 966068
rect 674834 966056 674840 966068
rect 674708 966028 674840 966056
rect 674708 966016 674714 966028
rect 674834 966016 674840 966028
rect 674892 966016 674898 966068
rect 673454 964316 673460 964368
rect 673512 964356 673518 964368
rect 675386 964356 675392 964368
rect 673512 964328 675392 964356
rect 673512 964316 673518 964328
rect 675386 964316 675392 964328
rect 675444 964316 675450 964368
rect 673546 963704 673552 963756
rect 673604 963744 673610 963756
rect 675386 963744 675392 963756
rect 673604 963716 675392 963744
rect 673604 963704 673610 963716
rect 675386 963704 675392 963716
rect 675444 963704 675450 963756
rect 41782 962412 41788 962464
rect 41840 962452 41846 962464
rect 42426 962452 42432 962464
rect 41840 962424 42432 962452
rect 41840 962412 41846 962424
rect 42426 962412 42432 962424
rect 42484 962412 42490 962464
rect 42334 960440 42340 960492
rect 42392 960480 42398 960492
rect 42610 960480 42616 960492
rect 42392 960452 42616 960480
rect 42392 960440 42398 960452
rect 42610 960440 42616 960452
rect 42668 960440 42674 960492
rect 41782 957040 41788 957092
rect 41840 957080 41846 957092
rect 42610 957080 42616 957092
rect 41840 957052 42616 957080
rect 41840 957040 41846 957052
rect 42260 956820 42288 957052
rect 42610 957040 42616 957052
rect 42668 957040 42674 957092
rect 42242 956768 42248 956820
rect 42300 956768 42306 956820
rect 673638 953844 673644 953896
rect 673696 953884 673702 953896
rect 675386 953884 675392 953896
rect 673696 953856 675392 953884
rect 673696 953844 673702 953856
rect 675386 953844 675392 953856
rect 675444 953844 675450 953896
rect 42518 946636 42524 946688
rect 42576 946676 42582 946688
rect 42702 946676 42708 946688
rect 42576 946648 42708 946676
rect 42576 946636 42582 946648
rect 42702 946636 42708 946648
rect 42760 946636 42766 946688
rect 674650 932832 674656 932884
rect 674708 932832 674714 932884
rect 674668 932804 674696 932832
rect 674834 932804 674840 932816
rect 674668 932776 674840 932804
rect 674834 932764 674840 932776
rect 674892 932764 674898 932816
rect 42518 927392 42524 927444
rect 42576 927432 42582 927444
rect 42702 927432 42708 927444
rect 42576 927404 42708 927432
rect 42576 927392 42582 927404
rect 42702 927392 42708 927404
rect 42760 927392 42766 927444
rect 39666 922904 39672 922956
rect 39724 922944 39730 922956
rect 42242 922944 42248 922956
rect 39724 922916 42248 922944
rect 39724 922904 39730 922916
rect 42242 922904 42248 922916
rect 42300 922904 42306 922956
rect 39850 915084 39856 915136
rect 39908 915124 39914 915136
rect 41414 915124 41420 915136
rect 39908 915096 41420 915124
rect 39908 915084 39914 915096
rect 41414 915084 41420 915096
rect 41472 915124 41478 915136
rect 42426 915124 42432 915136
rect 41472 915096 42432 915124
rect 41472 915084 41478 915096
rect 42426 915084 42432 915096
rect 42484 915084 42490 915136
rect 673546 910732 673552 910784
rect 673604 910772 673610 910784
rect 677870 910772 677876 910784
rect 673604 910744 677876 910772
rect 673604 910732 673610 910744
rect 677870 910732 677876 910744
rect 677928 910732 677934 910784
rect 675294 908080 675300 908132
rect 675352 908120 675358 908132
rect 677502 908120 677508 908132
rect 675352 908092 677508 908120
rect 675352 908080 675358 908092
rect 677502 908080 677508 908092
rect 677560 908080 677566 908132
rect 42518 908012 42524 908064
rect 42576 908052 42582 908064
rect 42702 908052 42708 908064
rect 42576 908024 42708 908052
rect 42576 908012 42582 908024
rect 42702 908012 42708 908024
rect 42760 908012 42766 908064
rect 41506 906652 41512 906704
rect 41564 906692 41570 906704
rect 42334 906692 42340 906704
rect 41564 906664 42340 906692
rect 41564 906652 41570 906664
rect 42334 906652 42340 906664
rect 42392 906652 42398 906704
rect 674834 902612 674840 902624
rect 674668 902584 674840 902612
rect 674668 902556 674696 902584
rect 674834 902572 674840 902584
rect 674892 902572 674898 902624
rect 674650 902504 674656 902556
rect 674708 902504 674714 902556
rect 674650 894208 674656 894260
rect 674708 894248 674714 894260
rect 674834 894248 674840 894260
rect 674708 894220 674840 894248
rect 674708 894208 674714 894220
rect 674834 894208 674840 894220
rect 674892 894208 674898 894260
rect 42518 888700 42524 888752
rect 42576 888740 42582 888752
rect 42702 888740 42708 888752
rect 42576 888712 42708 888740
rect 42576 888700 42582 888712
rect 42702 888700 42708 888712
rect 42760 888700 42766 888752
rect 41414 875848 41420 875900
rect 41472 875888 41478 875900
rect 42426 875888 42432 875900
rect 41472 875860 42432 875888
rect 41472 875848 41478 875860
rect 42426 875848 42432 875860
rect 42484 875848 42490 875900
rect 673454 875780 673460 875832
rect 673512 875820 673518 875832
rect 675386 875820 675392 875832
rect 673512 875792 675392 875820
rect 673512 875780 673518 875792
rect 675386 875780 675392 875792
rect 675444 875780 675450 875832
rect 673546 874828 673552 874880
rect 673604 874868 673610 874880
rect 675386 874868 675392 874880
rect 673604 874840 675392 874868
rect 673604 874828 673610 874840
rect 675386 874828 675392 874840
rect 675444 874828 675450 874880
rect 675202 870136 675208 870188
rect 675260 870176 675266 870188
rect 675386 870176 675392 870188
rect 675260 870148 675392 870176
rect 675260 870136 675266 870148
rect 675386 870136 675392 870148
rect 675444 870136 675450 870188
rect 673638 864968 673644 865020
rect 673696 865008 673702 865020
rect 675386 865008 675392 865020
rect 673696 864980 675392 865008
rect 673696 864968 673702 864980
rect 675386 864968 675392 864980
rect 675444 864968 675450 865020
rect 675294 862792 675300 862844
rect 675352 862792 675358 862844
rect 675312 862640 675340 862792
rect 675294 862588 675300 862640
rect 675352 862588 675358 862640
rect 42518 850076 42524 850128
rect 42576 850116 42582 850128
rect 42702 850116 42708 850128
rect 42576 850088 42708 850116
rect 42576 850076 42582 850088
rect 42702 850076 42708 850088
rect 42760 850076 42766 850128
rect 44174 836272 44180 836324
rect 44232 836312 44238 836324
rect 44358 836312 44364 836324
rect 44232 836284 44364 836312
rect 44232 836272 44238 836284
rect 44358 836272 44364 836284
rect 44416 836272 44422 836324
rect 674926 836272 674932 836324
rect 674984 836312 674990 836324
rect 675110 836312 675116 836324
rect 674984 836284 675116 836312
rect 674984 836272 674990 836284
rect 675110 836272 675116 836284
rect 675168 836272 675174 836324
rect 674926 827908 674932 827960
rect 674984 827948 674990 827960
rect 677594 827948 677600 827960
rect 674984 827920 677600 827948
rect 674984 827908 674990 827920
rect 677594 827908 677600 827920
rect 677652 827908 677658 827960
rect 39758 827500 39764 827552
rect 39816 827540 39822 827552
rect 44542 827540 44548 827552
rect 39816 827512 44548 827540
rect 39816 827500 39822 827512
rect 44542 827500 44548 827512
rect 44600 827500 44606 827552
rect 674742 823420 674748 823472
rect 674800 823460 674806 823472
rect 676122 823460 676128 823472
rect 674800 823432 676128 823460
rect 674800 823420 674806 823432
rect 676122 823420 676128 823432
rect 676180 823420 676186 823472
rect 675202 818660 675208 818712
rect 675260 818700 675266 818712
rect 676122 818700 676128 818712
rect 675260 818672 676128 818700
rect 675260 818660 675266 818672
rect 676122 818660 676128 818672
rect 676180 818700 676186 818712
rect 677410 818700 677416 818712
rect 676180 818672 677416 818700
rect 676180 818660 676186 818672
rect 677410 818660 677416 818672
rect 677468 818660 677474 818712
rect 44358 805944 44364 805996
rect 44416 805984 44422 805996
rect 44542 805984 44548 805996
rect 44416 805956 44548 805984
rect 44416 805944 44422 805956
rect 44542 805944 44548 805956
rect 44600 805944 44606 805996
rect 41782 799552 41788 799604
rect 41840 799592 41846 799604
rect 42426 799592 42432 799604
rect 41840 799564 42432 799592
rect 41840 799552 41846 799564
rect 42426 799552 42432 799564
rect 42484 799552 42490 799604
rect 41782 798668 41788 798720
rect 41840 798708 41846 798720
rect 42702 798708 42708 798720
rect 41840 798680 42708 798708
rect 41840 798668 41846 798680
rect 42702 798668 42708 798680
rect 42760 798668 42766 798720
rect 41782 792548 41788 792600
rect 41840 792588 41846 792600
rect 42426 792588 42432 792600
rect 41840 792560 42432 792588
rect 41840 792548 41846 792560
rect 42426 792548 42432 792560
rect 42484 792548 42490 792600
rect 42886 792072 42892 792124
rect 42944 792112 42950 792124
rect 43070 792112 43076 792124
rect 42944 792084 43076 792112
rect 42944 792072 42950 792084
rect 43070 792072 43076 792084
rect 43128 792072 43134 792124
rect 674834 792072 674840 792124
rect 674892 792112 674898 792124
rect 675110 792112 675116 792124
rect 674892 792084 675116 792112
rect 674892 792072 674898 792084
rect 675110 792072 675116 792084
rect 675168 792072 675174 792124
rect 41782 787856 41788 787908
rect 41840 787896 41846 787908
rect 42426 787896 42432 787908
rect 41840 787868 42432 787896
rect 41840 787856 41846 787868
rect 42426 787856 42432 787868
rect 42484 787896 42490 787908
rect 42610 787896 42616 787908
rect 42484 787868 42616 787896
rect 42484 787856 42490 787868
rect 42610 787856 42616 787868
rect 42668 787856 42674 787908
rect 673454 786904 673460 786956
rect 673512 786944 673518 786956
rect 673730 786944 673736 786956
rect 673512 786916 673736 786944
rect 673512 786904 673518 786916
rect 673730 786904 673736 786916
rect 673788 786944 673794 786956
rect 675386 786944 675392 786956
rect 673788 786916 675392 786944
rect 673788 786904 673794 786916
rect 675386 786904 675392 786916
rect 675444 786904 675450 786956
rect 41782 786632 41788 786684
rect 41840 786672 41846 786684
rect 42610 786672 42616 786684
rect 41840 786644 42616 786672
rect 41840 786632 41846 786644
rect 42610 786632 42616 786644
rect 42668 786632 42674 786684
rect 673546 786360 673552 786412
rect 673604 786400 673610 786412
rect 675386 786400 675392 786412
rect 673604 786372 675392 786400
rect 673604 786360 673610 786372
rect 675386 786360 675392 786372
rect 675444 786360 675450 786412
rect 675018 780988 675024 781040
rect 675076 781028 675082 781040
rect 675386 781028 675392 781040
rect 675076 781000 675392 781028
rect 675076 780988 675082 781000
rect 675386 780988 675392 781000
rect 675444 780988 675450 781040
rect 673638 774868 673644 774920
rect 673696 774908 673702 774920
rect 673914 774908 673920 774920
rect 673696 774880 673920 774908
rect 673696 774868 673702 774880
rect 673914 774868 673920 774880
rect 673972 774908 673978 774920
rect 675386 774908 675392 774920
rect 673972 774880 675392 774908
rect 673972 774868 673978 774880
rect 675386 774868 675392 774880
rect 675444 774868 675450 774920
rect 675018 773984 675024 774036
rect 675076 774024 675082 774036
rect 675386 774024 675392 774036
rect 675076 773996 675392 774024
rect 675076 773984 675082 773996
rect 675386 773984 675392 773996
rect 675444 773984 675450 774036
rect 42794 772828 42800 772880
rect 42852 772868 42858 772880
rect 43070 772868 43076 772880
rect 42852 772840 43076 772868
rect 42852 772828 42858 772840
rect 43070 772828 43076 772840
rect 43128 772828 43134 772880
rect 44358 767320 44364 767372
rect 44416 767360 44422 767372
rect 44542 767360 44548 767372
rect 44416 767332 44548 767360
rect 44416 767320 44422 767332
rect 44542 767320 44548 767332
rect 44600 767320 44606 767372
rect 42426 756508 42432 756560
rect 42484 756548 42490 756560
rect 42794 756548 42800 756560
rect 42484 756520 42800 756548
rect 42484 756508 42490 756520
rect 42794 756508 42800 756520
rect 42852 756508 42858 756560
rect 41782 756372 41788 756424
rect 41840 756412 41846 756424
rect 42426 756412 42432 756424
rect 41840 756384 42432 756412
rect 41840 756372 41846 756384
rect 42426 756372 42432 756384
rect 42484 756372 42490 756424
rect 41782 754468 41788 754520
rect 41840 754468 41846 754520
rect 41800 754440 41828 754468
rect 42702 754440 42708 754452
rect 41800 754412 42708 754440
rect 42702 754400 42708 754412
rect 42760 754400 42766 754452
rect 41782 749368 41788 749420
rect 41840 749408 41846 749420
rect 42426 749408 42432 749420
rect 41840 749380 42432 749408
rect 41840 749368 41846 749380
rect 42426 749368 42432 749380
rect 42484 749368 42490 749420
rect 673546 746512 673552 746564
rect 673604 746552 673610 746564
rect 674006 746552 674012 746564
rect 673604 746524 674012 746552
rect 673604 746512 673610 746524
rect 674006 746512 674012 746524
rect 674064 746512 674070 746564
rect 41782 745084 41788 745136
rect 41840 745124 41846 745136
rect 42426 745124 42432 745136
rect 41840 745096 42432 745124
rect 41840 745084 41846 745096
rect 42426 745084 42432 745096
rect 42484 745124 42490 745136
rect 42794 745124 42800 745136
rect 42484 745096 42800 745124
rect 42484 745084 42490 745096
rect 42794 745084 42800 745096
rect 42852 745084 42858 745136
rect 41782 744404 41788 744456
rect 41840 744444 41846 744456
rect 42610 744444 42616 744456
rect 41840 744416 42616 744444
rect 41840 744404 41846 744416
rect 42610 744404 42616 744416
rect 42668 744404 42674 744456
rect 673730 741888 673736 741940
rect 673788 741928 673794 741940
rect 675386 741928 675392 741940
rect 673788 741900 675392 741928
rect 673788 741888 673794 741900
rect 675386 741888 675392 741900
rect 675444 741888 675450 741940
rect 674006 740664 674012 740716
rect 674064 740704 674070 740716
rect 675386 740704 675392 740716
rect 674064 740676 675392 740704
rect 674064 740664 674070 740676
rect 675386 740664 675392 740676
rect 675444 740664 675450 740716
rect 44174 739576 44180 739628
rect 44232 739616 44238 739628
rect 44450 739616 44456 739628
rect 44232 739588 44456 739616
rect 44232 739576 44238 739588
rect 44450 739576 44456 739588
rect 44508 739576 44514 739628
rect 674834 739576 674840 739628
rect 674892 739616 674898 739628
rect 674926 739616 674932 739628
rect 674892 739588 674932 739616
rect 674892 739576 674898 739588
rect 674926 739576 674932 739588
rect 674984 739576 674990 739628
rect 675018 735972 675024 736024
rect 675076 736012 675082 736024
rect 675386 736012 675392 736024
rect 675076 735984 675392 736012
rect 675076 735972 675082 735984
rect 675386 735972 675392 735984
rect 675444 735972 675450 736024
rect 674834 734068 674840 734120
rect 674892 734108 674898 734120
rect 674926 734108 674932 734120
rect 674892 734080 674932 734108
rect 674892 734068 674898 734080
rect 674926 734068 674932 734080
rect 674984 734068 674990 734120
rect 42426 730804 42432 730856
rect 42484 730844 42490 730856
rect 42794 730844 42800 730856
rect 42484 730816 42800 730844
rect 42484 730804 42490 730816
rect 42794 730804 42800 730816
rect 42852 730804 42858 730856
rect 673546 730124 673552 730176
rect 673604 730164 673610 730176
rect 673914 730164 673920 730176
rect 673604 730136 673920 730164
rect 673604 730124 673610 730136
rect 673914 730124 673920 730136
rect 673972 730164 673978 730176
rect 675386 730164 675392 730176
rect 673972 730136 675392 730164
rect 673972 730124 673978 730136
rect 675386 730124 675392 730136
rect 675444 730124 675450 730176
rect 673638 729988 673644 730040
rect 673696 730028 673702 730040
rect 674006 730028 674012 730040
rect 673696 730000 674012 730028
rect 673696 729988 673702 730000
rect 674006 729988 674012 730000
rect 674064 729988 674070 730040
rect 675018 729036 675024 729088
rect 675076 729076 675082 729088
rect 675386 729076 675392 729088
rect 675076 729048 675392 729076
rect 675076 729036 675082 729048
rect 675386 729036 675392 729048
rect 675444 729036 675450 729088
rect 44174 720400 44180 720452
rect 44232 720440 44238 720452
rect 44450 720440 44456 720452
rect 44232 720412 44456 720440
rect 44232 720400 44238 720412
rect 44450 720400 44456 720412
rect 44508 720400 44514 720452
rect 674834 714756 674840 714808
rect 674892 714796 674898 714808
rect 675018 714796 675024 714808
rect 674892 714768 675024 714796
rect 674892 714756 674898 714768
rect 675018 714756 675024 714768
rect 675076 714756 675082 714808
rect 41782 713124 41788 713176
rect 41840 713164 41846 713176
rect 42426 713164 42432 713176
rect 41840 713136 42432 713164
rect 41840 713124 41846 713136
rect 42426 713124 42432 713136
rect 42484 713124 42490 713176
rect 41782 711288 41788 711340
rect 41840 711288 41846 711340
rect 41800 711260 41828 711288
rect 42886 711260 42892 711272
rect 41800 711232 42892 711260
rect 42886 711220 42892 711232
rect 42944 711220 42950 711272
rect 42518 708704 42524 708756
rect 42576 708744 42582 708756
rect 42794 708744 42800 708756
rect 42576 708716 42800 708744
rect 42576 708704 42582 708716
rect 42794 708704 42800 708716
rect 42852 708704 42858 708756
rect 41782 706188 41788 706240
rect 41840 706228 41846 706240
rect 42426 706228 42432 706240
rect 41840 706200 42432 706228
rect 41840 706188 41846 706200
rect 42426 706188 42432 706200
rect 42484 706188 42490 706240
rect 41782 700884 41788 700936
rect 41840 700924 41846 700936
rect 42518 700924 42524 700936
rect 41840 700896 42524 700924
rect 41840 700884 41846 700896
rect 42518 700884 42524 700896
rect 42576 700924 42582 700936
rect 42702 700924 42708 700936
rect 42576 700896 42708 700924
rect 42576 700884 42582 700896
rect 42702 700884 42708 700896
rect 42760 700884 42766 700936
rect 41782 700544 41788 700596
rect 41840 700584 41846 700596
rect 42610 700584 42616 700596
rect 41840 700556 42616 700584
rect 41840 700544 41846 700556
rect 42610 700544 42616 700556
rect 42668 700544 42674 700596
rect 673454 695920 673460 695972
rect 673512 695960 673518 695972
rect 673730 695960 673736 695972
rect 673512 695932 673736 695960
rect 673512 695920 673518 695932
rect 673730 695920 673736 695932
rect 673788 695960 673794 695972
rect 675386 695960 675392 695972
rect 673788 695932 675392 695960
rect 673788 695920 673794 695932
rect 675386 695920 675392 695932
rect 675444 695920 675450 695972
rect 674834 695512 674840 695564
rect 674892 695552 674898 695564
rect 675110 695552 675116 695564
rect 674892 695524 675116 695552
rect 674892 695512 674898 695524
rect 675110 695512 675116 695524
rect 675168 695512 675174 695564
rect 42886 695444 42892 695496
rect 42944 695484 42950 695496
rect 43070 695484 43076 695496
rect 42944 695456 43076 695484
rect 42944 695444 42950 695456
rect 43070 695444 43076 695456
rect 43128 695444 43134 695496
rect 673638 695308 673644 695360
rect 673696 695348 673702 695360
rect 675386 695348 675392 695360
rect 673696 695320 675392 695348
rect 673696 695308 673702 695320
rect 675386 695308 675392 695320
rect 675444 695308 675450 695360
rect 675018 691636 675024 691688
rect 675076 691676 675082 691688
rect 675386 691676 675392 691688
rect 675076 691648 675392 691676
rect 675076 691636 675082 691648
rect 675386 691636 675392 691648
rect 675444 691636 675450 691688
rect 673546 685176 673552 685228
rect 673604 685216 673610 685228
rect 675386 685216 675392 685228
rect 673604 685188 675392 685216
rect 673604 685176 673610 685188
rect 675386 685176 675392 685188
rect 675444 685176 675450 685228
rect 675018 684020 675024 684072
rect 675076 684060 675082 684072
rect 675386 684060 675392 684072
rect 675076 684032 675392 684060
rect 675076 684020 675082 684032
rect 675386 684020 675392 684032
rect 675444 684020 675450 684072
rect 44174 681708 44180 681760
rect 44232 681748 44238 681760
rect 44450 681748 44456 681760
rect 44232 681720 44456 681748
rect 44232 681708 44238 681720
rect 44450 681708 44456 681720
rect 44508 681708 44514 681760
rect 674834 676132 674840 676184
rect 674892 676172 674898 676184
rect 675018 676172 675024 676184
rect 674892 676144 675024 676172
rect 674892 676132 674898 676144
rect 675018 676132 675024 676144
rect 675076 676132 675082 676184
rect 41782 669944 41788 669996
rect 41840 669984 41846 669996
rect 42426 669984 42432 669996
rect 41840 669956 42432 669984
rect 41840 669944 41846 669956
rect 42426 669944 42432 669956
rect 42484 669944 42490 669996
rect 41782 669060 41788 669112
rect 41840 669100 41846 669112
rect 42610 669100 42616 669112
rect 41840 669072 42616 669100
rect 41840 669060 41846 669072
rect 42610 669060 42616 669072
rect 42668 669100 42674 669112
rect 42886 669100 42892 669112
rect 42668 669072 42892 669100
rect 42668 669060 42674 669072
rect 42886 669060 42892 669072
rect 42944 669060 42950 669112
rect 41782 663008 41788 663060
rect 41840 663048 41846 663060
rect 42426 663048 42432 663060
rect 41840 663020 42432 663048
rect 41840 663008 41846 663020
rect 42426 663008 42432 663020
rect 42484 663008 42490 663060
rect 41782 657636 41788 657688
rect 41840 657676 41846 657688
rect 42702 657676 42708 657688
rect 41840 657648 42708 657676
rect 41840 657636 41846 657648
rect 42702 657636 42708 657648
rect 42760 657676 42766 657688
rect 42978 657676 42984 657688
rect 42760 657648 42984 657676
rect 42760 657636 42766 657648
rect 42978 657636 42984 657648
rect 43036 657636 43042 657688
rect 41782 657092 41788 657144
rect 41840 657132 41846 657144
rect 42518 657132 42524 657144
rect 41840 657104 42524 657132
rect 41840 657092 41846 657104
rect 42518 657092 42524 657104
rect 42576 657132 42582 657144
rect 42702 657132 42708 657144
rect 42576 657104 42708 657132
rect 42576 657092 42582 657104
rect 42702 657092 42708 657104
rect 42760 657092 42766 657144
rect 674834 656888 674840 656940
rect 674892 656928 674898 656940
rect 675110 656928 675116 656940
rect 674892 656900 675116 656928
rect 674892 656888 674898 656900
rect 675110 656888 675116 656900
rect 675168 656888 675174 656940
rect 673454 651720 673460 651772
rect 673512 651760 673518 651772
rect 675386 651760 675392 651772
rect 673512 651732 675392 651760
rect 673512 651720 673518 651732
rect 675386 651720 675392 651732
rect 675444 651720 675450 651772
rect 673638 651108 673644 651160
rect 673696 651148 673702 651160
rect 675386 651148 675392 651160
rect 673696 651120 675392 651148
rect 673696 651108 673702 651120
rect 675386 651108 675392 651120
rect 675444 651108 675450 651160
rect 675018 645736 675024 645788
rect 675076 645776 675082 645788
rect 675386 645776 675392 645788
rect 675076 645748 675392 645776
rect 675076 645736 675082 645748
rect 675386 645736 675392 645748
rect 675444 645736 675450 645788
rect 44174 643084 44180 643136
rect 44232 643124 44238 643136
rect 44450 643124 44456 643136
rect 44232 643096 44456 643124
rect 44232 643084 44238 643096
rect 44450 643084 44456 643096
rect 44508 643084 44514 643136
rect 673546 639684 673552 639736
rect 673604 639724 673610 639736
rect 675386 639724 675392 639736
rect 673604 639696 675392 639724
rect 673604 639684 673610 639696
rect 675386 639684 675392 639696
rect 675444 639684 675450 639736
rect 675018 638800 675024 638852
rect 675076 638840 675082 638852
rect 675386 638840 675392 638852
rect 675076 638812 675392 638840
rect 675076 638800 675082 638812
rect 675386 638800 675392 638812
rect 675444 638800 675450 638852
rect 674742 637576 674748 637628
rect 674800 637616 674806 637628
rect 675110 637616 675116 637628
rect 674800 637588 675116 637616
rect 674800 637576 674806 637588
rect 675110 637576 675116 637588
rect 675168 637576 675174 637628
rect 42518 633360 42524 633412
rect 42576 633400 42582 633412
rect 42702 633400 42708 633412
rect 42576 633372 42708 633400
rect 42576 633360 42582 633372
rect 42702 633360 42708 633372
rect 42760 633360 42766 633412
rect 41782 626764 41788 626816
rect 41840 626804 41846 626816
rect 42426 626804 42432 626816
rect 41840 626776 42432 626804
rect 41840 626764 41846 626776
rect 42426 626764 42432 626776
rect 42484 626764 42490 626816
rect 41782 625880 41788 625932
rect 41840 625920 41846 625932
rect 42702 625920 42708 625932
rect 41840 625892 42708 625920
rect 41840 625880 41846 625892
rect 42702 625880 42708 625892
rect 42760 625880 42766 625932
rect 674742 623772 674748 623824
rect 674800 623772 674806 623824
rect 673546 623704 673552 623756
rect 673604 623704 673610 623756
rect 44174 623636 44180 623688
rect 44232 623676 44238 623688
rect 44450 623676 44456 623688
rect 44232 623648 44456 623676
rect 44232 623636 44238 623648
rect 44450 623636 44456 623648
rect 44508 623636 44514 623688
rect 673564 623676 673592 623704
rect 673822 623676 673828 623688
rect 673564 623648 673828 623676
rect 673822 623636 673828 623648
rect 673880 623636 673886 623688
rect 674760 623676 674788 623772
rect 674926 623676 674932 623688
rect 674760 623648 674932 623676
rect 674926 623636 674932 623648
rect 674984 623636 674990 623688
rect 41782 619760 41788 619812
rect 41840 619800 41846 619812
rect 42426 619800 42432 619812
rect 41840 619772 42432 619800
rect 41840 619760 41846 619772
rect 42426 619760 42432 619772
rect 42484 619760 42490 619812
rect 42702 618196 42708 618248
rect 42760 618236 42766 618248
rect 42978 618236 42984 618248
rect 42760 618208 42984 618236
rect 42760 618196 42766 618208
rect 42978 618196 42984 618208
rect 43036 618196 43042 618248
rect 674558 618196 674564 618248
rect 674616 618236 674622 618248
rect 674926 618236 674932 618248
rect 674616 618208 674932 618236
rect 674616 618196 674622 618208
rect 674926 618196 674932 618208
rect 674984 618196 674990 618248
rect 41782 614388 41788 614440
rect 41840 614428 41846 614440
rect 42426 614428 42432 614440
rect 41840 614400 42432 614428
rect 41840 614388 41846 614400
rect 42426 614388 42432 614400
rect 42484 614428 42490 614440
rect 42794 614428 42800 614440
rect 42484 614400 42800 614428
rect 42484 614388 42490 614400
rect 42794 614388 42800 614400
rect 42852 614388 42858 614440
rect 41782 614048 41788 614100
rect 41840 614088 41846 614100
rect 42610 614088 42616 614100
rect 41840 614060 42616 614088
rect 41840 614048 41846 614060
rect 42610 614048 42616 614060
rect 42668 614048 42674 614100
rect 673454 606704 673460 606756
rect 673512 606744 673518 606756
rect 674742 606744 674748 606756
rect 673512 606716 674748 606744
rect 673512 606704 673518 606716
rect 674742 606704 674748 606716
rect 674800 606744 674806 606756
rect 675386 606744 675392 606756
rect 674800 606716 675392 606744
rect 674800 606704 674806 606716
rect 675386 606704 675392 606716
rect 675444 606704 675450 606756
rect 673638 605480 673644 605532
rect 673696 605520 673702 605532
rect 675386 605520 675392 605532
rect 673696 605492 675392 605520
rect 673696 605480 673702 605492
rect 675386 605480 675392 605492
rect 675444 605480 675450 605532
rect 44174 604460 44180 604512
rect 44232 604500 44238 604512
rect 44450 604500 44456 604512
rect 44232 604472 44456 604500
rect 44232 604460 44238 604472
rect 44450 604460 44456 604472
rect 44508 604460 44514 604512
rect 673638 604460 673644 604512
rect 673696 604500 673702 604512
rect 673914 604500 673920 604512
rect 673696 604472 673920 604500
rect 673696 604460 673702 604472
rect 673914 604460 673920 604472
rect 673972 604460 673978 604512
rect 675110 600788 675116 600840
rect 675168 600828 675174 600840
rect 675386 600828 675392 600840
rect 675168 600800 675392 600828
rect 675168 600788 675174 600800
rect 675386 600788 675392 600800
rect 675444 600788 675450 600840
rect 674558 599020 674564 599072
rect 674616 599060 674622 599072
rect 674834 599060 674840 599072
rect 674616 599032 674840 599060
rect 674616 599020 674622 599032
rect 674834 599020 674840 599032
rect 674892 599020 674898 599072
rect 674650 598884 674656 598936
rect 674708 598924 674714 598936
rect 674742 598924 674748 598936
rect 674708 598896 674748 598924
rect 674708 598884 674714 598896
rect 674742 598884 674748 598896
rect 674800 598884 674806 598936
rect 674834 598884 674840 598936
rect 674892 598924 674898 598936
rect 675018 598924 675024 598936
rect 674892 598896 675024 598924
rect 674892 598884 674898 598896
rect 675018 598884 675024 598896
rect 675076 598884 675082 598936
rect 673638 594872 673644 594924
rect 673696 594912 673702 594924
rect 673822 594912 673828 594924
rect 673696 594884 673828 594912
rect 673696 594872 673702 594884
rect 673822 594872 673828 594884
rect 673880 594912 673886 594924
rect 675386 594912 675392 594924
rect 673880 594884 675392 594912
rect 673880 594872 673886 594884
rect 675386 594872 675392 594884
rect 675444 594872 675450 594924
rect 675110 593784 675116 593836
rect 675168 593824 675174 593836
rect 675386 593824 675392 593836
rect 675168 593796 675392 593824
rect 675168 593784 675174 593796
rect 675386 593784 675392 593796
rect 675444 593784 675450 593836
rect 44174 585012 44180 585064
rect 44232 585052 44238 585064
rect 44450 585052 44456 585064
rect 44232 585024 44456 585052
rect 44232 585012 44238 585024
rect 44450 585012 44456 585024
rect 44508 585012 44514 585064
rect 42426 583652 42432 583704
rect 42484 583692 42490 583704
rect 42794 583692 42800 583704
rect 42484 583664 42800 583692
rect 42484 583652 42490 583664
rect 42794 583652 42800 583664
rect 42852 583652 42858 583704
rect 41782 583516 41788 583568
rect 41840 583556 41846 583568
rect 42426 583556 42432 583568
rect 41840 583528 42432 583556
rect 41840 583516 41846 583528
rect 42426 583516 42432 583528
rect 42484 583516 42490 583568
rect 41782 581680 41788 581732
rect 41840 581680 41846 581732
rect 41800 581652 41828 581680
rect 42702 581652 42708 581664
rect 41800 581624 42708 581652
rect 42702 581612 42708 581624
rect 42760 581652 42766 581664
rect 42978 581652 42984 581664
rect 42760 581624 42984 581652
rect 42760 581612 42766 581624
rect 42978 581612 42984 581624
rect 43036 581612 43042 581664
rect 674650 579572 674656 579624
rect 674708 579612 674714 579624
rect 675018 579612 675024 579624
rect 674708 579584 675024 579612
rect 674708 579572 674714 579584
rect 675018 579572 675024 579584
rect 675076 579572 675082 579624
rect 41782 576580 41788 576632
rect 41840 576620 41846 576632
rect 42426 576620 42432 576632
rect 41840 576592 42432 576620
rect 41840 576580 41846 576592
rect 42426 576580 42432 576592
rect 42484 576580 42490 576632
rect 41782 572228 41788 572280
rect 41840 572268 41846 572280
rect 42426 572268 42432 572280
rect 41840 572240 42432 572268
rect 41840 572228 41846 572240
rect 42426 572228 42432 572240
rect 42484 572268 42490 572280
rect 42794 572268 42800 572280
rect 42484 572240 42800 572268
rect 42484 572228 42490 572240
rect 42794 572228 42800 572240
rect 42852 572228 42858 572280
rect 41782 571616 41788 571668
rect 41840 571656 41846 571668
rect 42610 571656 42616 571668
rect 41840 571628 42616 571656
rect 41840 571616 41846 571628
rect 42610 571616 42616 571628
rect 42668 571616 42674 571668
rect 44174 565836 44180 565888
rect 44232 565876 44238 565888
rect 44450 565876 44456 565888
rect 44232 565848 44456 565876
rect 44232 565836 44238 565848
rect 44450 565836 44456 565848
rect 44508 565836 44514 565888
rect 44174 564272 44180 564324
rect 44232 564312 44238 564324
rect 44450 564312 44456 564324
rect 44232 564284 44456 564312
rect 44232 564272 44238 564284
rect 44450 564272 44456 564284
rect 44508 564272 44514 564324
rect 673822 561212 673828 561264
rect 673880 561252 673886 561264
rect 674742 561252 674748 561264
rect 673880 561224 674748 561252
rect 673880 561212 673886 561224
rect 674742 561212 674748 561224
rect 674800 561252 674806 561264
rect 675386 561252 675392 561264
rect 674800 561224 675392 561252
rect 674800 561212 674806 561224
rect 675386 561212 675392 561224
rect 675444 561212 675450 561264
rect 673914 560940 673920 560992
rect 673972 560980 673978 560992
rect 675386 560980 675392 560992
rect 673972 560952 675392 560980
rect 673972 560940 673978 560952
rect 675386 560940 675392 560952
rect 675444 560940 675450 560992
rect 674650 560260 674656 560312
rect 674708 560300 674714 560312
rect 674834 560300 674840 560312
rect 674708 560272 674840 560300
rect 674708 560260 674714 560272
rect 674834 560260 674840 560272
rect 674892 560260 674898 560312
rect 42426 556112 42432 556164
rect 42484 556152 42490 556164
rect 42794 556152 42800 556164
rect 42484 556124 42800 556152
rect 42484 556112 42490 556124
rect 42794 556112 42800 556124
rect 42852 556112 42858 556164
rect 675110 555568 675116 555620
rect 675168 555608 675174 555620
rect 675386 555608 675392 555620
rect 675168 555580 675392 555608
rect 675168 555568 675174 555580
rect 675386 555568 675392 555580
rect 675444 555568 675450 555620
rect 673638 550468 673644 550520
rect 673696 550508 673702 550520
rect 675386 550508 675392 550520
rect 673696 550480 675392 550508
rect 673696 550468 673702 550480
rect 675386 550468 675392 550480
rect 675444 550468 675450 550520
rect 675110 548632 675116 548684
rect 675168 548672 675174 548684
rect 675386 548672 675392 548684
rect 675168 548644 675392 548672
rect 675168 548632 675174 548644
rect 675386 548632 675392 548644
rect 675444 548632 675450 548684
rect 674834 540948 674840 541000
rect 674892 540988 674898 541000
rect 675018 540988 675024 541000
rect 674892 540960 675024 540988
rect 674892 540948 674898 540960
rect 675018 540948 675024 540960
rect 675076 540948 675082 541000
rect 41782 540336 41788 540388
rect 41840 540376 41846 540388
rect 42426 540376 42432 540388
rect 41840 540348 42432 540376
rect 41840 540336 41846 540348
rect 42426 540336 42432 540348
rect 42484 540336 42490 540388
rect 41782 538500 41788 538552
rect 41840 538540 41846 538552
rect 42702 538540 42708 538552
rect 41840 538512 42708 538540
rect 41840 538500 41846 538512
rect 42702 538500 42708 538512
rect 42760 538500 42766 538552
rect 41782 533400 41788 533452
rect 41840 533440 41846 533452
rect 42426 533440 42432 533452
rect 41840 533412 42432 533440
rect 41840 533400 41846 533412
rect 42426 533400 42432 533412
rect 42484 533400 42490 533452
rect 41782 529048 41788 529100
rect 41840 529088 41846 529100
rect 42426 529088 42432 529100
rect 41840 529060 42432 529088
rect 41840 529048 41846 529060
rect 42426 529048 42432 529060
rect 42484 529088 42490 529100
rect 42794 529088 42800 529100
rect 42484 529060 42800 529088
rect 42484 529048 42490 529060
rect 42794 529048 42800 529060
rect 42852 529048 42858 529100
rect 41782 527756 41788 527808
rect 41840 527796 41846 527808
rect 42610 527796 42616 527808
rect 41840 527768 42616 527796
rect 41840 527756 41846 527768
rect 42610 527756 42616 527768
rect 42668 527756 42674 527808
rect 44174 527144 44180 527196
rect 44232 527184 44238 527196
rect 44450 527184 44456 527196
rect 44232 527156 44456 527184
rect 44232 527144 44238 527156
rect 44450 527144 44456 527156
rect 44508 527144 44514 527196
rect 674926 514020 674932 514072
rect 674984 514060 674990 514072
rect 676030 514060 676036 514072
rect 674984 514032 676036 514060
rect 674984 514020 674990 514032
rect 676030 514020 676036 514032
rect 676088 514060 676094 514072
rect 677410 514060 677416 514072
rect 676088 514032 677416 514060
rect 676088 514020 676094 514032
rect 677410 514020 677416 514032
rect 677468 514020 677474 514072
rect 675202 513748 675208 513800
rect 675260 513788 675266 513800
rect 676122 513788 676128 513800
rect 675260 513760 676128 513788
rect 675260 513748 675266 513760
rect 676122 513748 676128 513760
rect 676180 513788 676186 513800
rect 677502 513788 677508 513800
rect 676180 513760 677508 513788
rect 676180 513748 676186 513760
rect 677502 513748 677508 513760
rect 677560 513748 677566 513800
rect 676122 507832 676128 507884
rect 676180 507872 676186 507884
rect 677410 507872 677416 507884
rect 676180 507844 677416 507872
rect 676180 507832 676186 507844
rect 677410 507832 677416 507844
rect 677468 507832 677474 507884
rect 44174 507696 44180 507748
rect 44232 507736 44238 507748
rect 44450 507736 44456 507748
rect 44232 507708 44456 507736
rect 44232 507696 44238 507708
rect 44450 507696 44456 507708
rect 44508 507696 44514 507748
rect 42150 498176 42156 498228
rect 42208 498216 42214 498228
rect 42426 498216 42432 498228
rect 42208 498188 42432 498216
rect 42208 498176 42214 498188
rect 42426 498176 42432 498188
rect 42484 498176 42490 498228
rect 44174 488520 44180 488572
rect 44232 488560 44238 488572
rect 44450 488560 44456 488572
rect 44232 488532 44456 488560
rect 44232 488520 44238 488532
rect 44450 488520 44456 488532
rect 44508 488520 44514 488572
rect 42150 478864 42156 478916
rect 42208 478904 42214 478916
rect 42426 478904 42432 478916
rect 42208 478876 42432 478904
rect 42208 478864 42214 478876
rect 42426 478864 42432 478876
rect 42484 478864 42490 478916
rect 42150 469140 42156 469192
rect 42208 469180 42214 469192
rect 42426 469180 42432 469192
rect 42208 469152 42432 469180
rect 42208 469140 42214 469152
rect 42426 469140 42432 469152
rect 42484 469140 42490 469192
rect 675294 467508 675300 467560
rect 675352 467548 675358 467560
rect 677502 467548 677508 467560
rect 675352 467520 677508 467548
rect 675352 467508 675358 467520
rect 677502 467508 677508 467520
rect 677560 467508 677566 467560
rect 39850 463632 39856 463684
rect 39908 463672 39914 463684
rect 42150 463672 42156 463684
rect 39908 463644 42156 463672
rect 39908 463632 39914 463644
rect 42150 463632 42156 463644
rect 42208 463632 42214 463684
rect 42610 463632 42616 463684
rect 42668 463672 42674 463684
rect 42886 463672 42892 463684
rect 42668 463644 42892 463672
rect 42668 463632 42674 463644
rect 42886 463632 42892 463644
rect 42944 463632 42950 463684
rect 673730 463632 673736 463684
rect 673788 463672 673794 463684
rect 673822 463672 673828 463684
rect 673788 463644 673828 463672
rect 673788 463632 673794 463644
rect 673822 463632 673828 463644
rect 673880 463632 673886 463684
rect 676214 459960 676220 460012
rect 676272 460000 676278 460012
rect 677686 460000 677692 460012
rect 676272 459972 677692 460000
rect 676272 459960 676278 459972
rect 677686 459960 677692 459972
rect 677744 459960 677750 460012
rect 39390 458192 39396 458244
rect 39448 458232 39454 458244
rect 42242 458232 42248 458244
rect 39448 458204 42248 458232
rect 39448 458192 39454 458204
rect 42242 458192 42248 458204
rect 42300 458192 42306 458244
rect 44174 449896 44180 449948
rect 44232 449936 44238 449948
rect 44358 449936 44364 449948
rect 44232 449908 44364 449936
rect 44232 449896 44238 449908
rect 44358 449896 44364 449908
rect 44416 449896 44422 449948
rect 673730 449828 673736 449880
rect 673788 449868 673794 449880
rect 673914 449868 673920 449880
rect 673788 449840 673920 449868
rect 673788 449828 673794 449840
rect 673914 449828 673920 449840
rect 673972 449828 673978 449880
rect 42058 442688 42064 442740
rect 42116 442728 42122 442740
rect 42334 442728 42340 442740
rect 42116 442700 42340 442728
rect 42116 442688 42122 442700
rect 42334 442688 42340 442700
rect 42392 442688 42398 442740
rect 42426 441532 42432 441584
rect 42484 441572 42490 441584
rect 42610 441572 42616 441584
rect 42484 441544 42616 441572
rect 42484 441532 42490 441544
rect 42610 441532 42616 441544
rect 42668 441532 42674 441584
rect 676306 440172 676312 440224
rect 676364 440212 676370 440224
rect 677686 440212 677692 440224
rect 676364 440184 677692 440212
rect 676364 440172 676370 440184
rect 677686 440172 677692 440184
rect 677744 440172 677750 440224
rect 674006 430652 674012 430704
rect 674064 430652 674070 430704
rect 673914 430516 673920 430568
rect 673972 430556 673978 430568
rect 674024 430556 674052 430652
rect 673972 430528 674052 430556
rect 673972 430516 673978 430528
rect 676030 427796 676036 427848
rect 676088 427836 676094 427848
rect 677502 427836 677508 427848
rect 676088 427808 677508 427836
rect 676088 427796 676094 427808
rect 677502 427796 677508 427808
rect 677560 427796 677566 427848
rect 42334 425008 42340 425060
rect 42392 425048 42398 425060
rect 42794 425048 42800 425060
rect 42392 425020 42800 425048
rect 42392 425008 42398 425020
rect 42794 425008 42800 425020
rect 42852 425008 42858 425060
rect 42426 422288 42432 422340
rect 42484 422328 42490 422340
rect 42518 422328 42524 422340
rect 42484 422300 42524 422328
rect 42484 422288 42490 422300
rect 42518 422288 42524 422300
rect 42576 422288 42582 422340
rect 676122 420724 676128 420776
rect 676180 420764 676186 420776
rect 677502 420764 677508 420776
rect 676180 420736 677508 420764
rect 676180 420724 676186 420736
rect 677502 420724 677508 420736
rect 677560 420724 677566 420776
rect 42518 411312 42524 411324
rect 42444 411284 42524 411312
rect 42444 411256 42472 411284
rect 42518 411272 42524 411284
rect 42576 411272 42582 411324
rect 44174 411272 44180 411324
rect 44232 411312 44238 411324
rect 44358 411312 44364 411324
rect 44232 411284 44364 411312
rect 44232 411272 44238 411284
rect 44358 411272 44364 411284
rect 44416 411272 44422 411324
rect 42426 411204 42432 411256
rect 42484 411204 42490 411256
rect 41782 411068 41788 411120
rect 41840 411108 41846 411120
rect 42702 411108 42708 411120
rect 41840 411080 42708 411108
rect 41840 411068 41846 411080
rect 42702 411068 42708 411080
rect 42760 411068 42766 411120
rect 673086 408484 673092 408536
rect 673144 408524 673150 408536
rect 676306 408524 676312 408536
rect 673144 408496 676312 408524
rect 673144 408484 673150 408496
rect 676306 408484 676312 408496
rect 676364 408484 676370 408536
rect 41782 401344 41788 401396
rect 41840 401384 41846 401396
rect 42794 401384 42800 401396
rect 41840 401356 42800 401384
rect 41840 401344 41846 401356
rect 42794 401344 42800 401356
rect 42852 401344 42858 401396
rect 42150 397808 42156 397860
rect 42208 397848 42214 397860
rect 42794 397848 42800 397860
rect 42208 397820 42800 397848
rect 42208 397808 42214 397820
rect 42794 397808 42800 397820
rect 42852 397808 42858 397860
rect 675294 388628 675300 388680
rect 675352 388668 675358 388680
rect 676214 388668 676220 388680
rect 675352 388640 676220 388668
rect 675352 388628 675358 388640
rect 676214 388628 676220 388640
rect 676272 388628 676278 388680
rect 673454 384004 673460 384056
rect 673512 384044 673518 384056
rect 675386 384044 675392 384056
rect 673512 384016 675392 384044
rect 673512 384004 673518 384016
rect 675386 384004 675392 384016
rect 675444 384004 675450 384056
rect 673638 382712 673644 382764
rect 673696 382752 673702 382764
rect 675386 382752 675392 382764
rect 673696 382724 675392 382752
rect 673696 382712 673702 382724
rect 675386 382712 675392 382724
rect 675444 382712 675450 382764
rect 44174 372580 44180 372632
rect 44232 372620 44238 372632
rect 44358 372620 44364 372632
rect 44232 372592 44364 372620
rect 44232 372580 44238 372592
rect 44358 372580 44364 372592
rect 44416 372580 44422 372632
rect 673546 372308 673552 372360
rect 673604 372348 673610 372360
rect 675386 372348 675392 372360
rect 673604 372320 675392 372348
rect 673604 372308 673610 372320
rect 675386 372308 675392 372320
rect 675444 372308 675450 372360
rect 42426 370336 42432 370388
rect 42484 370376 42490 370388
rect 42702 370376 42708 370388
rect 42484 370348 42708 370376
rect 42484 370336 42490 370348
rect 42702 370336 42708 370348
rect 42760 370336 42766 370388
rect 42150 370200 42156 370252
rect 42208 370240 42214 370252
rect 42426 370240 42432 370252
rect 42208 370212 42432 370240
rect 42208 370200 42214 370212
rect 42426 370200 42432 370212
rect 42484 370200 42490 370252
rect 41782 367684 41788 367736
rect 41840 367724 41846 367736
rect 42518 367724 42524 367736
rect 41840 367696 42524 367724
rect 41840 367684 41846 367696
rect 42518 367684 42524 367696
rect 42576 367684 42582 367736
rect 41782 358232 41788 358284
rect 41840 358272 41846 358284
rect 42426 358272 42432 358284
rect 41840 358244 42432 358272
rect 41840 358232 41846 358244
rect 42426 358232 42432 358244
rect 42484 358272 42490 358284
rect 42610 358272 42616 358284
rect 42484 358244 42616 358272
rect 42484 358232 42490 358244
rect 42610 358232 42616 358244
rect 42668 358232 42674 358284
rect 41782 357280 41788 357332
rect 41840 357320 41846 357332
rect 42702 357320 42708 357332
rect 41840 357292 42708 357320
rect 41840 357280 41846 357292
rect 42702 357280 42708 357292
rect 42760 357280 42766 357332
rect 42426 356600 42432 356652
rect 42484 356640 42490 356652
rect 42702 356640 42708 356652
rect 42484 356612 42708 356640
rect 42484 356600 42490 356612
rect 42702 356600 42708 356612
rect 42760 356600 42766 356652
rect 42518 353200 42524 353252
rect 42576 353240 42582 353252
rect 42702 353240 42708 353252
rect 42576 353212 42708 353240
rect 42576 353200 42582 353212
rect 42702 353200 42708 353212
rect 42760 353200 42766 353252
rect 42334 339600 42340 339652
rect 42392 339640 42398 339652
rect 42610 339640 42616 339652
rect 42392 339612 42616 339640
rect 42392 339600 42398 339612
rect 42610 339600 42616 339612
rect 42668 339600 42674 339652
rect 673454 338104 673460 338156
rect 673512 338144 673518 338156
rect 673730 338144 673736 338156
rect 673512 338116 673736 338144
rect 673512 338104 673518 338116
rect 673730 338104 673736 338116
rect 673788 338144 673794 338156
rect 675386 338144 675392 338156
rect 673788 338116 675392 338144
rect 673788 338104 673794 338116
rect 675386 338104 675392 338116
rect 675444 338104 675450 338156
rect 673638 337492 673644 337544
rect 673696 337532 673702 337544
rect 675386 337532 675392 337544
rect 673696 337504 675392 337532
rect 673696 337492 673702 337504
rect 675386 337492 675392 337504
rect 675444 337492 675450 337544
rect 44174 333956 44180 334008
rect 44232 333996 44238 334008
rect 44358 333996 44364 334008
rect 44232 333968 44364 333996
rect 44232 333956 44238 333968
rect 44358 333956 44364 333968
rect 44416 333956 44422 334008
rect 673546 328040 673552 328092
rect 673604 328080 673610 328092
rect 675386 328080 675392 328092
rect 673604 328052 675392 328080
rect 673604 328040 673610 328052
rect 675386 328040 675392 328052
rect 675444 328040 675450 328092
rect 41782 324504 41788 324556
rect 41840 324544 41846 324556
rect 42702 324544 42708 324556
rect 41840 324516 42708 324544
rect 41840 324504 41846 324516
rect 42702 324504 42708 324516
rect 42760 324504 42766 324556
rect 41782 313488 41788 313540
rect 41840 313528 41846 313540
rect 42426 313528 42432 313540
rect 41840 313500 42432 313528
rect 41840 313488 41846 313500
rect 42426 313488 42432 313500
rect 42484 313528 42490 313540
rect 42610 313528 42616 313540
rect 42484 313500 42616 313528
rect 42484 313488 42490 313500
rect 42610 313488 42616 313500
rect 42668 313488 42674 313540
rect 673730 293836 673736 293888
rect 673788 293876 673794 293888
rect 674006 293876 674012 293888
rect 673788 293848 674012 293876
rect 673788 293836 673794 293848
rect 674006 293836 674012 293848
rect 674064 293876 674070 293888
rect 675386 293876 675392 293888
rect 674064 293848 675392 293876
rect 674064 293836 674070 293848
rect 675386 293836 675392 293848
rect 675444 293836 675450 293888
rect 673454 293564 673460 293616
rect 673512 293604 673518 293616
rect 673638 293604 673644 293616
rect 673512 293576 673644 293604
rect 673512 293564 673518 293576
rect 673638 293564 673644 293576
rect 673696 293604 673702 293616
rect 675386 293604 675392 293616
rect 673696 293576 675392 293604
rect 673696 293564 673702 293576
rect 675386 293564 675392 293576
rect 675444 293564 675450 293616
rect 42518 286628 42524 286680
rect 42576 286668 42582 286680
rect 42794 286668 42800 286680
rect 42576 286640 42800 286668
rect 42576 286628 42582 286640
rect 42794 286628 42800 286640
rect 42852 286628 42858 286680
rect 41782 282276 41788 282328
rect 41840 282316 41846 282328
rect 42426 282316 42432 282328
rect 41840 282288 42432 282316
rect 41840 282276 41846 282288
rect 42426 282276 42432 282288
rect 42484 282316 42490 282328
rect 42702 282316 42708 282328
rect 42484 282288 42708 282316
rect 42484 282276 42490 282288
rect 42702 282276 42708 282288
rect 42760 282276 42766 282328
rect 673546 282140 673552 282192
rect 673604 282140 673610 282192
rect 673564 282112 673592 282140
rect 675018 282112 675024 282124
rect 673564 282084 675024 282112
rect 675018 282072 675024 282084
rect 675076 282112 675082 282124
rect 675386 282112 675392 282124
rect 675076 282084 675392 282112
rect 675076 282072 675082 282084
rect 675386 282072 675392 282084
rect 675444 282072 675450 282124
rect 41782 270784 41788 270836
rect 41840 270824 41846 270836
rect 42794 270824 42800 270836
rect 41840 270796 42800 270824
rect 41840 270784 41846 270796
rect 42794 270784 42800 270796
rect 42852 270784 42858 270836
rect 42334 270716 42340 270768
rect 42392 270756 42398 270768
rect 42610 270756 42616 270768
rect 42392 270728 42616 270756
rect 42392 270716 42398 270728
rect 42610 270716 42616 270728
rect 42668 270716 42674 270768
rect 44266 270444 44272 270496
rect 44324 270484 44330 270496
rect 44358 270484 44364 270496
rect 44324 270456 44364 270484
rect 44324 270444 44330 270456
rect 44358 270444 44364 270456
rect 44416 270444 44422 270496
rect 675018 265044 675024 265056
rect 673748 265016 675024 265044
rect 673748 264988 673776 265016
rect 675018 265004 675024 265016
rect 675076 265004 675082 265056
rect 673730 264936 673736 264988
rect 673788 264936 673794 264988
rect 673822 264936 673828 264988
rect 673880 264976 673886 264988
rect 674006 264976 674012 264988
rect 673880 264948 674012 264976
rect 673880 264936 673886 264948
rect 674006 264936 674012 264948
rect 674064 264936 674070 264988
rect 44266 256708 44272 256760
rect 44324 256708 44330 256760
rect 44284 256624 44312 256708
rect 44266 256572 44272 256624
rect 44324 256572 44330 256624
rect 673546 249092 673552 249144
rect 673604 249132 673610 249144
rect 673822 249132 673828 249144
rect 673604 249104 673828 249132
rect 673604 249092 673610 249104
rect 673822 249092 673828 249104
rect 673880 249132 673886 249144
rect 675386 249132 675392 249144
rect 673880 249104 675392 249132
rect 673880 249092 673886 249104
rect 675386 249092 675392 249104
rect 675444 249092 675450 249144
rect 673454 248548 673460 248600
rect 673512 248588 673518 248600
rect 673638 248588 673644 248600
rect 673512 248560 673644 248588
rect 673512 248548 673518 248560
rect 673638 248548 673644 248560
rect 673696 248588 673702 248600
rect 675386 248588 675392 248600
rect 673696 248560 675392 248588
rect 673696 248548 673702 248560
rect 675386 248548 675392 248560
rect 675444 248548 675450 248600
rect 42334 246984 42340 247036
rect 42392 247024 42398 247036
rect 42702 247024 42708 247036
rect 42392 246996 42708 247024
rect 42392 246984 42398 246996
rect 42702 246984 42708 246996
rect 42760 246984 42766 247036
rect 41782 239028 41788 239080
rect 41840 239068 41846 239080
rect 42426 239068 42432 239080
rect 41840 239040 42432 239068
rect 41840 239028 41846 239040
rect 42426 239028 42432 239040
rect 42484 239068 42490 239080
rect 42610 239068 42616 239080
rect 42484 239040 42616 239068
rect 42484 239028 42490 239040
rect 42610 239028 42616 239040
rect 42668 239028 42674 239080
rect 673454 237668 673460 237720
rect 673512 237708 673518 237720
rect 673730 237708 673736 237720
rect 673512 237680 673736 237708
rect 673512 237668 673518 237680
rect 673730 237668 673736 237680
rect 673788 237708 673794 237720
rect 675386 237708 675392 237720
rect 673788 237680 675392 237708
rect 673788 237668 673794 237680
rect 675386 237668 675392 237680
rect 675444 237668 675450 237720
rect 42518 237396 42524 237448
rect 42576 237436 42582 237448
rect 42794 237436 42800 237448
rect 42576 237408 42800 237436
rect 42576 237396 42582 237408
rect 42794 237396 42800 237408
rect 42852 237396 42858 237448
rect 41782 227604 41788 227656
rect 41840 227644 41846 227656
rect 42426 227644 42432 227656
rect 41840 227616 42432 227644
rect 41840 227604 41846 227616
rect 42426 227604 42432 227616
rect 42484 227644 42490 227656
rect 42702 227644 42708 227656
rect 42484 227616 42708 227644
rect 42484 227604 42490 227616
rect 42702 227604 42708 227616
rect 42760 227604 42766 227656
rect 44174 218016 44180 218068
rect 44232 218056 44238 218068
rect 44358 218056 44364 218068
rect 44232 218028 44364 218056
rect 44232 218016 44238 218028
rect 44358 218016 44364 218028
rect 44416 218016 44422 218068
rect 673638 206932 673644 206984
rect 673696 206972 673702 206984
rect 675294 206972 675300 206984
rect 673696 206944 675300 206972
rect 673696 206932 673702 206944
rect 675294 206932 675300 206944
rect 675352 206932 675358 206984
rect 673546 202920 673552 202972
rect 673604 202960 673610 202972
rect 675386 202960 675392 202972
rect 673604 202932 675392 202960
rect 673604 202920 673610 202932
rect 675386 202920 675392 202932
rect 675444 202920 675450 202972
rect 42242 197344 42248 197396
rect 42300 197384 42306 197396
rect 42702 197384 42708 197396
rect 42300 197356 42708 197384
rect 42300 197344 42306 197356
rect 42702 197344 42708 197356
rect 42760 197344 42766 197396
rect 41782 195848 41788 195900
rect 41840 195888 41846 195900
rect 42610 195888 42616 195900
rect 41840 195860 42616 195888
rect 41840 195848 41846 195860
rect 42610 195848 42616 195860
rect 42668 195888 42674 195900
rect 44634 195888 44640 195900
rect 42668 195860 44640 195888
rect 42668 195848 42674 195860
rect 44634 195848 44640 195860
rect 44692 195848 44698 195900
rect 673454 191904 673460 191956
rect 673512 191944 673518 191956
rect 675386 191944 675392 191956
rect 673512 191916 675392 191944
rect 673512 191904 673518 191916
rect 675386 191904 675392 191916
rect 675444 191904 675450 191956
rect 41782 185444 41788 185496
rect 41840 185484 41846 185496
rect 42702 185484 42708 185496
rect 41840 185456 42708 185484
rect 41840 185444 41846 185456
rect 42702 185444 42708 185456
rect 42760 185444 42766 185496
rect 41782 184832 41788 184884
rect 41840 184872 41846 184884
rect 42242 184872 42248 184884
rect 41840 184844 42248 184872
rect 41840 184832 41846 184844
rect 42242 184832 42248 184844
rect 42300 184872 42306 184884
rect 42426 184872 42432 184884
rect 42300 184844 42432 184872
rect 42300 184832 42306 184844
rect 42426 184832 42432 184844
rect 42484 184832 42490 184884
rect 673730 184424 673736 184476
rect 673788 184464 673794 184476
rect 675202 184464 675208 184476
rect 673788 184436 675208 184464
rect 673788 184424 673794 184436
rect 675202 184424 675208 184436
rect 675260 184424 675266 184476
rect 42334 179392 42340 179444
rect 42392 179432 42398 179444
rect 42702 179432 42708 179444
rect 42392 179404 42708 179432
rect 42392 179392 42398 179404
rect 42702 179392 42708 179404
rect 42760 179392 42766 179444
rect 44174 179392 44180 179444
rect 44232 179432 44238 179444
rect 44358 179432 44364 179444
rect 44232 179404 44364 179432
rect 44232 179392 44238 179404
rect 44358 179392 44364 179404
rect 44416 179392 44422 179444
rect 673454 177964 673460 178016
rect 673512 178004 673518 178016
rect 673914 178004 673920 178016
rect 673512 177976 673920 178004
rect 673512 177964 673518 177976
rect 673914 177964 673920 177976
rect 673972 177964 673978 178016
rect 44450 173884 44456 173936
rect 44508 173924 44514 173936
rect 44726 173924 44732 173936
rect 44508 173896 44732 173924
rect 44508 173884 44514 173896
rect 44726 173884 44732 173896
rect 44784 173884 44790 173936
rect 673546 168308 673552 168360
rect 673604 168308 673610 168360
rect 673730 168308 673736 168360
rect 673788 168348 673794 168360
rect 675202 168348 675208 168360
rect 673788 168320 675208 168348
rect 673788 168308 673794 168320
rect 675202 168308 675208 168320
rect 675260 168308 675266 168360
rect 673564 168280 673592 168308
rect 675294 168280 675300 168292
rect 673564 168252 675300 168280
rect 675294 168240 675300 168252
rect 675352 168240 675358 168292
rect 44726 160188 44732 160200
rect 44652 160160 44732 160188
rect 44652 160064 44680 160160
rect 44726 160148 44732 160160
rect 44784 160148 44790 160200
rect 44634 160012 44640 160064
rect 44692 160012 44698 160064
rect 673454 157904 673460 157956
rect 673512 157944 673518 157956
rect 675386 157944 675392 157956
rect 673512 157916 675392 157944
rect 673512 157904 673518 157916
rect 675386 157904 675392 157916
rect 675444 157904 675450 157956
rect 673822 157292 673828 157344
rect 673880 157332 673886 157344
rect 675386 157332 675392 157344
rect 673880 157304 675392 157332
rect 673880 157292 673886 157304
rect 675386 157292 675392 157304
rect 675444 157292 675450 157344
rect 44634 154504 44640 154556
rect 44692 154544 44698 154556
rect 44818 154544 44824 154556
rect 44692 154516 44824 154544
rect 44692 154504 44698 154516
rect 44818 154504 44824 154516
rect 44876 154504 44882 154556
rect 673638 147840 673644 147892
rect 673696 147880 673702 147892
rect 673914 147880 673920 147892
rect 673696 147852 673920 147880
rect 673696 147840 673702 147852
rect 673914 147840 673920 147852
rect 673972 147880 673978 147892
rect 675386 147880 675392 147892
rect 673972 147852 675392 147880
rect 673972 147840 673978 147852
rect 675386 147840 675392 147852
rect 675444 147840 675450 147892
rect 44174 140768 44180 140820
rect 44232 140808 44238 140820
rect 44358 140808 44364 140820
rect 44232 140780 44364 140808
rect 44232 140768 44238 140780
rect 44358 140768 44364 140780
rect 44416 140768 44422 140820
rect 673454 129684 673460 129736
rect 673512 129724 673518 129736
rect 673730 129724 673736 129736
rect 673512 129696 673736 129724
rect 673512 129684 673518 129696
rect 673730 129684 673736 129696
rect 673788 129684 673794 129736
rect 673822 129684 673828 129736
rect 673880 129724 673886 129736
rect 675294 129724 675300 129736
rect 673880 129696 675300 129724
rect 673880 129684 673886 129696
rect 675294 129684 675300 129696
rect 675352 129684 675358 129736
rect 39850 125128 39856 125180
rect 39908 125168 39914 125180
rect 44174 125168 44180 125180
rect 39908 125140 44180 125168
rect 39908 125128 39914 125140
rect 44174 125128 44180 125140
rect 44232 125128 44238 125180
rect 39850 120164 39856 120216
rect 39908 120204 39914 120216
rect 44726 120204 44732 120216
rect 39908 120176 44732 120204
rect 39908 120164 39914 120176
rect 44726 120164 44732 120176
rect 44784 120164 44790 120216
rect 673454 112752 673460 112804
rect 673512 112792 673518 112804
rect 673730 112792 673736 112804
rect 673512 112764 673736 112792
rect 673512 112752 673518 112764
rect 673730 112752 673736 112764
rect 673788 112792 673794 112804
rect 675386 112792 675392 112804
rect 673788 112764 675392 112792
rect 673788 112752 673794 112764
rect 675386 112752 675392 112764
rect 675444 112752 675450 112804
rect 673546 112072 673552 112124
rect 673604 112112 673610 112124
rect 675386 112112 675392 112124
rect 673604 112084 675392 112112
rect 673604 112072 673610 112084
rect 675386 112072 675392 112084
rect 675444 112072 675450 112124
rect 673638 101668 673644 101720
rect 673696 101708 673702 101720
rect 675386 101708 675392 101720
rect 673696 101680 675392 101708
rect 673696 101668 673702 101680
rect 675386 101668 675392 101680
rect 675444 101668 675450 101720
rect 44266 96568 44272 96620
rect 44324 96608 44330 96620
rect 44450 96608 44456 96620
rect 44324 96580 44456 96608
rect 44324 96568 44330 96580
rect 44450 96568 44456 96580
rect 44508 96568 44514 96620
rect 44266 77256 44272 77308
rect 44324 77296 44330 77308
rect 44358 77296 44364 77308
rect 44324 77268 44364 77296
rect 44324 77256 44330 77268
rect 44358 77256 44364 77268
rect 44416 77256 44422 77308
rect 39666 74876 39672 74928
rect 39724 74916 39730 74928
rect 39850 74916 39856 74928
rect 39724 74888 39856 74916
rect 39724 74876 39730 74888
rect 39850 74876 39856 74888
rect 39908 74876 39914 74928
rect 44174 71748 44180 71800
rect 44232 71788 44238 71800
rect 44358 71788 44364 71800
rect 44232 71760 44364 71788
rect 44232 71748 44238 71760
rect 44358 71748 44364 71760
rect 44416 71748 44422 71800
rect 39574 67940 39580 67992
rect 39632 67980 39638 67992
rect 41414 67980 41420 67992
rect 39632 67952 41420 67980
rect 39632 67940 39638 67952
rect 41414 67940 41420 67952
rect 41472 67940 41478 67992
rect 41414 64472 41420 64524
rect 41472 64512 41478 64524
rect 42702 64512 42708 64524
rect 41472 64484 42708 64512
rect 41472 64472 41478 64484
rect 42702 64472 42708 64484
rect 42760 64472 42766 64524
rect 39666 52368 39672 52420
rect 39724 52408 39730 52420
rect 39850 52408 39856 52420
rect 39724 52380 39856 52408
rect 39724 52368 39730 52380
rect 39850 52368 39856 52380
rect 39908 52368 39914 52420
rect 42242 45840 42248 45892
rect 42300 45880 42306 45892
rect 145098 45880 145104 45892
rect 42300 45852 145104 45880
rect 42300 45840 42306 45852
rect 145098 45840 145104 45852
rect 145156 45840 145162 45892
rect 42702 45772 42708 45824
rect 42760 45812 42766 45824
rect 140958 45812 140964 45824
rect 42760 45784 140964 45812
rect 42760 45772 42766 45784
rect 140958 45772 140964 45784
rect 141016 45772 141022 45824
rect 578786 45704 578792 45756
rect 578844 45744 578850 45756
rect 673546 45744 673552 45756
rect 578844 45716 673552 45744
rect 578844 45704 578850 45716
rect 673546 45704 673552 45716
rect 673604 45704 673610 45756
rect 44174 45636 44180 45688
rect 44232 45676 44238 45688
rect 145834 45676 145840 45688
rect 44232 45648 145840 45676
rect 44232 45636 44238 45648
rect 145834 45636 145840 45648
rect 145892 45636 145898 45688
rect 528646 45636 528652 45688
rect 528704 45676 528710 45688
rect 673086 45676 673092 45688
rect 528704 45648 673092 45676
rect 528704 45636 528710 45648
rect 673086 45636 673092 45648
rect 673144 45636 673150 45688
rect 39850 45568 39856 45620
rect 39908 45608 39914 45620
rect 189258 45608 189264 45620
rect 39908 45580 189264 45608
rect 39908 45568 39914 45580
rect 189258 45568 189264 45580
rect 189316 45568 189322 45620
rect 529842 45568 529848 45620
rect 529900 45608 529906 45620
rect 673454 45608 673460 45620
rect 529900 45580 673460 45608
rect 529900 45568 529906 45580
rect 673454 45568 673460 45580
rect 673512 45568 673518 45620
rect 44910 45500 44916 45552
rect 44968 45540 44974 45552
rect 195974 45540 195980 45552
rect 44968 45512 195980 45540
rect 44968 45500 44974 45512
rect 195974 45500 195980 45512
rect 196032 45500 196038 45552
rect 516318 45500 516324 45552
rect 516376 45540 516382 45552
rect 673638 45540 673644 45552
rect 516376 45512 673644 45540
rect 516376 45500 516382 45512
rect 673638 45500 673644 45512
rect 673696 45500 673702 45552
rect 289814 44820 289820 44872
rect 289872 44860 289878 44872
rect 313182 44860 313188 44872
rect 289872 44832 313188 44860
rect 289872 44820 289878 44832
rect 313182 44820 313188 44832
rect 313240 44820 313246 44872
rect 458174 44820 458180 44872
rect 458232 44860 458238 44872
rect 458232 44832 531268 44860
rect 458232 44820 458238 44832
rect 250990 44752 250996 44804
rect 251048 44792 251054 44804
rect 252094 44792 252100 44804
rect 251048 44764 252100 44792
rect 251048 44752 251054 44764
rect 252094 44752 252100 44764
rect 252152 44792 252158 44804
rect 276014 44792 276020 44804
rect 252152 44764 276020 44792
rect 252152 44752 252158 44764
rect 276014 44752 276020 44764
rect 276072 44752 276078 44804
rect 380894 44752 380900 44804
rect 380952 44792 380958 44804
rect 400122 44792 400128 44804
rect 380952 44764 400128 44792
rect 380952 44752 380958 44764
rect 400122 44752 400128 44764
rect 400180 44752 400186 44804
rect 406746 44752 406752 44804
rect 406804 44792 406810 44804
rect 461486 44792 461492 44804
rect 406804 44764 461492 44792
rect 406804 44752 406810 44764
rect 461486 44752 461492 44764
rect 461544 44752 461550 44804
rect 231854 44724 231860 44736
rect 198752 44696 231860 44724
rect 193122 44616 193128 44668
rect 193180 44656 193186 44668
rect 198752 44656 198780 44696
rect 231854 44684 231860 44696
rect 231912 44684 231918 44736
rect 308214 44684 308220 44736
rect 308272 44724 308278 44736
rect 358722 44724 358728 44736
rect 308272 44696 358728 44724
rect 308272 44684 308278 44696
rect 358722 44684 358728 44696
rect 358780 44684 358786 44736
rect 362402 44684 362408 44736
rect 362460 44724 362466 44736
rect 362460 44696 367048 44724
rect 362460 44684 362466 44696
rect 193180 44628 198780 44656
rect 193180 44616 193186 44628
rect 247678 44616 247684 44668
rect 247736 44656 247742 44668
rect 307570 44656 307576 44668
rect 247736 44628 307576 44656
rect 247736 44616 247742 44628
rect 307570 44616 307576 44628
rect 307628 44616 307634 44668
rect 308306 44616 308312 44668
rect 308364 44656 308370 44668
rect 309134 44656 309140 44668
rect 308364 44628 309140 44656
rect 308364 44616 308370 44628
rect 309134 44616 309140 44628
rect 309192 44616 309198 44668
rect 328362 44616 328368 44668
rect 328420 44656 328426 44668
rect 347774 44656 347780 44668
rect 328420 44628 347780 44656
rect 328420 44616 328426 44628
rect 347774 44616 347780 44628
rect 347832 44616 347838 44668
rect 367020 44656 367048 44696
rect 488534 44684 488540 44736
rect 488592 44724 488598 44736
rect 499574 44724 499580 44736
rect 488592 44696 499580 44724
rect 488592 44684 488598 44696
rect 499574 44684 499580 44696
rect 499632 44684 499638 44736
rect 526806 44724 526812 44736
rect 521672 44696 526812 44724
rect 386414 44656 386420 44668
rect 367020 44628 386420 44656
rect 386414 44616 386420 44628
rect 386472 44616 386478 44668
rect 405642 44616 405648 44668
rect 405700 44656 405706 44668
rect 417234 44656 417240 44668
rect 405700 44628 417240 44656
rect 405700 44616 405706 44628
rect 417234 44616 417240 44628
rect 417292 44656 417298 44668
rect 425054 44656 425060 44668
rect 417292 44628 425060 44656
rect 417292 44616 417298 44628
rect 425054 44616 425060 44628
rect 425112 44616 425118 44668
rect 444282 44616 444288 44668
rect 444340 44656 444346 44668
rect 471974 44656 471980 44668
rect 444340 44628 471980 44656
rect 444340 44616 444346 44628
rect 471974 44616 471980 44628
rect 472032 44616 472038 44668
rect 472066 44616 472072 44668
rect 472124 44656 472130 44668
rect 472342 44656 472348 44668
rect 472124 44628 472348 44656
rect 472124 44616 472130 44628
rect 472342 44616 472348 44628
rect 472400 44656 472406 44668
rect 488442 44656 488448 44668
rect 472400 44628 488448 44656
rect 472400 44616 472406 44628
rect 488442 44616 488448 44628
rect 488500 44616 488506 44668
rect 518802 44616 518808 44668
rect 518860 44656 518866 44668
rect 521672 44656 521700 44696
rect 526806 44684 526812 44696
rect 526864 44684 526870 44736
rect 531240 44724 531268 44832
rect 546586 44820 546592 44872
rect 546644 44860 546650 44872
rect 560294 44860 560300 44872
rect 546644 44832 560300 44860
rect 546644 44820 546650 44832
rect 560294 44820 560300 44832
rect 560352 44820 560358 44872
rect 546402 44724 546408 44736
rect 531240 44696 546408 44724
rect 546402 44684 546408 44696
rect 546460 44684 546466 44736
rect 518860 44628 521700 44656
rect 518860 44616 518866 44628
rect 173894 44588 173900 44600
rect 160112 44560 173900 44588
rect 140958 44480 140964 44532
rect 141016 44520 141022 44532
rect 160112 44520 160140 44560
rect 173894 44548 173900 44560
rect 173952 44548 173958 44600
rect 289814 44548 289820 44600
rect 289872 44548 289878 44600
rect 309410 44548 309416 44600
rect 309468 44588 309474 44600
rect 309468 44560 310836 44588
rect 309468 44548 309474 44560
rect 141016 44492 160140 44520
rect 141016 44480 141022 44492
rect 199654 44480 199660 44532
rect 199712 44520 199718 44532
rect 212534 44520 212540 44532
rect 199712 44492 212540 44520
rect 199712 44480 199718 44492
rect 212534 44480 212540 44492
rect 212592 44480 212598 44532
rect 218054 44480 218060 44532
rect 218112 44520 218118 44532
rect 218112 44492 221320 44520
rect 218112 44480 218118 44492
rect 195974 44412 195980 44464
rect 196032 44452 196038 44464
rect 200758 44452 200764 44464
rect 196032 44424 200764 44452
rect 196032 44412 196038 44424
rect 200758 44412 200764 44424
rect 200816 44412 200822 44464
rect 200850 44412 200856 44464
rect 200908 44452 200914 44464
rect 217870 44452 217876 44464
rect 200908 44424 217876 44452
rect 200908 44412 200914 44424
rect 217870 44412 217876 44424
rect 217928 44412 217934 44464
rect 221292 44452 221320 44492
rect 276014 44480 276020 44532
rect 276072 44520 276078 44532
rect 289832 44520 289860 44548
rect 276072 44492 289860 44520
rect 276072 44480 276078 44492
rect 299566 44480 299572 44532
rect 299624 44520 299630 44532
rect 305730 44520 305736 44532
rect 299624 44492 305736 44520
rect 299624 44480 299630 44492
rect 305730 44480 305736 44492
rect 305788 44520 305794 44532
rect 310808 44520 310836 44560
rect 313182 44548 313188 44600
rect 313240 44588 313246 44600
rect 380894 44588 380900 44600
rect 313240 44560 380900 44588
rect 313240 44548 313246 44560
rect 380894 44548 380900 44560
rect 380952 44548 380958 44600
rect 400122 44548 400128 44600
rect 400180 44588 400186 44600
rect 419534 44588 419540 44600
rect 400180 44560 419540 44588
rect 400180 44548 400186 44560
rect 419534 44548 419540 44560
rect 419592 44548 419598 44600
rect 438762 44548 438768 44600
rect 438820 44588 438826 44600
rect 458174 44588 458180 44600
rect 438820 44560 458180 44588
rect 438820 44548 438826 44560
rect 458174 44548 458180 44560
rect 458232 44548 458238 44600
rect 352558 44520 352564 44532
rect 305788 44492 310744 44520
rect 310808 44492 352564 44520
rect 305788 44480 305794 44492
rect 242894 44452 242900 44464
rect 221292 44424 242900 44452
rect 242894 44412 242900 44424
rect 242952 44452 242958 44464
rect 297726 44452 297732 44464
rect 242952 44424 297732 44452
rect 242952 44412 242958 44424
rect 297726 44412 297732 44424
rect 297784 44452 297790 44464
rect 300762 44452 300768 44464
rect 297784 44424 300768 44452
rect 297784 44412 297790 44424
rect 300762 44412 300768 44424
rect 300820 44452 300826 44464
rect 306374 44452 306380 44464
rect 300820 44424 306380 44452
rect 300820 44412 300826 44424
rect 306374 44412 306380 44424
rect 306432 44412 306438 44464
rect 310716 44452 310744 44492
rect 352558 44480 352564 44492
rect 352616 44520 352622 44532
rect 355594 44520 355600 44532
rect 352616 44492 355600 44520
rect 352616 44480 352622 44492
rect 355594 44480 355600 44492
rect 355652 44520 355658 44532
rect 359918 44520 359924 44532
rect 355652 44492 359924 44520
rect 355652 44480 355658 44492
rect 359918 44480 359924 44492
rect 359976 44480 359982 44532
rect 364150 44480 364156 44532
rect 364208 44520 364214 44532
rect 407390 44520 407396 44532
rect 364208 44492 407396 44520
rect 364208 44480 364214 44492
rect 407390 44480 407396 44492
rect 407448 44520 407454 44532
rect 410426 44520 410432 44532
rect 407448 44492 410432 44520
rect 407448 44480 407454 44492
rect 410426 44480 410432 44492
rect 410484 44480 410490 44532
rect 419074 44480 419080 44532
rect 419132 44520 419138 44532
rect 462130 44520 462136 44532
rect 419132 44492 462136 44520
rect 419132 44480 419138 44492
rect 462130 44480 462136 44492
rect 462188 44520 462194 44532
rect 465166 44520 465172 44532
rect 462188 44492 465172 44520
rect 462188 44480 462194 44492
rect 465166 44480 465172 44492
rect 465224 44480 465230 44532
rect 473814 44480 473820 44532
rect 473872 44520 473878 44532
rect 516962 44520 516968 44532
rect 473872 44492 516968 44520
rect 473872 44480 473878 44492
rect 516962 44480 516968 44492
rect 517020 44480 517026 44532
rect 351914 44452 351920 44464
rect 310716 44424 351920 44452
rect 351914 44412 351920 44424
rect 351972 44452 351978 44464
rect 354398 44452 354404 44464
rect 351972 44424 354404 44452
rect 351972 44412 351978 44424
rect 354398 44412 354404 44424
rect 354456 44452 354462 44464
rect 360562 44452 360568 44464
rect 354456 44424 360568 44452
rect 354456 44412 354462 44424
rect 360562 44412 360568 44424
rect 360620 44412 360626 44464
rect 363046 44412 363052 44464
rect 363104 44452 363110 44464
rect 413554 44452 413560 44464
rect 363104 44424 413560 44452
rect 363104 44412 363110 44424
rect 413554 44412 413560 44424
rect 413612 44452 413618 44464
rect 417878 44452 417884 44464
rect 413612 44424 417884 44452
rect 413612 44412 413618 44424
rect 417878 44412 417884 44424
rect 417936 44452 417942 44464
rect 468294 44452 468300 44464
rect 417936 44424 468300 44452
rect 417936 44412 417942 44424
rect 468294 44412 468300 44424
rect 468352 44452 468358 44464
rect 472618 44452 472624 44464
rect 468352 44424 472624 44452
rect 468352 44412 468358 44424
rect 472618 44412 472624 44424
rect 472676 44452 472682 44464
rect 523126 44452 523132 44464
rect 472676 44424 523132 44452
rect 472676 44412 472682 44424
rect 523126 44412 523132 44424
rect 523184 44412 523190 44464
rect 199010 44344 199016 44396
rect 199068 44384 199074 44396
rect 217962 44384 217968 44396
rect 199068 44356 217968 44384
rect 199068 44344 199074 44356
rect 217962 44344 217968 44356
rect 218020 44344 218026 44396
rect 218146 44344 218152 44396
rect 218204 44384 218210 44396
rect 247402 44384 247408 44396
rect 218204 44356 247408 44384
rect 218204 44344 218210 44356
rect 247402 44344 247408 44356
rect 247460 44384 247466 44396
rect 247678 44384 247684 44396
rect 247460 44356 247684 44384
rect 247460 44344 247466 44356
rect 247678 44344 247684 44356
rect 247736 44344 247742 44396
rect 289814 44344 289820 44396
rect 289872 44344 289878 44396
rect 359366 44384 359372 44396
rect 304552 44356 359372 44384
rect 248322 44276 248328 44328
rect 248380 44316 248386 44328
rect 267734 44316 267740 44328
rect 248380 44288 267740 44316
rect 248380 44276 248386 44288
rect 267734 44276 267740 44288
rect 267792 44276 267798 44328
rect 286962 44276 286968 44328
rect 287020 44316 287026 44328
rect 289832 44316 289860 44344
rect 287020 44288 289860 44316
rect 287020 44276 287026 44288
rect 304552 44260 304580 44356
rect 359366 44344 359372 44356
rect 359424 44384 359430 44396
rect 414198 44384 414204 44396
rect 359424 44356 414204 44384
rect 359424 44344 359430 44356
rect 414198 44344 414204 44356
rect 414256 44384 414262 44396
rect 468938 44384 468944 44396
rect 414256 44356 468944 44384
rect 414256 44344 414262 44356
rect 468938 44344 468944 44356
rect 468996 44384 469002 44396
rect 523770 44384 523776 44396
rect 468996 44356 523776 44384
rect 468996 44344 469002 44356
rect 523770 44344 523776 44356
rect 523828 44344 523834 44396
rect 360562 44276 360568 44328
rect 360620 44316 360626 44328
rect 406746 44316 406752 44328
rect 360620 44288 406752 44316
rect 360620 44276 360626 44288
rect 406746 44276 406752 44288
rect 406804 44276 406810 44328
rect 411070 44276 411076 44328
rect 411128 44316 411134 44328
rect 411128 44288 413048 44316
rect 411128 44276 411134 44288
rect 145098 44208 145104 44260
rect 145156 44248 145162 44260
rect 195330 44248 195336 44260
rect 145156 44220 195336 44248
rect 145156 44208 145162 44220
rect 195330 44208 195336 44220
rect 195388 44248 195394 44260
rect 199654 44248 199660 44260
rect 195388 44220 199660 44248
rect 195388 44208 195394 44220
rect 199654 44208 199660 44220
rect 199712 44208 199718 44260
rect 200758 44208 200764 44260
rect 200816 44248 200822 44260
rect 304534 44248 304540 44260
rect 200816 44220 304540 44248
rect 200816 44208 200822 44220
rect 304534 44208 304540 44220
rect 304592 44208 304598 44260
rect 307570 44208 307576 44260
rect 307628 44248 307634 44260
rect 308306 44248 308312 44260
rect 307628 44220 308312 44248
rect 307628 44208 307634 44220
rect 308306 44208 308312 44220
rect 308364 44208 308370 44260
rect 186682 44140 186688 44192
rect 186740 44180 186746 44192
rect 194686 44180 194692 44192
rect 186740 44152 194692 44180
rect 186740 44140 186746 44152
rect 194686 44140 194692 44152
rect 194744 44140 194750 44192
rect 295242 44140 295248 44192
rect 295300 44180 295306 44192
rect 303246 44180 303252 44192
rect 295300 44152 303252 44180
rect 295300 44140 295306 44152
rect 303246 44140 303252 44152
rect 303304 44140 303310 44192
rect 306374 44140 306380 44192
rect 306432 44180 306438 44192
rect 309410 44180 309416 44192
rect 306432 44152 309416 44180
rect 306432 44140 306438 44152
rect 309410 44140 309416 44152
rect 309468 44140 309474 44192
rect 350074 44140 350080 44192
rect 350132 44180 350138 44192
rect 358078 44180 358084 44192
rect 350132 44152 358084 44180
rect 350132 44140 350138 44152
rect 358078 44140 358084 44152
rect 358136 44140 358142 44192
rect 404906 44140 404912 44192
rect 404964 44180 404970 44192
rect 412910 44180 412916 44192
rect 404964 44152 412916 44180
rect 404964 44140 404970 44152
rect 412910 44140 412916 44152
rect 412968 44140 412974 44192
rect 413020 44180 413048 44288
rect 419534 44276 419540 44328
rect 419592 44316 419598 44328
rect 438762 44316 438768 44328
rect 419592 44288 438768 44316
rect 419592 44276 419598 44288
rect 438762 44276 438768 44288
rect 438820 44276 438826 44328
rect 461486 44276 461492 44328
rect 461544 44316 461550 44328
rect 516318 44316 516324 44328
rect 461544 44288 516324 44316
rect 461544 44276 461550 44288
rect 516318 44276 516324 44288
rect 516376 44276 516382 44328
rect 465810 44208 465816 44260
rect 465868 44248 465874 44260
rect 474458 44248 474464 44260
rect 465868 44220 474464 44248
rect 465868 44208 465874 44220
rect 474458 44208 474464 44220
rect 474516 44208 474522 44260
rect 514478 44208 514484 44260
rect 514536 44248 514542 44260
rect 522482 44248 522488 44260
rect 514536 44220 522488 44248
rect 514536 44208 514542 44220
rect 522482 44208 522488 44220
rect 522540 44208 522546 44260
rect 523126 44208 523132 44260
rect 523184 44248 523190 44260
rect 527450 44248 527456 44260
rect 523184 44220 527456 44248
rect 523184 44208 523190 44220
rect 527450 44208 527456 44220
rect 527508 44248 527514 44260
rect 529842 44248 529848 44260
rect 527508 44220 529848 44248
rect 527508 44208 527514 44220
rect 529842 44208 529848 44220
rect 529900 44208 529906 44260
rect 419718 44180 419724 44192
rect 413020 44152 419724 44180
rect 419718 44140 419724 44152
rect 419776 44140 419782 44192
rect 459646 44140 459652 44192
rect 459704 44180 459710 44192
rect 467650 44180 467656 44192
rect 459704 44152 467656 44180
rect 459704 44140 459710 44152
rect 467650 44140 467656 44152
rect 467708 44140 467714 44192
rect 518802 44140 518808 44192
rect 518860 44180 518866 44192
rect 524966 44180 524972 44192
rect 518860 44152 524972 44180
rect 518860 44140 518866 44152
rect 524966 44140 524972 44152
rect 525024 44140 525030 44192
rect 525610 44140 525616 44192
rect 525668 44180 525674 44192
rect 528646 44180 528652 44192
rect 525668 44152 528652 44180
rect 525668 44140 525674 44152
rect 528646 44140 528652 44152
rect 528704 44140 528710 44192
rect 39758 44072 39764 44124
rect 39816 44112 39822 44124
rect 78950 44112 78956 44124
rect 39816 44084 78956 44112
rect 39816 44072 39822 44084
rect 78950 44072 78956 44084
rect 79008 44072 79014 44124
rect 347774 43664 347780 43716
rect 347832 43704 347838 43716
rect 362402 43704 362408 43716
rect 347832 43676 362408 43704
rect 347832 43664 347838 43676
rect 362402 43664 362408 43676
rect 362460 43664 362466 43716
rect 303890 42236 303896 42288
rect 303948 42276 303954 42288
rect 308214 42276 308220 42288
rect 303948 42248 308220 42276
rect 303948 42236 303954 42248
rect 308214 42236 308220 42248
rect 308272 42236 308278 42288
rect 189258 41896 189264 41948
rect 189316 41936 189322 41948
rect 191098 41936 191104 41948
rect 189316 41908 191104 41936
rect 189316 41896 189322 41908
rect 191098 41896 191104 41908
rect 191156 41936 191162 41948
rect 192294 41936 192300 41948
rect 191156 41908 192300 41936
rect 191156 41896 191162 41908
rect 192294 41896 192300 41908
rect 192352 41936 192358 41948
rect 193582 41936 193588 41948
rect 192352 41908 193588 41936
rect 192352 41896 192358 41908
rect 193582 41896 193588 41908
rect 193640 41936 193646 41948
rect 196434 41936 196440 41948
rect 193640 41908 196440 41936
rect 193640 41896 193646 41908
rect 196434 41896 196440 41908
rect 196492 41896 196498 41948
rect 198458 41896 198464 41948
rect 198516 41936 198522 41948
rect 200114 41936 200120 41948
rect 198516 41908 200120 41936
rect 198516 41896 198522 41908
rect 200114 41896 200120 41908
rect 200172 41896 200178 41948
rect 363506 41936 363512 41948
rect 361132 41908 363512 41936
rect 361132 41880 361160 41908
rect 363506 41896 363512 41908
rect 363564 41896 363570 41948
rect 188614 41868 188620 41880
rect 188540 41840 188620 41868
rect 135346 41692 135352 41744
rect 135404 41732 135410 41744
rect 154482 41732 154488 41744
rect 135404 41704 154488 41732
rect 135404 41692 135410 41704
rect 154482 41692 154488 41704
rect 154540 41692 154546 41744
rect 168282 41732 168288 41744
rect 160020 41704 168288 41732
rect 91278 41556 91284 41608
rect 91336 41596 91342 41608
rect 91336 41568 96660 41596
rect 91336 41556 91342 41568
rect 96632 41528 96660 41568
rect 102134 41556 102140 41608
rect 102192 41596 102198 41608
rect 102192 41568 115888 41596
rect 102192 41556 102198 41568
rect 102042 41528 102048 41540
rect 96632 41500 102048 41528
rect 102042 41488 102048 41500
rect 102100 41488 102106 41540
rect 115860 41528 115888 41568
rect 154482 41556 154488 41608
rect 154540 41596 154546 41608
rect 160020 41596 160048 41704
rect 168282 41692 168288 41704
rect 168340 41692 168346 41744
rect 188540 41732 188568 41840
rect 188614 41828 188620 41840
rect 188672 41868 188678 41880
rect 192938 41868 192944 41880
rect 188672 41840 192944 41868
rect 188672 41828 188678 41840
rect 192938 41828 192944 41840
rect 192996 41868 193002 41880
rect 201586 41868 201592 41880
rect 192996 41840 201592 41868
rect 192996 41828 193002 41840
rect 201586 41828 201592 41840
rect 201644 41868 201650 41880
rect 202506 41868 202512 41880
rect 201644 41840 202512 41868
rect 201644 41828 201650 41840
rect 202506 41828 202512 41840
rect 202564 41828 202570 41880
rect 299474 41868 299480 41880
rect 296916 41840 299480 41868
rect 296916 41812 296944 41840
rect 299474 41828 299480 41840
rect 299532 41828 299538 41880
rect 360010 41828 360016 41880
rect 360068 41868 360074 41880
rect 361114 41868 361120 41880
rect 360068 41840 361120 41868
rect 360068 41828 360074 41840
rect 361114 41828 361120 41840
rect 361172 41828 361178 41880
rect 409322 41828 409328 41880
rect 409380 41868 409386 41880
rect 412358 41868 412364 41880
rect 409380 41840 412364 41868
rect 409380 41828 409386 41840
rect 412358 41828 412364 41840
rect 412416 41868 412422 41880
rect 415210 41868 415216 41880
rect 412416 41840 415216 41868
rect 412416 41828 412422 41840
rect 415210 41828 415216 41840
rect 415268 41828 415274 41880
rect 465350 41828 465356 41880
rect 465408 41868 465414 41880
rect 466362 41868 466368 41880
rect 465408 41840 466368 41868
rect 465408 41828 465414 41840
rect 466362 41828 466368 41840
rect 466420 41868 466426 41880
rect 469398 41868 469404 41880
rect 466420 41840 469404 41868
rect 466420 41828 466426 41840
rect 469398 41828 469404 41840
rect 469456 41868 469462 41880
rect 470686 41868 470692 41880
rect 469456 41840 470692 41868
rect 469456 41828 469462 41840
rect 470686 41828 470692 41840
rect 470744 41868 470750 41880
rect 473078 41868 473084 41880
rect 470744 41840 473084 41868
rect 470744 41828 470750 41840
rect 473078 41828 473084 41840
rect 473136 41828 473142 41880
rect 517054 41828 517060 41880
rect 517112 41868 517118 41880
rect 520090 41868 520096 41880
rect 517112 41840 520096 41868
rect 517112 41828 517118 41840
rect 520090 41828 520096 41840
rect 520148 41868 520154 41880
rect 521378 41868 521384 41880
rect 520148 41840 521384 41868
rect 520148 41828 520154 41840
rect 521378 41828 521384 41840
rect 521436 41868 521442 41880
rect 524414 41868 524420 41880
rect 521436 41840 524420 41868
rect 521436 41828 521442 41840
rect 524414 41828 524420 41840
rect 524472 41868 524478 41880
rect 525518 41868 525524 41880
rect 524472 41840 525524 41868
rect 524472 41828 524478 41840
rect 525518 41828 525524 41840
rect 525576 41828 525582 41880
rect 525628 41840 527036 41868
rect 198918 41760 198924 41812
rect 198976 41760 198982 41812
rect 296898 41760 296904 41812
rect 296956 41760 296962 41812
rect 305270 41760 305276 41812
rect 305328 41800 305334 41812
rect 306282 41800 306288 41812
rect 305328 41772 306288 41800
rect 305328 41760 305334 41772
rect 306282 41760 306288 41772
rect 306340 41760 306346 41812
rect 358814 41760 358820 41812
rect 358872 41800 358878 41812
rect 362954 41800 362960 41812
rect 358872 41772 362960 41800
rect 358872 41760 358878 41772
rect 362954 41760 362960 41772
rect 363012 41760 363018 41812
rect 410518 41760 410524 41812
rect 410576 41800 410582 41812
rect 411530 41800 411536 41812
rect 410576 41772 411536 41800
rect 410576 41760 410582 41772
rect 411530 41760 411536 41772
rect 411588 41800 411594 41812
rect 414566 41800 414572 41812
rect 411588 41772 414572 41800
rect 411588 41760 411594 41772
rect 414566 41760 414572 41772
rect 414624 41800 414630 41812
rect 415854 41800 415860 41812
rect 414624 41772 415860 41800
rect 414624 41760 414630 41772
rect 415854 41760 415860 41772
rect 415912 41800 415918 41812
rect 418246 41800 418252 41812
rect 415912 41772 418252 41800
rect 415912 41760 415918 41772
rect 418246 41760 418252 41772
rect 418304 41760 418310 41812
rect 464154 41760 464160 41812
rect 464212 41800 464218 41812
rect 467190 41800 467196 41812
rect 464212 41772 467196 41800
rect 464212 41760 464218 41772
rect 467190 41760 467196 41772
rect 467248 41800 467254 41812
rect 470042 41800 470048 41812
rect 467248 41772 470048 41800
rect 467248 41760 467254 41772
rect 470042 41760 470048 41772
rect 470100 41760 470106 41812
rect 523862 41760 523868 41812
rect 523920 41800 523926 41812
rect 525628 41800 525656 41840
rect 523920 41772 525656 41800
rect 523920 41760 523926 41772
rect 526898 41760 526904 41812
rect 526956 41760 526962 41812
rect 198936 41732 198964 41760
rect 296916 41732 296944 41760
rect 171980 41704 188568 41732
rect 197832 41704 198964 41732
rect 296824 41704 296944 41732
rect 171980 41596 172008 41704
rect 154540 41568 160048 41596
rect 168392 41568 172008 41596
rect 154540 41556 154546 41568
rect 121362 41528 121368 41540
rect 115860 41500 121368 41528
rect 121362 41488 121368 41500
rect 121420 41488 121426 41540
rect 121454 41488 121460 41540
rect 121512 41528 121518 41540
rect 168392 41528 168420 41568
rect 121512 41500 125548 41528
rect 121512 41488 121518 41500
rect 125520 41460 125548 41500
rect 168208 41500 168420 41528
rect 135254 41460 135260 41472
rect 125520 41432 135260 41460
rect 135254 41420 135260 41432
rect 135312 41420 135318 41472
rect 149974 41420 149980 41472
rect 150032 41460 150038 41472
rect 168208 41460 168236 41500
rect 197832 41460 197860 41704
rect 253934 41556 253940 41608
rect 253992 41596 253998 41608
rect 253992 41568 256740 41596
rect 253992 41556 253998 41568
rect 256712 41528 256740 41568
rect 256712 41500 275968 41528
rect 150032 41432 168236 41460
rect 168484 41432 197860 41460
rect 150032 41420 150038 41432
rect 168282 41352 168288 41404
rect 168340 41392 168346 41404
rect 168484 41392 168512 41432
rect 202506 41420 202512 41472
rect 202564 41460 202570 41472
rect 240134 41460 240140 41472
rect 202564 41432 240140 41460
rect 202564 41420 202570 41432
rect 240134 41420 240140 41432
rect 240192 41420 240198 41472
rect 275940 41460 275968 41500
rect 296824 41460 296852 41704
rect 275940 41432 296852 41460
rect 526916 41460 526944 41760
rect 527008 41528 527036 41840
rect 569126 41528 569132 41540
rect 527008 41500 569132 41528
rect 569126 41488 569132 41500
rect 569184 41488 569190 41540
rect 629294 41460 629300 41472
rect 526916 41432 629300 41460
rect 629294 41420 629300 41432
rect 629352 41420 629358 41472
rect 168340 41364 168512 41392
rect 168340 41352 168346 41364
rect 78950 40196 78956 40248
rect 79008 40236 79014 40248
rect 86494 40236 86500 40248
rect 79008 40208 86500 40236
rect 79008 40196 79014 40208
rect 86494 40196 86500 40208
rect 86552 40236 86558 40248
rect 91278 40236 91284 40248
rect 86552 40208 91284 40236
rect 86552 40196 86558 40208
rect 91278 40196 91284 40208
rect 91336 40196 91342 40248
rect 133092 40196 133098 40248
rect 133150 40236 133156 40248
rect 143810 40236 143816 40248
rect 133150 40208 143816 40236
rect 133150 40196 133156 40208
rect 143810 40196 143816 40208
rect 143868 40196 143874 40248
rect 140990 40060 140996 40112
rect 141048 40100 141054 40112
rect 143066 40100 143072 40112
rect 141048 40072 143072 40100
rect 141048 40060 141054 40072
rect 142586 39950 142614 40072
rect 143066 40060 143072 40072
rect 143124 40100 143130 40112
rect 143350 40100 143356 40112
rect 143124 40072 143356 40100
rect 143124 40060 143130 40072
rect 143350 40060 143356 40072
rect 143408 40100 143414 40112
rect 143408 40072 144684 40100
rect 143408 40060 143414 40072
rect 144656 39984 144684 40072
<< via1 >>
rect 84016 995596 84068 995648
rect 91744 995596 91796 995648
rect 531964 995596 532016 995648
rect 539692 995596 539744 995648
rect 135352 995460 135404 995512
rect 143172 995460 143224 995512
rect 633808 995460 633860 995512
rect 641536 995460 641588 995512
rect 238208 995392 238260 995444
rect 245936 995392 245988 995444
rect 289636 995256 289688 995308
rect 297640 995256 297692 995308
rect 391480 995256 391532 995308
rect 399484 995256 399536 995308
rect 480444 995256 480496 995308
rect 488448 995256 488500 995308
rect 589556 992264 589608 992316
rect 674748 992264 674800 992316
rect 44088 992196 44140 992248
rect 329564 992196 329616 992248
rect 585048 992196 585100 992248
rect 675208 992196 675260 992248
rect 78864 990768 78916 990820
rect 130292 990768 130344 990820
rect 132408 990768 132460 990820
rect 181720 990768 181772 990820
rect 233056 990768 233108 990820
rect 79508 990700 79560 990752
rect 130936 990700 130988 990752
rect 182364 990700 182416 990752
rect 187700 990700 187752 990752
rect 206928 990700 206980 990752
rect 226340 990700 226392 990752
rect 88340 990632 88392 990684
rect 89996 990632 90048 990684
rect 141424 990632 141476 990684
rect 192852 990632 192904 990684
rect 132408 990564 132460 990616
rect 181720 990564 181772 990616
rect 186688 990564 186740 990616
rect 194692 990564 194744 990616
rect 233608 990564 233660 990616
rect 256608 990700 256660 990752
rect 285312 990768 285364 990820
rect 295708 990768 295760 990820
rect 246948 990632 247000 990684
rect 295524 990700 295576 990752
rect 314660 990700 314712 990752
rect 324228 990768 324280 990820
rect 333888 990768 333940 990820
rect 343640 990768 343692 990820
rect 353300 990768 353352 990820
rect 324320 990700 324372 990752
rect 333980 990700 334032 990752
rect 357808 990700 357860 990752
rect 372344 990700 372396 990752
rect 387156 990768 387208 990820
rect 475384 990768 475436 990820
rect 475476 990768 475528 990820
rect 526904 990768 526956 990820
rect 545948 990768 546000 990820
rect 546408 990768 546460 990820
rect 628656 990768 628708 990820
rect 353300 990632 353352 990684
rect 233056 990496 233108 990548
rect 244372 990564 244424 990616
rect 256700 990564 256752 990616
rect 256608 990496 256660 990548
rect 284576 990564 284628 990616
rect 284668 990564 284720 990616
rect 289820 990564 289872 990616
rect 309048 990564 309100 990616
rect 315948 990564 316000 990616
rect 187700 990428 187752 990480
rect 206928 990428 206980 990480
rect 295800 990428 295852 990480
rect 309048 990428 309100 990480
rect 314660 990428 314712 990480
rect 324228 990428 324280 990480
rect 324320 990428 324372 990480
rect 343640 990564 343692 990616
rect 343732 990564 343784 990616
rect 357992 990632 358044 990684
rect 372252 990632 372304 990684
rect 488448 990700 488500 990752
rect 527548 990700 527600 990752
rect 629300 990700 629352 990752
rect 372344 990564 372396 990616
rect 372252 990496 372304 990548
rect 386512 990564 386564 990616
rect 475476 990632 475528 990684
rect 546316 990632 546368 990684
rect 563060 990632 563112 990684
rect 486700 990564 486752 990616
rect 475384 990496 475436 990548
rect 476120 990496 476172 990548
rect 488356 990496 488408 990548
rect 582288 990564 582340 990616
rect 587992 990564 588044 990616
rect 623688 990564 623740 990616
rect 537852 990496 537904 990548
rect 585140 990496 585192 990548
rect 623872 990496 623924 990548
rect 639788 990496 639840 990548
rect 353208 990428 353260 990480
rect 353392 990428 353444 990480
rect 364340 990428 364392 990480
rect 397644 990428 397696 990480
rect 405648 990428 405700 990480
rect 546316 990428 546368 990480
rect 226340 990360 226392 990412
rect 233700 990360 233752 990412
rect 246948 990360 247000 990412
rect 285312 990360 285364 990412
rect 295708 990360 295760 990412
rect 233608 990292 233660 990344
rect 244372 990292 244424 990344
rect 256700 990292 256752 990344
rect 424968 990360 425020 990412
rect 430488 990360 430540 990412
rect 430580 990360 430632 990412
rect 383568 990292 383620 990344
rect 397644 990292 397696 990344
rect 405648 990292 405700 990344
rect 463608 990360 463660 990412
rect 469128 990360 469180 990412
rect 469220 990360 469272 990412
rect 471980 990360 472032 990412
rect 444380 990292 444432 990344
rect 315948 990224 316000 990276
rect 325700 990224 325752 990276
rect 405740 990224 405792 990276
rect 471980 990224 472032 990276
rect 486700 990224 486752 990276
rect 42340 990156 42392 990208
rect 79508 990156 79560 990208
rect 639788 990156 639840 990208
rect 673644 990156 673696 990208
rect 42248 990088 42300 990140
rect 78864 990088 78916 990140
rect 88340 990088 88392 990140
rect 325700 990088 325752 990140
rect 343732 990088 343784 990140
rect 628656 990088 628708 990140
rect 629300 990088 629352 990140
rect 673552 990088 673604 990140
rect 42524 990020 42576 990072
rect 673460 990020 673512 990072
rect 674840 985260 674892 985312
rect 675116 985260 675168 985312
rect 41788 969348 41840 969400
rect 42432 969348 42484 969400
rect 42524 968532 42576 968584
rect 41788 968464 41840 968516
rect 42708 968464 42760 968516
rect 42524 966016 42576 966068
rect 42708 966016 42760 966068
rect 674656 966016 674708 966068
rect 674840 966016 674892 966068
rect 673460 964316 673512 964368
rect 675392 964316 675444 964368
rect 673552 963704 673604 963756
rect 675392 963704 675444 963756
rect 41788 962412 41840 962464
rect 42432 962412 42484 962464
rect 42340 960440 42392 960492
rect 42616 960440 42668 960492
rect 41788 957040 41840 957092
rect 42616 957040 42668 957092
rect 42248 956768 42300 956820
rect 673644 953844 673696 953896
rect 675392 953844 675444 953896
rect 42524 946636 42576 946688
rect 42708 946636 42760 946688
rect 674656 932832 674708 932884
rect 674840 932764 674892 932816
rect 42524 927392 42576 927444
rect 42708 927392 42760 927444
rect 39672 922904 39724 922956
rect 42248 922904 42300 922956
rect 39856 915084 39908 915136
rect 41420 915084 41472 915136
rect 42432 915084 42484 915136
rect 673552 910732 673604 910784
rect 677876 910732 677928 910784
rect 675300 908080 675352 908132
rect 677508 908080 677560 908132
rect 42524 908012 42576 908064
rect 42708 908012 42760 908064
rect 41512 906652 41564 906704
rect 42340 906652 42392 906704
rect 674840 902572 674892 902624
rect 674656 902504 674708 902556
rect 674656 894208 674708 894260
rect 674840 894208 674892 894260
rect 42524 888700 42576 888752
rect 42708 888700 42760 888752
rect 41420 875848 41472 875900
rect 42432 875848 42484 875900
rect 673460 875780 673512 875832
rect 675392 875780 675444 875832
rect 673552 874828 673604 874880
rect 675392 874828 675444 874880
rect 675208 870136 675260 870188
rect 675392 870136 675444 870188
rect 673644 864968 673696 865020
rect 675392 864968 675444 865020
rect 675300 862792 675352 862844
rect 675300 862588 675352 862640
rect 42524 850076 42576 850128
rect 42708 850076 42760 850128
rect 44180 836272 44232 836324
rect 44364 836272 44416 836324
rect 674932 836272 674984 836324
rect 675116 836272 675168 836324
rect 674932 827908 674984 827960
rect 677600 827908 677652 827960
rect 39764 827500 39816 827552
rect 44548 827500 44600 827552
rect 674748 823420 674800 823472
rect 676128 823420 676180 823472
rect 675208 818660 675260 818712
rect 676128 818660 676180 818712
rect 677416 818660 677468 818712
rect 44364 805944 44416 805996
rect 44548 805944 44600 805996
rect 41788 799552 41840 799604
rect 42432 799552 42484 799604
rect 41788 798668 41840 798720
rect 42708 798668 42760 798720
rect 41788 792548 41840 792600
rect 42432 792548 42484 792600
rect 42892 792072 42944 792124
rect 43076 792072 43128 792124
rect 674840 792072 674892 792124
rect 675116 792072 675168 792124
rect 41788 787856 41840 787908
rect 42432 787856 42484 787908
rect 42616 787856 42668 787908
rect 673460 786904 673512 786956
rect 673736 786904 673788 786956
rect 675392 786904 675444 786956
rect 41788 786632 41840 786684
rect 42616 786632 42668 786684
rect 673552 786360 673604 786412
rect 675392 786360 675444 786412
rect 675024 780988 675076 781040
rect 675392 780988 675444 781040
rect 673644 774868 673696 774920
rect 673920 774868 673972 774920
rect 675392 774868 675444 774920
rect 675024 773984 675076 774036
rect 675392 773984 675444 774036
rect 42800 772828 42852 772880
rect 43076 772828 43128 772880
rect 44364 767320 44416 767372
rect 44548 767320 44600 767372
rect 42432 756508 42484 756560
rect 42800 756508 42852 756560
rect 41788 756372 41840 756424
rect 42432 756372 42484 756424
rect 41788 754468 41840 754520
rect 42708 754400 42760 754452
rect 41788 749368 41840 749420
rect 42432 749368 42484 749420
rect 673552 746512 673604 746564
rect 674012 746512 674064 746564
rect 41788 745084 41840 745136
rect 42432 745084 42484 745136
rect 42800 745084 42852 745136
rect 41788 744404 41840 744456
rect 42616 744404 42668 744456
rect 673736 741888 673788 741940
rect 675392 741888 675444 741940
rect 674012 740664 674064 740716
rect 675392 740664 675444 740716
rect 44180 739576 44232 739628
rect 44456 739576 44508 739628
rect 674840 739576 674892 739628
rect 674932 739576 674984 739628
rect 675024 735972 675076 736024
rect 675392 735972 675444 736024
rect 674840 734068 674892 734120
rect 674932 734068 674984 734120
rect 42432 730804 42484 730856
rect 42800 730804 42852 730856
rect 673552 730124 673604 730176
rect 673920 730124 673972 730176
rect 675392 730124 675444 730176
rect 673644 729988 673696 730040
rect 674012 729988 674064 730040
rect 675024 729036 675076 729088
rect 675392 729036 675444 729088
rect 44180 720400 44232 720452
rect 44456 720400 44508 720452
rect 674840 714756 674892 714808
rect 675024 714756 675076 714808
rect 41788 713124 41840 713176
rect 42432 713124 42484 713176
rect 41788 711288 41840 711340
rect 42892 711220 42944 711272
rect 42524 708704 42576 708756
rect 42800 708704 42852 708756
rect 41788 706188 41840 706240
rect 42432 706188 42484 706240
rect 41788 700884 41840 700936
rect 42524 700884 42576 700936
rect 42708 700884 42760 700936
rect 41788 700544 41840 700596
rect 42616 700544 42668 700596
rect 673460 695920 673512 695972
rect 673736 695920 673788 695972
rect 675392 695920 675444 695972
rect 674840 695512 674892 695564
rect 675116 695512 675168 695564
rect 42892 695444 42944 695496
rect 43076 695444 43128 695496
rect 673644 695308 673696 695360
rect 675392 695308 675444 695360
rect 675024 691636 675076 691688
rect 675392 691636 675444 691688
rect 673552 685176 673604 685228
rect 675392 685176 675444 685228
rect 675024 684020 675076 684072
rect 675392 684020 675444 684072
rect 44180 681708 44232 681760
rect 44456 681708 44508 681760
rect 674840 676132 674892 676184
rect 675024 676132 675076 676184
rect 41788 669944 41840 669996
rect 42432 669944 42484 669996
rect 41788 669060 41840 669112
rect 42616 669060 42668 669112
rect 42892 669060 42944 669112
rect 41788 663008 41840 663060
rect 42432 663008 42484 663060
rect 41788 657636 41840 657688
rect 42708 657636 42760 657688
rect 42984 657636 43036 657688
rect 41788 657092 41840 657144
rect 42524 657092 42576 657144
rect 42708 657092 42760 657144
rect 674840 656888 674892 656940
rect 675116 656888 675168 656940
rect 673460 651720 673512 651772
rect 675392 651720 675444 651772
rect 673644 651108 673696 651160
rect 675392 651108 675444 651160
rect 675024 645736 675076 645788
rect 675392 645736 675444 645788
rect 44180 643084 44232 643136
rect 44456 643084 44508 643136
rect 673552 639684 673604 639736
rect 675392 639684 675444 639736
rect 675024 638800 675076 638852
rect 675392 638800 675444 638852
rect 674748 637576 674800 637628
rect 675116 637576 675168 637628
rect 42524 633360 42576 633412
rect 42708 633360 42760 633412
rect 41788 626764 41840 626816
rect 42432 626764 42484 626816
rect 41788 625880 41840 625932
rect 42708 625880 42760 625932
rect 674748 623772 674800 623824
rect 673552 623704 673604 623756
rect 44180 623636 44232 623688
rect 44456 623636 44508 623688
rect 673828 623636 673880 623688
rect 674932 623636 674984 623688
rect 41788 619760 41840 619812
rect 42432 619760 42484 619812
rect 42708 618196 42760 618248
rect 42984 618196 43036 618248
rect 674564 618196 674616 618248
rect 674932 618196 674984 618248
rect 41788 614388 41840 614440
rect 42432 614388 42484 614440
rect 42800 614388 42852 614440
rect 41788 614048 41840 614100
rect 42616 614048 42668 614100
rect 673460 606704 673512 606756
rect 674748 606704 674800 606756
rect 675392 606704 675444 606756
rect 673644 605480 673696 605532
rect 675392 605480 675444 605532
rect 44180 604460 44232 604512
rect 44456 604460 44508 604512
rect 673644 604460 673696 604512
rect 673920 604460 673972 604512
rect 675116 600788 675168 600840
rect 675392 600788 675444 600840
rect 674564 599020 674616 599072
rect 674840 599020 674892 599072
rect 674656 598884 674708 598936
rect 674748 598884 674800 598936
rect 674840 598884 674892 598936
rect 675024 598884 675076 598936
rect 673644 594872 673696 594924
rect 673828 594872 673880 594924
rect 675392 594872 675444 594924
rect 675116 593784 675168 593836
rect 675392 593784 675444 593836
rect 44180 585012 44232 585064
rect 44456 585012 44508 585064
rect 42432 583652 42484 583704
rect 42800 583652 42852 583704
rect 41788 583516 41840 583568
rect 42432 583516 42484 583568
rect 41788 581680 41840 581732
rect 42708 581612 42760 581664
rect 42984 581612 43036 581664
rect 674656 579572 674708 579624
rect 675024 579572 675076 579624
rect 41788 576580 41840 576632
rect 42432 576580 42484 576632
rect 41788 572228 41840 572280
rect 42432 572228 42484 572280
rect 42800 572228 42852 572280
rect 41788 571616 41840 571668
rect 42616 571616 42668 571668
rect 44180 565836 44232 565888
rect 44456 565836 44508 565888
rect 44180 564272 44232 564324
rect 44456 564272 44508 564324
rect 673828 561212 673880 561264
rect 674748 561212 674800 561264
rect 675392 561212 675444 561264
rect 673920 560940 673972 560992
rect 675392 560940 675444 560992
rect 674656 560260 674708 560312
rect 674840 560260 674892 560312
rect 42432 556112 42484 556164
rect 42800 556112 42852 556164
rect 675116 555568 675168 555620
rect 675392 555568 675444 555620
rect 673644 550468 673696 550520
rect 675392 550468 675444 550520
rect 675116 548632 675168 548684
rect 675392 548632 675444 548684
rect 674840 540948 674892 541000
rect 675024 540948 675076 541000
rect 41788 540336 41840 540388
rect 42432 540336 42484 540388
rect 41788 538500 41840 538552
rect 42708 538500 42760 538552
rect 41788 533400 41840 533452
rect 42432 533400 42484 533452
rect 41788 529048 41840 529100
rect 42432 529048 42484 529100
rect 42800 529048 42852 529100
rect 41788 527756 41840 527808
rect 42616 527756 42668 527808
rect 44180 527144 44232 527196
rect 44456 527144 44508 527196
rect 674932 514020 674984 514072
rect 676036 514020 676088 514072
rect 677416 514020 677468 514072
rect 675208 513748 675260 513800
rect 676128 513748 676180 513800
rect 677508 513748 677560 513800
rect 676128 507832 676180 507884
rect 677416 507832 677468 507884
rect 44180 507696 44232 507748
rect 44456 507696 44508 507748
rect 42156 498176 42208 498228
rect 42432 498176 42484 498228
rect 44180 488520 44232 488572
rect 44456 488520 44508 488572
rect 42156 478864 42208 478916
rect 42432 478864 42484 478916
rect 42156 469140 42208 469192
rect 42432 469140 42484 469192
rect 675300 467508 675352 467560
rect 677508 467508 677560 467560
rect 39856 463632 39908 463684
rect 42156 463632 42208 463684
rect 42616 463632 42668 463684
rect 42892 463632 42944 463684
rect 673736 463632 673788 463684
rect 673828 463632 673880 463684
rect 676220 459960 676272 460012
rect 677692 459960 677744 460012
rect 39396 458192 39448 458244
rect 42248 458192 42300 458244
rect 44180 449896 44232 449948
rect 44364 449896 44416 449948
rect 673736 449828 673788 449880
rect 673920 449828 673972 449880
rect 42064 442688 42116 442740
rect 42340 442688 42392 442740
rect 42432 441532 42484 441584
rect 42616 441532 42668 441584
rect 676312 440172 676364 440224
rect 677692 440172 677744 440224
rect 674012 430652 674064 430704
rect 673920 430516 673972 430568
rect 676036 427796 676088 427848
rect 677508 427796 677560 427848
rect 42340 425008 42392 425060
rect 42800 425008 42852 425060
rect 42432 422288 42484 422340
rect 42524 422288 42576 422340
rect 676128 420724 676180 420776
rect 677508 420724 677560 420776
rect 42524 411272 42576 411324
rect 44180 411272 44232 411324
rect 44364 411272 44416 411324
rect 42432 411204 42484 411256
rect 41788 411068 41840 411120
rect 42708 411068 42760 411120
rect 673092 408484 673144 408536
rect 676312 408484 676364 408536
rect 41788 401344 41840 401396
rect 42800 401344 42852 401396
rect 42156 397808 42208 397860
rect 42800 397808 42852 397860
rect 675300 388628 675352 388680
rect 676220 388628 676272 388680
rect 673460 384004 673512 384056
rect 675392 384004 675444 384056
rect 673644 382712 673696 382764
rect 675392 382712 675444 382764
rect 44180 372580 44232 372632
rect 44364 372580 44416 372632
rect 673552 372308 673604 372360
rect 675392 372308 675444 372360
rect 42432 370336 42484 370388
rect 42708 370336 42760 370388
rect 42156 370200 42208 370252
rect 42432 370200 42484 370252
rect 41788 367684 41840 367736
rect 42524 367684 42576 367736
rect 41788 358232 41840 358284
rect 42432 358232 42484 358284
rect 42616 358232 42668 358284
rect 41788 357280 41840 357332
rect 42708 357280 42760 357332
rect 42432 356600 42484 356652
rect 42708 356600 42760 356652
rect 42524 353200 42576 353252
rect 42708 353200 42760 353252
rect 42340 339600 42392 339652
rect 42616 339600 42668 339652
rect 673460 338104 673512 338156
rect 673736 338104 673788 338156
rect 675392 338104 675444 338156
rect 673644 337492 673696 337544
rect 675392 337492 675444 337544
rect 44180 333956 44232 334008
rect 44364 333956 44416 334008
rect 673552 328040 673604 328092
rect 675392 328040 675444 328092
rect 41788 324504 41840 324556
rect 42708 324504 42760 324556
rect 41788 313488 41840 313540
rect 42432 313488 42484 313540
rect 42616 313488 42668 313540
rect 673736 293836 673788 293888
rect 674012 293836 674064 293888
rect 675392 293836 675444 293888
rect 673460 293564 673512 293616
rect 673644 293564 673696 293616
rect 675392 293564 675444 293616
rect 42524 286628 42576 286680
rect 42800 286628 42852 286680
rect 41788 282276 41840 282328
rect 42432 282276 42484 282328
rect 42708 282276 42760 282328
rect 673552 282140 673604 282192
rect 675024 282072 675076 282124
rect 675392 282072 675444 282124
rect 41788 270784 41840 270836
rect 42800 270784 42852 270836
rect 42340 270716 42392 270768
rect 42616 270716 42668 270768
rect 44272 270444 44324 270496
rect 44364 270444 44416 270496
rect 675024 265004 675076 265056
rect 673736 264936 673788 264988
rect 673828 264936 673880 264988
rect 674012 264936 674064 264988
rect 44272 256708 44324 256760
rect 44272 256572 44324 256624
rect 673552 249092 673604 249144
rect 673828 249092 673880 249144
rect 675392 249092 675444 249144
rect 673460 248548 673512 248600
rect 673644 248548 673696 248600
rect 675392 248548 675444 248600
rect 42340 246984 42392 247036
rect 42708 246984 42760 247036
rect 41788 239028 41840 239080
rect 42432 239028 42484 239080
rect 42616 239028 42668 239080
rect 673460 237668 673512 237720
rect 673736 237668 673788 237720
rect 675392 237668 675444 237720
rect 42524 237396 42576 237448
rect 42800 237396 42852 237448
rect 41788 227604 41840 227656
rect 42432 227604 42484 227656
rect 42708 227604 42760 227656
rect 44180 218016 44232 218068
rect 44364 218016 44416 218068
rect 673644 206932 673696 206984
rect 675300 206932 675352 206984
rect 673552 202920 673604 202972
rect 675392 202920 675444 202972
rect 42248 197344 42300 197396
rect 42708 197344 42760 197396
rect 41788 195848 41840 195900
rect 42616 195848 42668 195900
rect 44640 195848 44692 195900
rect 673460 191904 673512 191956
rect 675392 191904 675444 191956
rect 41788 185444 41840 185496
rect 42708 185444 42760 185496
rect 41788 184832 41840 184884
rect 42248 184832 42300 184884
rect 42432 184832 42484 184884
rect 673736 184424 673788 184476
rect 675208 184424 675260 184476
rect 42340 179392 42392 179444
rect 42708 179392 42760 179444
rect 44180 179392 44232 179444
rect 44364 179392 44416 179444
rect 673460 177964 673512 178016
rect 673920 177964 673972 178016
rect 44456 173884 44508 173936
rect 44732 173884 44784 173936
rect 673552 168308 673604 168360
rect 673736 168308 673788 168360
rect 675208 168308 675260 168360
rect 675300 168240 675352 168292
rect 44732 160148 44784 160200
rect 44640 160012 44692 160064
rect 673460 157904 673512 157956
rect 675392 157904 675444 157956
rect 673828 157292 673880 157344
rect 675392 157292 675444 157344
rect 44640 154504 44692 154556
rect 44824 154504 44876 154556
rect 673644 147840 673696 147892
rect 673920 147840 673972 147892
rect 675392 147840 675444 147892
rect 44180 140768 44232 140820
rect 44364 140768 44416 140820
rect 673460 129684 673512 129736
rect 673736 129684 673788 129736
rect 673828 129684 673880 129736
rect 675300 129684 675352 129736
rect 39856 125128 39908 125180
rect 44180 125128 44232 125180
rect 39856 120164 39908 120216
rect 44732 120164 44784 120216
rect 673460 112752 673512 112804
rect 673736 112752 673788 112804
rect 675392 112752 675444 112804
rect 673552 112072 673604 112124
rect 675392 112072 675444 112124
rect 673644 101668 673696 101720
rect 675392 101668 675444 101720
rect 44272 96568 44324 96620
rect 44456 96568 44508 96620
rect 44272 77256 44324 77308
rect 44364 77256 44416 77308
rect 39672 74876 39724 74928
rect 39856 74876 39908 74928
rect 44180 71748 44232 71800
rect 44364 71748 44416 71800
rect 39580 67940 39632 67992
rect 41420 67940 41472 67992
rect 41420 64472 41472 64524
rect 42708 64472 42760 64524
rect 39672 52368 39724 52420
rect 39856 52368 39908 52420
rect 42248 45840 42300 45892
rect 145104 45840 145156 45892
rect 42708 45772 42760 45824
rect 140964 45772 141016 45824
rect 578792 45704 578844 45756
rect 673552 45704 673604 45756
rect 44180 45636 44232 45688
rect 145840 45636 145892 45688
rect 528652 45636 528704 45688
rect 673092 45636 673144 45688
rect 39856 45568 39908 45620
rect 189264 45568 189316 45620
rect 529848 45568 529900 45620
rect 673460 45568 673512 45620
rect 44916 45500 44968 45552
rect 195980 45500 196032 45552
rect 516324 45500 516376 45552
rect 673644 45500 673696 45552
rect 289820 44820 289872 44872
rect 313188 44820 313240 44872
rect 458180 44820 458232 44872
rect 250996 44752 251048 44804
rect 252100 44752 252152 44804
rect 276020 44752 276072 44804
rect 380900 44752 380952 44804
rect 400128 44752 400180 44804
rect 406752 44752 406804 44804
rect 461492 44752 461544 44804
rect 193128 44616 193180 44668
rect 231860 44684 231912 44736
rect 308220 44684 308272 44736
rect 358728 44684 358780 44736
rect 362408 44684 362460 44736
rect 247684 44616 247736 44668
rect 307576 44616 307628 44668
rect 308312 44616 308364 44668
rect 309140 44616 309192 44668
rect 328368 44616 328420 44668
rect 347780 44616 347832 44668
rect 488540 44684 488592 44736
rect 499580 44684 499632 44736
rect 386420 44616 386472 44668
rect 405648 44616 405700 44668
rect 417240 44616 417292 44668
rect 425060 44616 425112 44668
rect 444288 44616 444340 44668
rect 471980 44616 472032 44668
rect 472072 44616 472124 44668
rect 472348 44616 472400 44668
rect 488448 44616 488500 44668
rect 518808 44616 518860 44668
rect 526812 44684 526864 44736
rect 546592 44820 546644 44872
rect 560300 44820 560352 44872
rect 546408 44684 546460 44736
rect 140964 44480 141016 44532
rect 173900 44548 173952 44600
rect 289820 44548 289872 44600
rect 309416 44548 309468 44600
rect 199660 44480 199712 44532
rect 212540 44480 212592 44532
rect 218060 44480 218112 44532
rect 195980 44412 196032 44464
rect 200764 44412 200816 44464
rect 200856 44412 200908 44464
rect 217876 44412 217928 44464
rect 276020 44480 276072 44532
rect 299572 44480 299624 44532
rect 305736 44480 305788 44532
rect 313188 44548 313240 44600
rect 380900 44548 380952 44600
rect 400128 44548 400180 44600
rect 419540 44548 419592 44600
rect 438768 44548 438820 44600
rect 458180 44548 458232 44600
rect 242900 44412 242952 44464
rect 297732 44412 297784 44464
rect 300768 44412 300820 44464
rect 306380 44412 306432 44464
rect 352564 44480 352616 44532
rect 355600 44480 355652 44532
rect 359924 44480 359976 44532
rect 364156 44480 364208 44532
rect 407396 44480 407448 44532
rect 410432 44480 410484 44532
rect 419080 44480 419132 44532
rect 462136 44480 462188 44532
rect 465172 44480 465224 44532
rect 473820 44480 473872 44532
rect 516968 44480 517020 44532
rect 351920 44412 351972 44464
rect 354404 44412 354456 44464
rect 360568 44412 360620 44464
rect 363052 44412 363104 44464
rect 413560 44412 413612 44464
rect 417884 44412 417936 44464
rect 468300 44412 468352 44464
rect 472624 44412 472676 44464
rect 523132 44412 523184 44464
rect 199016 44344 199068 44396
rect 217968 44344 218020 44396
rect 218152 44344 218204 44396
rect 247408 44344 247460 44396
rect 247684 44344 247736 44396
rect 289820 44344 289872 44396
rect 248328 44276 248380 44328
rect 267740 44276 267792 44328
rect 286968 44276 287020 44328
rect 359372 44344 359424 44396
rect 414204 44344 414256 44396
rect 468944 44344 468996 44396
rect 523776 44344 523828 44396
rect 360568 44276 360620 44328
rect 406752 44276 406804 44328
rect 411076 44276 411128 44328
rect 145104 44208 145156 44260
rect 195336 44208 195388 44260
rect 199660 44208 199712 44260
rect 200764 44208 200816 44260
rect 304540 44208 304592 44260
rect 307576 44208 307628 44260
rect 308312 44208 308364 44260
rect 186688 44140 186740 44192
rect 194692 44140 194744 44192
rect 295248 44140 295300 44192
rect 303252 44140 303304 44192
rect 306380 44140 306432 44192
rect 309416 44140 309468 44192
rect 350080 44140 350132 44192
rect 358084 44140 358136 44192
rect 404912 44140 404964 44192
rect 412916 44140 412968 44192
rect 419540 44276 419592 44328
rect 438768 44276 438820 44328
rect 461492 44276 461544 44328
rect 516324 44276 516376 44328
rect 465816 44208 465868 44260
rect 474464 44208 474516 44260
rect 514484 44208 514536 44260
rect 522488 44208 522540 44260
rect 523132 44208 523184 44260
rect 527456 44208 527508 44260
rect 529848 44208 529900 44260
rect 419724 44140 419776 44192
rect 459652 44140 459704 44192
rect 467656 44140 467708 44192
rect 518808 44140 518860 44192
rect 524972 44140 525024 44192
rect 525616 44140 525668 44192
rect 528652 44140 528704 44192
rect 39764 44072 39816 44124
rect 78956 44072 79008 44124
rect 347780 43664 347832 43716
rect 362408 43664 362460 43716
rect 303896 42236 303948 42288
rect 308220 42236 308272 42288
rect 189264 41896 189316 41948
rect 191104 41896 191156 41948
rect 192300 41896 192352 41948
rect 193588 41896 193640 41948
rect 196440 41896 196492 41948
rect 198464 41896 198516 41948
rect 200120 41896 200172 41948
rect 363512 41896 363564 41948
rect 135352 41692 135404 41744
rect 154488 41692 154540 41744
rect 91284 41556 91336 41608
rect 102140 41556 102192 41608
rect 102048 41488 102100 41540
rect 154488 41556 154540 41608
rect 168288 41692 168340 41744
rect 188620 41828 188672 41880
rect 192944 41828 192996 41880
rect 201592 41828 201644 41880
rect 202512 41828 202564 41880
rect 299480 41828 299532 41880
rect 360016 41828 360068 41880
rect 361120 41828 361172 41880
rect 409328 41828 409380 41880
rect 412364 41828 412416 41880
rect 415216 41828 415268 41880
rect 465356 41828 465408 41880
rect 466368 41828 466420 41880
rect 469404 41828 469456 41880
rect 470692 41828 470744 41880
rect 473084 41828 473136 41880
rect 517060 41828 517112 41880
rect 520096 41828 520148 41880
rect 521384 41828 521436 41880
rect 524420 41828 524472 41880
rect 525524 41828 525576 41880
rect 198924 41760 198976 41812
rect 296904 41760 296956 41812
rect 305276 41760 305328 41812
rect 306288 41760 306340 41812
rect 358820 41760 358872 41812
rect 362960 41760 363012 41812
rect 410524 41760 410576 41812
rect 411536 41760 411588 41812
rect 414572 41760 414624 41812
rect 415860 41760 415912 41812
rect 418252 41760 418304 41812
rect 464160 41760 464212 41812
rect 467196 41760 467248 41812
rect 470048 41760 470100 41812
rect 523868 41760 523920 41812
rect 526904 41760 526956 41812
rect 121368 41488 121420 41540
rect 121460 41488 121512 41540
rect 135260 41420 135312 41472
rect 149980 41420 150032 41472
rect 253940 41556 253992 41608
rect 168288 41352 168340 41404
rect 202512 41420 202564 41472
rect 240140 41420 240192 41472
rect 569132 41488 569184 41540
rect 629300 41420 629352 41472
rect 78956 40196 79008 40248
rect 86500 40196 86552 40248
rect 91284 40196 91336 40248
rect 133098 40196 133150 40248
rect 143816 40196 143868 40248
rect 140996 40060 141048 40112
rect 143072 40060 143124 40112
rect 143356 40060 143408 40112
<< metal2 >>
rect 585704 997529 585732 997628
rect 585046 997520 585102 997529
rect 585046 997455 585102 997464
rect 585690 997520 585746 997529
rect 585690 997455 585746 997464
rect 589554 997520 589610 997529
rect 589554 997455 589610 997464
rect 343638 997112 343694 997121
rect 343638 997047 343694 997056
rect 77049 995407 77105 995887
rect 77693 995407 77749 995887
rect 78337 995407 78393 995887
rect 44088 992248 44140 992254
rect 44088 992190 44140 992196
rect 42340 990208 42392 990214
rect 42340 990150 42392 990156
rect 42248 990140 42300 990146
rect 42248 990082 42300 990088
rect 41722 969870 41828 969898
rect 41800 969406 41828 969870
rect 41788 969400 41840 969406
rect 41788 969342 41840 969348
rect 41713 969217 42193 969273
rect 41788 968516 41840 968522
rect 41788 968458 41840 968464
rect 41800 968063 41828 968458
rect 41722 968035 41828 968063
rect 41713 967377 42193 967433
rect 41713 966733 42193 966789
rect 41713 965537 42193 965593
rect 41713 964341 42193 964397
rect 41713 963697 42193 963753
rect 41713 963053 42193 963109
rect 41713 962501 42193 962557
rect 41788 962464 41840 962470
rect 41788 962406 41840 962412
rect 41800 961874 41828 962406
rect 41722 961846 41828 961874
rect 41713 961213 42193 961269
rect 41713 960569 42193 960625
rect 41713 960017 42193 960073
rect 41713 959373 42193 959429
rect 41713 958729 42193 958785
rect 41713 958177 42193 958233
rect 41722 957547 41828 957575
rect 41800 957098 41828 957547
rect 41788 957092 41840 957098
rect 41788 957034 41840 957040
rect 42260 956931 42288 990082
rect 42352 960498 42380 990150
rect 42524 990072 42576 990078
rect 42524 990014 42576 990020
rect 42432 969400 42484 969406
rect 42432 969342 42484 969348
rect 42444 962470 42472 969342
rect 42536 968590 42564 990014
rect 42524 968584 42576 968590
rect 42524 968526 42576 968532
rect 42708 968516 42760 968522
rect 42708 968458 42760 968464
rect 42720 966074 42748 968458
rect 42524 966068 42576 966074
rect 42524 966010 42576 966016
rect 42708 966068 42760 966074
rect 42708 966010 42760 966016
rect 42432 962464 42484 962470
rect 42432 962406 42484 962412
rect 42340 960492 42392 960498
rect 42340 960434 42392 960440
rect 41722 956903 42288 956931
rect 42248 956820 42300 956826
rect 42248 956762 42300 956768
rect 41713 956337 42193 956393
rect 41713 955693 42193 955749
rect 41713 955049 42193 955105
rect 42260 941202 42288 956762
rect 42536 946694 42564 966010
rect 42616 960492 42668 960498
rect 42616 960434 42668 960440
rect 42628 957098 42656 960434
rect 42616 957092 42668 957098
rect 42616 957034 42668 957040
rect 42524 946688 42576 946694
rect 42524 946630 42576 946636
rect 42708 946688 42760 946694
rect 42708 946630 42760 946636
rect 42260 941174 42472 941202
rect 39486 928160 39542 928169
rect 39486 928095 39542 928104
rect 39500 922978 39528 928095
rect 39330 922962 39712 922978
rect 39330 922956 39724 922962
rect 39330 922950 39672 922956
rect 39672 922898 39724 922904
rect 42248 922956 42300 922962
rect 42248 922898 42300 922904
rect 41510 919728 41566 919737
rect 41510 919663 41566 919672
rect 39567 919006 39896 919034
rect 39868 915142 39896 919006
rect 41524 917289 41552 919663
rect 41510 917280 41566 917289
rect 41510 917215 41566 917224
rect 39856 915136 39908 915142
rect 39856 915078 39908 915084
rect 41420 915136 41472 915142
rect 41420 915078 41472 915084
rect 39330 912206 39620 912234
rect 39592 908177 39620 912206
rect 39578 908168 39634 908177
rect 39578 908103 39634 908112
rect 40038 908032 40094 908041
rect 40038 907967 40094 907976
rect 40052 889001 40080 907967
rect 40038 888992 40094 889001
rect 40038 888927 40094 888936
rect 40130 877568 40186 877577
rect 40130 877503 40186 877512
rect 40144 870097 40172 877503
rect 41432 875906 41460 915078
rect 41524 912257 41552 917215
rect 41510 912248 41566 912257
rect 41510 912183 41566 912192
rect 41524 906710 41552 912183
rect 41512 906704 41564 906710
rect 41512 906646 41564 906652
rect 41420 875900 41472 875906
rect 41420 875842 41472 875848
rect 41432 875129 41460 875842
rect 41418 875120 41474 875129
rect 41418 875055 41474 875064
rect 40130 870088 40186 870097
rect 40130 870023 40186 870032
rect 39854 869408 39910 869417
rect 39854 869343 39910 869352
rect 39868 850377 39896 869343
rect 39854 850368 39910 850377
rect 39854 850303 39910 850312
rect 39606 827750 39804 827778
rect 39776 827558 39804 827750
rect 39764 827552 39816 827558
rect 39762 827520 39764 827529
rect 39816 827520 39818 827529
rect 39762 827455 39818 827464
rect 41722 800075 41828 800103
rect 41800 799610 41828 800075
rect 41788 799604 41840 799610
rect 41788 799546 41840 799552
rect 41713 799417 42193 799473
rect 41788 798720 41840 798726
rect 41788 798662 41840 798668
rect 41800 798266 41828 798662
rect 41722 798238 41828 798266
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 41788 792600 41840 792606
rect 41788 792542 41840 792548
rect 41800 792099 41828 792542
rect 41722 792071 41828 792099
rect 41713 791413 42193 791469
rect 41713 790769 42193 790825
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 41788 787908 41840 787914
rect 41788 787850 41840 787856
rect 41800 787794 41828 787850
rect 41722 787766 41828 787794
rect 41722 787086 41828 787114
rect 41800 786690 41828 787086
rect 41788 786684 41840 786690
rect 41788 786626 41840 786632
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 41722 756894 41828 756922
rect 41800 756430 41828 756894
rect 41788 756424 41840 756430
rect 41788 756366 41840 756372
rect 41713 756217 42193 756273
rect 41722 755035 41828 755063
rect 41800 754526 41828 755035
rect 41788 754520 41840 754526
rect 41788 754462 41840 754468
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 41788 749420 41840 749426
rect 41788 749362 41840 749368
rect 41800 748898 41828 749362
rect 41722 748870 41828 748898
rect 41713 748213 42193 748269
rect 41713 747569 42193 747625
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 41788 745136 41840 745142
rect 41788 745078 41840 745084
rect 41800 744575 41828 745078
rect 41722 744547 41828 744575
rect 41788 744456 41840 744462
rect 41788 744398 41840 744404
rect 41800 743931 41828 744398
rect 41722 743903 41828 743931
rect 41713 743337 42193 743393
rect 41713 742693 42193 742749
rect 41713 742049 42193 742105
rect 41722 713675 41828 713703
rect 41800 713182 41828 713675
rect 41788 713176 41840 713182
rect 41788 713118 41840 713124
rect 41713 713017 42193 713073
rect 41722 711835 41828 711863
rect 41800 711346 41828 711835
rect 41788 711340 41840 711346
rect 41788 711282 41840 711288
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 41788 706240 41840 706246
rect 41788 706182 41840 706188
rect 41800 705699 41828 706182
rect 41722 705671 41828 705699
rect 41713 705013 42193 705069
rect 41713 704369 42193 704425
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 41722 701347 41828 701375
rect 41800 700942 41828 701347
rect 41788 700936 41840 700942
rect 41788 700878 41840 700884
rect 41722 700726 41828 700754
rect 41800 700602 41828 700726
rect 41788 700596 41840 700602
rect 41788 700538 41840 700544
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 41722 670475 41828 670503
rect 41800 670002 41828 670475
rect 41788 669996 41840 670002
rect 41788 669938 41840 669944
rect 41713 669817 42193 669873
rect 41788 669112 41840 669118
rect 41788 669054 41840 669060
rect 41800 668658 41828 669054
rect 41722 668630 41828 668658
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 41788 663060 41840 663066
rect 41788 663002 41840 663008
rect 41800 662499 41828 663002
rect 41722 662471 41828 662499
rect 41713 661813 42193 661869
rect 41713 661169 42193 661225
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 41722 658158 41828 658186
rect 41800 657694 41828 658158
rect 41788 657688 41840 657694
rect 41788 657630 41840 657636
rect 41722 657478 41828 657506
rect 41800 657150 41828 657478
rect 41788 657144 41840 657150
rect 41788 657086 41840 657092
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 41722 627286 41828 627314
rect 41800 626822 41828 627286
rect 41788 626816 41840 626822
rect 41788 626758 41840 626764
rect 41713 626617 42193 626673
rect 41788 625932 41840 625938
rect 41788 625874 41840 625880
rect 41800 625463 41828 625874
rect 41722 625435 41828 625463
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 41788 619812 41840 619818
rect 41788 619754 41840 619760
rect 41800 619290 41828 619754
rect 41722 619262 41828 619290
rect 41713 618613 42193 618669
rect 41713 617969 42193 618025
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41722 614947 41828 614975
rect 41800 614446 41828 614947
rect 41788 614440 41840 614446
rect 41788 614382 41840 614388
rect 41722 614303 41828 614331
rect 41800 614106 41828 614303
rect 41788 614100 41840 614106
rect 41788 614042 41840 614048
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 41722 584075 41828 584103
rect 41800 583574 41828 584075
rect 41788 583568 41840 583574
rect 41788 583510 41840 583516
rect 41713 583417 42193 583473
rect 41722 582235 41828 582263
rect 41800 581738 41828 582235
rect 41788 581732 41840 581738
rect 41788 581674 41840 581680
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 41788 576632 41840 576638
rect 41788 576574 41840 576580
rect 41800 576099 41828 576574
rect 41722 576071 41828 576099
rect 41713 575413 42193 575469
rect 41713 574769 42193 574825
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 41788 572280 41840 572286
rect 41788 572222 41840 572228
rect 41800 571775 41828 572222
rect 41722 571747 41828 571775
rect 41788 571668 41840 571674
rect 41788 571610 41840 571616
rect 41800 571146 41828 571610
rect 41722 571118 41828 571146
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 41722 540875 41828 540903
rect 41800 540394 41828 540875
rect 41788 540388 41840 540394
rect 41788 540330 41840 540336
rect 41713 540217 42193 540273
rect 41722 539022 41828 539050
rect 41800 538558 41828 539022
rect 41788 538552 41840 538558
rect 41788 538494 41840 538500
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 41788 533452 41840 533458
rect 41788 533394 41840 533400
rect 41800 532899 41828 533394
rect 41722 532871 41828 532899
rect 41713 532213 42193 532269
rect 41713 531569 42193 531625
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 41788 529100 41840 529106
rect 41788 529042 41840 529048
rect 41800 528578 41828 529042
rect 41722 528550 41828 528578
rect 41722 527903 41828 527931
rect 41800 527814 41828 527903
rect 41788 527808 41840 527814
rect 41788 527750 41840 527756
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 40222 516080 40278 516089
rect 40222 516015 40278 516024
rect 40236 497049 40264 516015
rect 42156 498228 42208 498234
rect 42156 498170 42208 498176
rect 40222 497040 40278 497049
rect 40222 496975 40278 496984
rect 39606 493190 39804 493218
rect 39776 492969 39804 493190
rect 39762 492960 39818 492969
rect 39762 492895 39818 492904
rect 39854 490512 39910 490521
rect 39854 490447 39910 490456
rect 39868 488073 39896 490447
rect 39854 488064 39910 488073
rect 39854 487999 39910 488008
rect 42168 478922 42196 498170
rect 42156 478916 42208 478922
rect 42156 478858 42208 478864
rect 40038 470656 40094 470665
rect 40038 470591 40094 470600
rect 39856 463684 39908 463690
rect 39856 463626 39908 463632
rect 39396 458244 39448 458250
rect 39396 458186 39448 458192
rect 39408 451874 39436 458186
rect 39670 451888 39726 451897
rect 39330 451846 39670 451874
rect 39670 451823 39726 451832
rect 39868 447794 39896 463626
rect 40052 461009 40080 470591
rect 42156 469192 42208 469198
rect 42156 469134 42208 469140
rect 42168 463690 42196 469134
rect 42156 463684 42208 463690
rect 42156 463626 42208 463632
rect 40038 461000 40094 461009
rect 40038 460935 40094 460944
rect 42260 458250 42288 922898
rect 42444 915142 42472 941174
rect 42720 927450 42748 946630
rect 42524 927444 42576 927450
rect 42524 927386 42576 927392
rect 42708 927444 42760 927450
rect 42708 927386 42760 927392
rect 42432 915136 42484 915142
rect 42432 915078 42484 915084
rect 42536 908070 42564 927386
rect 42524 908064 42576 908070
rect 42524 908006 42576 908012
rect 42708 908064 42760 908070
rect 42708 908006 42760 908012
rect 42340 906704 42392 906710
rect 42340 906646 42392 906652
rect 42248 458244 42300 458250
rect 42248 458186 42300 458192
rect 39946 455424 40002 455433
rect 39946 455359 40002 455368
rect 39567 447766 39896 447794
rect 39868 444417 39896 447766
rect 39854 444408 39910 444417
rect 39854 444343 39910 444352
rect 39670 441008 39726 441017
rect 39330 440966 39620 440994
rect 39592 440858 39620 440966
rect 39670 440943 39726 440952
rect 39684 440858 39712 440943
rect 39960 440858 39988 455359
rect 42352 448633 42380 906646
rect 42720 888758 42748 908006
rect 42524 888752 42576 888758
rect 42524 888694 42576 888700
rect 42708 888752 42760 888758
rect 42708 888694 42760 888700
rect 42432 875900 42484 875906
rect 42432 875842 42484 875848
rect 42444 807378 42472 875842
rect 42536 869417 42564 888694
rect 44100 877577 44128 992190
rect 78876 990826 78904 995452
rect 78864 990820 78916 990826
rect 78864 990762 78916 990768
rect 78876 990146 78904 990762
rect 79520 990758 79548 995452
rect 80177 995407 80233 995887
rect 80729 995407 80785 995887
rect 81373 995407 81429 995887
rect 82017 995407 82073 995887
rect 82569 995407 82625 995887
rect 83213 995407 83269 995887
rect 84016 995648 84068 995654
rect 84016 995590 84068 995596
rect 84028 995466 84056 995590
rect 83858 995438 84056 995466
rect 84501 995407 84557 995887
rect 85053 995407 85109 995887
rect 85697 995407 85753 995887
rect 86341 995407 86397 995887
rect 87537 995407 87593 995887
rect 88733 995407 88789 995887
rect 89377 995407 89433 995887
rect 79508 990752 79560 990758
rect 79508 990694 79560 990700
rect 79520 990214 79548 990694
rect 90008 990690 90036 995452
rect 91217 995407 91273 995887
rect 91744 995648 91796 995654
rect 91744 995590 91796 995596
rect 91756 995466 91784 995590
rect 91756 995438 91862 995466
rect 128449 995407 128505 995887
rect 129093 995407 129149 995887
rect 129737 995407 129793 995887
rect 130304 990826 130332 995452
rect 130292 990820 130344 990826
rect 130292 990762 130344 990768
rect 130948 990758 130976 995452
rect 131577 995407 131633 995887
rect 132129 995407 132185 995887
rect 132773 995407 132829 995887
rect 133417 995407 133473 995887
rect 133969 995407 134025 995887
rect 134613 995407 134669 995887
rect 135352 995512 135404 995518
rect 135286 995460 135352 995466
rect 135286 995454 135404 995460
rect 135286 995438 135392 995454
rect 135901 995407 135957 995887
rect 136453 995407 136509 995887
rect 137097 995407 137153 995887
rect 137741 995407 137797 995887
rect 138937 995407 138993 995887
rect 140133 995407 140189 995887
rect 140777 995407 140833 995887
rect 132408 990820 132460 990826
rect 132408 990762 132460 990768
rect 130936 990752 130988 990758
rect 130936 990694 130988 990700
rect 88340 990684 88392 990690
rect 88340 990626 88392 990632
rect 89996 990684 90048 990690
rect 89996 990626 90048 990632
rect 79508 990208 79560 990214
rect 79508 990150 79560 990156
rect 88352 990146 88380 990626
rect 132420 990622 132448 990762
rect 141436 990690 141464 995452
rect 142617 995407 142673 995887
rect 143172 995512 143224 995518
rect 143224 995460 143290 995466
rect 143172 995454 143290 995460
rect 143184 995438 143290 995454
rect 179849 995407 179905 995887
rect 180493 995407 180549 995887
rect 181137 995407 181193 995887
rect 181717 995438 181760 995466
rect 182361 995438 182404 995466
rect 181732 990826 181760 995438
rect 181720 990820 181772 990826
rect 181720 990762 181772 990768
rect 141424 990684 141476 990690
rect 141424 990626 141476 990632
rect 181732 990622 181760 990762
rect 182376 990758 182404 995438
rect 182977 995407 183033 995887
rect 183529 995407 183585 995887
rect 184173 995407 184229 995887
rect 184817 995407 184873 995887
rect 185369 995407 185425 995887
rect 186013 995407 186069 995887
rect 186685 995438 186728 995466
rect 182364 990752 182416 990758
rect 182364 990694 182416 990700
rect 186700 990622 186728 995438
rect 187301 995407 187357 995887
rect 187853 995407 187909 995887
rect 188497 995407 188553 995887
rect 189141 995407 189197 995887
rect 190337 995407 190393 995887
rect 191533 995407 191589 995887
rect 192177 995407 192233 995887
rect 192849 995438 192892 995466
rect 187700 990752 187752 990758
rect 187700 990694 187752 990700
rect 132408 990616 132460 990622
rect 132408 990558 132460 990564
rect 181720 990616 181772 990622
rect 181720 990558 181772 990564
rect 186688 990616 186740 990622
rect 186688 990558 186740 990564
rect 187712 990486 187740 990694
rect 192864 990690 192892 995438
rect 194017 995407 194073 995887
rect 194689 995438 194732 995466
rect 192852 990684 192904 990690
rect 192852 990626 192904 990632
rect 194704 990622 194732 995438
rect 231249 995407 231305 995887
rect 231893 995407 231949 995887
rect 232537 995407 232593 995887
rect 233068 995438 233117 995466
rect 233712 995438 233761 995466
rect 233068 990826 233096 995438
rect 233056 990820 233108 990826
rect 233056 990762 233108 990768
rect 206928 990752 206980 990758
rect 206928 990694 206980 990700
rect 226340 990752 226392 990758
rect 226340 990694 226392 990700
rect 194692 990616 194744 990622
rect 194692 990558 194744 990564
rect 206940 990486 206968 990694
rect 187700 990480 187752 990486
rect 187700 990422 187752 990428
rect 206928 990480 206980 990486
rect 206928 990422 206980 990428
rect 226352 990418 226380 990694
rect 233068 990554 233096 990762
rect 233608 990616 233660 990622
rect 233608 990558 233660 990564
rect 233056 990548 233108 990554
rect 233056 990490 233108 990496
rect 226340 990412 226392 990418
rect 226340 990354 226392 990360
rect 233620 990350 233648 990558
rect 233712 990418 233740 995438
rect 234377 995407 234433 995887
rect 234929 995407 234985 995887
rect 235573 995407 235629 995887
rect 236217 995407 236273 995887
rect 236769 995407 236825 995887
rect 237413 995407 237469 995887
rect 238085 995450 238248 995466
rect 238085 995444 238260 995450
rect 238085 995438 238208 995444
rect 238701 995407 238757 995887
rect 239253 995407 239309 995887
rect 239897 995407 239953 995887
rect 240541 995407 240597 995887
rect 241737 995407 241793 995887
rect 242933 995407 242989 995887
rect 243577 995407 243633 995887
rect 244200 995574 244412 995602
rect 244200 995466 244228 995574
rect 244200 995438 244249 995466
rect 238208 995386 238260 995392
rect 244384 990622 244412 995574
rect 245417 995407 245473 995887
rect 245948 995450 246089 995466
rect 245936 995444 246089 995450
rect 245988 995438 246089 995444
rect 282849 995407 282905 995887
rect 283493 995407 283549 995887
rect 284137 995407 284193 995887
rect 245936 995386 245988 995392
rect 256608 990752 256660 990758
rect 256608 990694 256660 990700
rect 246948 990684 247000 990690
rect 246948 990626 247000 990632
rect 244372 990616 244424 990622
rect 244372 990558 244424 990564
rect 233700 990412 233752 990418
rect 233700 990354 233752 990360
rect 244384 990350 244412 990558
rect 246960 990418 246988 990626
rect 256620 990554 256648 990694
rect 284680 990622 284708 995452
rect 285324 990826 285352 995452
rect 285977 995407 286033 995887
rect 286529 995407 286585 995887
rect 287173 995407 287229 995887
rect 287817 995407 287873 995887
rect 288369 995407 288425 995887
rect 289013 995407 289069 995887
rect 289648 995314 289676 995452
rect 290301 995407 290357 995887
rect 290853 995407 290909 995887
rect 291497 995407 291553 995887
rect 292141 995407 292197 995887
rect 293337 995407 293393 995887
rect 294533 995407 294589 995887
rect 295177 995407 295233 995887
rect 289636 995308 289688 995314
rect 289636 995250 289688 995256
rect 285312 990820 285364 990826
rect 285312 990762 285364 990768
rect 295708 990820 295760 990826
rect 295708 990762 295760 990768
rect 256700 990616 256752 990622
rect 256700 990558 256752 990564
rect 284576 990616 284628 990622
rect 284668 990616 284720 990622
rect 284628 990576 284668 990604
rect 284576 990558 284628 990564
rect 284668 990558 284720 990564
rect 256608 990548 256660 990554
rect 256608 990490 256660 990496
rect 246948 990412 247000 990418
rect 246948 990354 247000 990360
rect 256712 990350 256740 990558
rect 285324 990418 285352 990762
rect 295524 990752 295576 990758
rect 295524 990694 295576 990700
rect 289820 990616 289872 990622
rect 289818 990584 289820 990593
rect 295536 990593 295564 990694
rect 289872 990584 289874 990593
rect 289818 990519 289874 990528
rect 295522 990584 295578 990593
rect 295522 990519 295578 990528
rect 295720 990418 295748 990762
rect 295812 990486 295840 995452
rect 297017 995407 297073 995887
rect 297652 995314 297680 995452
rect 297640 995308 297692 995314
rect 297640 995250 297692 995256
rect 329562 992352 329618 992361
rect 329562 992287 329618 992296
rect 329576 992254 329604 992287
rect 329564 992248 329616 992254
rect 329564 992190 329616 992196
rect 333900 990826 334020 990842
rect 343652 990826 343680 997047
rect 384649 995407 384705 995887
rect 385293 995407 385349 995887
rect 385937 995407 385993 995887
rect 324228 990820 324280 990826
rect 324228 990762 324280 990768
rect 333888 990820 334020 990826
rect 333940 990814 334020 990820
rect 333888 990762 333940 990768
rect 314660 990752 314712 990758
rect 314660 990694 314712 990700
rect 309048 990616 309100 990622
rect 309048 990558 309100 990564
rect 309060 990486 309088 990558
rect 314672 990486 314700 990694
rect 315948 990616 316000 990622
rect 315948 990558 316000 990564
rect 295800 990480 295852 990486
rect 295800 990422 295852 990428
rect 309048 990480 309100 990486
rect 309048 990422 309100 990428
rect 314660 990480 314712 990486
rect 314660 990422 314712 990428
rect 285312 990412 285364 990418
rect 285312 990354 285364 990360
rect 295708 990412 295760 990418
rect 295708 990354 295760 990360
rect 233608 990344 233660 990350
rect 233608 990286 233660 990292
rect 244372 990344 244424 990350
rect 244372 990286 244424 990292
rect 256700 990344 256752 990350
rect 256700 990286 256752 990292
rect 315960 990282 315988 990558
rect 324240 990486 324268 990762
rect 333992 990758 334020 990814
rect 343640 990820 343692 990826
rect 343640 990762 343692 990768
rect 353300 990820 353352 990826
rect 353300 990762 353352 990768
rect 324320 990752 324372 990758
rect 324320 990694 324372 990700
rect 333980 990752 334032 990758
rect 333980 990694 334032 990700
rect 324332 990486 324360 990694
rect 343652 990622 343680 990762
rect 353312 990690 353340 990762
rect 357808 990752 357860 990758
rect 372344 990752 372396 990758
rect 357860 990700 358032 990706
rect 357808 990694 358032 990700
rect 372344 990694 372396 990700
rect 357820 990690 358032 990694
rect 353300 990684 353352 990690
rect 357820 990684 358044 990690
rect 357820 990678 357992 990684
rect 353300 990626 353352 990632
rect 357992 990626 358044 990632
rect 372252 990684 372304 990690
rect 372252 990626 372304 990632
rect 343640 990616 343692 990622
rect 343640 990558 343692 990564
rect 343732 990616 343784 990622
rect 343732 990558 343784 990564
rect 324228 990480 324280 990486
rect 324228 990422 324280 990428
rect 324320 990480 324372 990486
rect 324320 990422 324372 990428
rect 315948 990276 316000 990282
rect 315948 990218 316000 990224
rect 325700 990276 325752 990282
rect 325700 990218 325752 990224
rect 325712 990146 325740 990218
rect 343744 990146 343772 990558
rect 372264 990554 372292 990626
rect 372356 990622 372384 990694
rect 386524 990622 386552 995452
rect 387168 990826 387196 995452
rect 387777 995407 387833 995887
rect 388329 995407 388385 995887
rect 388973 995407 389029 995887
rect 389617 995407 389673 995887
rect 390169 995407 390225 995887
rect 390813 995407 390869 995887
rect 391492 995314 391520 995452
rect 392101 995407 392157 995887
rect 392653 995407 392709 995887
rect 393297 995407 393353 995887
rect 393941 995407 393997 995887
rect 395137 995407 395193 995887
rect 396333 995407 396389 995887
rect 396977 995407 397033 995887
rect 391480 995308 391532 995314
rect 391480 995250 391532 995256
rect 387156 990820 387208 990826
rect 387156 990762 387208 990768
rect 372344 990616 372396 990622
rect 372344 990558 372396 990564
rect 386512 990616 386564 990622
rect 386512 990558 386564 990564
rect 372252 990548 372304 990554
rect 372252 990490 372304 990496
rect 397656 990486 397684 995452
rect 398817 995407 398873 995887
rect 399496 995314 399524 995452
rect 473649 995407 473705 995887
rect 474293 995407 474349 995887
rect 474937 995407 474993 995887
rect 399484 995308 399536 995314
rect 399484 995250 399536 995256
rect 475488 990826 475516 995452
rect 475384 990820 475436 990826
rect 475384 990762 475436 990768
rect 475476 990820 475528 990826
rect 475476 990762 475528 990768
rect 475396 990554 475424 990762
rect 475488 990690 475516 990762
rect 475476 990684 475528 990690
rect 475476 990626 475528 990632
rect 476132 990554 476160 995452
rect 476777 995407 476833 995887
rect 477329 995407 477385 995887
rect 477973 995407 478029 995887
rect 478617 995407 478673 995887
rect 479169 995407 479225 995887
rect 479813 995407 479869 995887
rect 480456 995314 480484 995452
rect 481101 995407 481157 995887
rect 481653 995407 481709 995887
rect 482297 995407 482353 995887
rect 482941 995407 482997 995887
rect 484137 995407 484193 995887
rect 485333 995407 485389 995887
rect 485977 995407 486033 995887
rect 486634 995438 486740 995466
rect 480444 995308 480496 995314
rect 480444 995250 480496 995256
rect 486712 990622 486740 995438
rect 487817 995407 487873 995887
rect 488460 995314 488488 995452
rect 525049 995407 525105 995887
rect 525693 995407 525749 995887
rect 526337 995407 526393 995887
rect 488448 995308 488500 995314
rect 488448 995250 488500 995256
rect 526916 990826 526944 995452
rect 526904 990820 526956 990826
rect 526904 990762 526956 990768
rect 527560 990758 527588 995452
rect 528177 995407 528233 995887
rect 528729 995407 528785 995887
rect 529373 995407 529429 995887
rect 530017 995407 530073 995887
rect 530569 995407 530625 995887
rect 531213 995407 531269 995887
rect 531964 995648 532016 995654
rect 531964 995590 532016 995596
rect 531976 995466 532004 995590
rect 531898 995438 532004 995466
rect 532501 995407 532557 995887
rect 533053 995407 533109 995887
rect 533697 995407 533753 995887
rect 534341 995407 534397 995887
rect 535537 995407 535593 995887
rect 536733 995407 536789 995887
rect 537377 995407 537433 995887
rect 537864 995438 538062 995466
rect 488448 990752 488500 990758
rect 488368 990700 488448 990706
rect 488368 990694 488500 990700
rect 527548 990752 527600 990758
rect 527548 990694 527600 990700
rect 488368 990678 488488 990694
rect 486700 990616 486752 990622
rect 486700 990558 486752 990564
rect 475384 990548 475436 990554
rect 475384 990490 475436 990496
rect 476120 990548 476172 990554
rect 476120 990490 476172 990496
rect 353208 990480 353260 990486
rect 353392 990480 353444 990486
rect 353260 990428 353392 990434
rect 364340 990480 364392 990486
rect 353208 990422 353444 990428
rect 364338 990448 364340 990457
rect 397644 990480 397696 990486
rect 364392 990448 364394 990457
rect 353220 990406 353432 990422
rect 364338 990383 364394 990392
rect 383566 990448 383622 990457
rect 397644 990422 397696 990428
rect 405648 990480 405700 990486
rect 405648 990422 405700 990428
rect 383566 990383 383622 990392
rect 383580 990350 383608 990383
rect 397656 990350 397684 990422
rect 405660 990350 405688 990422
rect 430500 990418 430620 990434
rect 469140 990418 469260 990434
rect 424968 990412 425020 990418
rect 424968 990354 425020 990360
rect 430488 990412 430632 990418
rect 430540 990406 430580 990412
rect 430488 990354 430540 990360
rect 430580 990354 430632 990360
rect 463608 990412 463660 990418
rect 463608 990354 463660 990360
rect 469128 990412 469272 990418
rect 469180 990406 469220 990412
rect 469128 990354 469180 990360
rect 469220 990354 469272 990360
rect 471980 990412 472032 990418
rect 471980 990354 472032 990360
rect 383568 990344 383620 990350
rect 383568 990286 383620 990292
rect 397644 990344 397696 990350
rect 397644 990286 397696 990292
rect 405648 990344 405700 990350
rect 424980 990321 425008 990354
rect 444380 990344 444432 990350
rect 405648 990286 405700 990292
rect 405738 990312 405794 990321
rect 405738 990247 405740 990256
rect 405792 990247 405794 990256
rect 424966 990312 425022 990321
rect 424966 990247 425022 990256
rect 444378 990312 444380 990321
rect 463620 990321 463648 990354
rect 444432 990312 444434 990321
rect 444378 990247 444434 990256
rect 463606 990312 463662 990321
rect 471992 990282 472020 990354
rect 486712 990282 486740 990558
rect 488368 990554 488396 990678
rect 537864 990554 537892 995438
rect 539217 995407 539273 995887
rect 539692 995648 539744 995654
rect 539692 995590 539744 995596
rect 539704 995466 539732 995590
rect 539704 995438 539902 995466
rect 585060 992254 585088 997455
rect 589568 992322 589596 997455
rect 626849 995407 626905 995887
rect 627493 995407 627549 995887
rect 628137 995407 628193 995887
rect 628668 995438 628717 995466
rect 629312 995438 629361 995466
rect 589556 992316 589608 992322
rect 589556 992258 589608 992264
rect 585048 992248 585100 992254
rect 585048 992190 585100 992196
rect 545960 990826 546448 990842
rect 628668 990826 628696 995438
rect 545948 990820 546460 990826
rect 546000 990814 546408 990820
rect 545948 990762 546000 990768
rect 546408 990762 546460 990768
rect 628656 990820 628708 990826
rect 628656 990762 628708 990768
rect 563058 990720 563114 990729
rect 546316 990684 546368 990690
rect 563058 990655 563060 990664
rect 546316 990626 546368 990632
rect 563112 990655 563114 990664
rect 582286 990720 582342 990729
rect 582286 990655 582342 990664
rect 563060 990626 563112 990632
rect 488356 990548 488408 990554
rect 488356 990490 488408 990496
rect 537852 990548 537904 990554
rect 537852 990490 537904 990496
rect 546328 990486 546356 990626
rect 582300 990622 582328 990655
rect 582288 990616 582340 990622
rect 587992 990616 588044 990622
rect 582288 990558 582340 990564
rect 585138 990584 585194 990593
rect 585138 990519 585140 990528
rect 585192 990519 585194 990528
rect 587990 990584 587992 990593
rect 623688 990616 623740 990622
rect 588044 990584 588046 990593
rect 623740 990564 623912 990570
rect 623688 990558 623912 990564
rect 623700 990554 623912 990558
rect 623700 990548 623924 990554
rect 623700 990542 623872 990548
rect 587990 990519 588046 990528
rect 585140 990490 585192 990496
rect 623872 990490 623924 990496
rect 546316 990480 546368 990486
rect 546316 990422 546368 990428
rect 463606 990247 463662 990256
rect 471980 990276 472032 990282
rect 405740 990218 405792 990224
rect 471980 990218 472032 990224
rect 486700 990276 486752 990282
rect 486700 990218 486752 990224
rect 628668 990146 628696 990762
rect 629312 990758 629340 995438
rect 629977 995407 630033 995887
rect 630529 995407 630585 995887
rect 631173 995407 631229 995887
rect 631817 995407 631873 995887
rect 632369 995407 632425 995887
rect 633013 995407 633069 995887
rect 633808 995512 633860 995518
rect 633685 995460 633808 995466
rect 633685 995454 633860 995460
rect 633685 995438 633848 995454
rect 634301 995407 634357 995887
rect 634853 995407 634909 995887
rect 635497 995407 635553 995887
rect 636141 995407 636197 995887
rect 637337 995407 637393 995887
rect 638533 995407 638589 995887
rect 639177 995407 639233 995887
rect 639800 995438 639849 995466
rect 629300 990752 629352 990758
rect 629300 990694 629352 990700
rect 629312 990146 629340 990694
rect 639800 990554 639828 995438
rect 641017 995407 641073 995887
rect 641536 995512 641588 995518
rect 641588 995460 641689 995466
rect 641536 995454 641689 995460
rect 641548 995438 641689 995454
rect 674748 992316 674800 992322
rect 674748 992258 674800 992264
rect 639788 990548 639840 990554
rect 639788 990490 639840 990496
rect 639800 990214 639828 990490
rect 639788 990208 639840 990214
rect 639788 990150 639840 990156
rect 673644 990208 673696 990214
rect 673644 990150 673696 990156
rect 78864 990140 78916 990146
rect 78864 990082 78916 990088
rect 88340 990140 88392 990146
rect 88340 990082 88392 990088
rect 325700 990140 325752 990146
rect 325700 990082 325752 990088
rect 343732 990140 343784 990146
rect 343732 990082 343784 990088
rect 628656 990140 628708 990146
rect 628656 990082 628708 990088
rect 629300 990140 629352 990146
rect 629300 990082 629352 990088
rect 673552 990140 673604 990146
rect 673552 990082 673604 990088
rect 673460 990072 673512 990078
rect 673460 990014 673512 990020
rect 673472 964374 673500 990014
rect 673460 964368 673512 964374
rect 673460 964310 673512 964316
rect 44086 877568 44142 877577
rect 44086 877503 44142 877512
rect 673472 875838 673500 964310
rect 673564 963762 673592 990082
rect 673552 963756 673604 963762
rect 673552 963698 673604 963704
rect 673564 910790 673592 963698
rect 673656 953902 673684 990150
rect 674656 966068 674708 966074
rect 674656 966010 674708 966016
rect 673644 953896 673696 953902
rect 673644 953838 673696 953844
rect 673552 910784 673604 910790
rect 673552 910726 673604 910732
rect 673460 875832 673512 875838
rect 673460 875774 673512 875780
rect 44362 870088 44418 870097
rect 44362 870023 44418 870032
rect 42522 869408 42578 869417
rect 42522 869343 42578 869352
rect 42706 869408 42762 869417
rect 42706 869343 42762 869352
rect 42720 850134 42748 869343
rect 42524 850128 42576 850134
rect 42524 850070 42576 850076
rect 42708 850128 42760 850134
rect 42708 850070 42760 850076
rect 42536 836210 42564 850070
rect 44376 836330 44404 870023
rect 44180 836324 44232 836330
rect 44180 836266 44232 836272
rect 44364 836324 44416 836330
rect 44364 836266 44416 836272
rect 42536 836182 42748 836210
rect 42444 807350 42656 807378
rect 42432 799604 42484 799610
rect 42432 799546 42484 799552
rect 42444 792606 42472 799546
rect 42432 792600 42484 792606
rect 42432 792542 42484 792548
rect 42628 787914 42656 807350
rect 42720 798726 42748 836182
rect 42708 798720 42760 798726
rect 42708 798662 42760 798668
rect 42720 798266 42748 798662
rect 42720 798238 42932 798266
rect 42904 792130 42932 798238
rect 42892 792124 42944 792130
rect 42892 792066 42944 792072
rect 43076 792124 43128 792130
rect 43076 792066 43128 792072
rect 42432 787908 42484 787914
rect 42432 787850 42484 787856
rect 42616 787908 42668 787914
rect 42616 787850 42668 787856
rect 42444 756566 42472 787850
rect 42616 786684 42668 786690
rect 42616 786626 42668 786632
rect 42432 756560 42484 756566
rect 42432 756502 42484 756508
rect 42432 756424 42484 756430
rect 42432 756366 42484 756372
rect 42444 749426 42472 756366
rect 42432 749420 42484 749426
rect 42432 749362 42484 749368
rect 42432 745136 42484 745142
rect 42432 745078 42484 745084
rect 42444 730862 42472 745078
rect 42628 744462 42656 786626
rect 43088 772886 43116 792066
rect 42800 772880 42852 772886
rect 42800 772822 42852 772828
rect 43076 772880 43128 772886
rect 43076 772822 43128 772828
rect 42812 758962 42840 772822
rect 42720 758934 42840 758962
rect 42720 754458 42748 758934
rect 42800 756560 42852 756566
rect 42800 756502 42852 756508
rect 42708 754452 42760 754458
rect 42708 754394 42760 754400
rect 42616 744456 42668 744462
rect 42616 744398 42668 744404
rect 42432 730856 42484 730862
rect 42432 730798 42484 730804
rect 42432 713176 42484 713182
rect 42432 713118 42484 713124
rect 42444 706246 42472 713118
rect 42524 708756 42576 708762
rect 42524 708698 42576 708704
rect 42432 706240 42484 706246
rect 42432 706182 42484 706188
rect 42536 700942 42564 708698
rect 42524 700936 42576 700942
rect 42524 700878 42576 700884
rect 42628 700602 42656 744398
rect 42720 731082 42748 754394
rect 42812 745142 42840 756502
rect 42800 745136 42852 745142
rect 42800 745078 42852 745084
rect 44192 739634 44220 836266
rect 44270 835272 44326 835281
rect 44270 835207 44326 835216
rect 44180 739628 44232 739634
rect 44180 739570 44232 739576
rect 42720 731054 43024 731082
rect 42800 730856 42852 730862
rect 42800 730798 42852 730804
rect 42812 708762 42840 730798
rect 42892 711272 42944 711278
rect 42996 711226 43024 731054
rect 44180 720452 44232 720458
rect 44180 720394 44232 720400
rect 42944 711220 43024 711226
rect 42892 711214 43024 711220
rect 42904 711198 43024 711214
rect 42800 708756 42852 708762
rect 42800 708698 42852 708704
rect 42708 700936 42760 700942
rect 42708 700878 42760 700884
rect 42616 700596 42668 700602
rect 42616 700538 42668 700544
rect 42628 698850 42656 700538
rect 42536 698822 42656 698850
rect 42432 669996 42484 670002
rect 42432 669938 42484 669944
rect 42444 663066 42472 669938
rect 42432 663060 42484 663066
rect 42432 663002 42484 663008
rect 42536 657150 42564 698822
rect 42616 669112 42668 669118
rect 42616 669054 42668 669060
rect 42524 657144 42576 657150
rect 42524 657086 42576 657092
rect 42524 633412 42576 633418
rect 42524 633354 42576 633360
rect 42432 626816 42484 626822
rect 42432 626758 42484 626764
rect 42444 619818 42472 626758
rect 42536 623642 42564 633354
rect 42628 630170 42656 669054
rect 42720 668794 42748 700878
rect 42904 695502 42932 711198
rect 44192 701049 44220 720394
rect 44178 701040 44234 701049
rect 44178 700975 44234 700984
rect 42892 695496 42944 695502
rect 42892 695438 42944 695444
rect 43076 695496 43128 695502
rect 43076 695438 43128 695444
rect 43088 681442 43116 695438
rect 44180 681760 44232 681766
rect 44180 681702 44232 681708
rect 42904 681414 43116 681442
rect 42904 669118 42932 681414
rect 42892 669112 42944 669118
rect 42892 669054 42944 669060
rect 42720 668766 43024 668794
rect 42996 657694 43024 668766
rect 44192 662425 44220 681702
rect 44178 662416 44234 662425
rect 44178 662351 44234 662360
rect 42708 657688 42760 657694
rect 42984 657688 43036 657694
rect 42760 657636 42840 657642
rect 42708 657630 42840 657636
rect 42984 657630 43036 657636
rect 42720 657614 42840 657630
rect 42708 657144 42760 657150
rect 42708 657086 42760 657092
rect 42720 633418 42748 657086
rect 42708 633412 42760 633418
rect 42708 633354 42760 633360
rect 42628 630142 42748 630170
rect 42720 625938 42748 630142
rect 42708 625932 42760 625938
rect 42708 625874 42760 625880
rect 42536 623614 42656 623642
rect 42432 619812 42484 619818
rect 42432 619754 42484 619760
rect 42432 614440 42484 614446
rect 42432 614382 42484 614388
rect 42444 583710 42472 614382
rect 42628 614106 42656 623614
rect 42720 618254 42748 625874
rect 42708 618248 42760 618254
rect 42708 618190 42760 618196
rect 42812 614446 42840 657614
rect 44180 643136 44232 643142
rect 44180 643078 44232 643084
rect 44192 623694 44220 643078
rect 44180 623688 44232 623694
rect 44180 623630 44232 623636
rect 42984 618248 43036 618254
rect 42984 618190 43036 618196
rect 42800 614440 42852 614446
rect 42800 614382 42852 614388
rect 42616 614100 42668 614106
rect 42616 614042 42668 614048
rect 42432 583704 42484 583710
rect 42432 583646 42484 583652
rect 42432 583568 42484 583574
rect 42432 583510 42484 583516
rect 42444 576638 42472 583510
rect 42432 576632 42484 576638
rect 42432 576574 42484 576580
rect 42432 572280 42484 572286
rect 42432 572222 42484 572228
rect 42444 556170 42472 572222
rect 42628 571674 42656 614042
rect 42800 583704 42852 583710
rect 42800 583646 42852 583652
rect 42708 581664 42760 581670
rect 42708 581606 42760 581612
rect 42616 571668 42668 571674
rect 42616 571610 42668 571616
rect 42432 556164 42484 556170
rect 42432 556106 42484 556112
rect 42432 540388 42484 540394
rect 42432 540330 42484 540336
rect 42444 533458 42472 540330
rect 42432 533452 42484 533458
rect 42432 533394 42484 533400
rect 42432 529100 42484 529106
rect 42432 529042 42484 529048
rect 42444 498234 42472 529042
rect 42628 527814 42656 571610
rect 42720 538558 42748 581606
rect 42812 572286 42840 583646
rect 42996 581670 43024 618190
rect 44180 604512 44232 604518
rect 44180 604454 44232 604460
rect 44192 585070 44220 604454
rect 44180 585064 44232 585070
rect 44180 585006 44232 585012
rect 42984 581664 43036 581670
rect 42984 581606 43036 581612
rect 42800 572280 42852 572286
rect 42800 572222 42852 572228
rect 44180 565888 44232 565894
rect 44180 565830 44232 565836
rect 44192 564330 44220 565830
rect 44180 564324 44232 564330
rect 44180 564266 44232 564272
rect 42800 556164 42852 556170
rect 42800 556106 42852 556112
rect 42708 538552 42760 538558
rect 42708 538494 42760 538500
rect 42616 527808 42668 527814
rect 42616 527750 42668 527756
rect 42432 498228 42484 498234
rect 42432 498170 42484 498176
rect 42432 478916 42484 478922
rect 42432 478858 42484 478864
rect 42444 469198 42472 478858
rect 42432 469192 42484 469198
rect 42432 469134 42484 469140
rect 42628 463690 42656 527750
rect 42616 463684 42668 463690
rect 42616 463626 42668 463632
rect 42338 448624 42394 448633
rect 42338 448559 42394 448568
rect 42062 444408 42118 444417
rect 42062 444343 42118 444352
rect 42614 444408 42670 444417
rect 42614 444343 42670 444352
rect 42076 442746 42104 444343
rect 42064 442740 42116 442746
rect 42064 442682 42116 442688
rect 42340 442740 42392 442746
rect 42340 442682 42392 442688
rect 39592 440830 39988 440858
rect 42352 425066 42380 442682
rect 42628 441590 42656 444343
rect 42432 441584 42484 441590
rect 42432 441526 42484 441532
rect 42616 441584 42668 441590
rect 42616 441526 42668 441532
rect 42340 425060 42392 425066
rect 42340 425002 42392 425008
rect 42444 422346 42472 441526
rect 42432 422340 42484 422346
rect 42432 422282 42484 422288
rect 42524 422340 42576 422346
rect 42524 422282 42576 422288
rect 41722 413275 42288 413303
rect 41713 412617 42193 412673
rect 41722 411454 41828 411482
rect 41800 411126 41828 411454
rect 41788 411120 41840 411126
rect 41788 411062 41840 411068
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 42260 405770 42288 413275
rect 42536 411330 42564 422282
rect 42524 411324 42576 411330
rect 42524 411266 42576 411272
rect 42432 411256 42484 411262
rect 42432 411198 42484 411204
rect 41892 405742 42288 405770
rect 41892 405299 41920 405742
rect 41722 405271 41920 405299
rect 41713 404613 42193 404669
rect 41713 403969 42193 404025
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41788 401396 41840 401402
rect 41788 401338 41840 401344
rect 41800 400975 41828 401338
rect 41722 400947 41828 400975
rect 42444 400466 42472 411198
rect 42720 411126 42748 538494
rect 42812 529106 42840 556106
rect 42800 529100 42852 529106
rect 42800 529042 42852 529048
rect 44180 527196 44232 527202
rect 44180 527138 44232 527144
rect 44192 507754 44220 527138
rect 44180 507748 44232 507754
rect 44180 507690 44232 507696
rect 44284 493241 44312 835207
rect 44548 827552 44600 827558
rect 44548 827494 44600 827500
rect 44560 806002 44588 827494
rect 44364 805996 44416 806002
rect 44364 805938 44416 805944
rect 44548 805996 44600 806002
rect 44548 805938 44600 805944
rect 44376 786570 44404 805938
rect 673472 786962 673500 875774
rect 673564 874886 673592 910726
rect 673552 874880 673604 874886
rect 673552 874822 673604 874828
rect 673460 786956 673512 786962
rect 673460 786898 673512 786904
rect 44376 786542 44588 786570
rect 44560 767378 44588 786542
rect 673564 786418 673592 874822
rect 673656 865026 673684 953838
rect 674668 932890 674696 966010
rect 674656 932884 674708 932890
rect 674656 932826 674708 932832
rect 674656 902556 674708 902562
rect 674656 902498 674708 902504
rect 674668 894266 674696 902498
rect 674656 894260 674708 894266
rect 674656 894202 674708 894208
rect 673644 865020 673696 865026
rect 673644 864962 673696 864968
rect 673552 786412 673604 786418
rect 673552 786354 673604 786360
rect 44364 767372 44416 767378
rect 44364 767314 44416 767320
rect 44548 767372 44600 767378
rect 44548 767314 44600 767320
rect 44270 493232 44326 493241
rect 44270 493167 44326 493176
rect 44376 488617 44404 767314
rect 673564 746570 673592 786354
rect 673656 774926 673684 864962
rect 674760 823478 674788 992258
rect 675208 992248 675260 992254
rect 675208 992190 675260 992196
rect 675220 990842 675248 992190
rect 675128 990814 675248 990842
rect 675128 985318 675156 990814
rect 674840 985312 674892 985318
rect 674840 985254 674892 985260
rect 675116 985312 675168 985318
rect 675116 985254 675168 985260
rect 674852 966074 674880 985254
rect 675407 966695 675887 966751
rect 674840 966068 674892 966074
rect 675407 966051 675887 966107
rect 674840 966010 674892 966016
rect 675407 965407 675887 965463
rect 675404 964374 675432 964883
rect 675392 964368 675444 964374
rect 675392 964310 675444 964316
rect 675404 963762 675432 964239
rect 675392 963756 675444 963762
rect 675392 963698 675444 963704
rect 675407 963567 675887 963623
rect 675407 963015 675887 963071
rect 675407 962371 675887 962427
rect 675407 961727 675887 961783
rect 675407 961175 675887 961231
rect 675407 960531 675887 960587
rect 675312 959901 675418 959929
rect 675312 951810 675340 959901
rect 675407 959243 675887 959299
rect 675407 958691 675887 958747
rect 675407 958047 675887 958103
rect 675407 957403 675887 957459
rect 675407 956207 675887 956263
rect 675407 955011 675887 955067
rect 675407 954367 675887 954423
rect 675392 953896 675444 953902
rect 675392 953838 675444 953844
rect 675404 953751 675432 953838
rect 675407 952527 675887 952583
rect 675404 951810 675432 951932
rect 675312 951782 675432 951810
rect 674840 932816 674892 932822
rect 674840 932758 674892 932764
rect 674852 902630 674880 932758
rect 677796 918598 678086 918626
rect 677690 918368 677746 918377
rect 677690 918303 677746 918312
rect 677506 915376 677562 915385
rect 677506 915311 677562 915320
rect 677520 912801 677548 915311
rect 677506 912792 677562 912801
rect 677506 912727 677562 912736
rect 677520 908177 677548 912727
rect 677506 908168 677562 908177
rect 675300 908132 675352 908138
rect 677506 908103 677508 908112
rect 675300 908074 675352 908080
rect 677560 908103 677562 908112
rect 677508 908074 677560 908080
rect 674840 902624 674892 902630
rect 674840 902566 674892 902572
rect 674840 894260 674892 894266
rect 674840 894202 674892 894208
rect 674852 874970 674880 894202
rect 674852 874942 674972 874970
rect 674944 874834 674972 874942
rect 674944 874806 675064 874834
rect 675036 855658 675064 874806
rect 675208 870188 675260 870194
rect 675208 870130 675260 870136
rect 675220 862730 675248 870130
rect 675312 862850 675340 908074
rect 677704 907746 677732 918303
rect 677796 909401 677824 918598
rect 677888 913838 678046 913866
rect 677888 910790 677916 913838
rect 678018 913716 678046 913838
rect 677876 910784 677928 910790
rect 677876 910726 677928 910732
rect 677782 909392 677838 909401
rect 677782 909327 677838 909336
rect 677704 907718 678086 907746
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675392 875832 675444 875838
rect 675392 875774 675444 875780
rect 675404 875683 675432 875774
rect 675404 874886 675432 875039
rect 675392 874880 675444 874886
rect 675392 874822 675444 874828
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 871975 675887 872031
rect 675407 871331 675887 871387
rect 675404 870194 675432 870740
rect 675392 870188 675444 870194
rect 675392 870130 675444 870136
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675392 865020 675444 865026
rect 675392 864962 675444 864968
rect 675404 864551 675432 864962
rect 675407 863327 675887 863383
rect 675300 862844 675352 862850
rect 675300 862786 675352 862792
rect 675220 862702 675418 862730
rect 675300 862640 675352 862646
rect 675300 862582 675352 862588
rect 675036 855630 675156 855658
rect 675128 836330 675156 855630
rect 674932 836324 674984 836330
rect 674932 836266 674984 836272
rect 675116 836324 675168 836330
rect 675116 836266 675168 836272
rect 674944 827966 674972 836266
rect 674932 827960 674984 827966
rect 674932 827902 674984 827908
rect 674748 823472 674800 823478
rect 674748 823414 674800 823420
rect 674944 816898 674972 827902
rect 675208 818712 675260 818718
rect 675208 818654 675260 818660
rect 674944 816870 675064 816898
rect 675036 797722 675064 816870
rect 675036 797694 675156 797722
rect 675128 792130 675156 797694
rect 674840 792124 674892 792130
rect 674840 792066 674892 792072
rect 675116 792124 675168 792130
rect 675116 792066 675168 792072
rect 673736 786956 673788 786962
rect 673736 786898 673788 786904
rect 673644 774920 673696 774926
rect 673644 774862 673696 774868
rect 673552 746564 673604 746570
rect 673552 746506 673604 746512
rect 673748 741946 673776 786898
rect 673920 774920 673972 774926
rect 673920 774862 673972 774868
rect 673736 741940 673788 741946
rect 673736 741882 673788 741888
rect 44456 739628 44508 739634
rect 44456 739570 44508 739576
rect 44468 720458 44496 739570
rect 673552 730176 673604 730182
rect 673552 730118 673604 730124
rect 44456 720452 44508 720458
rect 44456 720394 44508 720400
rect 44454 701040 44510 701049
rect 44454 700975 44510 700984
rect 44468 681766 44496 700975
rect 673460 695972 673512 695978
rect 673460 695914 673512 695920
rect 44456 681760 44508 681766
rect 44456 681702 44508 681708
rect 44454 662416 44510 662425
rect 44454 662351 44510 662360
rect 44468 643142 44496 662351
rect 673472 651778 673500 695914
rect 673564 685234 673592 730118
rect 673644 730040 673696 730046
rect 673644 729982 673696 729988
rect 673656 695366 673684 729982
rect 673748 695978 673776 741882
rect 673932 730182 673960 774862
rect 674852 772834 674880 792066
rect 675024 781040 675076 781046
rect 675024 780982 675076 780988
rect 675036 774042 675064 780982
rect 675024 774036 675076 774042
rect 675024 773978 675076 773984
rect 674760 772806 674880 772834
rect 674760 758962 674788 772806
rect 674760 758934 675064 758962
rect 674012 746564 674064 746570
rect 674012 746506 674064 746512
rect 674024 740722 674052 746506
rect 675036 741497 675064 758934
rect 674944 741469 675064 741497
rect 674012 740716 674064 740722
rect 674012 740658 674064 740664
rect 673920 730176 673972 730182
rect 673920 730118 673972 730124
rect 674024 730046 674052 740658
rect 674944 739634 674972 741469
rect 674840 739628 674892 739634
rect 674840 739570 674892 739576
rect 674932 739628 674984 739634
rect 674932 739570 674984 739576
rect 674852 734126 674880 739570
rect 675024 736024 675076 736030
rect 675024 735966 675076 735972
rect 674840 734120 674892 734126
rect 674840 734062 674892 734068
rect 674932 734120 674984 734126
rect 674932 734062 674984 734068
rect 674012 730040 674064 730046
rect 674012 729982 674064 729988
rect 674944 728634 674972 734062
rect 675036 729094 675064 735966
rect 675024 729088 675076 729094
rect 675024 729030 675076 729036
rect 674944 728606 675064 728634
rect 675036 714814 675064 728606
rect 674840 714808 674892 714814
rect 674840 714750 674892 714756
rect 675024 714808 675076 714814
rect 675024 714750 675076 714756
rect 673736 695972 673788 695978
rect 673736 695914 673788 695920
rect 674852 695570 674880 714750
rect 674840 695564 674892 695570
rect 674840 695506 674892 695512
rect 675116 695564 675168 695570
rect 675116 695506 675168 695512
rect 673644 695360 673696 695366
rect 673644 695302 673696 695308
rect 673552 685228 673604 685234
rect 673552 685170 673604 685176
rect 673460 651772 673512 651778
rect 673460 651714 673512 651720
rect 44456 643136 44508 643142
rect 44456 643078 44508 643084
rect 44456 623688 44508 623694
rect 44456 623630 44508 623636
rect 44468 604518 44496 623630
rect 673472 606762 673500 651714
rect 673564 639742 673592 685170
rect 673656 651166 673684 695302
rect 675024 691688 675076 691694
rect 675024 691630 675076 691636
rect 675036 684078 675064 691630
rect 675024 684072 675076 684078
rect 675024 684014 675076 684020
rect 675128 681850 675156 695506
rect 674944 681822 675156 681850
rect 674944 681714 674972 681822
rect 674944 681686 675064 681714
rect 675036 676190 675064 681686
rect 674840 676184 674892 676190
rect 674840 676126 674892 676132
rect 675024 676184 675076 676190
rect 675024 676126 675076 676132
rect 674852 656946 674880 676126
rect 674840 656940 674892 656946
rect 674840 656882 674892 656888
rect 675116 656940 675168 656946
rect 675116 656882 675168 656888
rect 673644 651160 673696 651166
rect 673644 651102 673696 651108
rect 673552 639736 673604 639742
rect 673552 639678 673604 639684
rect 673564 623762 673592 639678
rect 673552 623756 673604 623762
rect 673552 623698 673604 623704
rect 673460 606756 673512 606762
rect 673460 606698 673512 606704
rect 673656 605538 673684 651102
rect 675024 645788 675076 645794
rect 675024 645730 675076 645736
rect 675036 638858 675064 645730
rect 675024 638852 675076 638858
rect 675024 638794 675076 638800
rect 675128 637634 675156 656882
rect 674748 637628 674800 637634
rect 674748 637570 674800 637576
rect 675116 637628 675168 637634
rect 675116 637570 675168 637576
rect 674760 623830 674788 637570
rect 674748 623824 674800 623830
rect 674748 623766 674800 623772
rect 673828 623688 673880 623694
rect 673828 623630 673880 623636
rect 674932 623688 674984 623694
rect 674932 623630 674984 623636
rect 673644 605532 673696 605538
rect 673644 605474 673696 605480
rect 673656 604518 673684 605474
rect 44456 604512 44508 604518
rect 44456 604454 44508 604460
rect 673644 604512 673696 604518
rect 673644 604454 673696 604460
rect 673840 594930 673868 623630
rect 674944 618254 674972 623630
rect 674564 618248 674616 618254
rect 674564 618190 674616 618196
rect 674932 618248 674984 618254
rect 674932 618190 674984 618196
rect 673920 604512 673972 604518
rect 673920 604454 673972 604460
rect 673644 594924 673696 594930
rect 673644 594866 673696 594872
rect 673828 594924 673880 594930
rect 673828 594866 673880 594872
rect 44456 585064 44508 585070
rect 44456 585006 44508 585012
rect 44468 565894 44496 585006
rect 44456 565888 44508 565894
rect 44456 565830 44508 565836
rect 44456 564324 44508 564330
rect 44456 564266 44508 564272
rect 44468 527202 44496 564266
rect 673656 550526 673684 594866
rect 673828 561264 673880 561270
rect 673828 561206 673880 561212
rect 673644 550520 673696 550526
rect 673644 550462 673696 550468
rect 44456 527196 44508 527202
rect 44456 527138 44508 527144
rect 673840 527082 673868 561206
rect 673932 560998 673960 604454
rect 674576 599078 674604 618190
rect 674748 606756 674800 606762
rect 674748 606698 674800 606704
rect 674564 599072 674616 599078
rect 674564 599014 674616 599020
rect 674760 598942 674788 606698
rect 675116 600840 675168 600846
rect 675116 600782 675168 600788
rect 674840 599072 674892 599078
rect 674840 599014 674892 599020
rect 674852 598942 674880 599014
rect 674656 598936 674708 598942
rect 674656 598878 674708 598884
rect 674748 598936 674800 598942
rect 674748 598878 674800 598884
rect 674840 598936 674892 598942
rect 674840 598878 674892 598884
rect 675024 598936 675076 598942
rect 675024 598878 675076 598884
rect 674668 589234 674696 598878
rect 675036 593586 675064 598878
rect 675128 593842 675156 600782
rect 675116 593836 675168 593842
rect 675116 593778 675168 593784
rect 675036 593558 675156 593586
rect 674668 589206 674788 589234
rect 674656 579624 674708 579630
rect 674656 579566 674708 579572
rect 673920 560992 673972 560998
rect 673920 560934 673972 560940
rect 674668 560318 674696 579566
rect 674760 561270 674788 589206
rect 675128 579714 675156 593558
rect 675036 579686 675156 579714
rect 675036 579630 675064 579686
rect 675024 579624 675076 579630
rect 675024 579566 675076 579572
rect 674748 561264 674800 561270
rect 674748 561206 674800 561212
rect 674656 560312 674708 560318
rect 674656 560254 674708 560260
rect 674840 560312 674892 560318
rect 674840 560254 674892 560260
rect 674852 541006 674880 560254
rect 675116 555620 675168 555626
rect 675116 555562 675168 555568
rect 675128 548690 675156 555562
rect 675116 548684 675168 548690
rect 675116 548626 675168 548632
rect 674840 541000 674892 541006
rect 674840 540942 674892 540948
rect 675024 541000 675076 541006
rect 675024 540942 675076 540948
rect 675036 531298 675064 540942
rect 674944 531270 675064 531298
rect 673840 527054 674052 527082
rect 44456 507748 44508 507754
rect 44456 507690 44508 507696
rect 44362 488608 44418 488617
rect 44180 488572 44232 488578
rect 44468 488578 44496 507690
rect 674024 492674 674052 527054
rect 674944 514078 674972 531270
rect 674932 514072 674984 514078
rect 674932 514014 674984 514020
rect 675220 513806 675248 818654
rect 675208 513800 675260 513806
rect 675208 513742 675260 513748
rect 673932 492646 674052 492674
rect 44362 488543 44418 488552
rect 44456 488572 44508 488578
rect 44180 488514 44232 488520
rect 44456 488514 44508 488520
rect 44192 488458 44220 488514
rect 44192 488430 44312 488458
rect 44284 488322 44312 488430
rect 44284 488294 44404 488322
rect 42892 463684 42944 463690
rect 42892 463626 42944 463632
rect 42904 444417 42932 463626
rect 44376 449954 44404 488294
rect 673932 469282 673960 492646
rect 673840 469254 673960 469282
rect 673840 463690 673868 469254
rect 675312 467566 675340 862582
rect 677612 827966 677640 828580
rect 677600 827960 677652 827966
rect 677600 827902 677652 827908
rect 676128 823472 676180 823478
rect 676128 823414 676180 823420
rect 676140 818718 676168 823414
rect 676128 818712 676180 818718
rect 676128 818654 676180 818660
rect 677416 818712 677468 818718
rect 677598 818680 677654 818689
rect 677468 818660 677598 818666
rect 677416 818654 677598 818660
rect 677428 818638 677598 818654
rect 677598 818615 677654 818624
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 675392 786956 675444 786962
rect 675392 786898 675444 786904
rect 675404 786483 675432 786898
rect 675392 786412 675444 786418
rect 675392 786354 675444 786360
rect 675404 785839 675432 786354
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 782775 675887 782831
rect 675407 782131 675887 782187
rect 675404 781046 675432 781524
rect 675392 781040 675444 781046
rect 675392 780982 675444 780988
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675404 774926 675432 775351
rect 675392 774920 675444 774926
rect 675392 774862 675444 774868
rect 675407 774127 675887 774183
rect 675392 774036 675444 774042
rect 675392 773978 675444 773984
rect 675404 773500 675432 773978
rect 675407 743295 675887 743351
rect 675407 742651 675887 742707
rect 675407 742007 675887 742063
rect 675392 741940 675444 741946
rect 675392 741882 675444 741888
rect 675404 741483 675432 741882
rect 675404 740722 675432 740860
rect 675392 740716 675444 740722
rect 675392 740658 675444 740664
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 737775 675887 737831
rect 675407 737131 675887 737187
rect 675404 736030 675432 736508
rect 675392 736024 675444 736030
rect 675392 735966 675444 735972
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675404 730182 675432 730351
rect 675392 730176 675444 730182
rect 675392 730118 675444 730124
rect 675407 729127 675887 729183
rect 675392 729088 675444 729094
rect 675392 729030 675444 729036
rect 675404 728484 675432 729030
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675404 695978 675432 696483
rect 675392 695972 675444 695978
rect 675392 695914 675444 695920
rect 675404 695366 675432 695844
rect 675392 695360 675444 695366
rect 675392 695302 675444 695308
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 692775 675887 692831
rect 675407 692131 675887 692187
rect 675392 691688 675444 691694
rect 675392 691630 675444 691636
rect 675404 691492 675432 691630
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675404 685234 675432 685372
rect 675392 685228 675444 685234
rect 675392 685170 675444 685176
rect 675407 684127 675887 684183
rect 675392 684072 675444 684078
rect 675392 684014 675444 684020
rect 675404 683511 675432 684014
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 675392 651772 675444 651778
rect 675392 651714 675444 651720
rect 675404 651283 675432 651714
rect 675392 651160 675444 651166
rect 675392 651102 675444 651108
rect 675404 650639 675432 651102
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 647575 675887 647631
rect 675407 646931 675887 646987
rect 675404 645794 675432 646340
rect 675392 645788 675444 645794
rect 675392 645730 675444 645736
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675404 639742 675432 640151
rect 675392 639736 675444 639742
rect 675392 639678 675444 639684
rect 675407 638927 675887 638983
rect 675392 638852 675444 638858
rect 675392 638794 675444 638800
rect 675404 638316 675432 638794
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 675392 606756 675444 606762
rect 675392 606698 675444 606704
rect 675404 606283 675432 606698
rect 675404 605538 675432 605639
rect 675392 605532 675444 605538
rect 675392 605474 675444 605480
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 602575 675887 602631
rect 675407 601931 675887 601987
rect 675404 600846 675432 601324
rect 675392 600840 675444 600846
rect 675392 600782 675444 600788
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675404 594930 675432 595151
rect 675392 594924 675444 594930
rect 675392 594866 675444 594872
rect 675407 593927 675887 593983
rect 675392 593836 675444 593842
rect 675392 593778 675444 593784
rect 675404 593300 675432 593778
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 675392 561264 675444 561270
rect 675392 561206 675444 561212
rect 675404 561068 675432 561206
rect 675392 560992 675444 560998
rect 675392 560934 675444 560940
rect 675404 560439 675432 560934
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675407 557375 675887 557431
rect 675407 556731 675887 556787
rect 675404 555626 675432 556115
rect 675392 555620 675444 555626
rect 675392 555562 675444 555568
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675392 550520 675444 550526
rect 675392 550462 675444 550468
rect 675404 549951 675432 550462
rect 675407 548727 675887 548783
rect 675392 548684 675444 548690
rect 675392 548626 675444 548632
rect 675404 548111 675432 548626
rect 676036 514072 676088 514078
rect 676036 514014 676088 514020
rect 677416 514072 677468 514078
rect 677468 514020 677626 514026
rect 677416 514014 677626 514020
rect 675300 467560 675352 467566
rect 675300 467502 675352 467508
rect 673736 463684 673788 463690
rect 673736 463626 673788 463632
rect 673828 463684 673880 463690
rect 673828 463626 673880 463632
rect 44180 449948 44232 449954
rect 44180 449890 44232 449896
rect 44364 449948 44416 449954
rect 44364 449890 44416 449896
rect 44192 449834 44220 449890
rect 673748 449886 673776 463626
rect 673736 449880 673788 449886
rect 44192 449806 44312 449834
rect 673736 449822 673788 449828
rect 673920 449880 673972 449886
rect 673920 449822 673972 449828
rect 42890 444408 42946 444417
rect 42890 444343 42946 444352
rect 44284 430658 44312 449806
rect 673932 444394 673960 449822
rect 673932 444366 674052 444394
rect 674024 430710 674052 444366
rect 674012 430704 674064 430710
rect 44284 430630 44404 430658
rect 674012 430646 674064 430652
rect 42800 425060 42852 425066
rect 42800 425002 42852 425008
rect 42708 411120 42760 411126
rect 42708 411062 42760 411068
rect 42720 404818 42748 411062
rect 41800 400438 42472 400466
rect 41800 400330 41828 400438
rect 41722 400302 41828 400330
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 42156 397860 42208 397866
rect 42156 397802 42208 397808
rect 42168 370258 42196 397802
rect 42444 370394 42472 400438
rect 42536 404790 42748 404818
rect 42432 370388 42484 370394
rect 42432 370330 42484 370336
rect 42156 370252 42208 370258
rect 42156 370194 42208 370200
rect 42432 370252 42484 370258
rect 42432 370194 42484 370200
rect 41722 370075 42288 370103
rect 41713 369417 42193 369473
rect 41722 368235 41828 368263
rect 41800 367742 41828 368235
rect 41788 367736 41840 367742
rect 41788 367678 41840 367684
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 42260 362250 42288 370075
rect 41800 362222 42288 362250
rect 41800 362114 41828 362222
rect 41722 362086 41828 362114
rect 41713 361413 42193 361469
rect 41713 360769 42193 360825
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 42444 358290 42472 370194
rect 42536 367742 42564 404790
rect 42812 401402 42840 425002
rect 44376 411330 44404 430630
rect 673920 430568 673972 430574
rect 673920 430510 673972 430516
rect 44180 411324 44232 411330
rect 44180 411266 44232 411272
rect 44364 411324 44416 411330
rect 44364 411266 44416 411272
rect 42800 401396 42852 401402
rect 42800 401338 42852 401344
rect 42812 397866 42840 401338
rect 42800 397860 42852 397866
rect 42800 397802 42852 397808
rect 44192 391898 44220 411266
rect 673932 411210 673960 430510
rect 676048 427854 676076 514014
rect 677428 513998 677626 514014
rect 676128 513800 676180 513806
rect 677508 513800 677560 513806
rect 676128 513742 676180 513748
rect 677506 513768 677508 513777
rect 677560 513768 677562 513777
rect 676140 507890 676168 513742
rect 677506 513703 677562 513712
rect 677428 507890 677626 507906
rect 676128 507884 676180 507890
rect 676128 507826 676180 507832
rect 677416 507884 677626 507890
rect 677468 507878 677626 507884
rect 677416 507826 677468 507832
rect 676036 427848 676088 427854
rect 676036 427790 676088 427796
rect 676140 420782 676168 507826
rect 678058 477592 678114 477601
rect 678058 477527 678114 477536
rect 678072 470778 678100 477527
rect 677888 470764 678100 470778
rect 677888 470750 678086 470764
rect 677888 469985 677916 470750
rect 677874 469976 677930 469985
rect 677874 469911 677930 469920
rect 677508 467560 677560 467566
rect 677506 467528 677508 467537
rect 677560 467528 677562 467537
rect 677506 467463 677562 467472
rect 677704 465990 678032 466018
rect 677704 460018 677732 465990
rect 676220 460012 676272 460018
rect 676220 459954 676272 459960
rect 677692 460012 677744 460018
rect 677692 459954 677744 459960
rect 676128 420776 676180 420782
rect 676128 420718 676180 420724
rect 673564 411182 673960 411210
rect 673092 408536 673144 408542
rect 673092 408478 673144 408484
rect 44192 391870 44404 391898
rect 44376 372638 44404 391870
rect 44180 372632 44232 372638
rect 44180 372574 44232 372580
rect 44364 372632 44416 372638
rect 44364 372574 44416 372580
rect 42708 370388 42760 370394
rect 42708 370330 42760 370336
rect 42524 367736 42576 367742
rect 42524 367678 42576 367684
rect 41788 358284 41840 358290
rect 41788 358226 41840 358232
rect 42432 358284 42484 358290
rect 42432 358226 42484 358232
rect 41800 357762 41828 358226
rect 41722 357734 41828 357762
rect 41788 357332 41840 357338
rect 41788 357274 41840 357280
rect 41800 357131 41828 357274
rect 41722 357103 41828 357131
rect 42432 356652 42484 356658
rect 42432 356594 42484 356600
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 42340 339652 42392 339658
rect 42340 339594 42392 339600
rect 41722 326862 42288 326890
rect 41713 326217 42193 326273
rect 41722 325035 41828 325063
rect 41800 324562 41828 325035
rect 41788 324556 41840 324562
rect 41788 324498 41840 324504
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 42260 318899 42288 326862
rect 41722 318871 42288 318899
rect 41713 318213 42193 318269
rect 41713 317569 42193 317625
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 42352 314575 42380 339594
rect 41722 314547 42380 314575
rect 41722 313903 41828 313931
rect 41800 313546 41828 313903
rect 41788 313540 41840 313546
rect 41788 313482 41840 313488
rect 42352 313426 42380 314547
rect 42444 313546 42472 356594
rect 42536 353258 42564 367678
rect 42616 358284 42668 358290
rect 42616 358226 42668 358232
rect 42524 353252 42576 353258
rect 42524 353194 42576 353200
rect 42628 339658 42656 358226
rect 42720 357338 42748 370330
rect 42708 357332 42760 357338
rect 42708 357274 42760 357280
rect 42720 356658 42748 357274
rect 42708 356652 42760 356658
rect 42708 356594 42760 356600
rect 44192 353274 44220 372574
rect 42708 353252 42760 353258
rect 44192 353246 44404 353274
rect 42708 353194 42760 353200
rect 42616 339652 42668 339658
rect 42616 339594 42668 339600
rect 42720 324562 42748 353194
rect 44376 334014 44404 353246
rect 44180 334008 44232 334014
rect 44180 333950 44232 333956
rect 44364 334008 44416 334014
rect 44364 333950 44416 333956
rect 42708 324556 42760 324562
rect 42708 324498 42760 324504
rect 42432 313540 42484 313546
rect 42432 313482 42484 313488
rect 42616 313540 42668 313546
rect 42616 313482 42668 313488
rect 42352 313398 42564 313426
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 42536 286686 42564 313398
rect 42524 286680 42576 286686
rect 42524 286622 42576 286628
rect 41722 283675 41920 283703
rect 41892 283234 41920 283675
rect 41892 283206 42288 283234
rect 41713 283017 42193 283073
rect 41788 282328 41840 282334
rect 41788 282270 41840 282276
rect 41800 281874 41828 282270
rect 41722 281846 41828 281874
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 41722 275671 41828 275699
rect 41800 275618 41828 275671
rect 42260 275618 42288 283206
rect 42432 282328 42484 282334
rect 42432 282270 42484 282276
rect 41800 275590 42288 275618
rect 41713 275013 42193 275069
rect 41713 274369 42193 274425
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 41722 271374 41828 271402
rect 41800 270842 41828 271374
rect 41788 270836 41840 270842
rect 41788 270778 41840 270784
rect 42352 270774 42380 270805
rect 42340 270768 42392 270774
rect 41722 270716 42340 270722
rect 41722 270710 42392 270716
rect 41722 270694 42380 270710
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 42352 247042 42380 270694
rect 42340 247036 42392 247042
rect 42340 246978 42392 246984
rect 41722 240502 42288 240530
rect 41713 239817 42193 239873
rect 41788 239080 41840 239086
rect 41788 239022 41840 239028
rect 41800 238663 41828 239022
rect 41722 238635 41828 238663
rect 41713 237977 42193 238033
rect 41713 237333 42193 237389
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 42260 232642 42288 240502
rect 42444 239086 42472 282270
rect 42628 270774 42656 313482
rect 42720 282334 42748 324498
rect 44192 314650 44220 333950
rect 44192 314622 44404 314650
rect 42800 286680 42852 286686
rect 42800 286622 42852 286628
rect 42708 282328 42760 282334
rect 42708 282270 42760 282276
rect 42812 270842 42840 286622
rect 42800 270836 42852 270842
rect 42800 270778 42852 270784
rect 42616 270768 42668 270774
rect 42616 270710 42668 270716
rect 42708 247036 42760 247042
rect 42708 246978 42760 246984
rect 42432 239080 42484 239086
rect 42432 239022 42484 239028
rect 42616 239080 42668 239086
rect 42616 239022 42668 239028
rect 42524 237448 42576 237454
rect 42524 237390 42576 237396
rect 41800 232614 42288 232642
rect 41800 232506 41828 232614
rect 41722 232478 41828 232506
rect 41713 231813 42193 231869
rect 41713 231169 42193 231225
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 41722 228126 41920 228154
rect 41892 227882 41920 228126
rect 42536 227882 42564 237390
rect 41892 227854 42564 227882
rect 41788 227656 41840 227662
rect 41788 227598 41840 227604
rect 41800 227531 41828 227598
rect 41722 227503 41828 227531
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 42260 197402 42288 227854
rect 42432 227656 42484 227662
rect 42432 227598 42484 227604
rect 42248 197396 42300 197402
rect 42248 197338 42300 197344
rect 41722 197254 42288 197282
rect 41713 196617 42193 196673
rect 41788 195900 41840 195906
rect 41788 195842 41840 195848
rect 41800 195463 41828 195842
rect 41722 195435 41828 195463
rect 41713 194777 42193 194833
rect 41713 194133 42193 194189
rect 41713 192937 42193 192993
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 42260 189394 42288 197254
rect 41800 189366 42288 189394
rect 41800 189299 41828 189366
rect 41722 189271 41828 189299
rect 41713 188613 42193 188669
rect 41713 187969 42193 188025
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 41788 185496 41840 185502
rect 41788 185438 41840 185444
rect 41800 184975 41828 185438
rect 41722 184947 41828 184975
rect 42444 184890 42472 227598
rect 42628 195906 42656 239022
rect 42720 227662 42748 246978
rect 42812 237454 42840 270778
rect 44376 270502 44404 314622
rect 44272 270496 44324 270502
rect 44272 270438 44324 270444
rect 44364 270496 44416 270502
rect 44364 270438 44416 270444
rect 44284 256766 44312 270438
rect 44272 256760 44324 256766
rect 44272 256702 44324 256708
rect 44272 256624 44324 256630
rect 44272 256566 44324 256572
rect 42800 237448 42852 237454
rect 42800 237390 42852 237396
rect 44284 237402 44312 256566
rect 44284 237374 44404 237402
rect 42708 227656 42760 227662
rect 42708 227598 42760 227604
rect 44376 218074 44404 237374
rect 44180 218068 44232 218074
rect 44180 218010 44232 218016
rect 44364 218068 44416 218074
rect 44364 218010 44416 218016
rect 44192 217954 44220 218010
rect 44192 217926 44312 217954
rect 44284 198778 44312 217926
rect 44284 198750 44404 198778
rect 42708 197396 42760 197402
rect 42708 197338 42760 197344
rect 42616 195900 42668 195906
rect 42616 195842 42668 195848
rect 42720 185502 42748 197338
rect 42708 185496 42760 185502
rect 42708 185438 42760 185444
rect 41788 184884 41840 184890
rect 41788 184826 41840 184832
rect 42248 184884 42300 184890
rect 42248 184826 42300 184832
rect 42432 184884 42484 184890
rect 42432 184826 42484 184832
rect 41800 184331 41828 184826
rect 41722 184303 41828 184331
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 39856 125180 39908 125186
rect 39856 125122 39908 125128
rect 39868 120306 39896 125122
rect 39606 120278 39896 120306
rect 39868 120222 39896 120278
rect 39856 120216 39908 120222
rect 39856 120158 39908 120164
rect 41418 115968 41474 115977
rect 41418 115903 41474 115912
rect 39394 83192 39450 83201
rect 39394 83127 39450 83136
rect 39408 79098 39436 83127
rect 39316 79070 39528 79098
rect 39316 78948 39344 79070
rect 39500 78962 39528 79070
rect 39500 78934 39896 78962
rect 39592 75126 39804 75154
rect 39592 75018 39620 75126
rect 39567 74990 39620 75018
rect 39672 74928 39724 74934
rect 39672 74870 39724 74876
rect 39330 68190 39620 68218
rect 39592 67998 39620 68190
rect 39580 67992 39632 67998
rect 39580 67934 39632 67940
rect 39684 52426 39712 74870
rect 39672 52420 39724 52426
rect 39672 52362 39724 52368
rect 39776 44130 39804 75126
rect 39868 74934 39896 78934
rect 39856 74928 39908 74934
rect 39856 74870 39908 74876
rect 41432 67998 41460 115903
rect 41420 67992 41472 67998
rect 41420 67934 41472 67940
rect 41432 64530 41460 67934
rect 41420 64524 41472 64530
rect 41420 64466 41472 64472
rect 39856 52420 39908 52426
rect 39856 52362 39908 52368
rect 39868 45626 39896 52362
rect 42260 45898 42288 184826
rect 42720 179450 42748 185438
rect 44376 179450 44404 198750
rect 44640 195900 44692 195906
rect 44640 195842 44692 195848
rect 44652 193225 44680 195842
rect 44454 193216 44510 193225
rect 44454 193151 44510 193160
rect 44638 193216 44694 193225
rect 44638 193151 44694 193160
rect 42340 179444 42392 179450
rect 42340 179386 42392 179392
rect 42708 179444 42760 179450
rect 42708 179386 42760 179392
rect 44180 179444 44232 179450
rect 44180 179386 44232 179392
rect 44364 179444 44416 179450
rect 44364 179386 44416 179392
rect 42352 115977 42380 179386
rect 44192 179330 44220 179386
rect 44192 179302 44312 179330
rect 44284 160154 44312 179302
rect 44468 173942 44496 193151
rect 44456 173936 44508 173942
rect 44456 173878 44508 173884
rect 44732 173936 44784 173942
rect 44732 173878 44784 173884
rect 44744 160206 44772 173878
rect 44732 160200 44784 160206
rect 44284 160126 44404 160154
rect 44732 160142 44784 160148
rect 44376 140826 44404 160126
rect 44640 160064 44692 160070
rect 44640 160006 44692 160012
rect 44652 154562 44680 160006
rect 44640 154556 44692 154562
rect 44640 154498 44692 154504
rect 44824 154556 44876 154562
rect 44824 154498 44876 154504
rect 44836 154442 44864 154498
rect 44836 154414 44956 154442
rect 44180 140820 44232 140826
rect 44180 140762 44232 140768
rect 44364 140820 44416 140826
rect 44364 140762 44416 140768
rect 44192 125186 44220 140762
rect 44180 125180 44232 125186
rect 44180 125122 44232 125128
rect 44928 121394 44956 154414
rect 44652 121366 44956 121394
rect 42338 115968 42394 115977
rect 42338 115903 42394 115912
rect 44652 102082 44680 121366
rect 44732 120216 44784 120222
rect 44732 120158 44784 120164
rect 44744 110650 44772 120158
rect 44744 110622 44956 110650
rect 44744 110537 44772 110622
rect 44730 110528 44786 110537
rect 44730 110463 44786 110472
rect 44468 102054 44680 102082
rect 44468 96626 44496 102054
rect 44272 96620 44324 96626
rect 44272 96562 44324 96568
rect 44456 96620 44508 96626
rect 44456 96562 44508 96568
rect 44284 77314 44312 96562
rect 44272 77308 44324 77314
rect 44272 77250 44324 77256
rect 44364 77308 44416 77314
rect 44364 77250 44416 77256
rect 44376 75993 44404 77250
rect 44362 75984 44418 75993
rect 44362 75919 44418 75928
rect 44376 73409 44404 75919
rect 44362 73400 44418 73409
rect 44362 73335 44418 73344
rect 44376 71806 44404 73335
rect 44180 71800 44232 71806
rect 44180 71742 44232 71748
rect 44364 71800 44416 71806
rect 44364 71742 44416 71748
rect 44192 68241 44220 71742
rect 44178 68232 44234 68241
rect 44178 68167 44234 68176
rect 42708 64524 42760 64530
rect 42708 64466 42760 64472
rect 42248 45892 42300 45898
rect 42248 45834 42300 45840
rect 42720 45830 42748 64466
rect 42708 45824 42760 45830
rect 42708 45766 42760 45772
rect 44192 45694 44220 68167
rect 44180 45688 44232 45694
rect 44180 45630 44232 45636
rect 39856 45620 39908 45626
rect 39856 45562 39908 45568
rect 44928 45558 44956 110622
rect 145104 45892 145156 45898
rect 145104 45834 145156 45840
rect 140964 45824 141016 45830
rect 140964 45766 141016 45772
rect 44916 45552 44968 45558
rect 44916 45494 44968 45500
rect 140976 44538 141004 45766
rect 140964 44532 141016 44538
rect 140964 44474 141016 44480
rect 39764 44124 39816 44130
rect 39764 44066 39816 44072
rect 78956 44124 79008 44130
rect 78956 44066 79008 44072
rect 78968 40254 78996 44066
rect 135352 41744 135404 41750
rect 135352 41686 135404 41692
rect 91284 41608 91336 41614
rect 102140 41608 102192 41614
rect 91284 41550 91336 41556
rect 102060 41556 102140 41562
rect 102060 41550 102192 41556
rect 91296 40254 91324 41550
rect 102060 41546 102180 41550
rect 121380 41546 121500 41562
rect 102048 41540 102180 41546
rect 102100 41534 102180 41540
rect 121368 41540 121512 41546
rect 102048 41482 102100 41488
rect 121420 41534 121460 41540
rect 121368 41482 121420 41488
rect 121460 41482 121512 41488
rect 135260 41472 135312 41478
rect 135364 41426 135392 41686
rect 135312 41420 135392 41426
rect 135260 41414 135392 41420
rect 135272 41398 135392 41414
rect 78956 40248 79008 40254
rect 78954 40216 78956 40225
rect 86500 40248 86552 40254
rect 79008 40216 79010 40225
rect 78954 40151 79010 40160
rect 86498 40216 86500 40225
rect 91284 40248 91336 40254
rect 86552 40216 86554 40225
rect 91284 40190 91336 40196
rect 133098 40248 133150 40254
rect 133098 40190 133150 40196
rect 140976 40202 141004 44474
rect 145116 44266 145144 45834
rect 578792 45756 578844 45762
rect 578792 45698 578844 45704
rect 145840 45688 145892 45694
rect 145840 45630 145892 45636
rect 528652 45688 528704 45694
rect 528652 45630 528704 45636
rect 145104 44260 145156 44266
rect 145104 44202 145156 44208
rect 143816 40248 143868 40254
rect 86498 40151 86554 40160
rect 78968 40125 78996 40151
rect 133110 39984 133138 40190
rect 140976 40174 141036 40202
rect 145116 40202 145144 44202
rect 145852 40361 145880 45630
rect 189264 45620 189316 45626
rect 189264 45562 189316 45568
rect 173900 44600 173952 44606
rect 173898 44568 173900 44577
rect 173952 44568 173954 44577
rect 173898 44503 173954 44512
rect 186688 44192 186740 44198
rect 186688 44134 186740 44140
rect 186700 41820 186728 44134
rect 154488 41744 154540 41750
rect 154488 41686 154540 41692
rect 168288 41744 168340 41750
rect 187327 41713 187383 42193
rect 189276 41954 189304 45562
rect 195980 45552 196032 45558
rect 195980 45494 196032 45500
rect 516324 45552 516376 45558
rect 516324 45494 516376 45500
rect 193128 44668 193180 44674
rect 193128 44610 193180 44616
rect 193140 44577 193168 44610
rect 193126 44568 193182 44577
rect 193126 44503 193182 44512
rect 195992 44470 196020 45494
rect 289820 44872 289872 44878
rect 289820 44814 289872 44820
rect 313188 44872 313240 44878
rect 313188 44814 313240 44820
rect 458180 44872 458232 44878
rect 458180 44814 458232 44820
rect 250996 44804 251048 44810
rect 250996 44746 251048 44752
rect 252100 44804 252152 44810
rect 252100 44746 252152 44752
rect 276020 44804 276072 44810
rect 276020 44746 276072 44752
rect 231860 44736 231912 44742
rect 231858 44704 231860 44713
rect 251008 44713 251036 44746
rect 231912 44704 231914 44713
rect 250994 44704 251050 44713
rect 231858 44639 231914 44648
rect 247684 44668 247736 44674
rect 250994 44639 251050 44648
rect 247684 44610 247736 44616
rect 212538 44568 212594 44577
rect 199660 44532 199712 44538
rect 212538 44503 212540 44512
rect 199660 44474 199712 44480
rect 212592 44503 212594 44512
rect 217888 44538 218100 44554
rect 217888 44532 218112 44538
rect 217888 44526 218060 44532
rect 212540 44474 212592 44480
rect 195980 44464 196032 44470
rect 195980 44406 196032 44412
rect 195336 44260 195388 44266
rect 195336 44202 195388 44208
rect 194692 44192 194744 44198
rect 194692 44134 194744 44140
rect 189264 41948 189316 41954
rect 189264 41890 189316 41896
rect 191104 41948 191156 41954
rect 191104 41890 191156 41896
rect 192300 41948 192352 41954
rect 192300 41890 192352 41896
rect 193588 41948 193640 41954
rect 193588 41890 193640 41896
rect 188620 41880 188672 41886
rect 188554 41828 188620 41834
rect 189276 41834 189304 41890
rect 191116 41834 191144 41890
rect 192312 41834 192340 41890
rect 192944 41880 192996 41886
rect 188554 41822 188672 41828
rect 188554 41806 188660 41822
rect 189198 41806 189304 41834
rect 191038 41806 191144 41834
rect 192234 41806 192340 41834
rect 192878 41828 192944 41834
rect 193600 41834 193628 41890
rect 192878 41822 192996 41828
rect 192878 41806 192984 41822
rect 193522 41806 193628 41834
rect 194043 41713 194099 42193
rect 194704 41820 194732 44134
rect 195348 41820 195376 44202
rect 195992 41820 196020 44406
rect 199016 44396 199068 44402
rect 199016 44338 199068 44344
rect 196440 41948 196492 41954
rect 196440 41890 196492 41896
rect 198464 41948 198516 41954
rect 198464 41890 198516 41896
rect 196452 41834 196480 41890
rect 198476 41834 198504 41890
rect 199028 41834 199056 44338
rect 199672 44266 199700 44474
rect 217888 44470 217916 44526
rect 218060 44474 218112 44480
rect 200764 44464 200816 44470
rect 200764 44406 200816 44412
rect 200856 44464 200908 44470
rect 200856 44406 200908 44412
rect 217876 44464 217928 44470
rect 242900 44464 242952 44470
rect 217876 44406 217928 44412
rect 200776 44266 200804 44406
rect 199660 44260 199712 44266
rect 199660 44202 199712 44208
rect 200764 44260 200816 44266
rect 200764 44202 200816 44208
rect 196452 41806 198504 41834
rect 198936 41820 199056 41834
rect 199672 41820 199700 44202
rect 200120 41948 200172 41954
rect 200120 41890 200172 41896
rect 200132 41834 200160 41890
rect 200868 41834 200896 44406
rect 217980 44402 218192 44418
rect 242900 44406 242952 44412
rect 217968 44396 218204 44402
rect 218020 44390 218152 44396
rect 217968 44338 218020 44344
rect 218152 44338 218204 44344
rect 201592 41880 201644 41886
rect 200132 41820 200896 41834
rect 201526 41828 201592 41834
rect 201526 41822 201644 41828
rect 202512 41880 202564 41886
rect 202512 41822 202564 41828
rect 198936 41818 199042 41820
rect 198924 41812 199042 41818
rect 198976 41806 199042 41812
rect 200132 41806 200882 41820
rect 201526 41806 201632 41822
rect 198924 41754 198976 41760
rect 168288 41686 168340 41692
rect 154500 41614 154528 41686
rect 154488 41608 154540 41614
rect 154488 41550 154540 41556
rect 149980 41472 150032 41478
rect 149980 41414 150032 41420
rect 149992 40361 150020 41414
rect 168300 41410 168328 41686
rect 202524 41478 202552 41822
rect 202512 41472 202564 41478
rect 202512 41414 202564 41420
rect 240140 41472 240192 41478
rect 240140 41414 240192 41420
rect 168288 41404 168340 41410
rect 168288 41346 168340 41352
rect 145838 40352 145894 40361
rect 145838 40287 145894 40296
rect 149978 40352 150034 40361
rect 149978 40287 150034 40296
rect 143816 40190 143868 40196
rect 141008 40118 141036 40174
rect 140996 40112 141048 40118
rect 140996 40054 141048 40060
rect 143072 40112 143124 40118
rect 143072 40054 143124 40060
rect 143356 40112 143408 40118
rect 143356 40054 143408 40060
rect 141008 39984 141036 40054
rect 143084 39984 143112 40054
rect 143368 39916 143396 40054
rect 143828 39916 143856 40190
rect 145103 40174 145144 40202
rect 145103 40000 145131 40174
rect 145091 39706 145143 40000
rect 240152 39953 240180 41414
rect 240138 39944 240194 39953
rect 240138 39879 240194 39888
rect 242912 39817 242940 44406
rect 247696 44402 247724 44610
rect 248326 44568 248382 44577
rect 248326 44503 248382 44512
rect 247408 44396 247460 44402
rect 247408 44338 247460 44344
rect 247684 44396 247736 44402
rect 247684 44338 247736 44344
rect 241242 39808 241298 39817
rect 241242 39743 241298 39752
rect 242898 39808 242954 39817
rect 242898 39743 242954 39752
rect 241256 39372 241284 39743
rect 247420 39581 247448 44338
rect 248340 44334 248368 44503
rect 248328 44328 248380 44334
rect 248328 44270 248380 44276
rect 247342 39553 247448 39581
rect 252112 39372 252140 44746
rect 276032 44538 276060 44746
rect 289832 44606 289860 44814
rect 308220 44736 308272 44742
rect 308220 44678 308272 44684
rect 307576 44668 307628 44674
rect 307576 44610 307628 44616
rect 289820 44600 289872 44606
rect 289820 44542 289872 44548
rect 276020 44532 276072 44538
rect 276020 44474 276072 44480
rect 299572 44532 299624 44538
rect 299572 44474 299624 44480
rect 305736 44532 305788 44538
rect 305736 44474 305788 44480
rect 297732 44464 297784 44470
rect 289818 44432 289874 44441
rect 286888 44390 287008 44418
rect 267740 44328 267792 44334
rect 267738 44296 267740 44305
rect 286888 44305 286916 44390
rect 286980 44334 287008 44390
rect 297732 44406 297784 44412
rect 289818 44367 289820 44376
rect 289872 44367 289874 44376
rect 289820 44338 289872 44344
rect 286968 44328 287020 44334
rect 267792 44296 267794 44305
rect 267738 44231 267794 44240
rect 286874 44296 286930 44305
rect 286968 44270 287020 44276
rect 286874 44231 286930 44240
rect 295248 44192 295300 44198
rect 295248 44134 295300 44140
rect 295260 41834 295288 44134
rect 297744 41834 297772 44406
rect 299480 41880 299532 41886
rect 295260 41806 295311 41834
rect 296916 41818 297151 41834
rect 296904 41812 297151 41818
rect 296956 41806 297151 41812
rect 297744 41806 297795 41834
rect 299584 41834 299612 44474
rect 300768 44464 300820 44470
rect 300768 44406 300820 44412
rect 303894 44432 303950 44441
rect 300780 41834 300808 44406
rect 303894 44367 303950 44376
rect 303252 44192 303304 44198
rect 303252 44134 303304 44140
rect 299532 41828 299635 41834
rect 299480 41822 299635 41828
rect 299492 41806 299635 41822
rect 300780 41806 302119 41834
rect 296904 41754 296956 41760
rect 302643 41713 302699 42193
rect 303264 41834 303292 44134
rect 303908 42294 303936 44367
rect 304540 44260 304592 44266
rect 304540 44202 304592 44208
rect 303896 42288 303948 42294
rect 303896 42230 303948 42236
rect 303908 41834 303936 42230
rect 304552 41834 304580 44202
rect 305748 41834 305776 44474
rect 306380 44464 306432 44470
rect 306380 44406 306432 44412
rect 306392 44198 306420 44406
rect 307588 44266 307616 44610
rect 307576 44260 307628 44266
rect 307576 44202 307628 44208
rect 306380 44192 306432 44198
rect 306380 44134 306432 44140
rect 306392 41834 306420 44134
rect 303264 41806 303315 41834
rect 303908 41806 303959 41834
rect 304552 41806 304603 41834
rect 305155 41818 305316 41834
rect 305155 41812 305328 41818
rect 305155 41806 305276 41812
rect 305748 41806 305799 41834
rect 306300 41818 306443 41834
rect 306288 41812 306443 41818
rect 305276 41754 305328 41760
rect 306340 41806 306443 41812
rect 306288 41754 306340 41760
rect 306967 41713 307023 42193
rect 307588 41834 307616 44202
rect 308232 42294 308260 44678
rect 308312 44668 308364 44674
rect 308312 44610 308364 44616
rect 309140 44668 309192 44674
rect 309140 44610 309192 44616
rect 308324 44266 308352 44610
rect 309152 44577 309180 44610
rect 313200 44606 313228 44814
rect 380900 44804 380952 44810
rect 380900 44746 380952 44752
rect 400128 44804 400180 44810
rect 400128 44746 400180 44752
rect 406752 44804 406804 44810
rect 406752 44746 406804 44752
rect 358728 44736 358780 44742
rect 358728 44678 358780 44684
rect 362408 44736 362460 44742
rect 362408 44678 362460 44684
rect 328368 44668 328420 44674
rect 328368 44610 328420 44616
rect 347780 44668 347832 44674
rect 347780 44610 347832 44616
rect 309416 44600 309468 44606
rect 309138 44568 309194 44577
rect 309416 44542 309468 44548
rect 313188 44600 313240 44606
rect 328380 44577 328408 44610
rect 313188 44542 313240 44548
rect 328366 44568 328422 44577
rect 309138 44503 309194 44512
rect 308312 44260 308364 44266
rect 308312 44202 308364 44208
rect 309428 44198 309456 44542
rect 328366 44503 328422 44512
rect 309416 44192 309468 44198
rect 309416 44134 309468 44140
rect 308220 42288 308272 42294
rect 308220 42230 308272 42236
rect 308232 41834 308260 42230
rect 309428 41834 309456 44134
rect 347792 43722 347820 44610
rect 352564 44532 352616 44538
rect 352564 44474 352616 44480
rect 355600 44532 355652 44538
rect 355600 44474 355652 44480
rect 351920 44464 351972 44470
rect 351920 44406 351972 44412
rect 350080 44192 350132 44198
rect 350080 44134 350132 44140
rect 347780 43716 347832 43722
rect 347780 43658 347832 43664
rect 307588 41806 307639 41834
rect 308232 41806 308283 41834
rect 308835 41806 309479 41834
rect 310095 41713 310151 42193
rect 350092 41820 350120 44134
rect 351932 41820 351960 44406
rect 352576 41820 352604 44474
rect 354404 44464 354456 44470
rect 354404 44406 354456 44412
rect 354416 41820 354444 44406
rect 355612 41834 355640 44474
rect 358084 44192 358136 44198
rect 358084 44134 358136 44140
rect 355612 41820 356914 41834
rect 355626 41806 356914 41820
rect 357443 41713 357499 42193
rect 358096 41820 358124 44134
rect 358740 41834 358768 44678
rect 359924 44532 359976 44538
rect 359924 44474 359976 44480
rect 359372 44396 359424 44402
rect 359372 44338 359424 44344
rect 358740 41820 358860 41834
rect 359384 41820 359412 44338
rect 359936 41834 359964 44474
rect 360568 44464 360620 44470
rect 360568 44406 360620 44412
rect 360580 44334 360608 44406
rect 360568 44328 360620 44334
rect 360568 44270 360620 44276
rect 360016 41880 360068 41886
rect 359936 41828 360016 41834
rect 359936 41822 360068 41828
rect 359936 41820 360056 41822
rect 360580 41820 360608 44270
rect 362420 43722 362448 44678
rect 380912 44606 380940 44746
rect 386420 44668 386472 44674
rect 386420 44610 386472 44616
rect 380900 44600 380952 44606
rect 386432 44577 386460 44610
rect 400140 44606 400168 44746
rect 405648 44668 405700 44674
rect 405648 44610 405700 44616
rect 400128 44600 400180 44606
rect 380900 44542 380952 44548
rect 386418 44568 386474 44577
rect 364156 44532 364208 44538
rect 405660 44577 405688 44610
rect 400128 44542 400180 44548
rect 405646 44568 405702 44577
rect 386418 44503 386474 44512
rect 405646 44503 405702 44512
rect 364156 44474 364208 44480
rect 363052 44464 363104 44470
rect 363052 44406 363104 44412
rect 362408 43716 362460 43722
rect 362408 43658 362460 43664
rect 361120 41880 361172 41886
rect 361172 41828 361238 41834
rect 361120 41822 361238 41828
rect 358754 41818 358860 41820
rect 358754 41812 358872 41818
rect 358754 41806 358820 41812
rect 359950 41806 360056 41820
rect 361132 41806 361238 41822
rect 358820 41754 358872 41760
rect 361767 41713 361823 42193
rect 362420 41820 362448 43658
rect 363064 41834 363092 44406
rect 363512 41948 363564 41954
rect 363512 41890 363564 41896
rect 362972 41820 363092 41834
rect 363524 41834 363552 41890
rect 364168 41834 364196 44474
rect 406764 44334 406792 44746
rect 417240 44668 417292 44674
rect 417240 44610 417292 44616
rect 425060 44668 425112 44674
rect 425060 44610 425112 44616
rect 444288 44668 444340 44674
rect 444288 44610 444340 44616
rect 407396 44532 407448 44538
rect 407396 44474 407448 44480
rect 410432 44532 410484 44538
rect 410432 44474 410484 44480
rect 406752 44328 406804 44334
rect 406752 44270 406804 44276
rect 404912 44192 404964 44198
rect 404912 44134 404964 44140
rect 362972 41818 363078 41820
rect 362960 41812 363078 41818
rect 363012 41806 363078 41812
rect 363524 41806 364274 41834
rect 362960 41754 363012 41760
rect 364895 41713 364951 42193
rect 404924 41820 404952 44134
rect 405527 41713 405583 42193
rect 406764 41820 406792 44270
rect 407408 41820 407436 44474
rect 409328 41880 409380 41886
rect 409262 41828 409328 41834
rect 409262 41822 409380 41828
rect 410444 41834 410472 44474
rect 413560 44464 413612 44470
rect 413560 44406 413612 44412
rect 411076 44328 411128 44334
rect 411076 44270 411128 44276
rect 409262 41806 409368 41822
rect 410444 41820 410564 41834
rect 411088 41820 411116 44270
rect 412916 44192 412968 44198
rect 412916 44134 412968 44140
rect 412243 41834 412299 42193
rect 412364 41880 412416 41886
rect 410458 41818 410564 41820
rect 411548 41818 411746 41834
rect 410458 41812 410576 41818
rect 410458 41806 410524 41812
rect 410524 41754 410576 41760
rect 411536 41812 411746 41818
rect 411588 41806 411746 41812
rect 412243 41828 412364 41834
rect 412243 41822 412416 41828
rect 412243 41806 412404 41822
rect 412928 41820 412956 44134
rect 413572 41820 413600 44406
rect 414204 44396 414256 44402
rect 414204 44338 414256 44344
rect 414216 41820 414244 44338
rect 415216 41880 415268 41886
rect 414584 41818 414782 41834
rect 415268 41828 415426 41834
rect 415216 41822 415426 41828
rect 414572 41812 414782 41818
rect 411536 41754 411588 41760
rect 412243 41713 412299 41806
rect 414624 41806 414782 41812
rect 415228 41806 415426 41822
rect 415872 41818 416070 41834
rect 415860 41812 416070 41818
rect 414572 41754 414624 41760
rect 415912 41806 416070 41812
rect 415860 41754 415912 41760
rect 416567 41713 416623 42193
rect 417252 41820 417280 44610
rect 419540 44600 419592 44606
rect 425072 44577 425100 44610
rect 438768 44600 438820 44606
rect 419540 44542 419592 44548
rect 425058 44568 425114 44577
rect 419080 44532 419132 44538
rect 419080 44474 419132 44480
rect 417884 44464 417936 44470
rect 417884 44406 417936 44412
rect 417896 41820 417924 44406
rect 419092 41834 419120 44474
rect 419552 44334 419580 44542
rect 444300 44577 444328 44610
rect 458192 44606 458220 44814
rect 461492 44804 461544 44810
rect 461492 44746 461544 44752
rect 458180 44600 458232 44606
rect 438768 44542 438820 44548
rect 444286 44568 444342 44577
rect 425058 44503 425114 44512
rect 438780 44334 438808 44542
rect 458180 44542 458232 44548
rect 444286 44503 444342 44512
rect 461504 44334 461532 44746
rect 488540 44736 488592 44742
rect 488460 44684 488540 44690
rect 488460 44678 488592 44684
rect 499580 44736 499632 44742
rect 499580 44678 499632 44684
rect 488460 44674 488580 44678
rect 471980 44668 472032 44674
rect 472072 44668 472124 44674
rect 472032 44628 472072 44656
rect 471980 44610 472032 44616
rect 472072 44610 472124 44616
rect 472348 44668 472400 44674
rect 472348 44610 472400 44616
rect 488448 44668 488580 44674
rect 488500 44662 488580 44668
rect 488448 44610 488500 44616
rect 462136 44532 462188 44538
rect 462136 44474 462188 44480
rect 465172 44532 465224 44538
rect 465172 44474 465224 44480
rect 419540 44328 419592 44334
rect 419540 44270 419592 44276
rect 438768 44328 438820 44334
rect 438768 44270 438820 44276
rect 461492 44328 461544 44334
rect 461492 44270 461544 44276
rect 419724 44192 419776 44198
rect 419724 44134 419776 44140
rect 459652 44192 459704 44198
rect 459652 44134 459704 44140
rect 419736 42193 419764 44134
rect 418264 41820 419120 41834
rect 419695 41820 419764 42193
rect 459664 41834 459692 44134
rect 418264 41818 419106 41820
rect 418252 41812 419106 41818
rect 418304 41806 419106 41812
rect 418252 41754 418304 41760
rect 419695 41713 419751 41820
rect 459664 41806 459711 41834
rect 460327 41713 460383 42193
rect 461504 41834 461532 44270
rect 462148 41834 462176 44474
rect 465184 41834 465212 44474
rect 468300 44464 468352 44470
rect 468300 44406 468352 44412
rect 465816 44260 465868 44266
rect 465816 44202 465868 44208
rect 465356 41880 465408 41886
rect 461504 41806 461551 41834
rect 462148 41806 462195 41834
rect 464035 41818 464200 41834
rect 465184 41828 465356 41834
rect 465184 41822 465408 41828
rect 465828 41834 465856 44202
rect 467656 44192 467708 44198
rect 467656 44134 467708 44140
rect 466368 41880 466420 41886
rect 464035 41812 464212 41818
rect 464035 41806 464160 41812
rect 465184 41806 465396 41822
rect 465828 41806 465875 41834
rect 467043 41834 467099 42193
rect 467668 41834 467696 44134
rect 468312 41834 468340 44406
rect 468944 44396 468996 44402
rect 468944 44338 468996 44344
rect 468956 41834 468984 44338
rect 469404 41880 469456 41886
rect 466420 41828 466519 41834
rect 466368 41822 466519 41828
rect 466380 41806 466519 41822
rect 467043 41818 467236 41834
rect 467043 41812 467248 41818
rect 467043 41806 467196 41812
rect 464160 41754 464212 41760
rect 467043 41713 467099 41806
rect 467668 41806 467715 41834
rect 468312 41806 468359 41834
rect 468956 41806 469003 41834
rect 470692 41880 470744 41886
rect 469456 41828 469555 41834
rect 469404 41822 469555 41828
rect 469416 41806 469555 41822
rect 470060 41818 470199 41834
rect 470744 41828 470843 41834
rect 470692 41822 470843 41828
rect 470048 41812 470199 41818
rect 467196 41754 467248 41760
rect 470100 41806 470199 41812
rect 470704 41806 470843 41822
rect 470048 41754 470100 41760
rect 471367 41713 471423 42193
rect 472360 41857 472388 44610
rect 499592 44577 499620 44678
rect 499578 44568 499634 44577
rect 473820 44532 473872 44538
rect 499578 44503 499634 44512
rect 473820 44474 473872 44480
rect 472624 44464 472676 44470
rect 472624 44406 472676 44412
rect 472011 41848 472067 41857
rect 472011 41783 472067 41792
rect 472346 41848 472402 41857
rect 472636 41834 472664 44406
rect 473084 41880 473136 41886
rect 472636 41806 472683 41834
rect 473832 41834 473860 44474
rect 516336 44334 516364 45494
rect 526812 44736 526864 44742
rect 526812 44678 526864 44684
rect 518808 44668 518860 44674
rect 518808 44610 518860 44616
rect 518820 44577 518848 44610
rect 518806 44568 518862 44577
rect 516968 44532 517020 44538
rect 518806 44503 518862 44512
rect 516968 44474 517020 44480
rect 516324 44328 516376 44334
rect 516324 44270 516376 44276
rect 474464 44260 474516 44266
rect 474464 44202 474516 44208
rect 514484 44260 514536 44266
rect 514484 44202 514536 44208
rect 474476 42193 474504 44202
rect 473136 41828 473879 41834
rect 473084 41822 473879 41828
rect 473096 41806 473879 41822
rect 474476 41806 474551 42193
rect 514496 41820 514524 44202
rect 472346 41783 472402 41792
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 516336 41820 516364 44270
rect 516980 41834 517008 44474
rect 523132 44464 523184 44470
rect 523132 44406 523184 44412
rect 523144 44266 523172 44406
rect 523776 44396 523828 44402
rect 523776 44338 523828 44344
rect 522488 44260 522540 44266
rect 522488 44202 522540 44208
rect 523132 44260 523184 44266
rect 523132 44202 523184 44208
rect 518808 44192 518860 44198
rect 518808 44134 518860 44140
rect 517060 41880 517112 41886
rect 516980 41828 517060 41834
rect 516980 41822 517112 41828
rect 516980 41820 517100 41822
rect 518820 41820 518848 44134
rect 520096 41880 520148 41886
rect 520030 41828 520096 41834
rect 520030 41822 520148 41828
rect 516994 41806 517100 41820
rect 520030 41806 520136 41822
rect 520647 41713 520703 42193
rect 521384 41880 521436 41886
rect 521318 41828 521384 41834
rect 521318 41822 521436 41828
rect 521318 41806 521424 41822
rect 521843 41713 521899 42193
rect 522500 41820 522528 44202
rect 523144 41820 523172 44202
rect 523788 41834 523816 44338
rect 524972 44192 525024 44198
rect 524972 44134 525024 44140
rect 525616 44192 525668 44198
rect 525616 44134 525668 44140
rect 524984 42193 525012 44134
rect 524420 41880 524472 41886
rect 523788 41820 523908 41834
rect 523802 41818 523908 41820
rect 524354 41828 524420 41834
rect 524354 41822 524472 41828
rect 523802 41812 523920 41818
rect 523802 41806 523868 41812
rect 524354 41806 524460 41822
rect 523868 41754 523920 41760
rect 524971 41713 525027 42193
rect 525524 41880 525576 41886
rect 525628 41834 525656 44134
rect 525576 41828 525656 41834
rect 525524 41822 525656 41828
rect 525536 41820 525656 41822
rect 525536 41806 525642 41820
rect 526167 41713 526223 42193
rect 526824 41834 526852 44678
rect 527456 44260 527508 44266
rect 527456 44202 527508 44208
rect 526824 41820 526944 41834
rect 527468 41820 527496 44202
rect 528664 44198 528692 45630
rect 529848 45620 529900 45626
rect 529848 45562 529900 45568
rect 529860 44266 529888 45562
rect 560312 44934 560524 44962
rect 560312 44878 560340 44934
rect 546592 44872 546644 44878
rect 546420 44820 546592 44826
rect 546420 44814 546644 44820
rect 560300 44872 560352 44878
rect 560300 44814 560352 44820
rect 546420 44798 546632 44814
rect 546420 44742 546448 44798
rect 546408 44736 546460 44742
rect 546408 44678 546460 44684
rect 529848 44260 529900 44266
rect 529848 44202 529900 44208
rect 528652 44192 528704 44198
rect 528652 44134 528704 44140
rect 528664 41834 528692 44134
rect 528034 41820 528692 41834
rect 526838 41818 526944 41820
rect 526838 41812 526956 41818
rect 526838 41806 526904 41812
rect 528034 41806 528678 41820
rect 526904 41754 526956 41760
rect 529295 41713 529351 42193
rect 253940 41608 253992 41614
rect 253940 41550 253992 41556
rect 253952 39953 253980 41550
rect 560496 40225 560524 44934
rect 569132 41540 569184 41546
rect 569132 41482 569184 41488
rect 560482 40216 560538 40225
rect 560482 40151 560538 40160
rect 253938 39944 253994 39953
rect 253938 39879 253994 39888
rect 569144 39644 569172 41482
rect 578804 40225 578832 45698
rect 673104 45694 673132 408478
rect 673564 392034 673592 411182
rect 673472 392006 673592 392034
rect 673472 384062 673500 392006
rect 676232 388686 676260 459954
rect 677704 459870 678086 459898
rect 677704 440230 677732 459870
rect 676312 440224 676364 440230
rect 676312 440166 676364 440172
rect 677692 440224 677744 440230
rect 677692 440166 677744 440172
rect 676324 408542 676352 440166
rect 677508 427848 677560 427854
rect 677508 427790 677560 427796
rect 677520 425762 677548 427790
rect 677598 425776 677654 425785
rect 677520 425734 677598 425762
rect 677598 425711 677654 425720
rect 677508 420776 677560 420782
rect 677506 420744 677508 420753
rect 677560 420744 677562 420753
rect 677506 420679 677562 420688
rect 676312 408536 676364 408542
rect 676312 408478 676364 408484
rect 675300 388680 675352 388686
rect 675300 388622 675352 388628
rect 676220 388680 676272 388686
rect 676220 388622 676272 388628
rect 673460 384056 673512 384062
rect 673460 383998 673512 384004
rect 673472 338162 673500 383998
rect 675312 383253 675340 388622
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 675392 384056 675444 384062
rect 675392 383998 675444 384004
rect 675404 383860 675432 383998
rect 675312 383239 675418 383253
rect 675312 383225 675432 383239
rect 675404 382770 675432 383225
rect 673644 382764 673696 382770
rect 673644 382706 673696 382712
rect 675392 382764 675444 382770
rect 675392 382706 675444 382712
rect 673552 372360 673604 372366
rect 673552 372302 673604 372308
rect 673460 338156 673512 338162
rect 673460 338098 673512 338104
rect 673564 328098 673592 372302
rect 673656 337550 673684 382706
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675407 380175 675887 380231
rect 675407 379531 675887 379587
rect 675312 378901 675418 378929
rect 675312 370925 675340 378901
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675404 372366 675432 372751
rect 675392 372360 675444 372366
rect 675392 372302 675444 372308
rect 675407 371527 675887 371583
rect 675312 370897 675418 370925
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675404 338162 675432 338708
rect 673736 338156 673788 338162
rect 673736 338098 673788 338104
rect 675392 338156 675444 338162
rect 675392 338098 675444 338104
rect 673644 337544 673696 337550
rect 673644 337486 673696 337492
rect 673552 328092 673604 328098
rect 673552 328034 673604 328040
rect 673460 293616 673512 293622
rect 673460 293558 673512 293564
rect 673472 248606 673500 293558
rect 673564 282198 673592 328034
rect 673656 293622 673684 337486
rect 673748 293894 673776 338098
rect 675404 337550 675432 338028
rect 675392 337544 675444 337550
rect 675392 337486 675444 337492
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 334975 675887 335031
rect 675407 334331 675887 334387
rect 675312 333701 675418 333729
rect 675312 325725 675340 333701
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675392 328092 675444 328098
rect 675392 328034 675444 328040
rect 675404 327556 675432 328034
rect 675407 326327 675887 326383
rect 675312 325697 675418 325725
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 673736 293888 673788 293894
rect 673736 293830 673788 293836
rect 674012 293888 674064 293894
rect 674012 293830 674064 293836
rect 675392 293888 675444 293894
rect 675392 293830 675444 293836
rect 673644 293616 673696 293622
rect 673644 293558 673696 293564
rect 673552 282192 673604 282198
rect 673552 282134 673604 282140
rect 674024 264994 674052 293830
rect 675404 293692 675432 293830
rect 675392 293616 675444 293622
rect 675392 293558 675444 293564
rect 675404 293012 675432 293558
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 289975 675887 290031
rect 675407 289331 675887 289387
rect 675312 288701 675418 288729
rect 675024 282124 675076 282130
rect 675024 282066 675076 282072
rect 675036 265062 675064 282066
rect 675312 280725 675340 288701
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 675404 282130 675432 282540
rect 675392 282124 675444 282130
rect 675392 282066 675444 282072
rect 675407 281327 675887 281383
rect 675312 280697 675418 280725
rect 675024 265056 675076 265062
rect 675024 264998 675076 265004
rect 673736 264988 673788 264994
rect 673736 264930 673788 264936
rect 673828 264988 673880 264994
rect 673828 264930 673880 264936
rect 674012 264988 674064 264994
rect 674012 264930 674064 264936
rect 673552 249144 673604 249150
rect 673552 249086 673604 249092
rect 673460 248600 673512 248606
rect 673460 248542 673512 248548
rect 673460 237720 673512 237726
rect 673460 237662 673512 237668
rect 673472 191962 673500 237662
rect 673564 202978 673592 249086
rect 673644 248600 673696 248606
rect 673644 248542 673696 248548
rect 673656 206990 673684 248542
rect 673748 237726 673776 264930
rect 673840 249150 673868 264930
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 673828 249144 673880 249150
rect 673828 249086 673880 249092
rect 675392 249144 675444 249150
rect 675392 249086 675444 249092
rect 675404 248676 675432 249086
rect 675392 248600 675444 248606
rect 675392 248542 675444 248548
rect 675404 248039 675432 248542
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 244975 675887 245031
rect 675407 244331 675887 244387
rect 675312 243701 675418 243729
rect 673736 237720 673788 237726
rect 673736 237662 673788 237668
rect 675312 235725 675340 243701
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 675407 238167 675887 238223
rect 675392 237720 675444 237726
rect 675392 237662 675444 237668
rect 675404 237524 675432 237662
rect 675407 236327 675887 236383
rect 675312 235697 675418 235725
rect 673644 206984 673696 206990
rect 673644 206926 673696 206932
rect 675300 206984 675352 206990
rect 675300 206926 675352 206932
rect 673552 202972 673604 202978
rect 673552 202914 673604 202920
rect 673460 191956 673512 191962
rect 673460 191898 673512 191904
rect 673472 178022 673500 191898
rect 673460 178016 673512 178022
rect 673460 177958 673512 177964
rect 673564 168366 673592 202914
rect 675312 202858 675340 206926
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 675404 202978 675432 203483
rect 675392 202972 675444 202978
rect 675392 202914 675444 202920
rect 675312 202844 675418 202858
rect 675312 202830 675432 202844
rect 675404 202314 675432 202830
rect 675220 202286 675432 202314
rect 675220 184482 675248 202286
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 199775 675887 199831
rect 675407 199131 675887 199187
rect 675312 198614 675432 198642
rect 675312 190525 675340 198614
rect 675404 198492 675432 198614
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 675407 194807 675887 194863
rect 675407 192967 675887 193023
rect 675404 191962 675432 192372
rect 675392 191956 675444 191962
rect 675392 191898 675444 191904
rect 675407 191127 675887 191183
rect 675312 190497 675418 190525
rect 673736 184476 673788 184482
rect 673736 184418 673788 184424
rect 675208 184476 675260 184482
rect 675208 184418 675260 184424
rect 673748 168366 673776 184418
rect 673920 178016 673972 178022
rect 673920 177958 673972 177964
rect 673552 168360 673604 168366
rect 673552 168302 673604 168308
rect 673736 168360 673788 168366
rect 673736 168302 673788 168308
rect 673460 157956 673512 157962
rect 673460 157898 673512 157904
rect 673472 129742 673500 157898
rect 673828 157344 673880 157350
rect 673828 157286 673880 157292
rect 673644 147892 673696 147898
rect 673644 147834 673696 147840
rect 673460 129736 673512 129742
rect 673460 129678 673512 129684
rect 673460 112804 673512 112810
rect 673460 112746 673512 112752
rect 673092 45688 673144 45694
rect 673092 45630 673144 45636
rect 673472 45626 673500 112746
rect 673552 112124 673604 112130
rect 673552 112066 673604 112072
rect 673564 45762 673592 112066
rect 673656 101726 673684 147834
rect 673840 129742 673868 157286
rect 673932 147898 673960 177958
rect 675208 168360 675260 168366
rect 675208 168302 675260 168308
rect 675220 157842 675248 168302
rect 675300 168292 675352 168298
rect 675300 168234 675352 168240
rect 675312 158386 675340 168234
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675404 158386 675432 158508
rect 675312 158358 675432 158386
rect 675404 157962 675432 158358
rect 675392 157956 675444 157962
rect 675392 157898 675444 157904
rect 675220 157828 675418 157842
rect 675220 157814 675432 157828
rect 675404 157350 675432 157814
rect 675392 157344 675444 157350
rect 675392 157286 675444 157292
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 154775 675887 154831
rect 675407 154131 675887 154187
rect 675312 153501 675418 153529
rect 673920 147892 673972 147898
rect 673920 147834 673972 147840
rect 675312 145525 675340 153501
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675392 147892 675444 147898
rect 675392 147834 675444 147840
rect 675404 147356 675432 147834
rect 675407 146127 675887 146183
rect 675312 145497 675418 145525
rect 673736 129736 673788 129742
rect 673736 129678 673788 129684
rect 673828 129736 673880 129742
rect 673828 129678 673880 129684
rect 675300 129736 675352 129742
rect 675300 129678 675352 129684
rect 673748 112810 673776 129678
rect 673736 112804 673788 112810
rect 673736 112746 673788 112752
rect 675312 112653 675340 129678
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675404 112810 675432 113283
rect 675392 112804 675444 112810
rect 675392 112746 675444 112752
rect 675312 112639 675418 112653
rect 675312 112625 675432 112639
rect 675404 112130 675432 112625
rect 675392 112124 675444 112130
rect 675392 112066 675444 112072
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675407 109575 675887 109631
rect 675407 108931 675887 108987
rect 675312 108310 675418 108338
rect 673644 101720 673696 101726
rect 673644 101662 673696 101668
rect 673552 45756 673604 45762
rect 673552 45698 673604 45704
rect 673460 45620 673512 45626
rect 673460 45562 673512 45568
rect 673656 45558 673684 101662
rect 675312 100314 675340 108310
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675404 101726 675432 102151
rect 675392 101720 675444 101726
rect 675392 101662 675444 101668
rect 675407 100927 675887 100983
rect 675312 100286 675418 100314
rect 673644 45552 673696 45558
rect 673644 45494 673696 45500
rect 629300 41472 629352 41478
rect 629300 41414 629352 41420
rect 622950 40488 623006 40497
rect 622950 40423 623006 40432
rect 578790 40216 578846 40225
rect 578790 40151 578846 40160
rect 622964 39681 622992 40423
rect 629312 40225 629340 41414
rect 629298 40216 629354 40225
rect 629298 40151 629354 40160
rect 622950 39672 623006 39681
rect 622950 39607 623006 39616
<< via2 >>
rect 585046 997464 585102 997520
rect 585690 997464 585746 997520
rect 589554 997464 589610 997520
rect 343638 997056 343694 997112
rect 39486 928104 39542 928160
rect 41510 919672 41566 919728
rect 41510 917224 41566 917280
rect 39578 908112 39634 908168
rect 40038 907976 40094 908032
rect 40038 888936 40094 888992
rect 40130 877512 40186 877568
rect 41510 912192 41566 912248
rect 41418 875064 41474 875120
rect 40130 870032 40186 870088
rect 39854 869352 39910 869408
rect 39854 850312 39910 850368
rect 39762 827500 39764 827520
rect 39764 827500 39816 827520
rect 39816 827500 39818 827520
rect 39762 827464 39818 827500
rect 40222 516024 40278 516080
rect 40222 496984 40278 497040
rect 39762 492904 39818 492960
rect 39854 490456 39910 490512
rect 39854 488008 39910 488064
rect 40038 470600 40094 470656
rect 39670 451832 39726 451888
rect 40038 460944 40094 461000
rect 39946 455368 40002 455424
rect 39854 444352 39910 444408
rect 39670 440952 39726 441008
rect 289818 990564 289820 990584
rect 289820 990564 289872 990584
rect 289872 990564 289874 990584
rect 289818 990528 289874 990564
rect 295522 990528 295578 990584
rect 329562 992296 329618 992352
rect 364338 990428 364340 990448
rect 364340 990428 364392 990448
rect 364392 990428 364394 990448
rect 364338 990392 364394 990428
rect 383566 990392 383622 990448
rect 405738 990276 405794 990312
rect 405738 990256 405740 990276
rect 405740 990256 405792 990276
rect 405792 990256 405794 990276
rect 424966 990256 425022 990312
rect 444378 990292 444380 990312
rect 444380 990292 444432 990312
rect 444432 990292 444434 990312
rect 444378 990256 444434 990292
rect 463606 990256 463662 990312
rect 563058 990684 563114 990720
rect 563058 990664 563060 990684
rect 563060 990664 563112 990684
rect 563112 990664 563114 990684
rect 582286 990664 582342 990720
rect 585138 990548 585194 990584
rect 585138 990528 585140 990548
rect 585140 990528 585192 990548
rect 585192 990528 585194 990548
rect 587990 990564 587992 990584
rect 587992 990564 588044 990584
rect 588044 990564 588046 990584
rect 587990 990528 588046 990564
rect 44086 877512 44142 877568
rect 44362 870032 44418 870088
rect 42522 869352 42578 869408
rect 42706 869352 42762 869408
rect 44270 835216 44326 835272
rect 44178 700984 44234 701040
rect 44178 662360 44234 662416
rect 42338 448568 42394 448624
rect 42062 444352 42118 444408
rect 42614 444352 42670 444408
rect 44270 493176 44326 493232
rect 677690 918312 677746 918368
rect 677506 915320 677562 915376
rect 677506 912736 677562 912792
rect 677506 908132 677562 908168
rect 677506 908112 677508 908132
rect 677508 908112 677560 908132
rect 677560 908112 677562 908132
rect 677782 909336 677838 909392
rect 44454 700984 44510 701040
rect 44454 662360 44510 662416
rect 44362 488552 44418 488608
rect 677598 818624 677654 818680
rect 42890 444352 42946 444408
rect 677506 513748 677508 513768
rect 677508 513748 677560 513768
rect 677560 513748 677562 513768
rect 677506 513712 677562 513748
rect 678058 477536 678114 477592
rect 677874 469920 677930 469976
rect 677506 467508 677508 467528
rect 677508 467508 677560 467528
rect 677560 467508 677562 467528
rect 677506 467472 677562 467508
rect 41418 115912 41474 115968
rect 39394 83136 39450 83192
rect 44454 193160 44510 193216
rect 44638 193160 44694 193216
rect 42338 115912 42394 115968
rect 44730 110472 44786 110528
rect 44362 75928 44418 75984
rect 44362 73344 44418 73400
rect 44178 68176 44234 68232
rect 78954 40196 78956 40216
rect 78956 40196 79008 40216
rect 79008 40196 79010 40216
rect 78954 40160 79010 40196
rect 86498 40196 86500 40216
rect 86500 40196 86552 40216
rect 86552 40196 86554 40216
rect 86498 40160 86554 40196
rect 173898 44548 173900 44568
rect 173900 44548 173952 44568
rect 173952 44548 173954 44568
rect 173898 44512 173954 44548
rect 193126 44512 193182 44568
rect 231858 44684 231860 44704
rect 231860 44684 231912 44704
rect 231912 44684 231914 44704
rect 231858 44648 231914 44684
rect 250994 44648 251050 44704
rect 212538 44532 212594 44568
rect 212538 44512 212540 44532
rect 212540 44512 212592 44532
rect 212592 44512 212594 44532
rect 145838 40296 145894 40352
rect 149978 40296 150034 40352
rect 240138 39888 240194 39944
rect 248326 44512 248382 44568
rect 241242 39752 241298 39808
rect 242898 39752 242954 39808
rect 289818 44396 289874 44432
rect 289818 44376 289820 44396
rect 289820 44376 289872 44396
rect 289872 44376 289874 44396
rect 267738 44276 267740 44296
rect 267740 44276 267792 44296
rect 267792 44276 267794 44296
rect 267738 44240 267794 44276
rect 286874 44240 286930 44296
rect 303894 44376 303950 44432
rect 309138 44512 309194 44568
rect 328366 44512 328422 44568
rect 386418 44512 386474 44568
rect 405646 44512 405702 44568
rect 425058 44512 425114 44568
rect 444286 44512 444342 44568
rect 499578 44512 499634 44568
rect 472011 41792 472067 41848
rect 472346 41792 472402 41848
rect 518806 44512 518862 44568
rect 560482 40160 560538 40216
rect 253938 39888 253994 39944
rect 677598 425720 677654 425776
rect 677506 420724 677508 420744
rect 677508 420724 677560 420744
rect 677560 420724 677562 420744
rect 677506 420688 677562 420724
rect 622950 40432 623006 40488
rect 578790 40160 578846 40216
rect 629298 40160 629354 40216
rect 622950 39616 623006 39672
<< metal3 >>
rect 338622 997522 338682 997628
rect 341006 997596 341012 997660
rect 341076 997596 341082 997660
rect 343590 997522 343650 997628
rect 580796 997598 581746 997658
rect 338622 997462 343650 997522
rect 581686 997522 581746 997598
rect 585550 997598 585764 997658
rect 585041 997522 585107 997525
rect 585550 997522 585610 997598
rect 581686 997520 585610 997522
rect 581686 997464 585046 997520
rect 585102 997464 585610 997520
rect 581686 997462 585610 997464
rect 585685 997522 585751 997525
rect 589549 997522 589615 997525
rect 585685 997520 589615 997522
rect 585685 997464 585690 997520
rect 585746 997464 589554 997520
rect 589610 997464 589615 997520
rect 585685 997462 589615 997464
rect 343590 997117 343650 997462
rect 585041 997459 585107 997462
rect 585685 997459 585751 997462
rect 589549 997459 589615 997462
rect 343590 997112 343699 997117
rect 343590 997056 343638 997112
rect 343694 997056 343699 997112
rect 343590 997054 343699 997056
rect 343633 997051 343699 997054
rect 329557 992354 329623 992357
rect 341006 992354 341012 992356
rect 329557 992352 341012 992354
rect 329557 992296 329562 992352
rect 329618 992296 341012 992352
rect 329557 992294 341012 992296
rect 329557 992291 329623 992294
rect 341006 992292 341012 992294
rect 341076 992292 341082 992356
rect 41270 990932 41276 990996
rect 41340 990994 41346 990996
rect 676254 990994 676260 990996
rect 41340 990934 676260 990994
rect 41340 990932 41346 990934
rect 676254 990932 676260 990934
rect 676324 990932 676330 990996
rect 563053 990722 563119 990725
rect 582281 990722 582347 990725
rect 563053 990720 582347 990722
rect 563053 990664 563058 990720
rect 563114 990664 582286 990720
rect 582342 990664 582347 990720
rect 563053 990662 582347 990664
rect 563053 990659 563119 990662
rect 582281 990659 582347 990662
rect 289813 990586 289879 990589
rect 295517 990586 295583 990589
rect 289813 990584 295583 990586
rect 289813 990528 289818 990584
rect 289874 990528 295522 990584
rect 295578 990528 295583 990584
rect 289813 990526 295583 990528
rect 289813 990523 289879 990526
rect 295517 990523 295583 990526
rect 585133 990586 585199 990589
rect 587985 990586 588051 990589
rect 585133 990584 588051 990586
rect 585133 990528 585138 990584
rect 585194 990528 587990 990584
rect 588046 990528 588051 990584
rect 585133 990526 588051 990528
rect 585133 990523 585199 990526
rect 587985 990523 588051 990526
rect 364333 990450 364399 990453
rect 383561 990450 383627 990453
rect 364333 990448 383627 990450
rect 364333 990392 364338 990448
rect 364394 990392 383566 990448
rect 383622 990392 383627 990448
rect 364333 990390 383627 990392
rect 364333 990387 364399 990390
rect 383561 990387 383627 990390
rect 405733 990314 405799 990317
rect 424961 990314 425027 990317
rect 405733 990312 425027 990314
rect 405733 990256 405738 990312
rect 405794 990256 424966 990312
rect 425022 990256 425027 990312
rect 405733 990254 425027 990256
rect 405733 990251 405799 990254
rect 424961 990251 425027 990254
rect 444373 990314 444439 990317
rect 463601 990314 463667 990317
rect 444373 990312 463667 990314
rect 444373 990256 444378 990312
rect 444434 990256 463606 990312
rect 463662 990256 463667 990312
rect 444373 990254 463667 990256
rect 444373 990251 444439 990254
rect 463601 990251 463667 990254
rect 39481 928162 39547 928165
rect 41270 928162 41276 928164
rect 39481 928160 41276 928162
rect 39481 928104 39486 928160
rect 39542 928104 41276 928160
rect 39481 928102 41276 928104
rect 39481 928099 39547 928102
rect 41270 928100 41276 928102
rect 41340 928100 41346 928164
rect 41505 919730 41571 919733
rect 39468 919728 41571 919730
rect 39468 919672 41510 919728
rect 41566 919672 41571 919728
rect 39468 919670 41571 919672
rect 41505 919667 41571 919670
rect 677542 918308 677548 918372
rect 677612 918370 677618 918372
rect 677685 918370 677751 918373
rect 677612 918368 677751 918370
rect 677612 918312 677690 918368
rect 677746 918312 677751 918368
rect 677612 918310 677751 918312
rect 677612 918308 677618 918310
rect 677685 918307 677751 918310
rect 41505 917282 41571 917285
rect 39468 917280 41571 917282
rect 39468 917224 41510 917280
rect 41566 917224 41571 917280
rect 39468 917222 41571 917224
rect 41505 917219 41571 917222
rect 677501 915378 677567 915381
rect 677501 915376 678132 915378
rect 677501 915320 677506 915376
rect 677562 915320 678132 915376
rect 677501 915318 678132 915320
rect 677501 915315 677567 915318
rect 677501 912794 677567 912797
rect 677501 912792 678132 912794
rect 677501 912736 677506 912792
rect 677562 912736 678132 912792
rect 677501 912734 678132 912736
rect 677501 912731 677567 912734
rect 41505 912250 41571 912253
rect 39468 912248 41571 912250
rect 39468 912192 41510 912248
rect 41566 912192 41571 912248
rect 39468 912190 41571 912192
rect 41505 912187 41571 912190
rect 677542 909332 677548 909396
rect 677612 909394 677618 909396
rect 677777 909394 677843 909397
rect 677612 909392 677843 909394
rect 677612 909336 677782 909392
rect 677838 909336 677843 909392
rect 677612 909334 677843 909336
rect 677612 909332 677618 909334
rect 677777 909331 677843 909334
rect 39573 908170 39639 908173
rect 40166 908170 40172 908172
rect 39573 908168 40172 908170
rect 39573 908112 39578 908168
rect 39634 908112 40172 908168
rect 39573 908110 40172 908112
rect 39573 908107 39639 908110
rect 40166 908108 40172 908110
rect 40236 908108 40242 908172
rect 677501 908170 677567 908173
rect 677501 908168 678162 908170
rect 677501 908112 677506 908168
rect 677562 908112 678162 908168
rect 677501 908110 678162 908112
rect 677501 908107 677567 908110
rect 40033 908034 40099 908037
rect 40166 908034 40172 908036
rect 40033 908032 40172 908034
rect 40033 907976 40038 908032
rect 40094 907976 40172 908032
rect 40033 907974 40172 907976
rect 40033 907971 40099 907974
rect 40166 907972 40172 907974
rect 40236 907972 40242 908036
rect 678102 907732 678162 908110
rect 40033 888994 40099 888997
rect 39806 888992 40099 888994
rect 39806 888936 40038 888992
rect 40094 888936 40099 888992
rect 39806 888934 40099 888936
rect 39806 888860 39866 888934
rect 40033 888931 40099 888934
rect 39798 888796 39804 888860
rect 39868 888796 39874 888860
rect 40125 877570 40191 877573
rect 44081 877570 44147 877573
rect 39622 877568 44147 877570
rect 39622 877512 40130 877568
rect 40186 877512 44086 877568
rect 44142 877512 44147 877568
rect 39622 877510 44147 877512
rect 39622 877404 39682 877510
rect 40125 877507 40191 877510
rect 44081 877507 44147 877510
rect 41413 875122 41479 875125
rect 39652 875120 41479 875122
rect 39652 875064 41418 875120
rect 41474 875064 41479 875120
rect 39652 875062 41479 875064
rect 41413 875059 41479 875062
rect 40125 870090 40191 870093
rect 44357 870090 44423 870093
rect 39622 870088 44423 870090
rect 39622 870032 40130 870088
rect 40186 870032 44362 870088
rect 44418 870032 44423 870088
rect 39622 870030 44423 870032
rect 39622 869924 39682 870030
rect 40125 870027 40191 870030
rect 44357 870027 44423 870030
rect 39849 869410 39915 869413
rect 40166 869410 40172 869412
rect 39849 869408 40172 869410
rect 39849 869352 39854 869408
rect 39910 869352 40172 869408
rect 39849 869350 40172 869352
rect 39849 869347 39915 869350
rect 40166 869348 40172 869350
rect 40236 869348 40242 869412
rect 42517 869410 42583 869413
rect 42701 869410 42767 869413
rect 42517 869408 42767 869410
rect 42517 869352 42522 869408
rect 42578 869352 42706 869408
rect 42762 869352 42767 869408
rect 42517 869350 42767 869352
rect 42517 869347 42583 869350
rect 42701 869347 42767 869350
rect 39849 850370 39915 850373
rect 39806 850368 39915 850370
rect 39806 850312 39854 850368
rect 39910 850312 39915 850368
rect 39806 850307 39915 850312
rect 39806 850236 39866 850307
rect 39798 850172 39804 850236
rect 39868 850172 39874 850236
rect 44265 835274 44331 835277
rect 39652 835272 44331 835274
rect 39652 835216 44270 835272
rect 44326 835216 44331 835272
rect 39652 835214 44331 835216
rect 44265 835211 44331 835214
rect 39652 827734 39866 827794
rect 39806 827525 39866 827734
rect 39757 827520 39866 827525
rect 39757 827464 39762 827520
rect 39818 827464 39866 827520
rect 39757 827462 39866 827464
rect 39757 827459 39823 827462
rect 677593 818682 677659 818685
rect 677593 818680 677764 818682
rect 677593 818624 677598 818680
rect 677654 818624 677764 818680
rect 677593 818622 677764 818624
rect 677593 818619 677659 818622
rect 44173 701042 44239 701045
rect 44449 701042 44515 701045
rect 44173 701040 44515 701042
rect 44173 700984 44178 701040
rect 44234 700984 44454 701040
rect 44510 700984 44515 701040
rect 44173 700982 44515 700984
rect 44173 700979 44239 700982
rect 44449 700979 44515 700982
rect 44173 662418 44239 662421
rect 44449 662418 44515 662421
rect 44173 662416 44515 662418
rect 44173 662360 44178 662416
rect 44234 662360 44454 662416
rect 44510 662360 44515 662416
rect 44173 662358 44515 662360
rect 44173 662355 44239 662358
rect 44449 662355 44515 662358
rect 40217 516084 40283 516085
rect 40166 516020 40172 516084
rect 40236 516082 40283 516084
rect 40236 516080 40328 516082
rect 40278 516024 40328 516080
rect 40236 516022 40328 516024
rect 40236 516020 40283 516022
rect 40217 516019 40283 516020
rect 677501 513770 677567 513773
rect 677734 513770 677794 514012
rect 677501 513768 677794 513770
rect 677501 513712 677506 513768
rect 677562 513712 677794 513768
rect 677501 513710 677794 513712
rect 677501 513707 677567 513710
rect 40217 497042 40283 497045
rect 40174 497040 40283 497042
rect 40174 496984 40222 497040
rect 40278 496984 40283 497040
rect 40174 496979 40283 496984
rect 40174 496908 40234 496979
rect 40166 496844 40172 496908
rect 40236 496844 40242 496908
rect 44265 493234 44331 493237
rect 39652 493232 44331 493234
rect 39652 493176 44270 493232
rect 44326 493176 44331 493232
rect 39652 493174 44331 493176
rect 39806 492965 39866 493174
rect 44265 493171 44331 493174
rect 39757 492960 39866 492965
rect 39757 492904 39762 492960
rect 39818 492904 39866 492960
rect 39757 492902 39866 492904
rect 39757 492899 39823 492902
rect 39849 490514 39915 490517
rect 40166 490514 40172 490516
rect 39849 490512 40172 490514
rect 39849 490456 39854 490512
rect 39910 490456 40172 490512
rect 39849 490454 40172 490456
rect 39849 490451 39915 490454
rect 40166 490452 40172 490454
rect 40236 490452 40242 490516
rect 44357 488610 44423 488613
rect 39806 488608 44423 488610
rect 39806 488552 44362 488608
rect 44418 488552 44423 488608
rect 39806 488550 44423 488552
rect 39806 488338 39866 488550
rect 44357 488547 44423 488550
rect 39652 488278 39866 488338
rect 39849 488068 39915 488069
rect 39798 488066 39804 488068
rect 39758 488006 39804 488066
rect 39868 488064 39915 488068
rect 39910 488008 39915 488064
rect 39798 488004 39804 488006
rect 39868 488004 39915 488008
rect 39849 488003 39915 488004
rect 677542 477532 677548 477596
rect 677612 477594 677618 477596
rect 678053 477594 678119 477597
rect 677612 477592 678119 477594
rect 677612 477536 678058 477592
rect 678114 477536 678119 477592
rect 677612 477534 678119 477536
rect 677612 477532 677618 477534
rect 678053 477531 678119 477534
rect 39798 470596 39804 470660
rect 39868 470658 39874 470660
rect 40033 470658 40099 470661
rect 39868 470656 40099 470658
rect 39868 470600 40038 470656
rect 40094 470600 40099 470656
rect 39868 470598 40099 470600
rect 39868 470596 39874 470598
rect 40033 470595 40099 470598
rect 677869 469978 677935 469981
rect 677869 469976 678132 469978
rect 677869 469920 677874 469976
rect 677930 469920 678132 469976
rect 677869 469918 678132 469920
rect 677869 469915 677935 469918
rect 677501 467530 677567 467533
rect 677501 467528 678132 467530
rect 677501 467472 677506 467528
rect 677562 467500 678132 467528
rect 677562 467472 678162 467500
rect 677501 467470 678162 467472
rect 677501 467467 677567 467470
rect 678102 465052 678162 467470
rect 40033 461004 40099 461005
rect 39982 460940 39988 461004
rect 40052 461002 40099 461004
rect 40052 461000 40144 461002
rect 40094 460944 40144 461000
rect 40052 460942 40144 460944
rect 40052 460940 40099 460942
rect 40033 460939 40099 460940
rect 39941 455428 40007 455429
rect 39941 455426 39988 455428
rect 39896 455424 39988 455426
rect 39896 455368 39946 455424
rect 39896 455366 39988 455368
rect 39941 455364 39988 455366
rect 40052 455364 40058 455428
rect 39941 455363 40007 455364
rect 39665 451890 39731 451893
rect 40166 451890 40172 451892
rect 39665 451888 40172 451890
rect 39665 451832 39670 451888
rect 39726 451832 40172 451888
rect 39665 451830 40172 451832
rect 39665 451827 39731 451830
rect 40166 451828 40172 451830
rect 40236 451828 40242 451892
rect 42333 448626 42399 448629
rect 39468 448624 42399 448626
rect 39468 448596 42338 448624
rect 39438 448568 42338 448596
rect 42394 448568 42399 448624
rect 39438 448566 42399 448568
rect 39438 446012 39498 448566
rect 42333 448563 42399 448566
rect 39849 444410 39915 444413
rect 42057 444410 42123 444413
rect 39849 444408 42123 444410
rect 39849 444352 39854 444408
rect 39910 444352 42062 444408
rect 42118 444352 42123 444408
rect 39849 444350 42123 444352
rect 39849 444347 39915 444350
rect 42057 444347 42123 444350
rect 42609 444410 42675 444413
rect 42885 444410 42951 444413
rect 42609 444408 42951 444410
rect 42609 444352 42614 444408
rect 42670 444352 42890 444408
rect 42946 444352 42951 444408
rect 42609 444350 42951 444352
rect 42609 444347 42675 444350
rect 42885 444347 42951 444350
rect 39665 441010 39731 441013
rect 39468 441008 39731 441010
rect 39468 440952 39670 441008
rect 39726 440952 39731 441008
rect 39468 440950 39731 440952
rect 39665 440947 39731 440950
rect 677593 425778 677659 425781
rect 677593 425776 677764 425778
rect 677593 425720 677598 425776
rect 677654 425720 677764 425776
rect 677593 425718 677764 425720
rect 677593 425715 677659 425718
rect 677501 420746 677567 420749
rect 677734 420746 677794 420852
rect 677501 420744 677794 420746
rect 677501 420688 677506 420744
rect 677562 420688 677794 420744
rect 677501 420686 677794 420688
rect 677501 420683 677567 420686
rect 44449 193218 44515 193221
rect 44633 193218 44699 193221
rect 44449 193216 44699 193218
rect 44449 193160 44454 193216
rect 44510 193160 44638 193216
rect 44694 193160 44699 193216
rect 44449 193158 44699 193160
rect 44449 193155 44515 193158
rect 44633 193155 44699 193158
rect 41413 115970 41479 115973
rect 42333 115970 42399 115973
rect 39806 115968 42399 115970
rect 39806 115912 41418 115968
rect 41474 115912 42338 115968
rect 42394 115912 42399 115968
rect 39806 115910 42399 115912
rect 39806 115562 39866 115910
rect 41413 115907 41479 115910
rect 42333 115907 42399 115910
rect 39622 115502 39866 115562
rect 39622 115396 39682 115502
rect 44725 110530 44791 110533
rect 39806 110528 44791 110530
rect 39806 110472 44730 110528
rect 44786 110472 44791 110528
rect 39806 110470 44791 110472
rect 39806 110430 39866 110470
rect 44725 110467 44791 110470
rect 39622 110370 39866 110430
rect 39622 110364 39682 110370
rect 39389 83194 39455 83197
rect 40166 83194 40172 83196
rect 39389 83192 40172 83194
rect 39389 83136 39394 83192
rect 39450 83136 40172 83192
rect 39389 83134 40172 83136
rect 39389 83131 39455 83134
rect 40166 83132 40172 83134
rect 40236 83132 40242 83196
rect 44357 75986 44423 75989
rect 39438 75984 44423 75986
rect 39438 75928 44362 75984
rect 44418 75928 44423 75984
rect 39438 75926 44423 75928
rect 39438 75684 39498 75926
rect 44357 75923 44423 75926
rect 44357 73402 44423 73405
rect 39438 73400 44423 73402
rect 39438 73344 44362 73400
rect 44418 73344 44423 73400
rect 39438 73342 44423 73344
rect 39438 73236 39498 73342
rect 44357 73339 44423 73342
rect 44173 68234 44239 68237
rect 39468 68232 44239 68234
rect 39468 68176 44178 68232
rect 44234 68176 44239 68232
rect 39468 68174 44239 68176
rect 44173 68171 44239 68174
rect 231853 44706 231919 44709
rect 250989 44706 251055 44709
rect 231853 44704 251055 44706
rect 231853 44648 231858 44704
rect 231914 44648 250994 44704
rect 251050 44648 251055 44704
rect 231853 44646 251055 44648
rect 231853 44643 231919 44646
rect 250989 44643 251055 44646
rect 173893 44570 173959 44573
rect 193121 44570 193187 44573
rect 173893 44568 193187 44570
rect 173893 44512 173898 44568
rect 173954 44512 193126 44568
rect 193182 44512 193187 44568
rect 173893 44510 193187 44512
rect 173893 44507 173959 44510
rect 193121 44507 193187 44510
rect 212533 44570 212599 44573
rect 248321 44570 248387 44573
rect 212533 44568 248387 44570
rect 212533 44512 212538 44568
rect 212594 44512 248326 44568
rect 248382 44512 248387 44568
rect 212533 44510 248387 44512
rect 212533 44507 212599 44510
rect 248321 44507 248387 44510
rect 309133 44570 309199 44573
rect 328361 44570 328427 44573
rect 309133 44568 328427 44570
rect 309133 44512 309138 44568
rect 309194 44512 328366 44568
rect 328422 44512 328427 44568
rect 309133 44510 328427 44512
rect 309133 44507 309199 44510
rect 328361 44507 328427 44510
rect 386413 44570 386479 44573
rect 405641 44570 405707 44573
rect 386413 44568 405707 44570
rect 386413 44512 386418 44568
rect 386474 44512 405646 44568
rect 405702 44512 405707 44568
rect 386413 44510 405707 44512
rect 386413 44507 386479 44510
rect 405641 44507 405707 44510
rect 425053 44570 425119 44573
rect 444281 44570 444347 44573
rect 425053 44568 444347 44570
rect 425053 44512 425058 44568
rect 425114 44512 444286 44568
rect 444342 44512 444347 44568
rect 425053 44510 444347 44512
rect 425053 44507 425119 44510
rect 444281 44507 444347 44510
rect 499573 44570 499639 44573
rect 518801 44570 518867 44573
rect 499573 44568 518867 44570
rect 499573 44512 499578 44568
rect 499634 44512 518806 44568
rect 518862 44512 518867 44568
rect 499573 44510 518867 44512
rect 499573 44507 499639 44510
rect 518801 44507 518867 44510
rect 289813 44434 289879 44437
rect 303889 44434 303955 44437
rect 289813 44432 303955 44434
rect 289813 44376 289818 44432
rect 289874 44376 303894 44432
rect 303950 44376 303955 44432
rect 289813 44374 303955 44376
rect 289813 44371 289879 44374
rect 303889 44371 303955 44374
rect 267733 44298 267799 44301
rect 286869 44298 286935 44301
rect 267733 44296 286935 44298
rect 267733 44240 267738 44296
rect 267794 44240 286874 44296
rect 286930 44240 286935 44296
rect 267733 44238 286935 44240
rect 267733 44235 267799 44238
rect 286869 44235 286935 44238
rect 472006 41850 472072 41853
rect 472341 41850 472407 41853
rect 472006 41848 472407 41850
rect 472006 41792 472011 41848
rect 472067 41792 472346 41848
rect 472402 41792 472407 41848
rect 472006 41790 472407 41792
rect 472006 41787 472072 41790
rect 472341 41787 472407 41790
rect 622945 40490 623011 40493
rect 84334 40488 623011 40490
rect 84334 40432 622950 40488
rect 623006 40432 623011 40488
rect 84334 40430 623011 40432
rect 78949 40218 79015 40221
rect 84334 40218 84394 40430
rect 622945 40427 623011 40430
rect 145833 40354 145899 40357
rect 149973 40354 150039 40357
rect 145708 40352 150039 40354
rect 145708 40296 145838 40352
rect 145894 40296 149978 40352
rect 150034 40296 150039 40352
rect 145708 40294 150039 40296
rect 145833 40291 145899 40294
rect 149973 40291 150039 40294
rect 78949 40216 79058 40218
rect 78949 40160 78954 40216
rect 79010 40160 79058 40216
rect 78949 40155 79058 40160
rect 78998 39644 79058 40155
rect 84150 40158 84394 40218
rect 86493 40218 86559 40221
rect 86493 40216 86602 40218
rect 86493 40160 86498 40216
rect 86554 40160 86602 40216
rect 84150 39644 84210 40158
rect 86493 40155 86602 40160
rect 86542 39644 86602 40155
rect 141667 38031 141813 39999
rect 145838 39967 145898 40291
rect 560477 40218 560543 40221
rect 578785 40218 578851 40221
rect 560477 40216 578851 40218
rect 560477 40160 560482 40216
rect 560538 40160 578790 40216
rect 578846 40160 578851 40216
rect 560477 40158 578851 40160
rect 560477 40155 560543 40158
rect 240133 39946 240199 39949
rect 253933 39946 253999 39949
rect 240133 39944 246498 39946
rect 240133 39888 240138 39944
rect 240194 39888 246498 39944
rect 240133 39886 246498 39888
rect 240133 39883 240199 39886
rect 241237 39810 241303 39813
rect 242893 39810 242959 39813
rect 241156 39808 242959 39810
rect 241156 39752 241242 39808
rect 241298 39752 242898 39808
rect 242954 39752 242959 39808
rect 241156 39750 242959 39752
rect 241237 39747 241346 39750
rect 242893 39747 242959 39750
rect 241286 39372 241346 39747
rect 246438 39538 246498 39886
rect 248830 39944 253999 39946
rect 248830 39888 253938 39944
rect 253994 39888 253999 39944
rect 248830 39886 253999 39888
rect 248830 39538 248890 39886
rect 253933 39883 253999 39886
rect 569174 39644 569234 40158
rect 576718 39644 576778 40158
rect 578785 40155 578851 40158
rect 629293 40218 629359 40221
rect 629293 40216 630506 40218
rect 629293 40160 629298 40216
rect 629354 40160 630506 40216
rect 629293 40158 630506 40160
rect 629293 40155 629359 40158
rect 622945 39674 623011 39677
rect 622945 39672 623116 39674
rect 622945 39616 622950 39672
rect 623006 39616 623116 39672
rect 630446 39644 630506 40158
rect 622945 39614 623116 39616
rect 622945 39611 623011 39614
rect 246438 39478 248890 39538
rect 246438 39372 246498 39478
rect 248830 39372 248890 39478
<< via3 >>
rect 341012 997596 341076 997660
rect 341012 992292 341076 992356
rect 41276 990932 41340 990996
rect 676260 990932 676324 990996
rect 41276 928100 41340 928164
rect 677548 918308 677612 918372
rect 677548 909332 677612 909396
rect 40172 908108 40236 908172
rect 40172 907972 40236 908036
rect 39804 888796 39868 888860
rect 40172 869348 40236 869412
rect 39804 850172 39868 850236
rect 40172 516080 40236 516084
rect 40172 516024 40222 516080
rect 40222 516024 40236 516080
rect 40172 516020 40236 516024
rect 40172 496844 40236 496908
rect 40172 490452 40236 490516
rect 39804 488064 39868 488068
rect 39804 488008 39854 488064
rect 39854 488008 39868 488064
rect 39804 488004 39868 488008
rect 677548 477532 677612 477596
rect 39804 470596 39868 470660
rect 39988 461000 40052 461004
rect 39988 460944 40038 461000
rect 40038 460944 40052 461000
rect 39988 460940 40052 460944
rect 39988 455424 40052 455428
rect 39988 455368 40002 455424
rect 40002 455368 40052 455424
rect 39988 455364 40052 455368
rect 40172 451828 40236 451892
rect 40172 83132 40236 83196
<< metal4 >>
rect 341011 997660 341077 997661
rect 341011 997596 341012 997660
rect 341076 997596 341077 997660
rect 341011 997595 341077 997596
rect 341014 992357 341074 997595
rect 341011 992356 341077 992357
rect 341011 992292 341012 992356
rect 341076 992292 341077 992356
rect 341011 992291 341077 992292
rect 41275 990996 41341 990997
rect 41275 990932 41276 990996
rect 41340 990932 41341 990996
rect 41275 990931 41341 990932
rect 676259 990996 676325 990997
rect 676259 990932 676260 990996
rect 676324 990932 676325 990996
rect 676259 990931 676325 990932
rect 41278 928165 41338 990931
rect 41275 928164 41341 928165
rect 41275 928100 41276 928164
rect 41340 928100 41341 928164
rect 41275 928099 41341 928100
rect 676262 918370 676322 990931
rect 677547 918372 677613 918373
rect 677547 918370 677548 918372
rect 676262 918310 677548 918370
rect 677547 918308 677548 918310
rect 677612 918308 677613 918372
rect 677547 918307 677613 918308
rect 677547 909396 677613 909397
rect 677547 909332 677548 909396
rect 677612 909332 677613 909396
rect 677547 909331 677613 909332
rect 40171 908172 40237 908173
rect 40171 908108 40172 908172
rect 40236 908108 40237 908172
rect 40171 908107 40237 908108
rect 40174 908037 40234 908107
rect 40171 908036 40237 908037
rect 40171 907972 40172 908036
rect 40236 907972 40237 908036
rect 40171 907971 40237 907972
rect 39803 888860 39869 888861
rect 39803 888796 39804 888860
rect 39868 888796 39869 888860
rect 39803 888795 39869 888796
rect 39806 874850 39866 888795
rect 39806 874790 40234 874850
rect 40174 869413 40234 874790
rect 40171 869412 40237 869413
rect 40171 869348 40172 869412
rect 40236 869348 40237 869412
rect 40171 869347 40237 869348
rect 39803 850236 39869 850237
rect 39803 850172 39804 850236
rect 39868 850172 39869 850236
rect 39803 850171 39869 850172
rect 39806 836090 39866 850171
rect 39806 836030 40050 836090
rect 39990 811610 40050 836030
rect 39990 811550 40418 811610
rect 40358 808210 40418 811550
rect 40358 808150 40602 808210
rect 40542 791890 40602 808150
rect 40542 791830 40786 791890
rect 40726 770130 40786 791830
rect 40358 770070 40786 770130
rect 40358 747098 40418 770070
rect 40174 731458 40234 746182
rect 40910 712330 40970 731222
rect 40358 712270 40970 712330
rect 40358 695330 40418 712270
rect 40358 695270 40602 695330
rect 40542 676290 40602 695270
rect 40358 676230 40602 676290
rect 40358 662778 40418 676230
rect 41462 651130 41522 662542
rect 41094 651070 41522 651130
rect 41094 632090 41154 651070
rect 40174 632030 41154 632090
rect 40174 628098 40234 632030
rect 41094 612370 41154 627862
rect 40542 612310 41154 612370
rect 40542 598770 40602 612310
rect 40358 598710 40602 598770
rect 40358 567490 40418 598710
rect 40358 567430 40602 567490
rect 40542 545050 40602 567430
rect 40358 544990 40602 545050
rect 40358 528730 40418 544990
rect 40174 528670 40418 528730
rect 40174 516085 40234 528670
rect 40171 516084 40237 516085
rect 40171 516020 40172 516084
rect 40236 516020 40237 516084
rect 40171 516019 40237 516020
rect 40171 496908 40237 496909
rect 40171 496844 40172 496908
rect 40236 496844 40237 496908
rect 40171 496843 40237 496844
rect 40174 490517 40234 496843
rect 40171 490516 40237 490517
rect 40171 490452 40172 490516
rect 40236 490452 40237 490516
rect 40171 490451 40237 490452
rect 39803 488068 39869 488069
rect 39803 488004 39804 488068
rect 39868 488004 39869 488068
rect 39803 488003 39869 488004
rect 39806 470661 39866 488003
rect 677550 477597 677610 909331
rect 677547 477596 677613 477597
rect 677547 477532 677548 477596
rect 677612 477532 677613 477596
rect 677547 477531 677613 477532
rect 39803 470660 39869 470661
rect 39803 470596 39804 470660
rect 39868 470596 39869 470660
rect 39803 470595 39869 470596
rect 39987 461004 40053 461005
rect 39987 460940 39988 461004
rect 40052 460940 40053 461004
rect 39987 460939 40053 460940
rect 39990 455429 40050 460939
rect 39987 455428 40053 455429
rect 39987 455364 39988 455428
rect 40052 455364 40053 455428
rect 39987 455363 40053 455364
rect 40171 451892 40237 451893
rect 40171 451828 40172 451892
rect 40236 451828 40237 451892
rect 40171 451827 40237 451828
rect 40174 83197 40234 451827
rect 40171 83196 40237 83197
rect 40171 83132 40172 83196
rect 40236 83132 40237 83196
rect 40171 83131 40237 83132
<< via4 >>
rect 40270 746862 40506 747098
rect 40086 746182 40322 746418
rect 40086 731222 40322 731458
rect 40822 731222 41058 731458
rect 40270 662542 40506 662778
rect 41374 662542 41610 662778
rect 40086 627862 40322 628098
rect 41006 627862 41242 628098
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334620 1018402 347160 1030924
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 576820 1018402 589360 1030924
rect 628240 1018512 640760 1031002
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6086 913863 19572 925191
rect 698028 909409 711514 920737
rect 698512 863640 711002 876160
rect 6675 828820 19197 841360
rect 698402 819640 710924 832180
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 40044 747098 40548 747140
rect 40044 746862 40270 747098
rect 40506 746862 40548 747098
rect 40044 746820 40548 746862
rect 40044 746418 40364 746820
rect 40044 746182 40086 746418
rect 40322 746182 40364 746418
rect 40044 746140 40364 746182
rect 40044 731458 41100 731500
rect 40044 731222 40086 731458
rect 40322 731222 40822 731458
rect 41058 731222 41100 731458
rect 40044 731180 41100 731222
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 40228 662778 41652 662820
rect 40228 662542 40270 662778
rect 40506 662542 41374 662778
rect 41610 662542 41652 662778
rect 40228 662500 41652 662542
rect 698512 639240 711002 651760
rect 40044 628098 41284 628140
rect 40044 627862 40086 628098
rect 40322 627862 41006 628098
rect 41242 627862 41284 628098
rect 40044 627820 41284 627862
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 6675 484220 19197 496760
rect 698028 461609 711514 472937
rect 6086 442663 19572 453991
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6675 111420 19197 123960
rect 698512 101240 711002 113760
rect 6086 69863 19572 81191
rect 80040 6675 92580 19197
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243009 6086 254337 19572
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 624040 6675 636580 19197
use sky130_ef_io__corner_pad  mgmt_corner\[0\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_177 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_381
timestamp 1607115945
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1607115945
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1
timestamp 1607115945
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_181 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_180
timestamp 1607115945
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_179 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_178 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_188
timestamp 1607115945
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1607115945
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1607115945
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1607115945
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_192
timestamp 1607115945
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_191
timestamp 1607115945
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_190
timestamp 1607115945
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_189
timestamp 1607115945
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__vssa_hvc_pad  mgmt_vssa_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 93800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_194
timestamp 1607115945
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_196
timestamp 1607115945
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_195
timestamp 1607115945
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1607115945
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_198
timestamp 1607115945
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_197
timestamp 1607115945
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1607115945
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1607115945
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1607115945
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1607115945
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1607115945
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_205
timestamp 1607115945
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_209
timestamp 1607115945
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_208
timestamp 1607115945
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_207
timestamp 1607115945
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_206
timestamp 1607115945
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_fd_io__top_xres4v2  resetb_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 147600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1607115945
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_215
timestamp 1607115945
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_214
timestamp 1607115945
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_213
timestamp 1607115945
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_212
timestamp 1607115945
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_211
timestamp 1607115945
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1607115945
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1607115945
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1607115945
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_224
timestamp 1607115945
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_223
timestamp 1607115945
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_222
timestamp 1607115945
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1607115945
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1607115945
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_226
timestamp 1607115945
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_225
timestamp 1607115945
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 202400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1607115945
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_232
timestamp 1607115945
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_231
timestamp 1607115945
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_230
timestamp 1607115945
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_229
timestamp 1607115945
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_228
timestamp 1607115945
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1607115945
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1607115945
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1607115945
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1607115945
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_242
timestamp 1607115945
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_241
timestamp 1607115945
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_240
timestamp 1607115945
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_239
timestamp 1607115945
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1607115945
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_243
timestamp 1607115945
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__vssd_lvc_pad  mgmt_vssd_lvclmap_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 256200 0 -1 39593
box 0 -7 15000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1607115945
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1607115945
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_249
timestamp 1607115945
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_248
timestamp 1607115945
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_247
timestamp 1607115945
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_246
timestamp 1607115945
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_245
timestamp 1607115945
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1607115945
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1607115945
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1607115945
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1607115945
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_260
timestamp 1607115945
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_259
timestamp 1607115945
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_258
timestamp 1607115945
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_257
timestamp 1607115945
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_256
timestamp 1607115945
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1607115945
transform -1 0 311000 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_262
timestamp 1607115945
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_263
timestamp 1607115945
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1607115945
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_266
timestamp 1607115945
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_265
timestamp 1607115945
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_264
timestamp 1607115945
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1607115945
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1607115945
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1607115945
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1607115945
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_277
timestamp 1607115945
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_276
timestamp 1607115945
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_275
timestamp 1607115945
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_274
timestamp 1607115945
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_273
timestamp 1607115945
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1607115945
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1607115945
transform -1 0 365800 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_280
timestamp 1607115945
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_279
timestamp 1607115945
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1607115945
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1607115945
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_283
timestamp 1607115945
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_282
timestamp 1607115945
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_281
timestamp 1607115945
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1607115945
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1607115945
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1607115945
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1607115945
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_294
timestamp 1607115945
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_293
timestamp 1607115945
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_292
timestamp 1607115945
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_291
timestamp 1607115945
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_290
timestamp 1607115945
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1607115945
transform -1 0 420600 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_296
timestamp 1607115945
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1607115945
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1607115945
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1607115945
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_300
timestamp 1607115945
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_299
timestamp 1607115945
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_298
timestamp 1607115945
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_297
timestamp 1607115945
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_307
timestamp 1607115945
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1607115945
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1607115945
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1607115945
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_311
timestamp 1607115945
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_310
timestamp 1607115945
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_309
timestamp 1607115945
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_308
timestamp 1607115945
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1607115945
transform -1 0 475400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_313
timestamp 1607115945
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_314
timestamp 1607115945
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1607115945
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_317
timestamp 1607115945
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_316
timestamp 1607115945
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_315
timestamp 1607115945
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1607115945
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1607115945
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1607115945
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1607115945
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1607115945
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_328
timestamp 1607115945
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_327
timestamp 1607115945
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_326
timestamp 1607115945
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_325
timestamp 1607115945
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_324
timestamp 1607115945
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1607115945
transform -1 0 530200 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1607115945
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_334
timestamp 1607115945
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_333
timestamp 1607115945
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_332
timestamp 1607115945
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_331
timestamp 1607115945
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_330
timestamp 1607115945
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1607115945
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1607115945
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_341
timestamp 1607115945
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1607115945
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1607115945
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1607115945
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_345
timestamp 1607115945
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_344
timestamp 1607115945
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_343
timestamp 1607115945
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_342
timestamp 1607115945
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__vssio_hvc_pad  mgmt_vssio_hvclamp_pad\[1\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 584000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_349
timestamp 1607115945
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_348
timestamp 1607115945
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_347
timestamp 1607115945
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1607115945
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1607115945
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1607115945
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1607115945
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_351
timestamp 1607115945
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_350
timestamp 1607115945
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_359
timestamp 1607115945
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_358
timestamp 1607115945
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1607115945
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1607115945
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_362
timestamp 1607115945
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_361
timestamp 1607115945
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_360
timestamp 1607115945
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__vdda_hvc_pad  mgmt_vdda_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_364
timestamp 1607115945
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_367
timestamp 1607115945
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_366
timestamp 1607115945
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_365
timestamp 1607115945
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1607115945
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_368
timestamp 1607115945
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1607115945
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1607115945
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1607115945
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1607115945
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1607115945
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1607115945
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_376
timestamp 1607115945
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1607115945
transform 0 1 676800 -1 0 40000
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_5um  FILLER_377
timestamp 1607115945
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_378
timestamp 1607115945
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_379
timestamp 1607115945
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_380
timestamp 1607115945
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_612
timestamp 1607115945
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_385
timestamp 1607115945
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1607115945
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_383
timestamp 1607115945
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_382
timestamp 1607115945
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_389
timestamp 1607115945
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_388
timestamp 1607115945
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_387
timestamp 1607115945
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_386
timestamp 1607115945
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  mgmt_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform 0 -1 39593 1 0 68000
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_391
timestamp 1607115945
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_613
timestamp 1607115945
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_614
timestamp 1607115945
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1607115945
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_616
timestamp 1607115945
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_617
timestamp 1607115945
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1607115945
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_1 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform 0 1 678007 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform 0 1 678007 -1 0 70000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_619
timestamp 1607115945
transform 0 1 678007 -1 0 69000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_622
timestamp 1607115945
transform 0 1 678007 -1 0 75000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_623
timestamp 1607115945
transform 0 1 678007 -1 0 79000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1607115945
transform 0 1 678007 -1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_625
timestamp 1607115945
transform 0 1 678007 -1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_395
timestamp 1607115945
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1607115945
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_393
timestamp 1607115945
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_392
timestamp 1607115945
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_399
timestamp 1607115945
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_398
timestamp 1607115945
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_397
timestamp 1607115945
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_396
timestamp 1607115945
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_pad  mgmt_vddio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1607115945
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_401
timestamp 1607115945
transform 0 -1 39593 1 0 125200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[0\]
timestamp 1607115945
transform 0 1 675407 -1 0 116000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_626
timestamp 1607115945
transform 0 1 678007 -1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_627
timestamp 1607115945
transform 0 1 678007 -1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1607115945
transform 0 1 678007 -1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_629
timestamp 1607115945
transform 0 1 678007 -1 0 100000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_631
timestamp 1607115945
transform 0 1 678007 -1 0 120000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_632
timestamp 1607115945
transform 0 1 678007 -1 0 124000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_633
timestamp 1607115945
transform 0 1 678007 -1 0 128000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_402
timestamp 1607115945
transform 0 -1 39593 1 0 129200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_403
timestamp 1607115945
transform 0 -1 39593 1 0 133200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_404
timestamp 1607115945
transform 0 -1 39593 1 0 137200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1607115945
transform 0 -1 39593 1 0 141200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_406
timestamp 1607115945
transform 0 -1 39593 1 0 145200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_407
timestamp 1607115945
transform 0 -1 39593 1 0 149200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_412
timestamp 1607115945
transform 0 -1 39593 1 0 154400
box 0 0 4000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_2
timestamp 1607115945
transform 0 -1 39593 1 0 153400
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1607115945
transform 0 -1 39593 1 0 152400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_409
timestamp 1607115945
transform 0 -1 39593 1 0 152200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_408
timestamp 1607115945
transform 0 -1 39593 1 0 151200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_413
timestamp 1607115945
transform 0 -1 39593 1 0 158400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_414
timestamp 1607115945
transform 0 -1 39593 1 0 162400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1607115945
transform 0 -1 39593 1 0 166400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[1\]
timestamp 1607115945
transform 0 1 675407 -1 0 161200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1607115945
transform 0 1 678007 -1 0 132000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_635
timestamp 1607115945
transform 0 1 678007 -1 0 136000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_636
timestamp 1607115945
transform 0 1 678007 -1 0 140000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1607115945
transform 0 1 678007 -1 0 144000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_638
timestamp 1607115945
transform 0 1 678007 -1 0 145000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_639
timestamp 1607115945
transform 0 1 678007 -1 0 145200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_641
timestamp 1607115945
transform 0 1 678007 -1 0 165200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_642
timestamp 1607115945
transform 0 1 678007 -1 0 169200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_420
timestamp 1607115945
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_419
timestamp 1607115945
transform 0 -1 39593 1 0 180400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_418
timestamp 1607115945
transform 0 -1 39593 1 0 178400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_417
timestamp 1607115945
transform 0 -1 39593 1 0 174400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1607115945
transform 0 -1 39593 1 0 170400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[19\]
timestamp 1607115945
transform 0 -1 42193 1 0 181600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_422
timestamp 1607115945
transform 0 -1 39593 1 0 197600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1607115945
transform 0 -1 39593 1 0 209600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_424
timestamp 1607115945
transform 0 -1 39593 1 0 205600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_423
timestamp 1607115945
transform 0 -1 39593 1 0 201600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[2\]
timestamp 1607115945
transform 0 1 675407 -1 0 206200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1607115945
transform 0 1 678007 -1 0 173200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_644
timestamp 1607115945
transform 0 1 678007 -1 0 177200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_645
timestamp 1607115945
transform 0 1 678007 -1 0 181200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1607115945
transform 0 1 678007 -1 0 185200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_647
timestamp 1607115945
transform 0 1 678007 -1 0 189200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_648
timestamp 1607115945
transform 0 1 678007 -1 0 190200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_650
timestamp 1607115945
transform 0 1 678007 -1 0 210200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_651
timestamp 1607115945
transform 0 1 678007 -1 0 214200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_430
timestamp 1607115945
transform 0 -1 39593 1 0 224600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_429
timestamp 1607115945
transform 0 -1 39593 1 0 223600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_428
timestamp 1607115945
transform 0 -1 39593 1 0 221600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_427
timestamp 1607115945
transform 0 -1 39593 1 0 217600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1607115945
transform 0 -1 39593 1 0 213600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[18\]
timestamp 1607115945
transform 0 -1 42193 1 0 224800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_432
timestamp 1607115945
transform 0 -1 39593 1 0 240800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1607115945
transform 0 -1 39593 1 0 252800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_434
timestamp 1607115945
transform 0 -1 39593 1 0 248800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_433
timestamp 1607115945
transform 0 -1 39593 1 0 244800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[3\]
timestamp 1607115945
transform 0 1 675407 -1 0 251400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_652
timestamp 1607115945
transform 0 1 678007 -1 0 218200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_653
timestamp 1607115945
transform 0 1 678007 -1 0 222200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_654
timestamp 1607115945
transform 0 1 678007 -1 0 226200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_655
timestamp 1607115945
transform 0 1 678007 -1 0 230200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1607115945
transform 0 1 678007 -1 0 234200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_657
timestamp 1607115945
transform 0 1 678007 -1 0 235200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_658
timestamp 1607115945
transform 0 1 678007 -1 0 235400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_660
timestamp 1607115945
transform 0 1 678007 -1 0 255400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[17\]
timestamp 1607115945
transform 0 -1 42193 1 0 268000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1607115945
transform 0 -1 39593 1 0 256800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_437
timestamp 1607115945
transform 0 -1 39593 1 0 260800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_438
timestamp 1607115945
transform 0 -1 39593 1 0 264800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_439
timestamp 1607115945
transform 0 -1 39593 1 0 266800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_440
timestamp 1607115945
transform 0 -1 39593 1 0 267800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_442
timestamp 1607115945
transform 0 -1 39593 1 0 284000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_443
timestamp 1607115945
transform 0 -1 39593 1 0 288000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_444
timestamp 1607115945
transform 0 -1 39593 1 0 292000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[4\]
timestamp 1607115945
transform 0 1 675407 -1 0 296400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_661
timestamp 1607115945
transform 0 1 678007 -1 0 259400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1607115945
transform 0 1 678007 -1 0 263400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_663
timestamp 1607115945
transform 0 1 678007 -1 0 267400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_664
timestamp 1607115945
transform 0 1 678007 -1 0 271400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1607115945
transform 0 1 678007 -1 0 275400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1607115945
transform 0 1 678007 -1 0 279400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_667
timestamp 1607115945
transform 0 1 678007 -1 0 280400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_450
timestamp 1607115945
transform 0 -1 39593 1 0 311000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_449
timestamp 1607115945
transform 0 -1 39593 1 0 310000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_448
timestamp 1607115945
transform 0 -1 39593 1 0 308000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_447
timestamp 1607115945
transform 0 -1 39593 1 0 304000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1607115945
transform 0 -1 39593 1 0 300000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1607115945
transform 0 -1 39593 1 0 296000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[16\]
timestamp 1607115945
transform 0 -1 42193 1 0 311200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_452
timestamp 1607115945
transform 0 -1 39593 1 0 327200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_454
timestamp 1607115945
transform 0 -1 39593 1 0 335200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_453
timestamp 1607115945
transform 0 -1 39593 1 0 331200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[5\]
timestamp 1607115945
transform 0 1 675407 -1 0 341400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_669
timestamp 1607115945
transform 0 1 678007 -1 0 300400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_670
timestamp 1607115945
transform 0 1 678007 -1 0 304400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1607115945
transform 0 1 678007 -1 0 308400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_672
timestamp 1607115945
transform 0 1 678007 -1 0 312400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_673
timestamp 1607115945
transform 0 1 678007 -1 0 316400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_674
timestamp 1607115945
transform 0 1 678007 -1 0 320400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1607115945
transform 0 1 678007 -1 0 324400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_676
timestamp 1607115945
transform 0 1 678007 -1 0 325400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_459
timestamp 1607115945
transform 0 -1 39593 1 0 353200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_458
timestamp 1607115945
transform 0 -1 39593 1 0 351200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_457
timestamp 1607115945
transform 0 -1 39593 1 0 347200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1607115945
transform 0 -1 39593 1 0 343200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1607115945
transform 0 -1 39593 1 0 339200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_460
timestamp 1607115945
transform 0 -1 39593 1 0 354200
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[15\]
timestamp 1607115945
transform 0 -1 42193 1 0 354400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_464
timestamp 1607115945
transform 0 -1 39593 1 0 378400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_463
timestamp 1607115945
transform 0 -1 39593 1 0 374400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_462
timestamp 1607115945
transform 0 -1 39593 1 0 370400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1607115945
transform 0 1 678007 -1 0 357400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_680
timestamp 1607115945
transform 0 1 678007 -1 0 353400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_679
timestamp 1607115945
transform 0 1 678007 -1 0 349400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_678
timestamp 1607115945
transform 0 1 678007 -1 0 345400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_685
timestamp 1607115945
transform 0 1 678007 -1 0 370400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1607115945
transform 0 1 678007 -1 0 369400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_683
timestamp 1607115945
transform 0 1 678007 -1 0 365400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_682
timestamp 1607115945
transform 0 1 678007 -1 0 361400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_686
timestamp 1607115945
transform 0 1 678007 -1 0 370600
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[6\]
timestamp 1607115945
transform 0 1 675407 -1 0 386600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_468
timestamp 1607115945
transform 0 -1 39593 1 0 394400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_467
timestamp 1607115945
transform 0 -1 39593 1 0 390400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1607115945
transform 0 -1 39593 1 0 386400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1607115945
transform 0 -1 39593 1 0 382400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_470
timestamp 1607115945
transform 0 -1 39593 1 0 397400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_469
timestamp 1607115945
transform 0 -1 39593 1 0 396400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[14\]
timestamp 1607115945
transform 0 -1 42193 1 0 397600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_474
timestamp 1607115945
transform 0 -1 39593 1 0 421600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_473
timestamp 1607115945
transform 0 -1 39593 1 0 417600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_472
timestamp 1607115945
transform 0 -1 39593 1 0 413600
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1607115945
transform 0 1 678007 -1 0 430600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_688
timestamp 1607115945
transform 0 1 678007 -1 0 390600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_689
timestamp 1607115945
transform 0 1 678007 -1 0 394600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1607115945
transform 0 1 678007 -1 0 398600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_691
timestamp 1607115945
transform 0 1 678007 -1 0 402600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_692
timestamp 1607115945
transform 0 1 678007 -1 0 406600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1607115945
transform 0 1 678007 -1 0 410600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1607115945
transform 0 1 678007 -1 0 414600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_695
timestamp 1607115945
transform 0 1 678007 -1 0 415600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_477
timestamp 1607115945
transform 0 -1 39593 1 0 433600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1607115945
transform 0 -1 39593 1 0 429600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1607115945
transform 0 -1 39593 1 0 425600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_480
timestamp 1607115945
transform 0 -1 39593 1 0 440600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_479
timestamp 1607115945
transform 0 -1 39593 1 0 439600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_478
timestamp 1607115945
transform 0 -1 39593 1 0 437600
box 0 0 2000 39593
use sky130_ef_io__vssd_lvc_pad  user2_vssd_lvclmap_pad
timestamp 1607115945
transform 0 -1 39593 1 0 440800
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_484
timestamp 1607115945
transform 0 -1 39593 1 0 463800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_483
timestamp 1607115945
transform 0 -1 39593 1 0 459800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_482
timestamp 1607115945
transform 0 -1 39593 1 0 455800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_698
timestamp 1607115945
transform 0 1 678007 -1 0 438600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_697
timestamp 1607115945
transform 0 1 678007 -1 0 434600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_702
timestamp 1607115945
transform 0 1 678007 -1 0 454600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_701
timestamp 1607115945
transform 0 1 678007 -1 0 450600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_700
timestamp 1607115945
transform 0 1 678007 -1 0 446600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_699
timestamp 1607115945
transform 0 1 678007 -1 0 442600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_705
timestamp 1607115945
transform 0 1 678007 -1 0 459800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_704
timestamp 1607115945
transform 0 1 678007 -1 0 459600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1607115945
transform 0 1 678007 -1 0 458600
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_pad  user1_vssd_lvclmap_pad
timestamp 1607115945
transform 0 1 678007 -1 0 474800
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_487
timestamp 1607115945
transform 0 -1 39593 1 0 475800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1607115945
transform 0 -1 39593 1 0 471800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1607115945
transform 0 -1 39593 1 0 467800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_490
timestamp 1607115945
transform 0 -1 39593 1 0 482800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_489
timestamp 1607115945
transform 0 -1 39593 1 0 481800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_488
timestamp 1607115945
transform 0 -1 39593 1 0 479800
box 0 0 2000 39593
use sky130_ef_io__vdda_hvc_pad  user2_vdda_hvclamp_pad
timestamp 1607115945
transform 0 -1 39593 1 0 483000
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_494
timestamp 1607115945
transform 0 -1 39593 1 0 506000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_493
timestamp 1607115945
transform 0 -1 39593 1 0 502000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_492
timestamp 1607115945
transform 0 -1 39593 1 0 498000
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1607115945
transform 0 1 678007 -1 0 518800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_707
timestamp 1607115945
transform 0 1 678007 -1 0 478800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_708
timestamp 1607115945
transform 0 1 678007 -1 0 482800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1607115945
transform 0 1 678007 -1 0 486800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_710
timestamp 1607115945
transform 0 1 678007 -1 0 490800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_711
timestamp 1607115945
transform 0 1 678007 -1 0 494800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1607115945
transform 0 1 678007 -1 0 498800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1607115945
transform 0 1 678007 -1 0 502800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_714
timestamp 1607115945
transform 0 1 678007 -1 0 503800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[13\]
timestamp 1607115945
transform 0 -1 42193 1 0 525200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1607115945
transform 0 -1 39593 1 0 510000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1607115945
transform 0 -1 39593 1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_497
timestamp 1607115945
transform 0 -1 39593 1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_498
timestamp 1607115945
transform 0 -1 39593 1 0 522000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_499
timestamp 1607115945
transform 0 -1 39593 1 0 524000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_500
timestamp 1607115945
transform 0 -1 39593 1 0 525000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_502
timestamp 1607115945
transform 0 -1 39593 1 0 541200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_503
timestamp 1607115945
transform 0 -1 39593 1 0 545200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[7\]
timestamp 1607115945
transform 0 1 675407 -1 0 563800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_716
timestamp 1607115945
transform 0 1 678007 -1 0 522800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_717
timestamp 1607115945
transform 0 1 678007 -1 0 526800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1607115945
transform 0 1 678007 -1 0 530800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_719
timestamp 1607115945
transform 0 1 678007 -1 0 534800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_720
timestamp 1607115945
transform 0 1 678007 -1 0 538800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_721
timestamp 1607115945
transform 0 1 678007 -1 0 542800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1607115945
transform 0 1 678007 -1 0 546800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_723
timestamp 1607115945
transform 0 1 678007 -1 0 547800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_507
timestamp 1607115945
transform 0 -1 39593 1 0 561200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1607115945
transform 0 -1 39593 1 0 557200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1607115945
transform 0 -1 39593 1 0 553200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_504
timestamp 1607115945
transform 0 -1 39593 1 0 549200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_510
timestamp 1607115945
transform 0 -1 39593 1 0 568200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_509
timestamp 1607115945
transform 0 -1 39593 1 0 567200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_508
timestamp 1607115945
transform 0 -1 39593 1 0 565200
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[12\]
timestamp 1607115945
transform 0 -1 42193 1 0 568400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_513
timestamp 1607115945
transform 0 -1 39593 1 0 588400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_512
timestamp 1607115945
transform 0 -1 39593 1 0 584400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_725
timestamp 1607115945
transform 0 1 678007 -1 0 567800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_726
timestamp 1607115945
transform 0 1 678007 -1 0 571800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_727
timestamp 1607115945
transform 0 1 678007 -1 0 575800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1607115945
transform 0 1 678007 -1 0 579800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_729
timestamp 1607115945
transform 0 1 678007 -1 0 583800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_730
timestamp 1607115945
transform 0 1 678007 -1 0 587800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1607115945
transform 0 1 678007 -1 0 591800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_517
timestamp 1607115945
transform 0 -1 39593 1 0 604400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1607115945
transform 0 -1 39593 1 0 600400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1607115945
transform 0 -1 39593 1 0 596400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_514
timestamp 1607115945
transform 0 -1 39593 1 0 592400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_520
timestamp 1607115945
transform 0 -1 39593 1 0 611400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_519
timestamp 1607115945
transform 0 -1 39593 1 0 610400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_518
timestamp 1607115945
transform 0 -1 39593 1 0 608400
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[11\]
timestamp 1607115945
transform 0 -1 42193 1 0 611600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_523
timestamp 1607115945
transform 0 -1 39593 1 0 631600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_522
timestamp 1607115945
transform 0 -1 39593 1 0 627600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[8\]
timestamp 1607115945
transform 0 1 675407 -1 0 609000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_732
timestamp 1607115945
transform 0 1 678007 -1 0 592800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_733
timestamp 1607115945
transform 0 1 678007 -1 0 593000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_735
timestamp 1607115945
transform 0 1 678007 -1 0 613000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_736
timestamp 1607115945
transform 0 1 678007 -1 0 617000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1607115945
transform 0 1 678007 -1 0 621000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_738
timestamp 1607115945
transform 0 1 678007 -1 0 625000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_739
timestamp 1607115945
transform 0 1 678007 -1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1607115945
transform 0 1 678007 -1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_527
timestamp 1607115945
transform 0 -1 39593 1 0 647600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1607115945
transform 0 -1 39593 1 0 643600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1607115945
transform 0 -1 39593 1 0 639600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_524
timestamp 1607115945
transform 0 -1 39593 1 0 635600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_530
timestamp 1607115945
transform 0 -1 39593 1 0 654600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_529
timestamp 1607115945
transform 0 -1 39593 1 0 653600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_528
timestamp 1607115945
transform 0 -1 39593 1 0 651600
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[10\]
timestamp 1607115945
transform 0 -1 42193 1 0 654800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_533
timestamp 1607115945
transform 0 -1 39593 1 0 674800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_532
timestamp 1607115945
transform 0 -1 39593 1 0 670800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[9\]
timestamp 1607115945
transform 0 1 675407 -1 0 654000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1607115945
transform 0 1 678007 -1 0 637000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_742
timestamp 1607115945
transform 0 1 678007 -1 0 638000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_744
timestamp 1607115945
transform 0 1 678007 -1 0 658000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_745
timestamp 1607115945
transform 0 1 678007 -1 0 662000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_746
timestamp 1607115945
transform 0 1 678007 -1 0 666000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_747
timestamp 1607115945
transform 0 1 678007 -1 0 670000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_748
timestamp 1607115945
transform 0 1 678007 -1 0 674000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_749
timestamp 1607115945
transform 0 1 678007 -1 0 678000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[9\]
timestamp 1607115945
transform 0 -1 42193 1 0 698000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_534
timestamp 1607115945
transform 0 -1 39593 1 0 678800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1607115945
transform 0 -1 39593 1 0 682800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1607115945
transform 0 -1 39593 1 0 686800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_537
timestamp 1607115945
transform 0 -1 39593 1 0 690800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_538
timestamp 1607115945
transform 0 -1 39593 1 0 694800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_539
timestamp 1607115945
transform 0 -1 39593 1 0 696800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_540
timestamp 1607115945
transform 0 -1 39593 1 0 697800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_542
timestamp 1607115945
transform 0 -1 39593 1 0 714000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[10\]
timestamp 1607115945
transform 0 1 675407 -1 0 699200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1607115945
transform 0 1 678007 -1 0 682000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_751
timestamp 1607115945
transform 0 1 678007 -1 0 683000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_752
timestamp 1607115945
transform 0 1 678007 -1 0 683200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_754
timestamp 1607115945
transform 0 1 678007 -1 0 703200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_755
timestamp 1607115945
transform 0 1 678007 -1 0 707200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1607115945
transform 0 1 678007 -1 0 711200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_757
timestamp 1607115945
transform 0 1 678007 -1 0 715200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_758
timestamp 1607115945
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1607115945
transform 0 -1 39593 1 0 730000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1607115945
transform 0 -1 39593 1 0 726000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_544
timestamp 1607115945
transform 0 -1 39593 1 0 722000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_543
timestamp 1607115945
transform 0 -1 39593 1 0 718000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_550
timestamp 1607115945
transform 0 -1 39593 1 0 741000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_549
timestamp 1607115945
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_548
timestamp 1607115945
transform 0 -1 39593 1 0 738000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_547
timestamp 1607115945
transform 0 -1 39593 1 0 734000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[8\]
timestamp 1607115945
transform 0 -1 42193 1 0 741200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_552
timestamp 1607115945
transform 0 -1 39593 1 0 757200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[11\]
timestamp 1607115945
transform 0 1 675407 -1 0 744200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1607115945
transform 0 1 678007 -1 0 723200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1607115945
transform 0 1 678007 -1 0 727200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_761
timestamp 1607115945
transform 0 1 678007 -1 0 728200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_763
timestamp 1607115945
transform 0 1 678007 -1 0 748200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_764
timestamp 1607115945
transform 0 1 678007 -1 0 752200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1607115945
transform 0 1 678007 -1 0 756200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_766
timestamp 1607115945
transform 0 1 678007 -1 0 760200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1607115945
transform 0 -1 39593 1 0 773200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1607115945
transform 0 -1 39593 1 0 769200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_554
timestamp 1607115945
transform 0 -1 39593 1 0 765200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_553
timestamp 1607115945
transform 0 -1 39593 1 0 761200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_560
timestamp 1607115945
transform 0 -1 39593 1 0 784200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_559
timestamp 1607115945
transform 0 -1 39593 1 0 783200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_558
timestamp 1607115945
transform 0 -1 39593 1 0 781200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_557
timestamp 1607115945
transform 0 -1 39593 1 0 777200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[7\]
timestamp 1607115945
transform 0 -1 42193 1 0 784400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_562
timestamp 1607115945
transform 0 -1 39593 1 0 800400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[12\]
timestamp 1607115945
transform 0 1 675407 -1 0 789200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_767
timestamp 1607115945
transform 0 1 678007 -1 0 764200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_768
timestamp 1607115945
transform 0 1 678007 -1 0 768200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1607115945
transform 0 1 678007 -1 0 772200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_770
timestamp 1607115945
transform 0 1 678007 -1 0 773200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_772
timestamp 1607115945
transform 0 1 678007 -1 0 793200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_773
timestamp 1607115945
transform 0 1 678007 -1 0 797200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_774
timestamp 1607115945
transform 0 1 678007 -1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1607115945
transform 0 1 678007 -1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1607115945
transform 0 -1 39593 1 0 816400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1607115945
transform 0 -1 39593 1 0 812400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_564
timestamp 1607115945
transform 0 -1 39593 1 0 808400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_563
timestamp 1607115945
transform 0 -1 39593 1 0 804400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_570
timestamp 1607115945
transform 0 -1 39593 1 0 827400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_569
timestamp 1607115945
transform 0 -1 39593 1 0 826400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_568
timestamp 1607115945
transform 0 -1 39593 1 0 824400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1607115945
transform 0 -1 39593 1 0 820400
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user2_vssa_hvclamp_pad
timestamp 1607115945
transform 0 -1 39593 1 0 827600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_572
timestamp 1607115945
transform 0 -1 39593 1 0 842600
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1607115945
transform 0 1 678007 -1 0 833400
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_776
timestamp 1607115945
transform 0 1 678007 -1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_777
timestamp 1607115945
transform 0 1 678007 -1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_778
timestamp 1607115945
transform 0 1 678007 -1 0 817200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_779
timestamp 1607115945
transform 0 1 678007 -1 0 818200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_780
timestamp 1607115945
transform 0 1 678007 -1 0 818400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_782
timestamp 1607115945
transform 0 1 678007 -1 0 837400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_783
timestamp 1607115945
transform 0 1 678007 -1 0 841400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1607115945
transform 0 1 678007 -1 0 845400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_576
timestamp 1607115945
transform 0 -1 39593 1 0 858600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1607115945
transform 0 -1 39593 1 0 854600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_574
timestamp 1607115945
transform 0 -1 39593 1 0 850600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_573
timestamp 1607115945
transform 0 -1 39593 1 0 846600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_580
timestamp 1607115945
transform 0 -1 39593 1 0 869600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_579
timestamp 1607115945
transform 0 -1 39593 1 0 868600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_578
timestamp 1607115945
transform 0 -1 39593 1 0 866600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_577
timestamp 1607115945
transform 0 -1 39593 1 0 862600
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1607115945
transform 0 -1 39593 1 0 869800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_582
timestamp 1607115945
transform 0 -1 39593 1 0 884800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[13\]
timestamp 1607115945
transform 0 1 675407 -1 0 878400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1607115945
transform 0 1 678007 -1 0 849400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_786
timestamp 1607115945
transform 0 1 678007 -1 0 853400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_787
timestamp 1607115945
transform 0 1 678007 -1 0 857400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_788
timestamp 1607115945
transform 0 1 678007 -1 0 861400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_789
timestamp 1607115945
transform 0 1 678007 -1 0 862400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_791
timestamp 1607115945
transform 0 1 678007 -1 0 882400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_792
timestamp 1607115945
transform 0 1 678007 -1 0 886400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1607115945
transform 0 -1 39593 1 0 900800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1607115945
transform 0 -1 39593 1 0 896800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_584
timestamp 1607115945
transform 0 -1 39593 1 0 892800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_583
timestamp 1607115945
transform 0 -1 39593 1 0 888800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_590
timestamp 1607115945
transform 0 -1 39593 1 0 911800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_589
timestamp 1607115945
transform 0 -1 39593 1 0 910800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_588
timestamp 1607115945
transform 0 -1 39593 1 0 908800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_587
timestamp 1607115945
transform 0 -1 39593 1 0 904800
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  user2_vccd_lvclamp_pad
timestamp 1607115945
transform 0 -1 39593 1 0 912000
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_592
timestamp 1607115945
transform 0 -1 39593 1 0 927000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_796
timestamp 1607115945
transform 0 1 678007 -1 0 902400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_795
timestamp 1607115945
transform 0 1 678007 -1 0 898400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_794
timestamp 1607115945
transform 0 1 678007 -1 0 894400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_793
timestamp 1607115945
transform 0 1 678007 -1 0 890400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_799
timestamp 1607115945
transform 0 1 678007 -1 0 907600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_798
timestamp 1607115945
transform 0 1 678007 -1 0 907400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_797
timestamp 1607115945
transform 0 1 678007 -1 0 906400
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  user1_vccd_lvclamp_pad
timestamp 1607115945
transform 0 1 678007 -1 0 922600
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_802
timestamp 1607115945
transform 0 1 678007 -1 0 930600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_801
timestamp 1607115945
transform 0 1 678007 -1 0 926600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1607115945
transform 0 -1 39593 1 0 943000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1607115945
transform 0 -1 39593 1 0 939000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_594
timestamp 1607115945
transform 0 -1 39593 1 0 935000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_593
timestamp 1607115945
transform 0 -1 39593 1 0 931000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_600
timestamp 1607115945
transform 0 -1 39593 1 0 954000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_599
timestamp 1607115945
transform 0 -1 39593 1 0 953000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_598
timestamp 1607115945
transform 0 -1 39593 1 0 951000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_597
timestamp 1607115945
transform 0 -1 39593 1 0 947000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[6\]
timestamp 1607115945
transform 0 -1 42193 1 0 954200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_602
timestamp 1607115945
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[14\]
timestamp 1607115945
transform 0 1 675407 -1 0 967600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_803
timestamp 1607115945
transform 0 1 678007 -1 0 934600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_804
timestamp 1607115945
transform 0 1 678007 -1 0 938600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_805
timestamp 1607115945
transform 0 1 678007 -1 0 942600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_806
timestamp 1607115945
transform 0 1 678007 -1 0 946600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_807
timestamp 1607115945
transform 0 1 678007 -1 0 950600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_808
timestamp 1607115945
transform 0 1 678007 -1 0 951600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_810
timestamp 1607115945
transform 0 1 678007 -1 0 971600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_607
timestamp 1607115945
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_606
timestamp 1607115945
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1607115945
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_604
timestamp 1607115945
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_603
timestamp 1607115945
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_611
timestamp 1607115945
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_610
timestamp 1607115945
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_609
timestamp 1607115945
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_608
timestamp 1607115945
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_5
timestamp 1607115945
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1607115945
transform 0 -1 40800 1 0 997600
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1607115945
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1607115945
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1607115945
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1607115945
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_13
timestamp 1607115945
transform 1 0 72800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1607115945
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1607115945
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1607115945
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_16
timestamp 1607115945
transform 1 0 76000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15
timestamp 1607115945
transform 1 0 75800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_14
timestamp 1607115945
transform 1 0 74800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[5\]
timestamp 1607115945
transform 1 0 76200 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1607115945
transform 1 0 92200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1607115945
transform 1 0 96200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1607115945
transform 1 0 100200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1607115945
transform 1 0 104200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1607115945
transform 1 0 108200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1607115945
transform 1 0 112200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1607115945
transform 1 0 116200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1607115945
transform 1 0 120200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_27
timestamp 1607115945
transform 1 0 126200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_26
timestamp 1607115945
transform 1 0 124200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_29
timestamp 1607115945
transform 1 0 127400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_28
timestamp 1607115945
transform 1 0 127200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[4\]
timestamp 1607115945
transform 1 0 127600 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1607115945
transform 1 0 155600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1607115945
transform 1 0 151600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1607115945
transform 1 0 147600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1607115945
transform 1 0 143600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1607115945
transform 1 0 167600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1607115945
transform 1 0 163600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1607115945
transform 1 0 159600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_42
timestamp 1607115945
transform 1 0 178800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_41
timestamp 1607115945
transform 1 0 178600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_40
timestamp 1607115945
transform 1 0 177600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_39
timestamp 1607115945
transform 1 0 175600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_38
timestamp 1607115945
transform 1 0 171600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[3\]
timestamp 1607115945
transform 1 0 179000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1607115945
transform 1 0 199000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1607115945
transform 1 0 195000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_47
timestamp 1607115945
transform 1 0 207000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1607115945
transform 1 0 203000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_52
timestamp 1607115945
transform 1 0 227000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1607115945
transform 1 0 223000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1607115945
transform 1 0 219000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1607115945
transform 1 0 215000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_48
timestamp 1607115945
transform 1 0 211000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1607115945
transform 1 0 230200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1607115945
transform 1 0 230000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_53
timestamp 1607115945
transform 1 0 229000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[2\]
timestamp 1607115945
transform 1 0 230400 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_58
timestamp 1607115945
transform 1 0 250400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_57
timestamp 1607115945
transform 1 0 246400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1607115945
transform 1 0 266400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1607115945
transform 1 0 262400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1607115945
transform 1 0 258400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_59
timestamp 1607115945
transform 1 0 254400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_69
timestamp 1607115945
transform 1 0 281800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_68
timestamp 1607115945
transform 1 0 281600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_67
timestamp 1607115945
transform 1 0 281400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_66
timestamp 1607115945
transform 1 0 280400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_65
timestamp 1607115945
transform 1 0 278400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1607115945
transform 1 0 274400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1607115945
transform 1 0 270400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[1\]
timestamp 1607115945
transform 1 0 282000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_74
timestamp 1607115945
transform 1 0 310000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1607115945
transform 1 0 306000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1607115945
transform 1 0 302000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1607115945
transform 1 0 298000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_77
timestamp 1607115945
transform 1 0 322000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_76
timestamp 1607115945
transform 1 0 318000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_75
timestamp 1607115945
transform 1 0 314000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_82
timestamp 1607115945
transform 1 0 333200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_81
timestamp 1607115945
transform 1 0 333000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_80
timestamp 1607115945
transform 1 0 332000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_79
timestamp 1607115945
transform 1 0 330000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1607115945
transform 1 0 326000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__vssio_hvc_pad  mgmt_vssio_hvclamp_pad\[0\]
timestamp 1607115945
transform 1 0 333400 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_84
timestamp 1607115945
transform 1 0 348400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_85
timestamp 1607115945
transform 1 0 352400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1607115945
transform 1 0 356400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1607115945
transform 1 0 360400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1607115945
transform 1 0 364400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1607115945
transform 1 0 368400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1607115945
transform 1 0 372400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1607115945
transform 1 0 376400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1607115945
transform 1 0 383600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_94
timestamp 1607115945
transform 1 0 383400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_93
timestamp 1607115945
transform 1 0 382400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_92
timestamp 1607115945
transform 1 0 380400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[0\]
timestamp 1607115945
transform 1 0 383800 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1607115945
transform 1 0 411800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_99
timestamp 1607115945
transform 1 0 407800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_98
timestamp 1607115945
transform 1 0 403800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_97
timestamp 1607115945
transform 1 0 399800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1607115945
transform 1 0 419800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1607115945
transform 1 0 415800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1607115945
transform 1 0 423800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1607115945
transform 1 0 427800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_106
timestamp 1607115945
transform 1 0 433800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_105
timestamp 1607115945
transform 1 0 431800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1607115945
transform 1 0 437200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_0
timestamp 1607115945
transform 1 0 436200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0
timestamp 1607115945
transform 1 0 435200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_108
timestamp 1607115945
transform 1 0 435000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_107
timestamp 1607115945
transform 1 0 434800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1607115945
transform 1 0 441200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1607115945
transform 1 0 445200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1607115945
transform 1 0 449200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1607115945
transform 1 0 453200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_116
timestamp 1607115945
transform 1 0 457200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_117
timestamp 1607115945
transform 1 0 461200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_123
timestamp 1607115945
transform 1 0 472600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_122
timestamp 1607115945
transform 1 0 472400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_121
timestamp 1607115945
transform 1 0 472200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_120
timestamp 1607115945
transform 1 0 471200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_119
timestamp 1607115945
transform 1 0 469200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_118
timestamp 1607115945
transform 1 0 465200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[17\]
timestamp 1607115945
transform 1 0 472800 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_126
timestamp 1607115945
transform 1 0 492800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1607115945
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_129
timestamp 1607115945
transform 1 0 504800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_128
timestamp 1607115945
transform 1 0 500800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_127
timestamp 1607115945
transform 1 0 496800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_133
timestamp 1607115945
transform 1 0 520800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_132
timestamp 1607115945
transform 1 0 516800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1607115945
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_130
timestamp 1607115945
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_136
timestamp 1607115945
transform 1 0 524000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_135
timestamp 1607115945
transform 1 0 523800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_134
timestamp 1607115945
transform 1 0 522800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[16\]
timestamp 1607115945
transform 1 0 524200 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_140
timestamp 1607115945
transform 1 0 548200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_139
timestamp 1607115945
transform 1 0 544200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_138
timestamp 1607115945
transform 1 0 540200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_143
timestamp 1607115945
transform 1 0 560200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_142
timestamp 1607115945
transform 1 0 556200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_141
timestamp 1607115945
transform 1 0 552200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_149
timestamp 1607115945
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_148
timestamp 1607115945
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_147
timestamp 1607115945
transform 1 0 574200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_146
timestamp 1607115945
transform 1 0 572200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_145
timestamp 1607115945
transform 1 0 568200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_144
timestamp 1607115945
transform 1 0 564200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1607115945
transform 1 0 575600 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_151
timestamp 1607115945
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_155
timestamp 1607115945
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_154
timestamp 1607115945
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_153
timestamp 1607115945
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_152
timestamp 1607115945
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_159
timestamp 1607115945
transform 1 0 622600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_158
timestamp 1607115945
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_157
timestamp 1607115945
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_156
timestamp 1607115945
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_162
timestamp 1607115945
transform 1 0 625800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_161
timestamp 1607115945
transform 1 0 625600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_160
timestamp 1607115945
transform 1 0 624600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[15\]
timestamp 1607115945
transform 1 0 626000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_164
timestamp 1607115945
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_165
timestamp 1607115945
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_166
timestamp 1607115945
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_167
timestamp 1607115945
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_168
timestamp 1607115945
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_169
timestamp 1607115945
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_170
timestamp 1607115945
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_171
timestamp 1607115945
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_172
timestamp 1607115945
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_815
timestamp 1607115945
transform 0 1 678007 -1 0 991600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_814
timestamp 1607115945
transform 0 1 678007 -1 0 987600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_813
timestamp 1607115945
transform 0 1 678007 -1 0 983600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_812
timestamp 1607115945
transform 0 1 678007 -1 0 979600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_811
timestamp 1607115945
transform 0 1 678007 -1 0 975600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_818
timestamp 1607115945
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_817
timestamp 1607115945
transform 0 1 678007 -1 0 996600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_816
timestamp 1607115945
transform 0 1 678007 -1 0 995600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_176
timestamp 1607115945
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_175
timestamp 1607115945
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_174
timestamp 1607115945
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_173
timestamp 1607115945
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__corner_pad  user1_corner
timestamp 1607115945
transform 1 0 677600 0 1 996800
box 0 0 40000 40800
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 1 nsew signal tristate
rlabel metal2 s 194043 41713 194099 42193 6 por
port 2 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 3 nsew signal tristate
rlabel metal2 s 361767 41713 361823 42193 6 flash_clk_core
port 4 nsew signal input
rlabel metal2 s 357443 41713 357499 42193 6 flash_clk_ieb_core
port 5 nsew signal input
rlabel metal2 s 364895 41713 364951 42193 6 flash_clk_oeb_core
port 6 nsew signal input
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 7 nsew signal tristate
rlabel metal2 s 306967 41713 307023 42193 6 flash_csb_core
port 8 nsew signal input
rlabel metal2 s 302643 41713 302699 42193 6 flash_csb_ieb_core
port 9 nsew signal input
rlabel metal2 s 310095 41713 310151 42193 6 flash_csb_oeb_core
port 10 nsew signal input
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 11 nsew signal bidirectional
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 12 nsew signal tristate
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 13 nsew signal input
rlabel metal2 s 412243 41713 412299 42193 6 flash_io0_ieb_core
port 14 nsew signal input
rlabel metal2 s 419695 41713 419751 42193 6 flash_io0_oeb_core
port 15 nsew signal input
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 16 nsew signal bidirectional
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 17 nsew signal tristate
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 18 nsew signal input
rlabel metal2 s 467043 41713 467099 42193 6 flash_io1_ieb_core
port 19 nsew signal input
rlabel metal2 s 474495 41713 474551 42193 6 flash_io1_oeb_core
port 20 nsew signal input
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 21 nsew signal bidirectional
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 22 nsew signal tristate
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 23 nsew signal input
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 24 nsew signal input
rlabel metal2 s 524971 41713 525027 42193 6 gpio_mode1_core
port 25 nsew signal input
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 26 nsew signal input
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 27 nsew signal input
rlabel metal5 s 6086 69863 19572 81191 6 vccd
port 28 nsew signal bidirectional
rlabel metal5 s 624040 6675 636580 19197 6 vdda
port 29 nsew signal bidirectional
rlabel metal5 s 6675 111420 19197 123960 6 vddio
port 30 nsew signal bidirectional
rlabel metal5 s 80040 6675 92580 19197 6 vssa
port 31 nsew signal bidirectional
rlabel metal5 s 243009 6086 254337 19572 6 vssd
port 32 nsew signal bidirectional
rlabel metal5 s 334620 1018402 347160 1030924 6 vssio
port 33 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 34 nsew signal bidirectional
rlabel metal2 s 675407 105803 675887 105859 6 mprj_io_analog_en[0]
port 35 nsew signal input
rlabel metal2 s 675407 107091 675887 107147 6 mprj_io_analog_pol[0]
port 36 nsew signal input
rlabel metal2 s 675407 110127 675887 110183 6 mprj_io_analog_sel[0]
port 37 nsew signal input
rlabel metal2 s 675407 106447 675887 106503 6 mprj_io_dm[0]
port 38 nsew signal input
rlabel metal2 s 675407 104607 675887 104663 6 mprj_io_dm[1]
port 39 nsew signal input
rlabel metal2 s 675407 110771 675887 110827 6 mprj_io_dm[2]
port 40 nsew signal input
rlabel metal2 s 675407 108931 675887 108987 6 mprj_io_enh[0]
port 41 nsew signal input
rlabel metal2 s 675407 109575 675887 109631 6 mprj_io_hldh_n[0]
port 42 nsew signal input
rlabel metal2 s 675407 111415 675887 111471 6 mprj_io_holdover[0]
port 43 nsew signal input
rlabel metal2 s 675407 114451 675887 114507 6 mprj_io_ib_mode_sel[0]
port 44 nsew signal input
rlabel metal2 s 675407 107643 675887 107699 6 mprj_io_inp_dis[0]
port 45 nsew signal input
rlabel metal2 s 675407 115095 675887 115151 6 mprj_io_oeb[0]
port 46 nsew signal input
rlabel metal2 s 675407 111967 675887 112023 6 mprj_io_out[0]
port 47 nsew signal input
rlabel metal2 s 675407 102767 675887 102823 6 mprj_io_slow_sel[0]
port 48 nsew signal input
rlabel metal2 s 675407 113807 675887 113863 6 mprj_io_vtrip_sel[0]
port 49 nsew signal input
rlabel metal2 s 675407 100927 675887 100983 6 mprj_io_in[0]
port 50 nsew signal tristate
rlabel metal2 s 675407 686611 675887 686667 6 mprj_analog_io[3]
port 51 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 52 nsew signal bidirectional
rlabel metal2 s 675407 689003 675887 689059 6 mprj_io_analog_en[10]
port 53 nsew signal input
rlabel metal2 s 675407 690291 675887 690347 6 mprj_io_analog_pol[10]
port 54 nsew signal input
rlabel metal2 s 675407 693327 675887 693383 6 mprj_io_analog_sel[10]
port 55 nsew signal input
rlabel metal2 s 675407 689647 675887 689703 6 mprj_io_dm[30]
port 56 nsew signal input
rlabel metal2 s 675407 687807 675887 687863 6 mprj_io_dm[31]
port 57 nsew signal input
rlabel metal2 s 675407 693971 675887 694027 6 mprj_io_dm[32]
port 58 nsew signal input
rlabel metal2 s 675407 692131 675887 692187 6 mprj_io_enh[10]
port 59 nsew signal input
rlabel metal2 s 675407 692775 675887 692831 6 mprj_io_hldh_n[10]
port 60 nsew signal input
rlabel metal2 s 675407 694615 675887 694671 6 mprj_io_holdover[10]
port 61 nsew signal input
rlabel metal2 s 675407 697651 675887 697707 6 mprj_io_ib_mode_sel[10]
port 62 nsew signal input
rlabel metal2 s 675407 690843 675887 690899 6 mprj_io_inp_dis[10]
port 63 nsew signal input
rlabel metal2 s 675407 698295 675887 698351 6 mprj_io_oeb[10]
port 64 nsew signal input
rlabel metal2 s 675407 695167 675887 695223 6 mprj_io_out[10]
port 65 nsew signal input
rlabel metal2 s 675407 685967 675887 686023 6 mprj_io_slow_sel[10]
port 66 nsew signal input
rlabel metal2 s 675407 697007 675887 697063 6 mprj_io_vtrip_sel[10]
port 67 nsew signal input
rlabel metal2 s 675407 684127 675887 684183 6 mprj_io_in[10]
port 68 nsew signal tristate
rlabel metal2 s 675407 731611 675887 731667 6 mprj_analog_io[4]
port 69 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 70 nsew signal bidirectional
rlabel metal2 s 675407 734003 675887 734059 6 mprj_io_analog_en[11]
port 71 nsew signal input
rlabel metal2 s 675407 735291 675887 735347 6 mprj_io_analog_pol[11]
port 72 nsew signal input
rlabel metal2 s 675407 738327 675887 738383 6 mprj_io_analog_sel[11]
port 73 nsew signal input
rlabel metal2 s 675407 734647 675887 734703 6 mprj_io_dm[33]
port 74 nsew signal input
rlabel metal2 s 675407 732807 675887 732863 6 mprj_io_dm[34]
port 75 nsew signal input
rlabel metal2 s 675407 738971 675887 739027 6 mprj_io_dm[35]
port 76 nsew signal input
rlabel metal2 s 675407 737131 675887 737187 6 mprj_io_enh[11]
port 77 nsew signal input
rlabel metal2 s 675407 737775 675887 737831 6 mprj_io_hldh_n[11]
port 78 nsew signal input
rlabel metal2 s 675407 739615 675887 739671 6 mprj_io_holdover[11]
port 79 nsew signal input
rlabel metal2 s 675407 742651 675887 742707 6 mprj_io_ib_mode_sel[11]
port 80 nsew signal input
rlabel metal2 s 675407 735843 675887 735899 6 mprj_io_inp_dis[11]
port 81 nsew signal input
rlabel metal2 s 675407 743295 675887 743351 6 mprj_io_oeb[11]
port 82 nsew signal input
rlabel metal2 s 675407 740167 675887 740223 6 mprj_io_out[11]
port 83 nsew signal input
rlabel metal2 s 675407 730967 675887 731023 6 mprj_io_slow_sel[11]
port 84 nsew signal input
rlabel metal2 s 675407 742007 675887 742063 6 mprj_io_vtrip_sel[11]
port 85 nsew signal input
rlabel metal2 s 675407 729127 675887 729183 6 mprj_io_in[11]
port 86 nsew signal tristate
rlabel metal2 s 675407 776611 675887 776667 6 mprj_analog_io[5]
port 87 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 88 nsew signal bidirectional
rlabel metal2 s 675407 779003 675887 779059 6 mprj_io_analog_en[12]
port 89 nsew signal input
rlabel metal2 s 675407 780291 675887 780347 6 mprj_io_analog_pol[12]
port 90 nsew signal input
rlabel metal2 s 675407 783327 675887 783383 6 mprj_io_analog_sel[12]
port 91 nsew signal input
rlabel metal2 s 675407 779647 675887 779703 6 mprj_io_dm[36]
port 92 nsew signal input
rlabel metal2 s 675407 777807 675887 777863 6 mprj_io_dm[37]
port 93 nsew signal input
rlabel metal2 s 675407 783971 675887 784027 6 mprj_io_dm[38]
port 94 nsew signal input
rlabel metal2 s 675407 782131 675887 782187 6 mprj_io_enh[12]
port 95 nsew signal input
rlabel metal2 s 675407 782775 675887 782831 6 mprj_io_hldh_n[12]
port 96 nsew signal input
rlabel metal2 s 675407 784615 675887 784671 6 mprj_io_holdover[12]
port 97 nsew signal input
rlabel metal2 s 675407 787651 675887 787707 6 mprj_io_ib_mode_sel[12]
port 98 nsew signal input
rlabel metal2 s 675407 780843 675887 780899 6 mprj_io_inp_dis[12]
port 99 nsew signal input
rlabel metal2 s 675407 788295 675887 788351 6 mprj_io_oeb[12]
port 100 nsew signal input
rlabel metal2 s 675407 785167 675887 785223 6 mprj_io_out[12]
port 101 nsew signal input
rlabel metal2 s 675407 775967 675887 776023 6 mprj_io_slow_sel[12]
port 102 nsew signal input
rlabel metal2 s 675407 787007 675887 787063 6 mprj_io_vtrip_sel[12]
port 103 nsew signal input
rlabel metal2 s 675407 774127 675887 774183 6 mprj_io_in[12]
port 104 nsew signal tristate
rlabel metal2 s 675407 865811 675887 865867 6 mprj_analog_io[6]
port 105 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 106 nsew signal bidirectional
rlabel metal2 s 675407 868203 675887 868259 6 mprj_io_analog_en[13]
port 107 nsew signal input
rlabel metal2 s 675407 869491 675887 869547 6 mprj_io_analog_pol[13]
port 108 nsew signal input
rlabel metal2 s 675407 872527 675887 872583 6 mprj_io_analog_sel[13]
port 109 nsew signal input
rlabel metal2 s 675407 868847 675887 868903 6 mprj_io_dm[39]
port 110 nsew signal input
rlabel metal2 s 675407 867007 675887 867063 6 mprj_io_dm[40]
port 111 nsew signal input
rlabel metal2 s 675407 873171 675887 873227 6 mprj_io_dm[41]
port 112 nsew signal input
rlabel metal2 s 675407 871331 675887 871387 6 mprj_io_enh[13]
port 113 nsew signal input
rlabel metal2 s 675407 871975 675887 872031 6 mprj_io_hldh_n[13]
port 114 nsew signal input
rlabel metal2 s 675407 873815 675887 873871 6 mprj_io_holdover[13]
port 115 nsew signal input
rlabel metal2 s 675407 876851 675887 876907 6 mprj_io_ib_mode_sel[13]
port 116 nsew signal input
rlabel metal2 s 675407 870043 675887 870099 6 mprj_io_inp_dis[13]
port 117 nsew signal input
rlabel metal2 s 675407 877495 675887 877551 6 mprj_io_oeb[13]
port 118 nsew signal input
rlabel metal2 s 675407 874367 675887 874423 6 mprj_io_out[13]
port 119 nsew signal input
rlabel metal2 s 675407 865167 675887 865223 6 mprj_io_slow_sel[13]
port 120 nsew signal input
rlabel metal2 s 675407 876207 675887 876263 6 mprj_io_vtrip_sel[13]
port 121 nsew signal input
rlabel metal2 s 675407 863327 675887 863383 6 mprj_io_in[13]
port 122 nsew signal tristate
rlabel metal2 s 675407 955011 675887 955067 6 mprj_analog_io[7]
port 123 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 124 nsew signal bidirectional
rlabel metal2 s 675407 957403 675887 957459 6 mprj_io_analog_en[14]
port 125 nsew signal input
rlabel metal2 s 675407 958691 675887 958747 6 mprj_io_analog_pol[14]
port 126 nsew signal input
rlabel metal2 s 675407 961727 675887 961783 6 mprj_io_analog_sel[14]
port 127 nsew signal input
rlabel metal2 s 675407 958047 675887 958103 6 mprj_io_dm[42]
port 128 nsew signal input
rlabel metal2 s 675407 956207 675887 956263 6 mprj_io_dm[43]
port 129 nsew signal input
rlabel metal2 s 675407 962371 675887 962427 6 mprj_io_dm[44]
port 130 nsew signal input
rlabel metal2 s 675407 960531 675887 960587 6 mprj_io_enh[14]
port 131 nsew signal input
rlabel metal2 s 675407 961175 675887 961231 6 mprj_io_hldh_n[14]
port 132 nsew signal input
rlabel metal2 s 675407 963015 675887 963071 6 mprj_io_holdover[14]
port 133 nsew signal input
rlabel metal2 s 675407 966051 675887 966107 6 mprj_io_ib_mode_sel[14]
port 134 nsew signal input
rlabel metal2 s 675407 959243 675887 959299 6 mprj_io_inp_dis[14]
port 135 nsew signal input
rlabel metal2 s 675407 966695 675887 966751 6 mprj_io_oeb[14]
port 136 nsew signal input
rlabel metal2 s 675407 963567 675887 963623 6 mprj_io_out[14]
port 137 nsew signal input
rlabel metal2 s 675407 954367 675887 954423 6 mprj_io_slow_sel[14]
port 138 nsew signal input
rlabel metal2 s 675407 965407 675887 965463 6 mprj_io_vtrip_sel[14]
port 139 nsew signal input
rlabel metal2 s 675407 952527 675887 952583 6 mprj_io_in[14]
port 140 nsew signal tristate
rlabel metal2 s 638533 995407 638589 995887 6 mprj_analog_io[8]
port 141 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 142 nsew signal bidirectional
rlabel metal2 s 636141 995407 636197 995887 6 mprj_io_analog_en[15]
port 143 nsew signal input
rlabel metal2 s 634853 995407 634909 995887 6 mprj_io_analog_pol[15]
port 144 nsew signal input
rlabel metal2 s 631817 995407 631873 995887 6 mprj_io_analog_sel[15]
port 145 nsew signal input
rlabel metal2 s 635497 995407 635553 995887 6 mprj_io_dm[45]
port 146 nsew signal input
rlabel metal2 s 637337 995407 637393 995887 6 mprj_io_dm[46]
port 147 nsew signal input
rlabel metal2 s 631173 995407 631229 995887 6 mprj_io_dm[47]
port 148 nsew signal input
rlabel metal2 s 633013 995407 633069 995887 6 mprj_io_enh[15]
port 149 nsew signal input
rlabel metal2 s 632369 995407 632425 995887 6 mprj_io_hldh_n[15]
port 150 nsew signal input
rlabel metal2 s 630529 995407 630585 995887 6 mprj_io_holdover[15]
port 151 nsew signal input
rlabel metal2 s 627493 995407 627549 995887 6 mprj_io_ib_mode_sel[15]
port 152 nsew signal input
rlabel metal2 s 634301 995407 634357 995887 6 mprj_io_inp_dis[15]
port 153 nsew signal input
rlabel metal2 s 626849 995407 626905 995887 6 mprj_io_oeb[15]
port 154 nsew signal input
rlabel metal2 s 629977 995407 630033 995887 6 mprj_io_out[15]
port 155 nsew signal input
rlabel metal2 s 639177 995407 639233 995887 6 mprj_io_slow_sel[15]
port 156 nsew signal input
rlabel metal2 s 628137 995407 628193 995887 6 mprj_io_vtrip_sel[15]
port 157 nsew signal input
rlabel metal2 s 641017 995407 641073 995887 6 mprj_io_in[15]
port 158 nsew signal tristate
rlabel metal2 s 536733 995407 536789 995887 6 mprj_analog_io[9]
port 159 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 160 nsew signal bidirectional
rlabel metal2 s 534341 995407 534397 995887 6 mprj_io_analog_en[16]
port 161 nsew signal input
rlabel metal2 s 533053 995407 533109 995887 6 mprj_io_analog_pol[16]
port 162 nsew signal input
rlabel metal2 s 530017 995407 530073 995887 6 mprj_io_analog_sel[16]
port 163 nsew signal input
rlabel metal2 s 533697 995407 533753 995887 6 mprj_io_dm[48]
port 164 nsew signal input
rlabel metal2 s 535537 995407 535593 995887 6 mprj_io_dm[49]
port 165 nsew signal input
rlabel metal2 s 529373 995407 529429 995887 6 mprj_io_dm[50]
port 166 nsew signal input
rlabel metal2 s 531213 995407 531269 995887 6 mprj_io_enh[16]
port 167 nsew signal input
rlabel metal2 s 530569 995407 530625 995887 6 mprj_io_hldh_n[16]
port 168 nsew signal input
rlabel metal2 s 528729 995407 528785 995887 6 mprj_io_holdover[16]
port 169 nsew signal input
rlabel metal2 s 525693 995407 525749 995887 6 mprj_io_ib_mode_sel[16]
port 170 nsew signal input
rlabel metal2 s 532501 995407 532557 995887 6 mprj_io_inp_dis[16]
port 171 nsew signal input
rlabel metal2 s 525049 995407 525105 995887 6 mprj_io_oeb[16]
port 172 nsew signal input
rlabel metal2 s 528177 995407 528233 995887 6 mprj_io_out[16]
port 173 nsew signal input
rlabel metal2 s 537377 995407 537433 995887 6 mprj_io_slow_sel[16]
port 174 nsew signal input
rlabel metal2 s 526337 995407 526393 995887 6 mprj_io_vtrip_sel[16]
port 175 nsew signal input
rlabel metal2 s 539217 995407 539273 995887 6 mprj_io_in[16]
port 176 nsew signal tristate
rlabel metal2 s 485333 995407 485389 995887 6 mprj_analog_io[10]
port 177 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 178 nsew signal bidirectional
rlabel metal2 s 482941 995407 482997 995887 6 mprj_io_analog_en[17]
port 179 nsew signal input
rlabel metal2 s 481653 995407 481709 995887 6 mprj_io_analog_pol[17]
port 180 nsew signal input
rlabel metal2 s 478617 995407 478673 995887 6 mprj_io_analog_sel[17]
port 181 nsew signal input
rlabel metal2 s 482297 995407 482353 995887 6 mprj_io_dm[51]
port 182 nsew signal input
rlabel metal2 s 484137 995407 484193 995887 6 mprj_io_dm[52]
port 183 nsew signal input
rlabel metal2 s 477973 995407 478029 995887 6 mprj_io_dm[53]
port 184 nsew signal input
rlabel metal2 s 479813 995407 479869 995887 6 mprj_io_enh[17]
port 185 nsew signal input
rlabel metal2 s 479169 995407 479225 995887 6 mprj_io_hldh_n[17]
port 186 nsew signal input
rlabel metal2 s 477329 995407 477385 995887 6 mprj_io_holdover[17]
port 187 nsew signal input
rlabel metal2 s 474293 995407 474349 995887 6 mprj_io_ib_mode_sel[17]
port 188 nsew signal input
rlabel metal2 s 481101 995407 481157 995887 6 mprj_io_inp_dis[17]
port 189 nsew signal input
rlabel metal2 s 473649 995407 473705 995887 6 mprj_io_oeb[17]
port 190 nsew signal input
rlabel metal2 s 476777 995407 476833 995887 6 mprj_io_out[17]
port 191 nsew signal input
rlabel metal2 s 485977 995407 486033 995887 6 mprj_io_slow_sel[17]
port 192 nsew signal input
rlabel metal2 s 474937 995407 474993 995887 6 mprj_io_vtrip_sel[17]
port 193 nsew signal input
rlabel metal2 s 487817 995407 487873 995887 6 mprj_io_in[17]
port 194 nsew signal tristate
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 195 nsew signal bidirectional
rlabel metal2 s 675407 151003 675887 151059 6 mprj_io_analog_en[1]
port 196 nsew signal input
rlabel metal2 s 675407 152291 675887 152347 6 mprj_io_analog_pol[1]
port 197 nsew signal input
rlabel metal2 s 675407 155327 675887 155383 6 mprj_io_analog_sel[1]
port 198 nsew signal input
rlabel metal2 s 675407 151647 675887 151703 6 mprj_io_dm[3]
port 199 nsew signal input
rlabel metal2 s 675407 149807 675887 149863 6 mprj_io_dm[4]
port 200 nsew signal input
rlabel metal2 s 675407 155971 675887 156027 6 mprj_io_dm[5]
port 201 nsew signal input
rlabel metal2 s 675407 154131 675887 154187 6 mprj_io_enh[1]
port 202 nsew signal input
rlabel metal2 s 675407 154775 675887 154831 6 mprj_io_hldh_n[1]
port 203 nsew signal input
rlabel metal2 s 675407 156615 675887 156671 6 mprj_io_holdover[1]
port 204 nsew signal input
rlabel metal2 s 675407 159651 675887 159707 6 mprj_io_ib_mode_sel[1]
port 205 nsew signal input
rlabel metal2 s 675407 152843 675887 152899 6 mprj_io_inp_dis[1]
port 206 nsew signal input
rlabel metal2 s 675407 160295 675887 160351 6 mprj_io_oeb[1]
port 207 nsew signal input
rlabel metal2 s 675407 157167 675887 157223 6 mprj_io_out[1]
port 208 nsew signal input
rlabel metal2 s 675407 147967 675887 148023 6 mprj_io_slow_sel[1]
port 209 nsew signal input
rlabel metal2 s 675407 159007 675887 159063 6 mprj_io_vtrip_sel[1]
port 210 nsew signal input
rlabel metal2 s 675407 146127 675887 146183 6 mprj_io_in[1]
port 211 nsew signal tristate
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 212 nsew signal bidirectional
rlabel metal2 s 675407 196003 675887 196059 6 mprj_io_analog_en[2]
port 213 nsew signal input
rlabel metal2 s 675407 197291 675887 197347 6 mprj_io_analog_pol[2]
port 214 nsew signal input
rlabel metal2 s 675407 200327 675887 200383 6 mprj_io_analog_sel[2]
port 215 nsew signal input
rlabel metal2 s 675407 196647 675887 196703 6 mprj_io_dm[6]
port 216 nsew signal input
rlabel metal2 s 675407 194807 675887 194863 6 mprj_io_dm[7]
port 217 nsew signal input
rlabel metal2 s 675407 200971 675887 201027 6 mprj_io_dm[8]
port 218 nsew signal input
rlabel metal2 s 675407 199131 675887 199187 6 mprj_io_enh[2]
port 219 nsew signal input
rlabel metal2 s 675407 199775 675887 199831 6 mprj_io_hldh_n[2]
port 220 nsew signal input
rlabel metal2 s 675407 201615 675887 201671 6 mprj_io_holdover[2]
port 221 nsew signal input
rlabel metal2 s 675407 204651 675887 204707 6 mprj_io_ib_mode_sel[2]
port 222 nsew signal input
rlabel metal2 s 675407 197843 675887 197899 6 mprj_io_inp_dis[2]
port 223 nsew signal input
rlabel metal2 s 675407 205295 675887 205351 6 mprj_io_oeb[2]
port 224 nsew signal input
rlabel metal2 s 675407 202167 675887 202223 6 mprj_io_out[2]
port 225 nsew signal input
rlabel metal2 s 675407 192967 675887 193023 6 mprj_io_slow_sel[2]
port 226 nsew signal input
rlabel metal2 s 675407 204007 675887 204063 6 mprj_io_vtrip_sel[2]
port 227 nsew signal input
rlabel metal2 s 675407 191127 675887 191183 6 mprj_io_in[2]
port 228 nsew signal tristate
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 229 nsew signal bidirectional
rlabel metal2 s 675407 241203 675887 241259 6 mprj_io_analog_en[3]
port 230 nsew signal input
rlabel metal2 s 675407 242491 675887 242547 6 mprj_io_analog_pol[3]
port 231 nsew signal input
rlabel metal2 s 675407 245527 675887 245583 6 mprj_io_analog_sel[3]
port 232 nsew signal input
rlabel metal2 s 675407 240007 675887 240063 6 mprj_io_dm[10]
port 233 nsew signal input
rlabel metal2 s 675407 246171 675887 246227 6 mprj_io_dm[11]
port 234 nsew signal input
rlabel metal2 s 675407 241847 675887 241903 6 mprj_io_dm[9]
port 235 nsew signal input
rlabel metal2 s 675407 244331 675887 244387 6 mprj_io_enh[3]
port 236 nsew signal input
rlabel metal2 s 675407 244975 675887 245031 6 mprj_io_hldh_n[3]
port 237 nsew signal input
rlabel metal2 s 675407 246815 675887 246871 6 mprj_io_holdover[3]
port 238 nsew signal input
rlabel metal2 s 675407 249851 675887 249907 6 mprj_io_ib_mode_sel[3]
port 239 nsew signal input
rlabel metal2 s 675407 243043 675887 243099 6 mprj_io_inp_dis[3]
port 240 nsew signal input
rlabel metal2 s 675407 250495 675887 250551 6 mprj_io_oeb[3]
port 241 nsew signal input
rlabel metal2 s 675407 247367 675887 247423 6 mprj_io_out[3]
port 242 nsew signal input
rlabel metal2 s 675407 238167 675887 238223 6 mprj_io_slow_sel[3]
port 243 nsew signal input
rlabel metal2 s 675407 249207 675887 249263 6 mprj_io_vtrip_sel[3]
port 244 nsew signal input
rlabel metal2 s 675407 236327 675887 236383 6 mprj_io_in[3]
port 245 nsew signal tristate
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 246 nsew signal bidirectional
rlabel metal2 s 675407 286203 675887 286259 6 mprj_io_analog_en[4]
port 247 nsew signal input
rlabel metal2 s 675407 287491 675887 287547 6 mprj_io_analog_pol[4]
port 248 nsew signal input
rlabel metal2 s 675407 290527 675887 290583 6 mprj_io_analog_sel[4]
port 249 nsew signal input
rlabel metal2 s 675407 286847 675887 286903 6 mprj_io_dm[12]
port 250 nsew signal input
rlabel metal2 s 675407 285007 675887 285063 6 mprj_io_dm[13]
port 251 nsew signal input
rlabel metal2 s 675407 291171 675887 291227 6 mprj_io_dm[14]
port 252 nsew signal input
rlabel metal2 s 675407 289331 675887 289387 6 mprj_io_enh[4]
port 253 nsew signal input
rlabel metal2 s 675407 289975 675887 290031 6 mprj_io_hldh_n[4]
port 254 nsew signal input
rlabel metal2 s 675407 291815 675887 291871 6 mprj_io_holdover[4]
port 255 nsew signal input
rlabel metal2 s 675407 294851 675887 294907 6 mprj_io_ib_mode_sel[4]
port 256 nsew signal input
rlabel metal2 s 675407 288043 675887 288099 6 mprj_io_inp_dis[4]
port 257 nsew signal input
rlabel metal2 s 675407 295495 675887 295551 6 mprj_io_oeb[4]
port 258 nsew signal input
rlabel metal2 s 675407 292367 675887 292423 6 mprj_io_out[4]
port 259 nsew signal input
rlabel metal2 s 675407 283167 675887 283223 6 mprj_io_slow_sel[4]
port 260 nsew signal input
rlabel metal2 s 675407 294207 675887 294263 6 mprj_io_vtrip_sel[4]
port 261 nsew signal input
rlabel metal2 s 675407 281327 675887 281383 6 mprj_io_in[4]
port 262 nsew signal tristate
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 263 nsew signal bidirectional
rlabel metal2 s 675407 331203 675887 331259 6 mprj_io_analog_en[5]
port 264 nsew signal input
rlabel metal2 s 675407 332491 675887 332547 6 mprj_io_analog_pol[5]
port 265 nsew signal input
rlabel metal2 s 675407 335527 675887 335583 6 mprj_io_analog_sel[5]
port 266 nsew signal input
rlabel metal2 s 675407 331847 675887 331903 6 mprj_io_dm[15]
port 267 nsew signal input
rlabel metal2 s 675407 330007 675887 330063 6 mprj_io_dm[16]
port 268 nsew signal input
rlabel metal2 s 675407 336171 675887 336227 6 mprj_io_dm[17]
port 269 nsew signal input
rlabel metal2 s 675407 334331 675887 334387 6 mprj_io_enh[5]
port 270 nsew signal input
rlabel metal2 s 675407 334975 675887 335031 6 mprj_io_hldh_n[5]
port 271 nsew signal input
rlabel metal2 s 675407 336815 675887 336871 6 mprj_io_holdover[5]
port 272 nsew signal input
rlabel metal2 s 675407 339851 675887 339907 6 mprj_io_ib_mode_sel[5]
port 273 nsew signal input
rlabel metal2 s 675407 333043 675887 333099 6 mprj_io_inp_dis[5]
port 274 nsew signal input
rlabel metal2 s 675407 340495 675887 340551 6 mprj_io_oeb[5]
port 275 nsew signal input
rlabel metal2 s 675407 337367 675887 337423 6 mprj_io_out[5]
port 276 nsew signal input
rlabel metal2 s 675407 328167 675887 328223 6 mprj_io_slow_sel[5]
port 277 nsew signal input
rlabel metal2 s 675407 339207 675887 339263 6 mprj_io_vtrip_sel[5]
port 278 nsew signal input
rlabel metal2 s 675407 326327 675887 326383 6 mprj_io_in[5]
port 279 nsew signal tristate
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 280 nsew signal bidirectional
rlabel metal2 s 675407 376403 675887 376459 6 mprj_io_analog_en[6]
port 281 nsew signal input
rlabel metal2 s 675407 377691 675887 377747 6 mprj_io_analog_pol[6]
port 282 nsew signal input
rlabel metal2 s 675407 380727 675887 380783 6 mprj_io_analog_sel[6]
port 283 nsew signal input
rlabel metal2 s 675407 377047 675887 377103 6 mprj_io_dm[18]
port 284 nsew signal input
rlabel metal2 s 675407 375207 675887 375263 6 mprj_io_dm[19]
port 285 nsew signal input
rlabel metal2 s 675407 381371 675887 381427 6 mprj_io_dm[20]
port 286 nsew signal input
rlabel metal2 s 675407 379531 675887 379587 6 mprj_io_enh[6]
port 287 nsew signal input
rlabel metal2 s 675407 380175 675887 380231 6 mprj_io_hldh_n[6]
port 288 nsew signal input
rlabel metal2 s 675407 382015 675887 382071 6 mprj_io_holdover[6]
port 289 nsew signal input
rlabel metal2 s 675407 385051 675887 385107 6 mprj_io_ib_mode_sel[6]
port 290 nsew signal input
rlabel metal2 s 675407 378243 675887 378299 6 mprj_io_inp_dis[6]
port 291 nsew signal input
rlabel metal2 s 675407 385695 675887 385751 6 mprj_io_oeb[6]
port 292 nsew signal input
rlabel metal2 s 675407 382567 675887 382623 6 mprj_io_out[6]
port 293 nsew signal input
rlabel metal2 s 675407 373367 675887 373423 6 mprj_io_slow_sel[6]
port 294 nsew signal input
rlabel metal2 s 675407 384407 675887 384463 6 mprj_io_vtrip_sel[6]
port 295 nsew signal input
rlabel metal2 s 675407 371527 675887 371583 6 mprj_io_in[6]
port 296 nsew signal tristate
rlabel metal2 s 675407 551211 675887 551267 6 mprj_analog_io[0]
port 297 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 298 nsew signal bidirectional
rlabel metal2 s 675407 553603 675887 553659 6 mprj_io_analog_en[7]
port 299 nsew signal input
rlabel metal2 s 675407 554891 675887 554947 6 mprj_io_analog_pol[7]
port 300 nsew signal input
rlabel metal2 s 675407 557927 675887 557983 6 mprj_io_analog_sel[7]
port 301 nsew signal input
rlabel metal2 s 675407 554247 675887 554303 6 mprj_io_dm[21]
port 302 nsew signal input
rlabel metal2 s 675407 552407 675887 552463 6 mprj_io_dm[22]
port 303 nsew signal input
rlabel metal2 s 675407 558571 675887 558627 6 mprj_io_dm[23]
port 304 nsew signal input
rlabel metal2 s 675407 556731 675887 556787 6 mprj_io_enh[7]
port 305 nsew signal input
rlabel metal2 s 675407 557375 675887 557431 6 mprj_io_hldh_n[7]
port 306 nsew signal input
rlabel metal2 s 675407 559215 675887 559271 6 mprj_io_holdover[7]
port 307 nsew signal input
rlabel metal2 s 675407 562251 675887 562307 6 mprj_io_ib_mode_sel[7]
port 308 nsew signal input
rlabel metal2 s 675407 555443 675887 555499 6 mprj_io_inp_dis[7]
port 309 nsew signal input
rlabel metal2 s 675407 562895 675887 562951 6 mprj_io_oeb[7]
port 310 nsew signal input
rlabel metal2 s 675407 559767 675887 559823 6 mprj_io_out[7]
port 311 nsew signal input
rlabel metal2 s 675407 550567 675887 550623 6 mprj_io_slow_sel[7]
port 312 nsew signal input
rlabel metal2 s 675407 561607 675887 561663 6 mprj_io_vtrip_sel[7]
port 313 nsew signal input
rlabel metal2 s 675407 548727 675887 548783 6 mprj_io_in[7]
port 314 nsew signal tristate
rlabel metal2 s 675407 596411 675887 596467 6 mprj_analog_io[1]
port 315 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 316 nsew signal bidirectional
rlabel metal2 s 675407 598803 675887 598859 6 mprj_io_analog_en[8]
port 317 nsew signal input
rlabel metal2 s 675407 600091 675887 600147 6 mprj_io_analog_pol[8]
port 318 nsew signal input
rlabel metal2 s 675407 603127 675887 603183 6 mprj_io_analog_sel[8]
port 319 nsew signal input
rlabel metal2 s 675407 599447 675887 599503 6 mprj_io_dm[24]
port 320 nsew signal input
rlabel metal2 s 675407 597607 675887 597663 6 mprj_io_dm[25]
port 321 nsew signal input
rlabel metal2 s 675407 603771 675887 603827 6 mprj_io_dm[26]
port 322 nsew signal input
rlabel metal2 s 675407 601931 675887 601987 6 mprj_io_enh[8]
port 323 nsew signal input
rlabel metal2 s 675407 602575 675887 602631 6 mprj_io_hldh_n[8]
port 324 nsew signal input
rlabel metal2 s 675407 604415 675887 604471 6 mprj_io_holdover[8]
port 325 nsew signal input
rlabel metal2 s 675407 607451 675887 607507 6 mprj_io_ib_mode_sel[8]
port 326 nsew signal input
rlabel metal2 s 675407 600643 675887 600699 6 mprj_io_inp_dis[8]
port 327 nsew signal input
rlabel metal2 s 675407 608095 675887 608151 6 mprj_io_oeb[8]
port 328 nsew signal input
rlabel metal2 s 675407 604967 675887 605023 6 mprj_io_out[8]
port 329 nsew signal input
rlabel metal2 s 675407 595767 675887 595823 6 mprj_io_slow_sel[8]
port 330 nsew signal input
rlabel metal2 s 675407 606807 675887 606863 6 mprj_io_vtrip_sel[8]
port 331 nsew signal input
rlabel metal2 s 675407 593927 675887 593983 6 mprj_io_in[8]
port 332 nsew signal tristate
rlabel metal2 s 675407 641411 675887 641467 6 mprj_analog_io[2]
port 333 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 334 nsew signal bidirectional
rlabel metal2 s 675407 643803 675887 643859 6 mprj_io_analog_en[9]
port 335 nsew signal input
rlabel metal2 s 675407 645091 675887 645147 6 mprj_io_analog_pol[9]
port 336 nsew signal input
rlabel metal2 s 675407 648127 675887 648183 6 mprj_io_analog_sel[9]
port 337 nsew signal input
rlabel metal2 s 675407 644447 675887 644503 6 mprj_io_dm[27]
port 338 nsew signal input
rlabel metal2 s 675407 642607 675887 642663 6 mprj_io_dm[28]
port 339 nsew signal input
rlabel metal2 s 675407 648771 675887 648827 6 mprj_io_dm[29]
port 340 nsew signal input
rlabel metal2 s 675407 646931 675887 646987 6 mprj_io_enh[9]
port 341 nsew signal input
rlabel metal2 s 675407 647575 675887 647631 6 mprj_io_hldh_n[9]
port 342 nsew signal input
rlabel metal2 s 675407 649415 675887 649471 6 mprj_io_holdover[9]
port 343 nsew signal input
rlabel metal2 s 675407 652451 675887 652507 6 mprj_io_ib_mode_sel[9]
port 344 nsew signal input
rlabel metal2 s 675407 645643 675887 645699 6 mprj_io_inp_dis[9]
port 345 nsew signal input
rlabel metal2 s 675407 653095 675887 653151 6 mprj_io_oeb[9]
port 346 nsew signal input
rlabel metal2 s 675407 649967 675887 650023 6 mprj_io_out[9]
port 347 nsew signal input
rlabel metal2 s 675407 640767 675887 640823 6 mprj_io_slow_sel[9]
port 348 nsew signal input
rlabel metal2 s 675407 651807 675887 651863 6 mprj_io_vtrip_sel[9]
port 349 nsew signal input
rlabel metal2 s 675407 638927 675887 638983 6 mprj_io_in[9]
port 350 nsew signal tristate
rlabel metal2 s 396333 995407 396389 995887 6 mprj_analog_io[11]
port 351 nsew signal bidirectional
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 352 nsew signal bidirectional
rlabel metal2 s 393941 995407 393997 995887 6 mprj_io_analog_en[18]
port 353 nsew signal input
rlabel metal2 s 392653 995407 392709 995887 6 mprj_io_analog_pol[18]
port 354 nsew signal input
rlabel metal2 s 389617 995407 389673 995887 6 mprj_io_analog_sel[18]
port 355 nsew signal input
rlabel metal2 s 393297 995407 393353 995887 6 mprj_io_dm[54]
port 356 nsew signal input
rlabel metal2 s 395137 995407 395193 995887 6 mprj_io_dm[55]
port 357 nsew signal input
rlabel metal2 s 388973 995407 389029 995887 6 mprj_io_dm[56]
port 358 nsew signal input
rlabel metal2 s 390813 995407 390869 995887 6 mprj_io_enh[18]
port 359 nsew signal input
rlabel metal2 s 390169 995407 390225 995887 6 mprj_io_hldh_n[18]
port 360 nsew signal input
rlabel metal2 s 388329 995407 388385 995887 6 mprj_io_holdover[18]
port 361 nsew signal input
rlabel metal2 s 385293 995407 385349 995887 6 mprj_io_ib_mode_sel[18]
port 362 nsew signal input
rlabel metal2 s 392101 995407 392157 995887 6 mprj_io_inp_dis[18]
port 363 nsew signal input
rlabel metal2 s 384649 995407 384705 995887 6 mprj_io_oeb[18]
port 364 nsew signal input
rlabel metal2 s 387777 995407 387833 995887 6 mprj_io_out[18]
port 365 nsew signal input
rlabel metal2 s 396977 995407 397033 995887 6 mprj_io_slow_sel[18]
port 366 nsew signal input
rlabel metal2 s 385937 995407 385993 995887 6 mprj_io_vtrip_sel[18]
port 367 nsew signal input
rlabel metal2 s 398817 995407 398873 995887 6 mprj_io_in[18]
port 368 nsew signal tristate
rlabel metal2 s 41713 667333 42193 667389 6 mprj_analog_io[21]
port 369 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 370 nsew signal bidirectional
rlabel metal2 s 41713 664941 42193 664997 6 mprj_io_analog_en[28]
port 371 nsew signal input
rlabel metal2 s 41713 663653 42193 663709 6 mprj_io_analog_pol[28]
port 372 nsew signal input
rlabel metal2 s 41713 660617 42193 660673 6 mprj_io_analog_sel[28]
port 373 nsew signal input
rlabel metal2 s 41713 664297 42193 664353 6 mprj_io_dm[84]
port 374 nsew signal input
rlabel metal2 s 41713 666137 42193 666193 6 mprj_io_dm[85]
port 375 nsew signal input
rlabel metal2 s 41713 659973 42193 660029 6 mprj_io_dm[86]
port 376 nsew signal input
rlabel metal2 s 41713 661813 42193 661869 6 mprj_io_enh[28]
port 377 nsew signal input
rlabel metal2 s 41713 661169 42193 661225 6 mprj_io_hldh_n[28]
port 378 nsew signal input
rlabel metal2 s 41713 659329 42193 659385 6 mprj_io_holdover[28]
port 379 nsew signal input
rlabel metal2 s 41713 656293 42193 656349 6 mprj_io_ib_mode_sel[28]
port 380 nsew signal input
rlabel metal2 s 41713 663101 42193 663157 6 mprj_io_inp_dis[28]
port 381 nsew signal input
rlabel metal2 s 41713 655649 42193 655705 6 mprj_io_oeb[28]
port 382 nsew signal input
rlabel metal2 s 41713 658777 42193 658833 6 mprj_io_out[28]
port 383 nsew signal input
rlabel metal2 s 41713 667977 42193 668033 6 mprj_io_slow_sel[28]
port 384 nsew signal input
rlabel metal2 s 41713 656937 42193 656993 6 mprj_io_vtrip_sel[28]
port 385 nsew signal input
rlabel metal2 s 41713 669817 42193 669873 6 mprj_io_in[28]
port 386 nsew signal tristate
rlabel metal2 s 41713 624133 42193 624189 6 mprj_analog_io[22]
port 387 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 388 nsew signal bidirectional
rlabel metal2 s 41713 621741 42193 621797 6 mprj_io_analog_en[29]
port 389 nsew signal input
rlabel metal2 s 41713 620453 42193 620509 6 mprj_io_analog_pol[29]
port 390 nsew signal input
rlabel metal2 s 41713 617417 42193 617473 6 mprj_io_analog_sel[29]
port 391 nsew signal input
rlabel metal2 s 41713 621097 42193 621153 6 mprj_io_dm[87]
port 392 nsew signal input
rlabel metal2 s 41713 622937 42193 622993 6 mprj_io_dm[88]
port 393 nsew signal input
rlabel metal2 s 41713 616773 42193 616829 6 mprj_io_dm[89]
port 394 nsew signal input
rlabel metal2 s 41713 618613 42193 618669 6 mprj_io_enh[29]
port 395 nsew signal input
rlabel metal2 s 41713 617969 42193 618025 6 mprj_io_hldh_n[29]
port 396 nsew signal input
rlabel metal2 s 41713 616129 42193 616185 6 mprj_io_holdover[29]
port 397 nsew signal input
rlabel metal2 s 41713 613093 42193 613149 6 mprj_io_ib_mode_sel[29]
port 398 nsew signal input
rlabel metal2 s 41713 619901 42193 619957 6 mprj_io_inp_dis[29]
port 399 nsew signal input
rlabel metal2 s 41713 612449 42193 612505 6 mprj_io_oeb[29]
port 400 nsew signal input
rlabel metal2 s 41713 615577 42193 615633 6 mprj_io_out[29]
port 401 nsew signal input
rlabel metal2 s 41713 624777 42193 624833 6 mprj_io_slow_sel[29]
port 402 nsew signal input
rlabel metal2 s 41713 613737 42193 613793 6 mprj_io_vtrip_sel[29]
port 403 nsew signal input
rlabel metal2 s 41713 626617 42193 626673 6 mprj_io_in[29]
port 404 nsew signal tristate
rlabel metal2 s 41713 580933 42193 580989 6 mprj_analog_io[23]
port 405 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 406 nsew signal bidirectional
rlabel metal2 s 41713 578541 42193 578597 6 mprj_io_analog_en[30]
port 407 nsew signal input
rlabel metal2 s 41713 577253 42193 577309 6 mprj_io_analog_pol[30]
port 408 nsew signal input
rlabel metal2 s 41713 574217 42193 574273 6 mprj_io_analog_sel[30]
port 409 nsew signal input
rlabel metal2 s 41713 577897 42193 577953 6 mprj_io_dm[90]
port 410 nsew signal input
rlabel metal2 s 41713 579737 42193 579793 6 mprj_io_dm[91]
port 411 nsew signal input
rlabel metal2 s 41713 573573 42193 573629 6 mprj_io_dm[92]
port 412 nsew signal input
rlabel metal2 s 41713 575413 42193 575469 6 mprj_io_enh[30]
port 413 nsew signal input
rlabel metal2 s 41713 574769 42193 574825 6 mprj_io_hldh_n[30]
port 414 nsew signal input
rlabel metal2 s 41713 572929 42193 572985 6 mprj_io_holdover[30]
port 415 nsew signal input
rlabel metal2 s 41713 569893 42193 569949 6 mprj_io_ib_mode_sel[30]
port 416 nsew signal input
rlabel metal2 s 41713 576701 42193 576757 6 mprj_io_inp_dis[30]
port 417 nsew signal input
rlabel metal2 s 41713 569249 42193 569305 6 mprj_io_oeb[30]
port 418 nsew signal input
rlabel metal2 s 41713 572377 42193 572433 6 mprj_io_out[30]
port 419 nsew signal input
rlabel metal2 s 41713 581577 42193 581633 6 mprj_io_slow_sel[30]
port 420 nsew signal input
rlabel metal2 s 41713 570537 42193 570593 6 mprj_io_vtrip_sel[30]
port 421 nsew signal input
rlabel metal2 s 41713 583417 42193 583473 6 mprj_io_in[30]
port 422 nsew signal tristate
rlabel metal2 s 41713 537733 42193 537789 6 mprj_analog_io[24]
port 423 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 424 nsew signal bidirectional
rlabel metal2 s 41713 535341 42193 535397 6 mprj_io_analog_en[31]
port 425 nsew signal input
rlabel metal2 s 41713 534053 42193 534109 6 mprj_io_analog_pol[31]
port 426 nsew signal input
rlabel metal2 s 41713 531017 42193 531073 6 mprj_io_analog_sel[31]
port 427 nsew signal input
rlabel metal2 s 41713 534697 42193 534753 6 mprj_io_dm[93]
port 428 nsew signal input
rlabel metal2 s 41713 536537 42193 536593 6 mprj_io_dm[94]
port 429 nsew signal input
rlabel metal2 s 41713 530373 42193 530429 6 mprj_io_dm[95]
port 430 nsew signal input
rlabel metal2 s 41713 532213 42193 532269 6 mprj_io_enh[31]
port 431 nsew signal input
rlabel metal2 s 41713 531569 42193 531625 6 mprj_io_hldh_n[31]
port 432 nsew signal input
rlabel metal2 s 41713 529729 42193 529785 6 mprj_io_holdover[31]
port 433 nsew signal input
rlabel metal2 s 41713 526693 42193 526749 6 mprj_io_ib_mode_sel[31]
port 434 nsew signal input
rlabel metal2 s 41713 533501 42193 533557 6 mprj_io_inp_dis[31]
port 435 nsew signal input
rlabel metal2 s 41713 526049 42193 526105 6 mprj_io_oeb[31]
port 436 nsew signal input
rlabel metal2 s 41713 529177 42193 529233 6 mprj_io_out[31]
port 437 nsew signal input
rlabel metal2 s 41713 538377 42193 538433 6 mprj_io_slow_sel[31]
port 438 nsew signal input
rlabel metal2 s 41713 527337 42193 527393 6 mprj_io_vtrip_sel[31]
port 439 nsew signal input
rlabel metal2 s 41713 540217 42193 540273 6 mprj_io_in[31]
port 440 nsew signal tristate
rlabel metal2 s 41713 410133 42193 410189 6 mprj_analog_io[25]
port 441 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 442 nsew signal bidirectional
rlabel metal2 s 41713 407741 42193 407797 6 mprj_io_analog_en[32]
port 443 nsew signal input
rlabel metal2 s 41713 406453 42193 406509 6 mprj_io_analog_pol[32]
port 444 nsew signal input
rlabel metal2 s 41713 403417 42193 403473 6 mprj_io_analog_sel[32]
port 445 nsew signal input
rlabel metal2 s 41713 407097 42193 407153 6 mprj_io_dm[96]
port 446 nsew signal input
rlabel metal2 s 41713 408937 42193 408993 6 mprj_io_dm[97]
port 447 nsew signal input
rlabel metal2 s 41713 402773 42193 402829 6 mprj_io_dm[98]
port 448 nsew signal input
rlabel metal2 s 41713 404613 42193 404669 6 mprj_io_enh[32]
port 449 nsew signal input
rlabel metal2 s 41713 403969 42193 404025 6 mprj_io_hldh_n[32]
port 450 nsew signal input
rlabel metal2 s 41713 402129 42193 402185 6 mprj_io_holdover[32]
port 451 nsew signal input
rlabel metal2 s 41713 399093 42193 399149 6 mprj_io_ib_mode_sel[32]
port 452 nsew signal input
rlabel metal2 s 41713 405901 42193 405957 6 mprj_io_inp_dis[32]
port 453 nsew signal input
rlabel metal2 s 41713 398449 42193 398505 6 mprj_io_oeb[32]
port 454 nsew signal input
rlabel metal2 s 41713 401577 42193 401633 6 mprj_io_out[32]
port 455 nsew signal input
rlabel metal2 s 41713 410777 42193 410833 6 mprj_io_slow_sel[32]
port 456 nsew signal input
rlabel metal2 s 41713 399737 42193 399793 6 mprj_io_vtrip_sel[32]
port 457 nsew signal input
rlabel metal2 s 41713 412617 42193 412673 6 mprj_io_in[32]
port 458 nsew signal tristate
rlabel metal2 s 41713 366933 42193 366989 6 mprj_analog_io[26]
port 459 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 460 nsew signal bidirectional
rlabel metal2 s 41713 364541 42193 364597 6 mprj_io_analog_en[33]
port 461 nsew signal input
rlabel metal2 s 41713 363253 42193 363309 6 mprj_io_analog_pol[33]
port 462 nsew signal input
rlabel metal2 s 41713 360217 42193 360273 6 mprj_io_analog_sel[33]
port 463 nsew signal input
rlabel metal2 s 41713 365737 42193 365793 6 mprj_io_dm[100]
port 464 nsew signal input
rlabel metal2 s 41713 359573 42193 359629 6 mprj_io_dm[101]
port 465 nsew signal input
rlabel metal2 s 41713 363897 42193 363953 6 mprj_io_dm[99]
port 466 nsew signal input
rlabel metal2 s 41713 361413 42193 361469 6 mprj_io_enh[33]
port 467 nsew signal input
rlabel metal2 s 41713 360769 42193 360825 6 mprj_io_hldh_n[33]
port 468 nsew signal input
rlabel metal2 s 41713 358929 42193 358985 6 mprj_io_holdover[33]
port 469 nsew signal input
rlabel metal2 s 41713 355893 42193 355949 6 mprj_io_ib_mode_sel[33]
port 470 nsew signal input
rlabel metal2 s 41713 362701 42193 362757 6 mprj_io_inp_dis[33]
port 471 nsew signal input
rlabel metal2 s 41713 355249 42193 355305 6 mprj_io_oeb[33]
port 472 nsew signal input
rlabel metal2 s 41713 358377 42193 358433 6 mprj_io_out[33]
port 473 nsew signal input
rlabel metal2 s 41713 367577 42193 367633 6 mprj_io_slow_sel[33]
port 474 nsew signal input
rlabel metal2 s 41713 356537 42193 356593 6 mprj_io_vtrip_sel[33]
port 475 nsew signal input
rlabel metal2 s 41713 369417 42193 369473 6 mprj_io_in[33]
port 476 nsew signal tristate
rlabel metal2 s 41713 323733 42193 323789 6 mprj_analog_io[27]
port 477 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 478 nsew signal bidirectional
rlabel metal2 s 41713 321341 42193 321397 6 mprj_io_analog_en[34]
port 479 nsew signal input
rlabel metal2 s 41713 320053 42193 320109 6 mprj_io_analog_pol[34]
port 480 nsew signal input
rlabel metal2 s 41713 317017 42193 317073 6 mprj_io_analog_sel[34]
port 481 nsew signal input
rlabel metal2 s 41713 320697 42193 320753 6 mprj_io_dm[102]
port 482 nsew signal input
rlabel metal2 s 41713 322537 42193 322593 6 mprj_io_dm[103]
port 483 nsew signal input
rlabel metal2 s 41713 316373 42193 316429 6 mprj_io_dm[104]
port 484 nsew signal input
rlabel metal2 s 41713 318213 42193 318269 6 mprj_io_enh[34]
port 485 nsew signal input
rlabel metal2 s 41713 317569 42193 317625 6 mprj_io_hldh_n[34]
port 486 nsew signal input
rlabel metal2 s 41713 315729 42193 315785 6 mprj_io_holdover[34]
port 487 nsew signal input
rlabel metal2 s 41713 312693 42193 312749 6 mprj_io_ib_mode_sel[34]
port 488 nsew signal input
rlabel metal2 s 41713 319501 42193 319557 6 mprj_io_inp_dis[34]
port 489 nsew signal input
rlabel metal2 s 41713 312049 42193 312105 6 mprj_io_oeb[34]
port 490 nsew signal input
rlabel metal2 s 41713 315177 42193 315233 6 mprj_io_out[34]
port 491 nsew signal input
rlabel metal2 s 41713 324377 42193 324433 6 mprj_io_slow_sel[34]
port 492 nsew signal input
rlabel metal2 s 41713 313337 42193 313393 6 mprj_io_vtrip_sel[34]
port 493 nsew signal input
rlabel metal2 s 41713 326217 42193 326273 6 mprj_io_in[34]
port 494 nsew signal tristate
rlabel metal2 s 41713 280533 42193 280589 6 mprj_analog_io[28]
port 495 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 496 nsew signal bidirectional
rlabel metal2 s 41713 278141 42193 278197 6 mprj_io_analog_en[35]
port 497 nsew signal input
rlabel metal2 s 41713 276853 42193 276909 6 mprj_io_analog_pol[35]
port 498 nsew signal input
rlabel metal2 s 41713 273817 42193 273873 6 mprj_io_analog_sel[35]
port 499 nsew signal input
rlabel metal2 s 41713 277497 42193 277553 6 mprj_io_dm[105]
port 500 nsew signal input
rlabel metal2 s 41713 279337 42193 279393 6 mprj_io_dm[106]
port 501 nsew signal input
rlabel metal2 s 41713 273173 42193 273229 6 mprj_io_dm[107]
port 502 nsew signal input
rlabel metal2 s 41713 275013 42193 275069 6 mprj_io_enh[35]
port 503 nsew signal input
rlabel metal2 s 41713 274369 42193 274425 6 mprj_io_hldh_n[35]
port 504 nsew signal input
rlabel metal2 s 41713 272529 42193 272585 6 mprj_io_holdover[35]
port 505 nsew signal input
rlabel metal2 s 41713 269493 42193 269549 6 mprj_io_ib_mode_sel[35]
port 506 nsew signal input
rlabel metal2 s 41713 276301 42193 276357 6 mprj_io_inp_dis[35]
port 507 nsew signal input
rlabel metal2 s 41713 268849 42193 268905 6 mprj_io_oeb[35]
port 508 nsew signal input
rlabel metal2 s 41713 271977 42193 272033 6 mprj_io_out[35]
port 509 nsew signal input
rlabel metal2 s 41713 281177 42193 281233 6 mprj_io_slow_sel[35]
port 510 nsew signal input
rlabel metal2 s 41713 270137 42193 270193 6 mprj_io_vtrip_sel[35]
port 511 nsew signal input
rlabel metal2 s 41713 283017 42193 283073 6 mprj_io_in[35]
port 512 nsew signal tristate
rlabel metal2 s 41713 237333 42193 237389 6 mprj_analog_io[29]
port 513 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 514 nsew signal bidirectional
rlabel metal2 s 41713 234941 42193 234997 6 mprj_io_analog_en[36]
port 515 nsew signal input
rlabel metal2 s 41713 233653 42193 233709 6 mprj_io_analog_pol[36]
port 516 nsew signal input
rlabel metal2 s 41713 230617 42193 230673 6 mprj_io_analog_sel[36]
port 517 nsew signal input
rlabel metal2 s 41713 234297 42193 234353 6 mprj_io_dm[108]
port 518 nsew signal input
rlabel metal2 s 41713 236137 42193 236193 6 mprj_io_dm[109]
port 519 nsew signal input
rlabel metal2 s 41713 229973 42193 230029 6 mprj_io_dm[110]
port 520 nsew signal input
rlabel metal2 s 41713 231813 42193 231869 6 mprj_io_enh[36]
port 521 nsew signal input
rlabel metal2 s 41713 231169 42193 231225 6 mprj_io_hldh_n[36]
port 522 nsew signal input
rlabel metal2 s 41713 229329 42193 229385 6 mprj_io_holdover[36]
port 523 nsew signal input
rlabel metal2 s 41713 226293 42193 226349 6 mprj_io_ib_mode_sel[36]
port 524 nsew signal input
rlabel metal2 s 41713 233101 42193 233157 6 mprj_io_inp_dis[36]
port 525 nsew signal input
rlabel metal2 s 41713 225649 42193 225705 6 mprj_io_oeb[36]
port 526 nsew signal input
rlabel metal2 s 41713 228777 42193 228833 6 mprj_io_out[36]
port 527 nsew signal input
rlabel metal2 s 41713 237977 42193 238033 6 mprj_io_slow_sel[36]
port 528 nsew signal input
rlabel metal2 s 41713 226937 42193 226993 6 mprj_io_vtrip_sel[36]
port 529 nsew signal input
rlabel metal2 s 41713 239817 42193 239873 6 mprj_io_in[36]
port 530 nsew signal tristate
rlabel metal2 s 41713 194133 42193 194189 6 mprj_analog_io[30]
port 531 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 532 nsew signal bidirectional
rlabel metal2 s 41713 191741 42193 191797 6 mprj_io_analog_en[37]
port 533 nsew signal input
rlabel metal2 s 41713 190453 42193 190509 6 mprj_io_analog_pol[37]
port 534 nsew signal input
rlabel metal2 s 41713 187417 42193 187473 6 mprj_io_analog_sel[37]
port 535 nsew signal input
rlabel metal2 s 41713 191097 42193 191153 6 mprj_io_dm[111]
port 536 nsew signal input
rlabel metal2 s 41713 192937 42193 192993 6 mprj_io_dm[112]
port 537 nsew signal input
rlabel metal2 s 41713 186773 42193 186829 6 mprj_io_dm[113]
port 538 nsew signal input
rlabel metal2 s 41713 188613 42193 188669 6 mprj_io_enh[37]
port 539 nsew signal input
rlabel metal2 s 41713 187969 42193 188025 6 mprj_io_hldh_n[37]
port 540 nsew signal input
rlabel metal2 s 41713 186129 42193 186185 6 mprj_io_holdover[37]
port 541 nsew signal input
rlabel metal2 s 41713 183093 42193 183149 6 mprj_io_ib_mode_sel[37]
port 542 nsew signal input
rlabel metal2 s 41713 189901 42193 189957 6 mprj_io_inp_dis[37]
port 543 nsew signal input
rlabel metal2 s 41713 182449 42193 182505 6 mprj_io_oeb[37]
port 544 nsew signal input
rlabel metal2 s 41713 185577 42193 185633 6 mprj_io_out[37]
port 545 nsew signal input
rlabel metal2 s 41713 194777 42193 194833 6 mprj_io_slow_sel[37]
port 546 nsew signal input
rlabel metal2 s 41713 183737 42193 183793 6 mprj_io_vtrip_sel[37]
port 547 nsew signal input
rlabel metal2 s 41713 196617 42193 196673 6 mprj_io_in[37]
port 548 nsew signal tristate
rlabel metal2 s 294533 995407 294589 995887 6 mprj_analog_io[12]
port 549 nsew signal bidirectional
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 550 nsew signal bidirectional
rlabel metal2 s 292141 995407 292197 995887 6 mprj_io_analog_en[19]
port 551 nsew signal input
rlabel metal2 s 290853 995407 290909 995887 6 mprj_io_analog_pol[19]
port 552 nsew signal input
rlabel metal2 s 287817 995407 287873 995887 6 mprj_io_analog_sel[19]
port 553 nsew signal input
rlabel metal2 s 291497 995407 291553 995887 6 mprj_io_dm[57]
port 554 nsew signal input
rlabel metal2 s 293337 995407 293393 995887 6 mprj_io_dm[58]
port 555 nsew signal input
rlabel metal2 s 287173 995407 287229 995887 6 mprj_io_dm[59]
port 556 nsew signal input
rlabel metal2 s 289013 995407 289069 995887 6 mprj_io_enh[19]
port 557 nsew signal input
rlabel metal2 s 288369 995407 288425 995887 6 mprj_io_hldh_n[19]
port 558 nsew signal input
rlabel metal2 s 286529 995407 286585 995887 6 mprj_io_holdover[19]
port 559 nsew signal input
rlabel metal2 s 283493 995407 283549 995887 6 mprj_io_ib_mode_sel[19]
port 560 nsew signal input
rlabel metal2 s 290301 995407 290357 995887 6 mprj_io_inp_dis[19]
port 561 nsew signal input
rlabel metal2 s 282849 995407 282905 995887 6 mprj_io_oeb[19]
port 562 nsew signal input
rlabel metal2 s 285977 995407 286033 995887 6 mprj_io_out[19]
port 563 nsew signal input
rlabel metal2 s 295177 995407 295233 995887 6 mprj_io_slow_sel[19]
port 564 nsew signal input
rlabel metal2 s 284137 995407 284193 995887 6 mprj_io_vtrip_sel[19]
port 565 nsew signal input
rlabel metal2 s 297017 995407 297073 995887 6 mprj_io_in[19]
port 566 nsew signal tristate
rlabel metal2 s 242933 995407 242989 995887 6 mprj_analog_io[13]
port 567 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 568 nsew signal bidirectional
rlabel metal2 s 240541 995407 240597 995887 6 mprj_io_analog_en[20]
port 569 nsew signal input
rlabel metal2 s 239253 995407 239309 995887 6 mprj_io_analog_pol[20]
port 570 nsew signal input
rlabel metal2 s 236217 995407 236273 995887 6 mprj_io_analog_sel[20]
port 571 nsew signal input
rlabel metal2 s 239897 995407 239953 995887 6 mprj_io_dm[60]
port 572 nsew signal input
rlabel metal2 s 241737 995407 241793 995887 6 mprj_io_dm[61]
port 573 nsew signal input
rlabel metal2 s 235573 995407 235629 995887 6 mprj_io_dm[62]
port 574 nsew signal input
rlabel metal2 s 237413 995407 237469 995887 6 mprj_io_enh[20]
port 575 nsew signal input
rlabel metal2 s 236769 995407 236825 995887 6 mprj_io_hldh_n[20]
port 576 nsew signal input
rlabel metal2 s 234929 995407 234985 995887 6 mprj_io_holdover[20]
port 577 nsew signal input
rlabel metal2 s 231893 995407 231949 995887 6 mprj_io_ib_mode_sel[20]
port 578 nsew signal input
rlabel metal2 s 238701 995407 238757 995887 6 mprj_io_inp_dis[20]
port 579 nsew signal input
rlabel metal2 s 231249 995407 231305 995887 6 mprj_io_oeb[20]
port 580 nsew signal input
rlabel metal2 s 234377 995407 234433 995887 6 mprj_io_out[20]
port 581 nsew signal input
rlabel metal2 s 243577 995407 243633 995887 6 mprj_io_slow_sel[20]
port 582 nsew signal input
rlabel metal2 s 232537 995407 232593 995887 6 mprj_io_vtrip_sel[20]
port 583 nsew signal input
rlabel metal2 s 245417 995407 245473 995887 6 mprj_io_in[20]
port 584 nsew signal tristate
rlabel metal2 s 191533 995407 191589 995887 6 mprj_analog_io[14]
port 585 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 586 nsew signal bidirectional
rlabel metal2 s 189141 995407 189197 995887 6 mprj_io_analog_en[21]
port 587 nsew signal input
rlabel metal2 s 187853 995407 187909 995887 6 mprj_io_analog_pol[21]
port 588 nsew signal input
rlabel metal2 s 184817 995407 184873 995887 6 mprj_io_analog_sel[21]
port 589 nsew signal input
rlabel metal2 s 188497 995407 188553 995887 6 mprj_io_dm[63]
port 590 nsew signal input
rlabel metal2 s 190337 995407 190393 995887 6 mprj_io_dm[64]
port 591 nsew signal input
rlabel metal2 s 184173 995407 184229 995887 6 mprj_io_dm[65]
port 592 nsew signal input
rlabel metal2 s 186013 995407 186069 995887 6 mprj_io_enh[21]
port 593 nsew signal input
rlabel metal2 s 185369 995407 185425 995887 6 mprj_io_hldh_n[21]
port 594 nsew signal input
rlabel metal2 s 183529 995407 183585 995887 6 mprj_io_holdover[21]
port 595 nsew signal input
rlabel metal2 s 180493 995407 180549 995887 6 mprj_io_ib_mode_sel[21]
port 596 nsew signal input
rlabel metal2 s 187301 995407 187357 995887 6 mprj_io_inp_dis[21]
port 597 nsew signal input
rlabel metal2 s 179849 995407 179905 995887 6 mprj_io_oeb[21]
port 598 nsew signal input
rlabel metal2 s 182977 995407 183033 995887 6 mprj_io_out[21]
port 599 nsew signal input
rlabel metal2 s 192177 995407 192233 995887 6 mprj_io_slow_sel[21]
port 600 nsew signal input
rlabel metal2 s 181137 995407 181193 995887 6 mprj_io_vtrip_sel[21]
port 601 nsew signal input
rlabel metal2 s 194017 995407 194073 995887 6 mprj_io_in[21]
port 602 nsew signal tristate
rlabel metal2 s 140133 995407 140189 995887 6 mprj_analog_io[15]
port 603 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 604 nsew signal bidirectional
rlabel metal2 s 137741 995407 137797 995887 6 mprj_io_analog_en[22]
port 605 nsew signal input
rlabel metal2 s 136453 995407 136509 995887 6 mprj_io_analog_pol[22]
port 606 nsew signal input
rlabel metal2 s 133417 995407 133473 995887 6 mprj_io_analog_sel[22]
port 607 nsew signal input
rlabel metal2 s 137097 995407 137153 995887 6 mprj_io_dm[66]
port 608 nsew signal input
rlabel metal2 s 138937 995407 138993 995887 6 mprj_io_dm[67]
port 609 nsew signal input
rlabel metal2 s 132773 995407 132829 995887 6 mprj_io_dm[68]
port 610 nsew signal input
rlabel metal2 s 134613 995407 134669 995887 6 mprj_io_enh[22]
port 611 nsew signal input
rlabel metal2 s 133969 995407 134025 995887 6 mprj_io_hldh_n[22]
port 612 nsew signal input
rlabel metal2 s 132129 995407 132185 995887 6 mprj_io_holdover[22]
port 613 nsew signal input
rlabel metal2 s 129093 995407 129149 995887 6 mprj_io_ib_mode_sel[22]
port 614 nsew signal input
rlabel metal2 s 135901 995407 135957 995887 6 mprj_io_inp_dis[22]
port 615 nsew signal input
rlabel metal2 s 128449 995407 128505 995887 6 mprj_io_oeb[22]
port 616 nsew signal input
rlabel metal2 s 131577 995407 131633 995887 6 mprj_io_out[22]
port 617 nsew signal input
rlabel metal2 s 140777 995407 140833 995887 6 mprj_io_slow_sel[22]
port 618 nsew signal input
rlabel metal2 s 129737 995407 129793 995887 6 mprj_io_vtrip_sel[22]
port 619 nsew signal input
rlabel metal2 s 142617 995407 142673 995887 6 mprj_io_in[22]
port 620 nsew signal tristate
rlabel metal2 s 88733 995407 88789 995887 6 mprj_analog_io[16]
port 621 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 622 nsew signal bidirectional
rlabel metal2 s 86341 995407 86397 995887 6 mprj_io_analog_en[23]
port 623 nsew signal input
rlabel metal2 s 85053 995407 85109 995887 6 mprj_io_analog_pol[23]
port 624 nsew signal input
rlabel metal2 s 82017 995407 82073 995887 6 mprj_io_analog_sel[23]
port 625 nsew signal input
rlabel metal2 s 85697 995407 85753 995887 6 mprj_io_dm[69]
port 626 nsew signal input
rlabel metal2 s 87537 995407 87593 995887 6 mprj_io_dm[70]
port 627 nsew signal input
rlabel metal2 s 81373 995407 81429 995887 6 mprj_io_dm[71]
port 628 nsew signal input
rlabel metal2 s 83213 995407 83269 995887 6 mprj_io_enh[23]
port 629 nsew signal input
rlabel metal2 s 82569 995407 82625 995887 6 mprj_io_hldh_n[23]
port 630 nsew signal input
rlabel metal2 s 80729 995407 80785 995887 6 mprj_io_holdover[23]
port 631 nsew signal input
rlabel metal2 s 77693 995407 77749 995887 6 mprj_io_ib_mode_sel[23]
port 632 nsew signal input
rlabel metal2 s 84501 995407 84557 995887 6 mprj_io_inp_dis[23]
port 633 nsew signal input
rlabel metal2 s 77049 995407 77105 995887 6 mprj_io_oeb[23]
port 634 nsew signal input
rlabel metal2 s 80177 995407 80233 995887 6 mprj_io_out[23]
port 635 nsew signal input
rlabel metal2 s 89377 995407 89433 995887 6 mprj_io_slow_sel[23]
port 636 nsew signal input
rlabel metal2 s 78337 995407 78393 995887 6 mprj_io_vtrip_sel[23]
port 637 nsew signal input
rlabel metal2 s 91217 995407 91273 995887 6 mprj_io_in[23]
port 638 nsew signal tristate
rlabel metal2 s 41713 966733 42193 966789 6 mprj_analog_io[17]
port 639 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 640 nsew signal bidirectional
rlabel metal2 s 41713 964341 42193 964397 6 mprj_io_analog_en[24]
port 641 nsew signal input
rlabel metal2 s 41713 963053 42193 963109 6 mprj_io_analog_pol[24]
port 642 nsew signal input
rlabel metal2 s 41713 960017 42193 960073 6 mprj_io_analog_sel[24]
port 643 nsew signal input
rlabel metal2 s 41713 963697 42193 963753 6 mprj_io_dm[72]
port 644 nsew signal input
rlabel metal2 s 41713 965537 42193 965593 6 mprj_io_dm[73]
port 645 nsew signal input
rlabel metal2 s 41713 959373 42193 959429 6 mprj_io_dm[74]
port 646 nsew signal input
rlabel metal2 s 41713 961213 42193 961269 6 mprj_io_enh[24]
port 647 nsew signal input
rlabel metal2 s 41713 960569 42193 960625 6 mprj_io_hldh_n[24]
port 648 nsew signal input
rlabel metal2 s 41713 958729 42193 958785 6 mprj_io_holdover[24]
port 649 nsew signal input
rlabel metal2 s 41713 955693 42193 955749 6 mprj_io_ib_mode_sel[24]
port 650 nsew signal input
rlabel metal2 s 41713 962501 42193 962557 6 mprj_io_inp_dis[24]
port 651 nsew signal input
rlabel metal2 s 41713 955049 42193 955105 6 mprj_io_oeb[24]
port 652 nsew signal input
rlabel metal2 s 41713 958177 42193 958233 6 mprj_io_out[24]
port 653 nsew signal input
rlabel metal2 s 41713 967377 42193 967433 6 mprj_io_slow_sel[24]
port 654 nsew signal input
rlabel metal2 s 41713 956337 42193 956393 6 mprj_io_vtrip_sel[24]
port 655 nsew signal input
rlabel metal2 s 41713 969217 42193 969273 6 mprj_io_in[24]
port 656 nsew signal tristate
rlabel metal2 s 41713 796933 42193 796989 6 mprj_analog_io[18]
port 657 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 658 nsew signal bidirectional
rlabel metal2 s 41713 794541 42193 794597 6 mprj_io_analog_en[25]
port 659 nsew signal input
rlabel metal2 s 41713 793253 42193 793309 6 mprj_io_analog_pol[25]
port 660 nsew signal input
rlabel metal2 s 41713 790217 42193 790273 6 mprj_io_analog_sel[25]
port 661 nsew signal input
rlabel metal2 s 41713 793897 42193 793953 6 mprj_io_dm[75]
port 662 nsew signal input
rlabel metal2 s 41713 795737 42193 795793 6 mprj_io_dm[76]
port 663 nsew signal input
rlabel metal2 s 41713 789573 42193 789629 6 mprj_io_dm[77]
port 664 nsew signal input
rlabel metal2 s 41713 791413 42193 791469 6 mprj_io_enh[25]
port 665 nsew signal input
rlabel metal2 s 41713 790769 42193 790825 6 mprj_io_hldh_n[25]
port 666 nsew signal input
rlabel metal2 s 41713 788929 42193 788985 6 mprj_io_holdover[25]
port 667 nsew signal input
rlabel metal2 s 41713 785893 42193 785949 6 mprj_io_ib_mode_sel[25]
port 668 nsew signal input
rlabel metal2 s 41713 792701 42193 792757 6 mprj_io_inp_dis[25]
port 669 nsew signal input
rlabel metal2 s 41713 785249 42193 785305 6 mprj_io_oeb[25]
port 670 nsew signal input
rlabel metal2 s 41713 788377 42193 788433 6 mprj_io_out[25]
port 671 nsew signal input
rlabel metal2 s 41713 797577 42193 797633 6 mprj_io_slow_sel[25]
port 672 nsew signal input
rlabel metal2 s 41713 786537 42193 786593 6 mprj_io_vtrip_sel[25]
port 673 nsew signal input
rlabel metal2 s 41713 799417 42193 799473 6 mprj_io_in[25]
port 674 nsew signal tristate
rlabel metal2 s 41713 753733 42193 753789 6 mprj_analog_io[19]
port 675 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 676 nsew signal bidirectional
rlabel metal2 s 41713 751341 42193 751397 6 mprj_io_analog_en[26]
port 677 nsew signal input
rlabel metal2 s 41713 750053 42193 750109 6 mprj_io_analog_pol[26]
port 678 nsew signal input
rlabel metal2 s 41713 747017 42193 747073 6 mprj_io_analog_sel[26]
port 679 nsew signal input
rlabel metal2 s 41713 750697 42193 750753 6 mprj_io_dm[78]
port 680 nsew signal input
rlabel metal2 s 41713 752537 42193 752593 6 mprj_io_dm[79]
port 681 nsew signal input
rlabel metal2 s 41713 746373 42193 746429 6 mprj_io_dm[80]
port 682 nsew signal input
rlabel metal2 s 41713 748213 42193 748269 6 mprj_io_enh[26]
port 683 nsew signal input
rlabel metal2 s 41713 747569 42193 747625 6 mprj_io_hldh_n[26]
port 684 nsew signal input
rlabel metal2 s 41713 745729 42193 745785 6 mprj_io_holdover[26]
port 685 nsew signal input
rlabel metal2 s 41713 742693 42193 742749 6 mprj_io_ib_mode_sel[26]
port 686 nsew signal input
rlabel metal2 s 41713 749501 42193 749557 6 mprj_io_inp_dis[26]
port 687 nsew signal input
rlabel metal2 s 41713 742049 42193 742105 6 mprj_io_oeb[26]
port 688 nsew signal input
rlabel metal2 s 41713 745177 42193 745233 6 mprj_io_out[26]
port 689 nsew signal input
rlabel metal2 s 41713 754377 42193 754433 6 mprj_io_slow_sel[26]
port 690 nsew signal input
rlabel metal2 s 41713 743337 42193 743393 6 mprj_io_vtrip_sel[26]
port 691 nsew signal input
rlabel metal2 s 41713 756217 42193 756273 6 mprj_io_in[26]
port 692 nsew signal tristate
rlabel metal2 s 41713 710533 42193 710589 6 mprj_analog_io[20]
port 693 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 694 nsew signal bidirectional
rlabel metal2 s 41713 708141 42193 708197 6 mprj_io_analog_en[27]
port 695 nsew signal input
rlabel metal2 s 41713 706853 42193 706909 6 mprj_io_analog_pol[27]
port 696 nsew signal input
rlabel metal2 s 41713 703817 42193 703873 6 mprj_io_analog_sel[27]
port 697 nsew signal input
rlabel metal2 s 41713 707497 42193 707553 6 mprj_io_dm[81]
port 698 nsew signal input
rlabel metal2 s 41713 709337 42193 709393 6 mprj_io_dm[82]
port 699 nsew signal input
rlabel metal2 s 41713 703173 42193 703229 6 mprj_io_dm[83]
port 700 nsew signal input
rlabel metal2 s 41713 705013 42193 705069 6 mprj_io_enh[27]
port 701 nsew signal input
rlabel metal2 s 41713 704369 42193 704425 6 mprj_io_hldh_n[27]
port 702 nsew signal input
rlabel metal2 s 41713 702529 42193 702585 6 mprj_io_holdover[27]
port 703 nsew signal input
rlabel metal2 s 41713 699493 42193 699549 6 mprj_io_ib_mode_sel[27]
port 704 nsew signal input
rlabel metal2 s 41713 706301 42193 706357 6 mprj_io_inp_dis[27]
port 705 nsew signal input
rlabel metal2 s 41713 698849 42193 698905 6 mprj_io_oeb[27]
port 706 nsew signal input
rlabel metal2 s 41713 701977 42193 702033 6 mprj_io_out[27]
port 707 nsew signal input
rlabel metal2 s 41713 711177 42193 711233 6 mprj_io_slow_sel[27]
port 708 nsew signal input
rlabel metal2 s 41713 700137 42193 700193 6 mprj_io_vtrip_sel[27]
port 709 nsew signal input
rlabel metal2 s 41713 713017 42193 713073 6 mprj_io_in[27]
port 710 nsew signal tristate
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 711 nsew signal input
rlabel metal5 s 136713 7143 144149 18309 6 resetb
port 712 nsew signal input
rlabel metal3 s 141667 38031 141813 39999 6 resetb_core_h
port 713 nsew signal tristate
rlabel metal5 s 698028 909409 711514 920737 6 vccd1
port 714 nsew signal bidirectional
rlabel metal5 s 698402 819640 710924 832180 6 vdda1
port 715 nsew signal bidirectional
rlabel metal5 s 576820 1018402 589360 1030924 6 vssa1
port 716 nsew signal bidirectional
rlabel metal5 s 698028 461609 711514 472937 6 vssd1
port 717 nsew signal bidirectional
rlabel metal5 s 6086 913863 19572 925191 6 vccd2
port 718 nsew signal bidirectional
rlabel metal5 s 6675 484220 19197 496760 6 vdda2
port 719 nsew signal bidirectional
rlabel metal5 s 6675 828820 19197 841360 6 vssa2
port 720 nsew signal bidirectional
rlabel metal5 s 6086 442663 19572 453991 6 vssd2
port 721 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
