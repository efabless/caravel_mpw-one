magic
tech sky130A
magscale 12 1
timestamp 1598786078
<< metal5 >>
rect 15 90 30 105
rect 10 85 45 90
rect 5 80 45 85
rect 0 75 45 80
rect 0 60 20 75
rect 0 55 35 60
rect 5 50 40 55
rect 10 45 45 50
rect 25 30 45 45
rect 0 25 45 30
rect 0 20 40 25
rect 0 15 35 20
rect 15 0 30 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
