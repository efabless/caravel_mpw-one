.subckt condiode  A C 
.ends
