magic
tech sky130A
magscale 1 2
timestamp 1625094921
<< metal1 >>
rect 181456 1002267 181462 1002319
rect 181514 1002307 181520 1002319
rect 184048 1002307 184054 1002319
rect 181514 1002279 184054 1002307
rect 181514 1002267 181520 1002279
rect 184048 1002267 184054 1002279
rect 184106 1002267 184112 1002319
rect 482608 1002267 482614 1002319
rect 482666 1002307 482672 1002319
rect 483856 1002307 483862 1002319
rect 482666 1002279 483862 1002307
rect 482666 1002267 482672 1002279
rect 483856 1002267 483862 1002279
rect 483914 1002267 483920 1002319
rect 181360 992203 181366 992255
rect 181418 992243 181424 992255
rect 184240 992243 184246 992255
rect 181418 992215 184246 992243
rect 181418 992203 181424 992215
rect 184240 992203 184246 992215
rect 184298 992203 184304 992255
rect 535696 992129 535702 992181
rect 535754 992169 535760 992181
rect 538576 992169 538582 992181
rect 535754 992141 538582 992169
rect 535754 992129 535760 992141
rect 538576 992129 538582 992141
rect 538634 992129 538640 992181
rect 394576 991463 394582 991515
rect 394634 991503 394640 991515
rect 397456 991503 397462 991515
rect 394634 991475 397462 991503
rect 394634 991463 394640 991475
rect 397456 991463 397462 991475
rect 397514 991463 397520 991515
rect 240880 982953 240886 983005
rect 240938 982993 240944 983005
rect 241936 982993 241942 983005
rect 240938 982965 241942 982993
rect 240938 982953 240944 982965
rect 241936 982953 241942 982965
rect 241994 982953 242000 983005
rect 656656 982993 656662 983005
rect 650866 982965 656662 982993
rect 391600 982879 391606 982931
rect 391658 982919 391664 982931
rect 649456 982919 649462 982931
rect 391658 982891 649462 982919
rect 391658 982879 391664 982891
rect 649456 982879 649462 982891
rect 649514 982879 649520 982931
rect 394576 982805 394582 982857
rect 394634 982845 394640 982857
rect 650866 982845 650894 982965
rect 656656 982953 656662 982965
rect 656714 982953 656720 983005
rect 394634 982817 650894 982845
rect 394634 982805 394640 982817
rect 649456 981991 649462 982043
rect 649514 982031 649520 982043
rect 652240 982031 652246 982043
rect 649514 982003 652246 982031
rect 649514 981991 649520 982003
rect 652240 981991 652246 982003
rect 652298 981991 652304 982043
rect 656656 979253 656662 979305
rect 656714 979293 656720 979305
rect 679696 979293 679702 979305
rect 656714 979265 679702 979293
rect 656714 979253 656720 979265
rect 679696 979253 679702 979265
rect 679754 979253 679760 979305
rect 652240 979179 652246 979231
rect 652298 979219 652304 979231
rect 677584 979219 677590 979231
rect 652298 979191 677590 979219
rect 652298 979179 652304 979191
rect 677584 979179 677590 979191
rect 677642 979179 677648 979231
rect 677488 967635 677494 967687
rect 677546 967675 677552 967687
rect 679696 967675 679702 967687
rect 677546 967647 679702 967675
rect 677546 967635 677552 967647
rect 679696 967635 679702 967647
rect 679754 967635 679760 967687
rect 40144 959051 40150 959103
rect 40202 959091 40208 959103
rect 60016 959091 60022 959103
rect 40202 959063 60022 959091
rect 40202 959051 40208 959063
rect 60016 959051 60022 959063
rect 60074 959051 60080 959103
rect 653776 950319 653782 950371
rect 653834 950359 653840 950371
rect 676816 950359 676822 950371
rect 653834 950331 676822 950359
rect 653834 950319 653840 950331
rect 676816 950319 676822 950331
rect 676874 950319 676880 950371
rect 655408 892969 655414 893021
rect 655466 893009 655472 893021
rect 676144 893009 676150 893021
rect 655466 892981 676150 893009
rect 655466 892969 655472 892981
rect 676144 892969 676150 892981
rect 676202 892969 676208 893021
rect 655216 892895 655222 892947
rect 655274 892935 655280 892947
rect 676240 892935 676246 892947
rect 655274 892907 676246 892935
rect 655274 892895 655280 892907
rect 676240 892895 676246 892907
rect 676298 892895 676304 892947
rect 655120 892821 655126 892873
rect 655178 892861 655184 892873
rect 676048 892861 676054 892873
rect 655178 892833 676054 892861
rect 655178 892821 655184 892833
rect 676048 892821 676054 892833
rect 676106 892821 676112 892873
rect 673360 892377 673366 892429
rect 673418 892417 673424 892429
rect 676048 892417 676054 892429
rect 673418 892389 676054 892417
rect 673418 892377 673424 892389
rect 676048 892377 676054 892389
rect 676106 892377 676112 892429
rect 670960 891415 670966 891467
rect 671018 891455 671024 891467
rect 676048 891455 676054 891467
rect 671018 891427 676054 891455
rect 671018 891415 671024 891427
rect 676048 891415 676054 891427
rect 676106 891415 676112 891467
rect 670864 890379 670870 890431
rect 670922 890419 670928 890431
rect 676048 890419 676054 890431
rect 670922 890391 676054 890419
rect 670922 890379 670928 890391
rect 676048 890379 676054 890391
rect 676106 890379 676112 890431
rect 673936 887863 673942 887915
rect 673994 887903 674000 887915
rect 676240 887903 676246 887915
rect 673994 887875 676246 887903
rect 673994 887863 674000 887875
rect 676240 887863 676246 887875
rect 676298 887863 676304 887915
rect 674128 887123 674134 887175
rect 674186 887163 674192 887175
rect 676048 887163 676054 887175
rect 674186 887135 676054 887163
rect 674186 887123 674192 887135
rect 676048 887123 676054 887135
rect 676106 887123 676112 887175
rect 674224 887049 674230 887101
rect 674282 887089 674288 887101
rect 676240 887089 676246 887101
rect 674282 887061 676246 887089
rect 674282 887049 674288 887061
rect 676240 887049 676246 887061
rect 676298 887049 676304 887101
rect 674032 885051 674038 885103
rect 674090 885091 674096 885103
rect 676048 885091 676054 885103
rect 674090 885063 676054 885091
rect 674090 885051 674096 885063
rect 676048 885051 676054 885063
rect 676106 885051 676112 885103
rect 674512 884237 674518 884289
rect 674570 884277 674576 884289
rect 676048 884277 676054 884289
rect 674570 884249 676054 884277
rect 674570 884237 674576 884249
rect 676048 884237 676054 884249
rect 676106 884237 676112 884289
rect 674416 883571 674422 883623
rect 674474 883611 674480 883623
rect 676048 883611 676054 883623
rect 674474 883583 676054 883611
rect 674474 883571 674480 883583
rect 676048 883571 676054 883583
rect 676106 883571 676112 883623
rect 675280 883201 675286 883253
rect 675338 883241 675344 883253
rect 679984 883241 679990 883253
rect 675338 883213 679990 883241
rect 675338 883201 675344 883213
rect 679984 883201 679990 883213
rect 680042 883201 680048 883253
rect 675088 883127 675094 883179
rect 675146 883167 675152 883179
rect 680176 883167 680182 883179
rect 675146 883139 680182 883167
rect 675146 883127 675152 883139
rect 680176 883127 680182 883139
rect 680234 883127 680240 883179
rect 674992 883053 674998 883105
rect 675050 883093 675056 883105
rect 676048 883093 676054 883105
rect 675050 883065 676054 883093
rect 675050 883053 675056 883065
rect 676048 883053 676054 883065
rect 676106 883053 676112 883105
rect 674992 882831 674998 882883
rect 675050 882871 675056 882883
rect 679696 882871 679702 882883
rect 675050 882843 679702 882871
rect 675050 882831 675056 882843
rect 679696 882831 679702 882843
rect 679754 882831 679760 882883
rect 649456 881425 649462 881477
rect 649514 881465 649520 881477
rect 679696 881465 679702 881477
rect 649514 881437 679702 881465
rect 649514 881425 649520 881437
rect 679696 881425 679702 881437
rect 679754 881425 679760 881477
rect 655312 881351 655318 881403
rect 655370 881391 655376 881403
rect 675472 881391 675478 881403
rect 655370 881363 675478 881391
rect 655370 881351 655376 881363
rect 675472 881351 675478 881363
rect 675530 881351 675536 881403
rect 674320 881203 674326 881255
rect 674378 881243 674384 881255
rect 680080 881243 680086 881255
rect 674378 881215 680086 881243
rect 674378 881203 674384 881215
rect 680080 881203 680086 881215
rect 680138 881203 680144 881255
rect 674608 880093 674614 880145
rect 674666 880133 674672 880145
rect 679792 880133 679798 880145
rect 674666 880105 679798 880133
rect 674666 880093 674672 880105
rect 679792 880093 679798 880105
rect 679850 880093 679856 880145
rect 675184 879501 675190 879553
rect 675242 879541 675248 879553
rect 679888 879541 679894 879553
rect 675242 879513 679894 879541
rect 675242 879501 675248 879513
rect 679888 879501 679894 879513
rect 679946 879501 679952 879553
rect 674896 878317 674902 878369
rect 674954 878357 674960 878369
rect 675760 878357 675766 878369
rect 674954 878329 675766 878357
rect 674954 878317 674960 878329
rect 675760 878317 675766 878329
rect 675818 878317 675824 878369
rect 674992 877207 674998 877259
rect 675050 877247 675056 877259
rect 675472 877247 675478 877259
rect 675050 877219 675478 877247
rect 675050 877207 675056 877219
rect 675472 877207 675478 877219
rect 675530 877207 675536 877259
rect 675184 876615 675190 876667
rect 675242 876615 675248 876667
rect 675202 876223 675230 876615
rect 675184 876171 675190 876223
rect 675242 876171 675248 876223
rect 674224 876097 674230 876149
rect 674282 876137 674288 876149
rect 675088 876137 675094 876149
rect 674282 876109 675094 876137
rect 674282 876097 674288 876109
rect 675088 876097 675094 876109
rect 675146 876097 675152 876149
rect 674512 875431 674518 875483
rect 674570 875471 674576 875483
rect 674992 875471 674998 875483
rect 674570 875443 674998 875471
rect 674570 875431 674576 875443
rect 674992 875431 674998 875443
rect 675050 875431 675056 875483
rect 673936 875209 673942 875261
rect 673994 875249 674000 875261
rect 674416 875249 674422 875261
rect 673994 875221 674422 875249
rect 673994 875209 674000 875221
rect 674416 875209 674422 875221
rect 674474 875209 674480 875261
rect 674320 874913 674326 874965
rect 674378 874953 674384 874965
rect 675472 874953 675478 874965
rect 674378 874925 675478 874953
rect 674378 874913 674384 874925
rect 675472 874913 675478 874925
rect 675530 874913 675536 874965
rect 674608 874247 674614 874299
rect 674666 874287 674672 874299
rect 675472 874287 675478 874299
rect 674666 874259 675478 874287
rect 674666 874247 674672 874259
rect 675472 874247 675478 874259
rect 675530 874247 675536 874299
rect 675184 873507 675190 873559
rect 675242 873547 675248 873559
rect 675376 873547 675382 873559
rect 675242 873519 675382 873547
rect 675242 873507 675248 873519
rect 675376 873507 675382 873519
rect 675434 873507 675440 873559
rect 674896 872915 674902 872967
rect 674954 872955 674960 872967
rect 675376 872955 675382 872967
rect 674954 872927 675382 872955
rect 674954 872915 674960 872927
rect 675376 872915 675382 872927
rect 675434 872915 675440 872967
rect 654160 872619 654166 872671
rect 654218 872659 654224 872671
rect 674608 872659 674614 872671
rect 654218 872631 674614 872659
rect 654218 872619 654224 872631
rect 674608 872619 674614 872631
rect 674666 872619 674672 872671
rect 674512 869807 674518 869859
rect 674570 869847 674576 869859
rect 675376 869847 675382 869859
rect 674570 869819 675382 869847
rect 674570 869807 674576 869819
rect 675376 869807 675382 869819
rect 675434 869807 675440 869859
rect 674128 868105 674134 868157
rect 674186 868145 674192 868157
rect 674992 868145 674998 868157
rect 674186 868117 674998 868145
rect 674186 868105 674192 868117
rect 674992 868105 674998 868117
rect 675050 868105 675056 868157
rect 674608 868031 674614 868083
rect 674666 868071 674672 868083
rect 675088 868071 675094 868083
rect 674666 868043 675094 868071
rect 674666 868031 674672 868043
rect 675088 868031 675094 868043
rect 675146 868031 675152 868083
rect 674032 867365 674038 867417
rect 674090 867405 674096 867417
rect 675472 867405 675478 867417
rect 674090 867377 675478 867405
rect 674090 867365 674096 867377
rect 675472 867365 675478 867377
rect 675530 867365 675536 867417
rect 674416 865737 674422 865789
rect 674474 865777 674480 865789
rect 675184 865777 675190 865789
rect 674474 865749 675190 865777
rect 674474 865737 674480 865749
rect 675184 865737 675190 865749
rect 675242 865737 675248 865789
rect 653776 863961 653782 864013
rect 653834 864001 653840 864013
rect 675088 864001 675094 864013
rect 653834 863973 675094 864001
rect 653834 863961 653840 863973
rect 675088 863961 675094 863973
rect 675146 863961 675152 864013
rect 41776 817933 41782 817985
rect 41834 817973 41840 817985
rect 47440 817973 47446 817985
rect 41834 817945 47446 817973
rect 41834 817933 41840 817945
rect 47440 817933 47446 817945
rect 47498 817933 47504 817985
rect 41776 817267 41782 817319
rect 41834 817307 41840 817319
rect 44848 817307 44854 817319
rect 41834 817279 44854 817307
rect 41834 817267 41840 817279
rect 44848 817267 44854 817279
rect 44906 817267 44912 817319
rect 41584 816527 41590 816579
rect 41642 816567 41648 816579
rect 44944 816567 44950 816579
rect 41642 816539 44950 816567
rect 41642 816527 41648 816539
rect 44944 816527 44950 816539
rect 45002 816527 45008 816579
rect 41776 815787 41782 815839
rect 41834 815827 41840 815839
rect 43216 815827 43222 815839
rect 41834 815799 43222 815827
rect 41834 815787 41840 815799
rect 43216 815787 43222 815799
rect 43274 815787 43280 815839
rect 41776 814825 41782 814877
rect 41834 814865 41840 814877
rect 44656 814865 44662 814877
rect 41834 814837 44662 814865
rect 41834 814825 41840 814837
rect 44656 814825 44662 814837
rect 44714 814825 44720 814877
rect 41584 813567 41590 813619
rect 41642 813607 41648 813619
rect 44752 813607 44758 813619
rect 41642 813579 44758 813607
rect 41642 813567 41648 813579
rect 44752 813567 44758 813579
rect 44810 813567 44816 813619
rect 41584 812383 41590 812435
rect 41642 812423 41648 812435
rect 42928 812423 42934 812435
rect 41642 812395 42934 812423
rect 41642 812383 41648 812395
rect 42928 812383 42934 812395
rect 42986 812383 42992 812435
rect 41584 809867 41590 809919
rect 41642 809907 41648 809919
rect 42832 809907 42838 809919
rect 41642 809879 42838 809907
rect 41642 809867 41648 809879
rect 42832 809867 42838 809879
rect 42890 809867 42896 809919
rect 41776 809793 41782 809845
rect 41834 809833 41840 809845
rect 42736 809833 42742 809845
rect 41834 809805 42742 809833
rect 41834 809793 41840 809805
rect 42736 809793 42742 809805
rect 42794 809793 42800 809845
rect 41776 808609 41782 808661
rect 41834 808649 41840 808661
rect 43120 808649 43126 808661
rect 41834 808621 43126 808649
rect 41834 808609 41840 808621
rect 43120 808609 43126 808621
rect 43178 808609 43184 808661
rect 41776 807351 41782 807403
rect 41834 807391 41840 807403
rect 42640 807391 42646 807403
rect 41834 807363 42646 807391
rect 41834 807351 41840 807363
rect 42640 807351 42646 807363
rect 42698 807351 42704 807403
rect 41584 806611 41590 806663
rect 41642 806651 41648 806663
rect 43024 806651 43030 806663
rect 41642 806623 43030 806651
rect 41642 806611 41648 806623
rect 43024 806611 43030 806623
rect 43082 806611 43088 806663
rect 41584 805131 41590 805183
rect 41642 805171 41648 805183
rect 44560 805171 44566 805183
rect 41642 805143 44566 805171
rect 41642 805131 41648 805143
rect 44560 805131 44566 805143
rect 44618 805131 44624 805183
rect 42832 800765 42838 800817
rect 42890 800805 42896 800817
rect 43504 800805 43510 800817
rect 42890 800777 43510 800805
rect 42890 800765 42896 800777
rect 43504 800765 43510 800777
rect 43562 800765 43568 800817
rect 42736 800691 42742 800743
rect 42794 800731 42800 800743
rect 57712 800731 57718 800743
rect 42794 800703 57718 800731
rect 42794 800691 42800 800703
rect 57712 800691 57718 800703
rect 57770 800691 57776 800743
rect 42832 800617 42838 800669
rect 42890 800657 42896 800669
rect 57616 800657 57622 800669
rect 42890 800629 57622 800657
rect 42890 800617 42896 800629
rect 57616 800617 57622 800629
rect 57674 800617 57680 800669
rect 41872 800173 41878 800225
rect 41930 800173 41936 800225
rect 42160 800173 42166 800225
rect 42218 800213 42224 800225
rect 43312 800213 43318 800225
rect 42218 800185 43318 800213
rect 42218 800173 42224 800185
rect 43312 800173 43318 800185
rect 43370 800173 43376 800225
rect 41890 800003 41918 800173
rect 41872 799951 41878 800003
rect 41930 799951 41936 800003
rect 42160 798101 42166 798153
rect 42218 798141 42224 798153
rect 42544 798141 42550 798153
rect 42218 798113 42550 798141
rect 42218 798101 42224 798113
rect 42544 798101 42550 798113
rect 42602 798101 42608 798153
rect 42640 797879 42646 797931
rect 42698 797919 42704 797931
rect 42698 797891 42878 797919
rect 42698 797879 42704 797891
rect 42064 797287 42070 797339
rect 42122 797327 42128 797339
rect 42736 797327 42742 797339
rect 42122 797299 42742 797327
rect 42122 797287 42128 797299
rect 42736 797287 42742 797299
rect 42794 797287 42800 797339
rect 42850 797253 42878 797891
rect 42754 797225 42878 797253
rect 42754 796895 42782 797225
rect 42736 796843 42742 796895
rect 42794 796843 42800 796895
rect 42160 796251 42166 796303
rect 42218 796291 42224 796303
rect 43120 796291 43126 796303
rect 42218 796263 43126 796291
rect 42218 796251 42224 796263
rect 43120 796251 43126 796263
rect 43178 796251 43184 796303
rect 43216 796251 43222 796303
rect 43274 796251 43280 796303
rect 43234 796081 43262 796251
rect 43216 796029 43222 796081
rect 43274 796029 43280 796081
rect 42064 795585 42070 795637
rect 42122 795625 42128 795637
rect 42832 795625 42838 795637
rect 42122 795597 42838 795625
rect 42122 795585 42128 795597
rect 42832 795585 42838 795597
rect 42890 795585 42896 795637
rect 42160 794771 42166 794823
rect 42218 794811 42224 794823
rect 43024 794811 43030 794823
rect 42218 794783 43030 794811
rect 42218 794771 42224 794783
rect 43024 794771 43030 794783
rect 43082 794771 43088 794823
rect 43024 794623 43030 794675
rect 43082 794663 43088 794675
rect 43504 794663 43510 794675
rect 43082 794635 43510 794663
rect 43082 794623 43088 794635
rect 43504 794623 43510 794635
rect 43562 794623 43568 794675
rect 42160 793587 42166 793639
rect 42218 793627 42224 793639
rect 42736 793627 42742 793639
rect 42218 793599 42742 793627
rect 42218 793587 42224 793599
rect 42736 793587 42742 793599
rect 42794 793587 42800 793639
rect 42928 792107 42934 792159
rect 42986 792147 42992 792159
rect 43504 792147 43510 792159
rect 42986 792119 43510 792147
rect 42986 792107 42992 792119
rect 43504 792107 43510 792119
rect 43562 792107 43568 792159
rect 655120 792033 655126 792085
rect 655178 792073 655184 792085
rect 675376 792073 675382 792085
rect 655178 792045 675382 792073
rect 655178 792033 655184 792045
rect 675376 792033 675382 792045
rect 675434 792033 675440 792085
rect 42160 790627 42166 790679
rect 42218 790667 42224 790679
rect 43120 790667 43126 790679
rect 42218 790639 43126 790667
rect 42218 790627 42224 790639
rect 43120 790627 43126 790639
rect 43178 790627 43184 790679
rect 43120 790479 43126 790531
rect 43178 790519 43184 790531
rect 43504 790519 43510 790531
rect 43178 790491 43510 790519
rect 43178 790479 43184 790491
rect 43504 790479 43510 790491
rect 43562 790479 43568 790531
rect 42160 789443 42166 789495
rect 42218 789483 42224 789495
rect 42736 789483 42742 789495
rect 42218 789455 42742 789483
rect 42218 789443 42224 789455
rect 42736 789443 42742 789455
rect 42794 789443 42800 789495
rect 42928 789147 42934 789199
rect 42986 789187 42992 789199
rect 58192 789187 58198 789199
rect 42986 789159 58198 789187
rect 42986 789147 42992 789159
rect 58192 789147 58198 789159
rect 58250 789147 58256 789199
rect 44944 789073 44950 789125
rect 45002 789113 45008 789125
rect 58384 789113 58390 789125
rect 45002 789085 58390 789113
rect 45002 789073 45008 789085
rect 58384 789073 58390 789085
rect 58442 789073 58448 789125
rect 42160 788703 42166 788755
rect 42218 788743 42224 788755
rect 43024 788743 43030 788755
rect 42218 788715 43030 788743
rect 42218 788703 42224 788715
rect 43024 788703 43030 788715
rect 43082 788703 43088 788755
rect 42160 786853 42166 786905
rect 42218 786893 42224 786905
rect 43120 786893 43126 786905
rect 42218 786865 43126 786893
rect 42218 786853 42224 786865
rect 43120 786853 43126 786865
rect 43178 786853 43184 786905
rect 42160 786409 42166 786461
rect 42218 786449 42224 786461
rect 42736 786449 42742 786461
rect 42218 786421 42742 786449
rect 42218 786409 42224 786421
rect 42736 786409 42742 786421
rect 42794 786409 42800 786461
rect 42064 785595 42070 785647
rect 42122 785635 42128 785647
rect 42832 785635 42838 785647
rect 42122 785607 42838 785635
rect 42122 785595 42128 785607
rect 42832 785595 42838 785607
rect 42890 785595 42896 785647
rect 44848 785521 44854 785573
rect 44906 785561 44912 785573
rect 59152 785561 59158 785573
rect 44906 785533 59158 785561
rect 44906 785521 44912 785533
rect 59152 785521 59158 785533
rect 59210 785521 59216 785573
rect 47440 785373 47446 785425
rect 47498 785413 47504 785425
rect 59632 785413 59638 785425
rect 47498 785385 59638 785413
rect 47498 785373 47504 785385
rect 59632 785373 59638 785385
rect 59690 785373 59696 785425
rect 42160 785003 42166 785055
rect 42218 785043 42224 785055
rect 42928 785043 42934 785055
rect 42218 785015 42934 785043
rect 42218 785003 42224 785015
rect 42928 785003 42934 785015
rect 42986 785003 42992 785055
rect 656560 783449 656566 783501
rect 656618 783489 656624 783501
rect 674992 783489 674998 783501
rect 656618 783461 674998 783489
rect 656618 783449 656624 783461
rect 674992 783449 674998 783461
rect 675050 783449 675056 783501
rect 654352 780489 654358 780541
rect 654410 780529 654416 780541
rect 675280 780529 675286 780541
rect 654410 780501 675286 780529
rect 654410 780489 654416 780501
rect 675280 780489 675286 780501
rect 675338 780489 675344 780541
rect 674992 778861 674998 778913
rect 675050 778901 675056 778913
rect 675376 778901 675382 778913
rect 675050 778873 675382 778901
rect 675050 778861 675056 778873
rect 675376 778861 675382 778873
rect 675434 778861 675440 778913
rect 673072 778713 673078 778765
rect 673130 778753 673136 778765
rect 675472 778753 675478 778765
rect 673130 778725 675478 778753
rect 673130 778713 673136 778725
rect 675472 778713 675478 778725
rect 675530 778713 675536 778765
rect 41776 774643 41782 774695
rect 41834 774683 41840 774695
rect 47536 774683 47542 774695
rect 41834 774655 47542 774683
rect 41834 774643 41840 774655
rect 47536 774643 47542 774655
rect 47594 774643 47600 774695
rect 41584 773903 41590 773955
rect 41642 773943 41648 773955
rect 44848 773943 44854 773955
rect 41642 773915 44854 773943
rect 41642 773903 41648 773915
rect 44848 773903 44854 773915
rect 44906 773903 44912 773955
rect 674512 773607 674518 773659
rect 674570 773647 674576 773659
rect 675280 773647 675286 773659
rect 674570 773619 675286 773647
rect 674570 773607 674576 773619
rect 675280 773607 675286 773619
rect 675338 773607 675344 773659
rect 41584 773311 41590 773363
rect 41642 773351 41648 773363
rect 44944 773351 44950 773363
rect 41642 773323 44950 773351
rect 41642 773311 41648 773323
rect 44944 773311 44950 773323
rect 45002 773311 45008 773363
rect 41776 773237 41782 773289
rect 41834 773277 41840 773289
rect 43408 773277 43414 773289
rect 41834 773249 43414 773277
rect 41834 773237 41840 773249
rect 43408 773237 43414 773249
rect 43466 773237 43472 773289
rect 41776 772571 41782 772623
rect 41834 772611 41840 772623
rect 43312 772611 43318 772623
rect 41834 772583 43318 772611
rect 41834 772571 41840 772583
rect 43312 772571 43318 772583
rect 43370 772571 43376 772623
rect 42736 771905 42742 771957
rect 42794 771945 42800 771957
rect 62032 771945 62038 771957
rect 42794 771917 62038 771945
rect 42794 771905 42800 771917
rect 62032 771905 62038 771917
rect 62090 771905 62096 771957
rect 41584 771831 41590 771883
rect 41642 771871 41648 771883
rect 61840 771871 61846 771883
rect 41642 771843 61846 771871
rect 41642 771831 41648 771843
rect 61840 771831 61846 771843
rect 61898 771831 61904 771883
rect 41776 768131 41782 768183
rect 41834 768171 41840 768183
rect 42832 768171 42838 768183
rect 41834 768143 42838 768171
rect 41834 768131 41840 768143
rect 42832 768131 42838 768143
rect 42890 768131 42896 768183
rect 41776 765097 41782 765149
rect 41834 765137 41840 765149
rect 42928 765137 42934 765149
rect 41834 765109 42934 765137
rect 41834 765097 41840 765109
rect 42928 765097 42934 765109
rect 42986 765097 42992 765149
rect 41776 764135 41782 764187
rect 41834 764175 41840 764187
rect 43024 764175 43030 764187
rect 41834 764147 43030 764175
rect 41834 764135 41840 764147
rect 43024 764135 43030 764147
rect 43082 764135 43088 764187
rect 41584 763395 41590 763447
rect 41642 763435 41648 763447
rect 43120 763435 43126 763447
rect 41642 763407 43126 763435
rect 41642 763395 41648 763407
rect 43120 763395 43126 763407
rect 43178 763395 43184 763447
rect 41776 762063 41782 762115
rect 41834 762103 41840 762115
rect 47440 762103 47446 762115
rect 41834 762075 47446 762103
rect 41834 762063 41840 762075
rect 47440 762063 47446 762075
rect 47498 762063 47504 762115
rect 42928 757623 42934 757675
rect 42986 757663 42992 757675
rect 43216 757663 43222 757675
rect 42986 757635 43222 757663
rect 42986 757623 42992 757635
rect 43216 757623 43222 757635
rect 43274 757623 43280 757675
rect 42928 757475 42934 757527
rect 42986 757515 42992 757527
rect 58672 757515 58678 757527
rect 42986 757487 58678 757515
rect 42986 757475 42992 757487
rect 58672 757475 58678 757487
rect 58730 757475 58736 757527
rect 41392 757327 41398 757379
rect 41450 757367 41456 757379
rect 43600 757367 43606 757379
rect 41450 757339 43606 757367
rect 41450 757327 41456 757339
rect 43600 757327 43606 757339
rect 43658 757327 43664 757379
rect 41488 757253 41494 757305
rect 41546 757293 41552 757305
rect 43504 757293 43510 757305
rect 41546 757265 43510 757293
rect 41546 757253 41552 757265
rect 43504 757253 43510 757265
rect 43562 757253 43568 757305
rect 41872 756957 41878 757009
rect 41930 756957 41936 757009
rect 41890 756787 41918 756957
rect 41872 756735 41878 756787
rect 41930 756735 41936 756787
rect 42160 754219 42166 754271
rect 42218 754259 42224 754271
rect 42928 754259 42934 754271
rect 42218 754231 42934 754259
rect 42218 754219 42224 754231
rect 42928 754219 42934 754231
rect 42986 754219 42992 754271
rect 42064 753035 42070 753087
rect 42122 753075 42128 753087
rect 42352 753075 42358 753087
rect 42122 753047 42358 753075
rect 42122 753035 42128 753047
rect 42352 753035 42358 753047
rect 42410 753035 42416 753087
rect 42352 752887 42358 752939
rect 42410 752927 42416 752939
rect 43024 752927 43030 752939
rect 42410 752899 43030 752927
rect 42410 752887 42416 752899
rect 43024 752887 43030 752899
rect 43082 752887 43088 752939
rect 42064 751777 42070 751829
rect 42122 751817 42128 751829
rect 43216 751817 43222 751829
rect 42122 751789 43222 751817
rect 42122 751777 42128 751789
rect 43216 751777 43222 751789
rect 43274 751777 43280 751829
rect 42064 751481 42070 751533
rect 42122 751521 42128 751533
rect 42928 751521 42934 751533
rect 42122 751493 42934 751521
rect 42122 751481 42128 751493
rect 42928 751481 42934 751493
rect 42986 751481 42992 751533
rect 42064 751111 42070 751163
rect 42122 751151 42128 751163
rect 43120 751151 43126 751163
rect 42122 751123 43126 751151
rect 42122 751111 42128 751123
rect 43120 751111 43126 751123
rect 43178 751111 43184 751163
rect 43120 750963 43126 751015
rect 43178 751003 43184 751015
rect 43504 751003 43510 751015
rect 43178 750975 43510 751003
rect 43178 750963 43184 750975
rect 43504 750963 43510 750975
rect 43562 750963 43568 751015
rect 42160 750593 42166 750645
rect 42218 750633 42224 750645
rect 42352 750633 42358 750645
rect 42218 750605 42358 750633
rect 42218 750593 42224 750605
rect 42352 750593 42358 750605
rect 42410 750593 42416 750645
rect 42064 749779 42070 749831
rect 42122 749819 42128 749831
rect 42928 749819 42934 749831
rect 42122 749791 42934 749819
rect 42122 749779 42128 749791
rect 42928 749779 42934 749791
rect 42986 749779 42992 749831
rect 42928 749631 42934 749683
rect 42986 749671 42992 749683
rect 43600 749671 43606 749683
rect 42986 749643 43606 749671
rect 42986 749631 42992 749643
rect 43600 749631 43606 749643
rect 43658 749631 43664 749683
rect 655696 748817 655702 748869
rect 655754 748857 655760 748869
rect 675376 748857 675382 748869
rect 655754 748829 675382 748857
rect 655754 748817 655760 748829
rect 675376 748817 675382 748829
rect 675434 748817 675440 748869
rect 42064 746079 42070 746131
rect 42122 746119 42128 746131
rect 43120 746119 43126 746131
rect 42122 746091 43126 746119
rect 42122 746079 42128 746091
rect 43120 746079 43126 746091
rect 43178 746079 43184 746131
rect 43120 745931 43126 745983
rect 43178 745971 43184 745983
rect 54640 745971 54646 745983
rect 43178 745943 54646 745971
rect 43178 745931 43184 745943
rect 54640 745931 54646 745943
rect 54698 745931 54704 745983
rect 54736 745931 54742 745983
rect 54794 745971 54800 745983
rect 57616 745971 57622 745983
rect 54794 745943 57622 745971
rect 54794 745931 54800 745943
rect 57616 745931 57622 745943
rect 57674 745931 57680 745983
rect 42160 745487 42166 745539
rect 42218 745527 42224 745539
rect 42448 745527 42454 745539
rect 42218 745499 42454 745527
rect 42218 745487 42224 745499
rect 42448 745487 42454 745499
rect 42506 745487 42512 745539
rect 43216 745265 43222 745317
rect 43274 745305 43280 745317
rect 59632 745305 59638 745317
rect 43274 745277 59638 745305
rect 43274 745265 43280 745277
rect 59632 745265 59638 745277
rect 59690 745265 59696 745317
rect 44944 745117 44950 745169
rect 45002 745157 45008 745169
rect 58192 745157 58198 745169
rect 45002 745129 58198 745157
rect 45002 745117 45008 745129
rect 58192 745117 58198 745129
rect 58250 745117 58256 745169
rect 42160 743563 42166 743615
rect 42218 743603 42224 743615
rect 43024 743603 43030 743615
rect 42218 743575 43030 743603
rect 42218 743563 42224 743575
rect 43024 743563 43030 743575
rect 43082 743563 43088 743615
rect 42064 743193 42070 743245
rect 42122 743233 42128 743245
rect 42928 743233 42934 743245
rect 42122 743205 42934 743233
rect 42122 743193 42128 743205
rect 42928 743193 42934 743205
rect 42986 743193 42992 743245
rect 47536 742971 47542 743023
rect 47594 743011 47600 743023
rect 59632 743011 59638 743023
rect 47594 742983 59638 743011
rect 47594 742971 47600 742983
rect 59632 742971 59638 742983
rect 59690 742971 59696 743023
rect 44848 742897 44854 742949
rect 44906 742937 44912 742949
rect 59728 742937 59734 742949
rect 44906 742909 59734 742937
rect 44906 742897 44912 742909
rect 59728 742897 59734 742909
rect 59786 742897 59792 742949
rect 42160 742601 42166 742653
rect 42218 742641 42224 742653
rect 42448 742641 42454 742653
rect 42218 742613 42454 742641
rect 42218 742601 42224 742613
rect 42448 742601 42454 742613
rect 42506 742601 42512 742653
rect 674416 742083 674422 742135
rect 674474 742123 674480 742135
rect 675184 742123 675190 742135
rect 674474 742095 675190 742123
rect 674474 742083 674480 742095
rect 675184 742083 675190 742095
rect 675242 742083 675248 742135
rect 42160 741935 42166 741987
rect 42218 741975 42224 741987
rect 43120 741975 43126 741987
rect 42218 741947 43126 741975
rect 42218 741935 42224 741947
rect 43120 741935 43126 741947
rect 43178 741935 43184 741987
rect 673168 738235 673174 738287
rect 673226 738275 673232 738287
rect 675376 738275 675382 738287
rect 673226 738247 675382 738275
rect 673226 738235 673232 738247
rect 675376 738235 675382 738247
rect 675434 738235 675440 738287
rect 672112 737569 672118 737621
rect 672170 737609 672176 737621
rect 675280 737609 675286 737621
rect 672170 737581 675286 737609
rect 672170 737569 672176 737581
rect 675280 737569 675286 737581
rect 675338 737569 675344 737621
rect 654064 737421 654070 737473
rect 654122 737461 654128 737473
rect 675280 737461 675286 737473
rect 654122 737433 675286 737461
rect 654122 737421 654128 737433
rect 675280 737421 675286 737433
rect 675338 737421 675344 737473
rect 654160 737347 654166 737399
rect 654218 737387 654224 737399
rect 674608 737387 674614 737399
rect 654218 737359 674614 737387
rect 654218 737347 654224 737359
rect 674608 737347 674614 737359
rect 674666 737347 674672 737399
rect 672880 734757 672886 734809
rect 672938 734797 672944 734809
rect 675376 734797 675382 734809
rect 672938 734769 675382 734797
rect 672938 734757 672944 734769
rect 675376 734757 675382 734769
rect 675434 734757 675440 734809
rect 672304 734387 672310 734439
rect 672362 734427 672368 734439
rect 675376 734427 675382 734439
rect 672362 734399 675382 734427
rect 672362 734387 672368 734399
rect 675376 734387 675382 734399
rect 675434 734387 675440 734439
rect 672400 734165 672406 734217
rect 672458 734205 672464 734217
rect 675376 734205 675382 734217
rect 672458 734177 675382 734205
rect 672458 734165 672464 734177
rect 675376 734165 675382 734177
rect 675434 734165 675440 734217
rect 675184 733869 675190 733921
rect 675242 733909 675248 733921
rect 675472 733909 675478 733921
rect 675242 733881 675478 733909
rect 675242 733869 675248 733881
rect 675472 733869 675478 733881
rect 675530 733869 675536 733921
rect 672784 732315 672790 732367
rect 672842 732355 672848 732367
rect 675472 732355 675478 732367
rect 672842 732327 675478 732355
rect 672842 732315 672848 732327
rect 675472 732315 675478 732327
rect 675530 732315 675536 732367
rect 674608 732019 674614 732071
rect 674666 732059 674672 732071
rect 675376 732059 675382 732071
rect 674666 732031 675382 732059
rect 674666 732019 674672 732031
rect 675376 732019 675382 732031
rect 675434 732019 675440 732071
rect 41776 731427 41782 731479
rect 41834 731467 41840 731479
rect 47632 731467 47638 731479
rect 41834 731439 47638 731467
rect 41834 731427 41840 731439
rect 47632 731427 47638 731439
rect 47690 731427 47696 731479
rect 41584 730687 41590 730739
rect 41642 730727 41648 730739
rect 44848 730727 44854 730739
rect 41642 730699 44854 730727
rect 41642 730687 41648 730699
rect 44848 730687 44854 730699
rect 44906 730687 44912 730739
rect 674416 730465 674422 730517
rect 674474 730505 674480 730517
rect 675472 730505 675478 730517
rect 674474 730477 675478 730505
rect 674474 730465 674480 730477
rect 675472 730465 675478 730477
rect 675530 730465 675536 730517
rect 41776 730317 41782 730369
rect 41834 730357 41840 730369
rect 44944 730357 44950 730369
rect 41834 730329 44950 730357
rect 41834 730317 41840 730329
rect 44944 730317 44950 730329
rect 45002 730317 45008 730369
rect 41584 730169 41590 730221
rect 41642 730209 41648 730221
rect 43312 730209 43318 730221
rect 41642 730181 43318 730209
rect 41642 730169 41648 730181
rect 43312 730169 43318 730181
rect 43370 730169 43376 730221
rect 41584 729207 41590 729259
rect 41642 729247 41648 729259
rect 43888 729247 43894 729259
rect 41642 729219 43894 729247
rect 41642 729207 41648 729219
rect 43888 729207 43894 729219
rect 43946 729207 43952 729259
rect 41776 728763 41782 728815
rect 41834 728803 41840 728815
rect 43792 728803 43798 728815
rect 41834 728775 43798 728803
rect 41834 728763 41840 728775
rect 43792 728763 43798 728775
rect 43850 728763 43856 728815
rect 40432 728689 40438 728741
rect 40490 728729 40496 728741
rect 62224 728729 62230 728741
rect 40490 728701 62230 728729
rect 40490 728689 40496 728701
rect 62224 728689 62230 728701
rect 62282 728689 62288 728741
rect 41392 728615 41398 728667
rect 41450 728655 41456 728667
rect 62416 728655 62422 728667
rect 41450 728627 62422 728655
rect 41450 728615 41456 728627
rect 62416 728615 62422 728627
rect 62474 728615 62480 728667
rect 674224 728615 674230 728667
rect 674282 728655 674288 728667
rect 675472 728655 675478 728667
rect 674282 728627 675478 728655
rect 674282 728615 674288 728627
rect 675472 728615 675478 728627
rect 675530 728615 675536 728667
rect 41776 727875 41782 727927
rect 41834 727915 41840 727927
rect 43696 727915 43702 727927
rect 41834 727887 43702 727915
rect 41834 727875 41840 727887
rect 43696 727875 43702 727887
rect 43754 727875 43760 727927
rect 41872 722917 41878 722969
rect 41930 722957 41936 722969
rect 42928 722957 42934 722969
rect 41930 722929 42934 722957
rect 41930 722917 41936 722929
rect 42928 722917 42934 722929
rect 42986 722917 42992 722969
rect 41584 720401 41590 720453
rect 41642 720441 41648 720453
rect 43024 720441 43030 720453
rect 41642 720413 43030 720441
rect 41642 720401 41648 720413
rect 43024 720401 43030 720413
rect 43082 720401 43088 720453
rect 41584 720179 41590 720231
rect 41642 720219 41648 720231
rect 43120 720219 43126 720231
rect 41642 720191 43126 720219
rect 41642 720179 41648 720191
rect 43120 720179 43126 720191
rect 43178 720179 43184 720231
rect 41584 718699 41590 718751
rect 41642 718739 41648 718751
rect 47536 718739 47542 718751
rect 41642 718711 47542 718739
rect 41642 718699 41648 718711
rect 47536 718699 47542 718711
rect 47594 718699 47600 718751
rect 655600 714703 655606 714755
rect 655658 714743 655664 714755
rect 676240 714743 676246 714755
rect 655658 714715 676246 714743
rect 655658 714703 655664 714715
rect 676240 714703 676246 714715
rect 676298 714703 676304 714755
rect 655408 714555 655414 714607
rect 655466 714595 655472 714607
rect 676336 714595 676342 714607
rect 655466 714567 676342 714595
rect 655466 714555 655472 714567
rect 676336 714555 676342 714567
rect 676394 714555 676400 714607
rect 655216 714407 655222 714459
rect 655274 714447 655280 714459
rect 676144 714447 676150 714459
rect 655274 714419 676150 714447
rect 655274 714407 655280 714419
rect 676144 714407 676150 714419
rect 676202 714407 676208 714459
rect 43216 714259 43222 714311
rect 43274 714299 43280 714311
rect 59632 714299 59638 714311
rect 43274 714271 59638 714299
rect 43274 714259 43280 714271
rect 59632 714259 59638 714271
rect 59690 714259 59696 714311
rect 673360 714185 673366 714237
rect 673418 714225 673424 714237
rect 676048 714225 676054 714237
rect 673418 714197 676054 714225
rect 673418 714185 673424 714197
rect 676048 714185 676054 714197
rect 676106 714185 676112 714237
rect 41680 714037 41686 714089
rect 41738 714077 41744 714089
rect 43504 714077 43510 714089
rect 41738 714049 43510 714077
rect 41738 714037 41744 714049
rect 43504 714037 43510 714049
rect 43562 714037 43568 714089
rect 42160 713889 42166 713941
rect 42218 713929 42224 713941
rect 43408 713929 43414 713941
rect 42218 713901 43414 713929
rect 42218 713889 42224 713901
rect 43408 713889 43414 713901
rect 43466 713889 43472 713941
rect 41776 713815 41782 713867
rect 41834 713815 41840 713867
rect 41794 713571 41822 713815
rect 41776 713519 41782 713571
rect 41834 713519 41840 713571
rect 672688 713371 672694 713423
rect 672746 713411 672752 713423
rect 676240 713411 676246 713423
rect 672746 713383 676246 713411
rect 672746 713371 672752 713383
rect 676240 713371 676246 713383
rect 676298 713371 676304 713423
rect 669712 713075 669718 713127
rect 669770 713115 669776 713127
rect 670960 713115 670966 713127
rect 669770 713087 670966 713115
rect 669770 713075 669776 713087
rect 670960 713075 670966 713087
rect 671018 713115 671024 713127
rect 676048 713115 676054 713127
rect 671018 713087 676054 713115
rect 671018 713075 671024 713087
rect 676048 713075 676054 713087
rect 676106 713075 676112 713127
rect 670672 712631 670678 712683
rect 670730 712671 670736 712683
rect 676048 712671 676054 712683
rect 670730 712643 676054 712671
rect 670730 712631 670736 712643
rect 676048 712631 676054 712643
rect 676106 712631 676112 712683
rect 42448 711965 42454 712017
rect 42506 712005 42512 712017
rect 43216 712005 43222 712017
rect 42506 711977 43222 712005
rect 42506 711965 42512 711977
rect 43216 711965 43222 711977
rect 43274 711965 43280 712017
rect 669520 711891 669526 711943
rect 669578 711931 669584 711943
rect 670864 711931 670870 711943
rect 669578 711903 670870 711931
rect 669578 711891 669584 711903
rect 670864 711891 670870 711903
rect 670922 711931 670928 711943
rect 676240 711931 676246 711943
rect 670922 711903 676246 711931
rect 670922 711891 670928 711903
rect 676240 711891 676246 711903
rect 676298 711891 676304 711943
rect 43216 711817 43222 711869
rect 43274 711857 43280 711869
rect 43792 711857 43798 711869
rect 43274 711829 43798 711857
rect 43274 711817 43280 711829
rect 43792 711817 43798 711829
rect 43850 711817 43856 711869
rect 43024 711521 43030 711573
rect 43082 711561 43088 711573
rect 43408 711561 43414 711573
rect 43082 711533 43414 711561
rect 43082 711521 43088 711533
rect 43408 711521 43414 711533
rect 43466 711521 43472 711573
rect 670768 711521 670774 711573
rect 670826 711561 670832 711573
rect 676048 711561 676054 711573
rect 670826 711533 676054 711561
rect 670826 711521 670832 711533
rect 676048 711521 676054 711533
rect 676106 711521 676112 711573
rect 43408 711373 43414 711425
rect 43466 711413 43472 711425
rect 43888 711413 43894 711425
rect 43466 711385 43894 711413
rect 43466 711373 43472 711385
rect 43888 711373 43894 711385
rect 43946 711373 43952 711425
rect 674896 711299 674902 711351
rect 674954 711339 674960 711351
rect 676048 711339 676054 711351
rect 674954 711311 676054 711339
rect 674954 711299 674960 711311
rect 676048 711299 676054 711311
rect 676106 711299 676112 711351
rect 43024 711151 43030 711203
rect 43082 711191 43088 711203
rect 43082 711163 43646 711191
rect 43082 711151 43088 711163
rect 43618 711129 43646 711163
rect 43600 711077 43606 711129
rect 43658 711077 43664 711129
rect 674512 711077 674518 711129
rect 674570 711117 674576 711129
rect 676048 711117 676054 711129
rect 674570 711089 676054 711117
rect 674570 711077 674576 711089
rect 676048 711077 676054 711089
rect 676106 711077 676112 711129
rect 42160 710855 42166 710907
rect 42218 710895 42224 710907
rect 42448 710895 42454 710907
rect 42218 710867 42454 710895
rect 42218 710855 42224 710867
rect 42448 710855 42454 710867
rect 42506 710855 42512 710907
rect 42160 709893 42166 709945
rect 42218 709933 42224 709945
rect 43504 709933 43510 709945
rect 42218 709905 43510 709933
rect 42218 709893 42224 709905
rect 43504 709893 43510 709905
rect 43562 709893 43568 709945
rect 42064 708487 42070 708539
rect 42122 708527 42128 708539
rect 43504 708527 43510 708539
rect 42122 708499 43510 708527
rect 42122 708487 42128 708499
rect 43504 708487 43510 708499
rect 43562 708487 43568 708539
rect 674992 708413 674998 708465
rect 675050 708453 675056 708465
rect 676048 708453 676054 708465
rect 675050 708425 676054 708453
rect 675050 708413 675056 708425
rect 676048 708413 676054 708425
rect 676106 708413 676112 708465
rect 42064 708339 42070 708391
rect 42122 708379 42128 708391
rect 43120 708379 43126 708391
rect 42122 708351 43126 708379
rect 42122 708339 42128 708351
rect 43120 708339 43126 708351
rect 43178 708339 43184 708391
rect 43120 708191 43126 708243
rect 43178 708231 43184 708243
rect 43600 708231 43606 708243
rect 43178 708203 43606 708231
rect 43178 708191 43184 708203
rect 43600 708191 43606 708203
rect 43658 708191 43664 708243
rect 42160 708043 42166 708095
rect 42218 708083 42224 708095
rect 42928 708083 42934 708095
rect 42218 708055 42934 708083
rect 42218 708043 42224 708055
rect 42928 708043 42934 708055
rect 42986 708043 42992 708095
rect 42160 706563 42166 706615
rect 42218 706603 42224 706615
rect 43120 706603 43126 706615
rect 42218 706575 43126 706603
rect 42218 706563 42224 706575
rect 43120 706563 43126 706575
rect 43178 706563 43184 706615
rect 42928 706415 42934 706467
rect 42986 706455 42992 706467
rect 43120 706455 43126 706467
rect 42986 706427 43126 706455
rect 42986 706415 42992 706427
rect 43120 706415 43126 706427
rect 43178 706415 43184 706467
rect 42448 704935 42454 704987
rect 42506 704935 42512 704987
rect 42160 704269 42166 704321
rect 42218 704309 42224 704321
rect 42466 704309 42494 704935
rect 673072 704861 673078 704913
rect 673130 704901 673136 704913
rect 676240 704901 676246 704913
rect 673130 704873 676246 704901
rect 673130 704861 673136 704873
rect 676240 704861 676246 704873
rect 676298 704861 676304 704913
rect 42218 704281 42494 704309
rect 42218 704269 42224 704281
rect 42064 703677 42070 703729
rect 42122 703717 42128 703729
rect 43024 703717 43030 703729
rect 42122 703689 43030 703717
rect 42122 703677 42128 703689
rect 43024 703677 43030 703689
rect 43082 703677 43088 703729
rect 653776 702789 653782 702841
rect 653834 702829 653840 702841
rect 675376 702829 675382 702841
rect 653834 702801 675382 702829
rect 653834 702789 653840 702801
rect 675376 702789 675382 702801
rect 675434 702789 675440 702841
rect 649456 702715 649462 702767
rect 649514 702755 649520 702767
rect 679984 702755 679990 702767
rect 649514 702727 679990 702755
rect 649514 702715 649520 702727
rect 679984 702715 679990 702727
rect 680042 702715 680048 702767
rect 42160 702641 42166 702693
rect 42218 702681 42224 702693
rect 42352 702681 42358 702693
rect 42218 702653 42358 702681
rect 42218 702641 42224 702653
rect 42352 702641 42358 702653
rect 42410 702641 42416 702693
rect 43504 702641 43510 702693
rect 43562 702681 43568 702693
rect 58768 702681 58774 702693
rect 43562 702653 58774 702681
rect 43562 702641 43568 702653
rect 58768 702641 58774 702653
rect 58826 702641 58832 702693
rect 44944 702567 44950 702619
rect 45002 702607 45008 702619
rect 58672 702607 58678 702619
rect 45002 702579 58678 702607
rect 45002 702567 45008 702579
rect 58672 702567 58678 702579
rect 58730 702567 58736 702619
rect 42160 702271 42166 702323
rect 42218 702311 42224 702323
rect 43120 702311 43126 702323
rect 42218 702283 43126 702311
rect 42218 702271 42224 702283
rect 43120 702271 43126 702283
rect 43178 702271 43184 702323
rect 42064 700495 42070 700547
rect 42122 700535 42128 700547
rect 43024 700535 43030 700547
rect 42122 700507 43030 700535
rect 42122 700495 42128 700507
rect 43024 700495 43030 700507
rect 43082 700495 43088 700547
rect 47632 699755 47638 699807
rect 47690 699795 47696 699807
rect 59248 699795 59254 699807
rect 47690 699767 59254 699795
rect 47690 699755 47696 699767
rect 59248 699755 59254 699767
rect 59306 699755 59312 699807
rect 44848 699681 44854 699733
rect 44906 699721 44912 699733
rect 58864 699721 58870 699733
rect 44906 699693 58870 699721
rect 44906 699681 44912 699693
rect 58864 699681 58870 699693
rect 58922 699681 58928 699733
rect 42160 699385 42166 699437
rect 42218 699425 42224 699437
rect 42928 699425 42934 699437
rect 42218 699397 42934 699425
rect 42218 699385 42224 699397
rect 42928 699385 42934 699397
rect 42986 699385 42992 699437
rect 42064 698719 42070 698771
rect 42122 698759 42128 698771
rect 45232 698759 45238 698771
rect 42122 698731 45238 698759
rect 42122 698719 42128 698731
rect 45232 698719 45238 698731
rect 45290 698719 45296 698771
rect 654160 694131 654166 694183
rect 654218 694171 654224 694183
rect 674992 694171 674998 694183
rect 654218 694143 674998 694171
rect 654218 694131 654224 694143
rect 674992 694131 674998 694143
rect 675050 694131 675056 694183
rect 672592 693613 672598 693665
rect 672650 693653 672656 693665
rect 675472 693653 675478 693665
rect 672650 693625 675478 693653
rect 672650 693613 672656 693625
rect 675472 693613 675478 693625
rect 675530 693613 675536 693665
rect 673072 692873 673078 692925
rect 673130 692913 673136 692925
rect 675376 692913 675382 692925
rect 673130 692885 675382 692913
rect 673130 692873 673136 692885
rect 675376 692873 675382 692885
rect 675434 692873 675440 692925
rect 654064 691319 654070 691371
rect 654122 691359 654128 691371
rect 675184 691359 675190 691371
rect 654122 691331 675190 691359
rect 654122 691319 654128 691331
rect 675184 691319 675190 691331
rect 675242 691319 675248 691371
rect 674896 690431 674902 690483
rect 674954 690471 674960 690483
rect 675472 690471 675478 690483
rect 674954 690443 675478 690471
rect 674954 690431 674960 690443
rect 675472 690431 675478 690443
rect 675530 690431 675536 690483
rect 672976 689765 672982 689817
rect 673034 689805 673040 689817
rect 675376 689805 675382 689817
rect 673034 689777 675382 689805
rect 673034 689765 673040 689777
rect 675376 689765 675382 689777
rect 675434 689765 675440 689817
rect 672016 689321 672022 689373
rect 672074 689361 672080 689373
rect 675376 689361 675382 689373
rect 672074 689333 675382 689361
rect 672074 689321 672080 689333
rect 675376 689321 675382 689333
rect 675434 689321 675440 689373
rect 672208 689099 672214 689151
rect 672266 689139 672272 689151
rect 675376 689139 675382 689151
rect 672266 689111 675382 689139
rect 672266 689099 672272 689111
rect 675376 689099 675382 689111
rect 675434 689099 675440 689151
rect 674992 688877 674998 688929
rect 675050 688917 675056 688929
rect 675472 688917 675478 688929
rect 675050 688889 675478 688917
rect 675050 688877 675056 688889
rect 675472 688877 675478 688889
rect 675530 688877 675536 688929
rect 41776 688211 41782 688263
rect 41834 688251 41840 688263
rect 50320 688251 50326 688263
rect 41834 688223 50326 688251
rect 41834 688211 41840 688223
rect 50320 688211 50326 688223
rect 50378 688211 50384 688263
rect 41584 687471 41590 687523
rect 41642 687511 41648 687523
rect 47728 687511 47734 687523
rect 41642 687483 47734 687511
rect 41642 687471 41648 687483
rect 47728 687471 47734 687483
rect 47786 687471 47792 687523
rect 672496 687323 672502 687375
rect 672554 687363 672560 687375
rect 675472 687363 675478 687375
rect 672554 687335 675478 687363
rect 672554 687323 672560 687335
rect 675472 687323 675478 687335
rect 675530 687323 675536 687375
rect 41776 687175 41782 687227
rect 41834 687215 41840 687227
rect 45040 687215 45046 687227
rect 41834 687187 45046 687215
rect 41834 687175 41840 687187
rect 45040 687175 45046 687187
rect 45098 687175 45104 687227
rect 675184 687027 675190 687079
rect 675242 687067 675248 687079
rect 675472 687067 675478 687079
rect 675242 687039 675478 687067
rect 675242 687027 675248 687039
rect 675472 687027 675478 687039
rect 675530 687027 675536 687079
rect 41584 686953 41590 687005
rect 41642 686993 41648 687005
rect 43408 686993 43414 687005
rect 41642 686965 43414 686993
rect 41642 686953 41648 686965
rect 43408 686953 43414 686965
rect 43466 686953 43472 687005
rect 41584 685991 41590 686043
rect 41642 686031 41648 686043
rect 43504 686031 43510 686043
rect 41642 686003 43510 686031
rect 41642 685991 41648 686003
rect 43504 685991 43510 686003
rect 43562 685991 43568 686043
rect 674320 685473 674326 685525
rect 674378 685513 674384 685525
rect 675472 685513 675478 685525
rect 674378 685485 675478 685513
rect 674378 685473 674384 685485
rect 675472 685473 675478 685485
rect 675530 685473 675536 685525
rect 41776 685325 41782 685377
rect 41834 685365 41840 685377
rect 43216 685365 43222 685377
rect 41834 685337 43222 685365
rect 41834 685325 41840 685337
rect 43216 685325 43222 685337
rect 43274 685365 43280 685377
rect 44944 685365 44950 685377
rect 43274 685337 44950 685365
rect 43274 685325 43280 685337
rect 44944 685325 44950 685337
rect 45002 685325 45008 685377
rect 41776 684141 41782 684193
rect 41834 684181 41840 684193
rect 43312 684181 43318 684193
rect 41834 684153 43318 684181
rect 41834 684141 41840 684153
rect 43312 684141 43318 684153
rect 43370 684181 43376 684193
rect 44848 684181 44854 684193
rect 43370 684153 44854 684181
rect 43370 684141 43376 684153
rect 44848 684141 44854 684153
rect 44906 684141 44912 684193
rect 674512 683623 674518 683675
rect 674570 683663 674576 683675
rect 675472 683663 675478 683675
rect 674570 683635 675478 683663
rect 674570 683623 674576 683635
rect 675472 683623 675478 683635
rect 675530 683623 675536 683675
rect 41776 683031 41782 683083
rect 41834 683071 41840 683083
rect 42928 683071 42934 683083
rect 41834 683043 42934 683071
rect 41834 683031 41840 683043
rect 42928 683031 42934 683043
rect 42986 683031 42992 683083
rect 41584 677259 41590 677311
rect 41642 677299 41648 677311
rect 43120 677299 43126 677311
rect 41642 677271 43126 677299
rect 41642 677259 41648 677271
rect 43120 677259 43126 677271
rect 43178 677259 43184 677311
rect 41584 676963 41590 677015
rect 41642 677003 41648 677015
rect 43024 677003 43030 677015
rect 41642 676975 43030 677003
rect 41642 676963 41648 676975
rect 43024 676963 43030 676975
rect 43082 676963 43088 677015
rect 41584 675483 41590 675535
rect 41642 675523 41648 675535
rect 47632 675523 47638 675535
rect 41642 675495 47638 675523
rect 41642 675483 41648 675495
rect 47632 675483 47638 675495
rect 47690 675483 47696 675535
rect 34480 672449 34486 672501
rect 34538 672489 34544 672501
rect 40336 672489 40342 672501
rect 34538 672461 40342 672489
rect 34538 672449 34544 672461
rect 40336 672449 40342 672461
rect 40394 672449 40400 672501
rect 37360 671265 37366 671317
rect 37418 671305 37424 671317
rect 43696 671305 43702 671317
rect 37418 671277 43702 671305
rect 37418 671265 37424 671277
rect 43696 671265 43702 671277
rect 43754 671265 43760 671317
rect 39856 671191 39862 671243
rect 39914 671231 39920 671243
rect 43600 671231 43606 671243
rect 39914 671203 43606 671231
rect 39914 671191 39920 671203
rect 43600 671191 43606 671203
rect 43658 671191 43664 671243
rect 40336 671117 40342 671169
rect 40394 671157 40400 671169
rect 43312 671157 43318 671169
rect 40394 671129 43318 671157
rect 40394 671117 40400 671129
rect 43312 671117 43318 671129
rect 43370 671117 43376 671169
rect 42736 671043 42742 671095
rect 42794 671083 42800 671095
rect 59632 671083 59638 671095
rect 42794 671055 59638 671083
rect 42794 671043 42800 671055
rect 59632 671043 59638 671055
rect 59690 671043 59696 671095
rect 43504 670969 43510 671021
rect 43562 670969 43568 671021
rect 41680 670821 41686 670873
rect 41738 670861 41744 670873
rect 42832 670861 42838 670873
rect 41738 670833 42838 670861
rect 41738 670821 41744 670833
rect 42832 670821 42838 670833
rect 42890 670821 42896 670873
rect 43024 670821 43030 670873
rect 43082 670861 43088 670873
rect 43312 670861 43318 670873
rect 43082 670833 43318 670861
rect 43082 670821 43088 670833
rect 43312 670821 43318 670833
rect 43370 670821 43376 670873
rect 42256 670747 42262 670799
rect 42314 670787 42320 670799
rect 42314 670759 43454 670787
rect 42314 670747 42320 670759
rect 43426 670725 43454 670759
rect 43522 670725 43550 670969
rect 42064 670673 42070 670725
rect 42122 670713 42128 670725
rect 43120 670713 43126 670725
rect 42122 670685 43126 670713
rect 42122 670673 42128 670685
rect 43120 670673 43126 670685
rect 43178 670673 43184 670725
rect 43408 670673 43414 670725
rect 43466 670673 43472 670725
rect 43504 670673 43510 670725
rect 43562 670673 43568 670725
rect 41776 670599 41782 670651
rect 41834 670599 41840 670651
rect 41872 670599 41878 670651
rect 41930 670639 41936 670651
rect 43024 670639 43030 670651
rect 41930 670611 43030 670639
rect 41930 670599 41936 670611
rect 43024 670599 43030 670611
rect 43082 670599 43088 670651
rect 41794 670355 41822 670599
rect 41776 670303 41782 670355
rect 41834 670303 41840 670355
rect 672688 669193 672694 669245
rect 672746 669233 672752 669245
rect 676048 669233 676054 669245
rect 672746 669205 676054 669233
rect 672746 669193 672752 669205
rect 676048 669193 676054 669205
rect 676106 669193 676112 669245
rect 42160 668527 42166 668579
rect 42218 668567 42224 668579
rect 42928 668567 42934 668579
rect 42218 668539 42934 668567
rect 42218 668527 42224 668539
rect 42928 668527 42934 668539
rect 42986 668527 42992 668579
rect 655504 668527 655510 668579
rect 655562 668567 655568 668579
rect 676144 668567 676150 668579
rect 655562 668539 676150 668567
rect 655562 668527 655568 668539
rect 676144 668527 676150 668539
rect 676202 668527 676208 668579
rect 673264 668453 673270 668505
rect 673322 668493 673328 668505
rect 676048 668493 676054 668505
rect 673322 668465 676054 668493
rect 673322 668453 673328 668465
rect 676048 668453 676054 668465
rect 676106 668453 676112 668505
rect 42928 668379 42934 668431
rect 42986 668419 42992 668431
rect 43216 668419 43222 668431
rect 42986 668391 43222 668419
rect 42986 668379 42992 668391
rect 43216 668379 43222 668391
rect 43274 668379 43280 668431
rect 655312 668379 655318 668431
rect 655370 668419 655376 668431
rect 676240 668419 676246 668431
rect 655370 668391 676246 668419
rect 655370 668379 655376 668391
rect 676240 668379 676246 668391
rect 676298 668379 676304 668431
rect 655120 668157 655126 668209
rect 655178 668197 655184 668209
rect 676336 668197 676342 668209
rect 655178 668169 676342 668197
rect 655178 668157 655184 668169
rect 676336 668157 676342 668169
rect 676394 668157 676400 668209
rect 674416 668083 674422 668135
rect 674474 668123 674480 668135
rect 676048 668123 676054 668135
rect 674474 668095 676054 668123
rect 674474 668083 674480 668095
rect 676048 668083 676054 668095
rect 676106 668083 676112 668135
rect 670672 668009 670678 668061
rect 670730 668049 670736 668061
rect 675952 668049 675958 668061
rect 670730 668021 675958 668049
rect 670730 668009 670736 668021
rect 675952 668009 675958 668021
rect 676010 668009 676016 668061
rect 42160 667861 42166 667913
rect 42218 667901 42224 667913
rect 42736 667901 42742 667913
rect 42218 667873 42742 667901
rect 42218 667861 42224 667873
rect 42736 667861 42742 667873
rect 42794 667861 42800 667913
rect 42736 667713 42742 667765
rect 42794 667753 42800 667765
rect 43312 667753 43318 667765
rect 42794 667725 43318 667753
rect 42794 667713 42800 667725
rect 43312 667713 43318 667725
rect 43370 667713 43376 667765
rect 670768 667639 670774 667691
rect 670826 667679 670832 667691
rect 675952 667679 675958 667691
rect 670826 667651 675958 667679
rect 670826 667639 670832 667651
rect 675952 667639 675958 667651
rect 676010 667639 676016 667691
rect 652240 666751 652246 666803
rect 652298 666791 652304 666803
rect 670864 666791 670870 666803
rect 652298 666763 670870 666791
rect 652298 666751 652304 666763
rect 670864 666751 670870 666763
rect 670922 666791 670928 666803
rect 676240 666791 676246 666803
rect 670922 666763 676246 666791
rect 670922 666751 670928 666763
rect 676240 666751 676246 666763
rect 676298 666751 676304 666803
rect 42160 666677 42166 666729
rect 42218 666717 42224 666729
rect 42928 666717 42934 666729
rect 42218 666689 42934 666717
rect 42218 666677 42224 666689
rect 42928 666677 42934 666689
rect 42986 666677 42992 666729
rect 649744 666677 649750 666729
rect 649802 666717 649808 666729
rect 670672 666717 670678 666729
rect 649802 666689 670678 666717
rect 649802 666677 649808 666689
rect 670672 666677 670678 666689
rect 670730 666677 670736 666729
rect 42928 666529 42934 666581
rect 42986 666569 42992 666581
rect 43408 666569 43414 666581
rect 42986 666541 43414 666569
rect 42986 666529 42992 666541
rect 43408 666529 43414 666541
rect 43466 666529 43472 666581
rect 670960 666307 670966 666359
rect 671018 666347 671024 666359
rect 676240 666347 676246 666359
rect 671018 666319 676246 666347
rect 671018 666307 671024 666319
rect 676240 666307 676246 666319
rect 676298 666307 676304 666359
rect 42160 665271 42166 665323
rect 42218 665311 42224 665323
rect 43216 665311 43222 665323
rect 42218 665283 43222 665311
rect 42218 665271 42224 665283
rect 43216 665271 43222 665283
rect 43274 665271 43280 665323
rect 674224 665197 674230 665249
rect 674282 665237 674288 665249
rect 676048 665237 676054 665249
rect 674282 665209 676054 665237
rect 674282 665197 674288 665209
rect 676048 665197 676054 665209
rect 676106 665197 676112 665249
rect 42160 665123 42166 665175
rect 42218 665163 42224 665175
rect 42736 665163 42742 665175
rect 42218 665135 42742 665163
rect 42218 665123 42224 665135
rect 42736 665123 42742 665135
rect 42794 665123 42800 665175
rect 42160 664827 42166 664879
rect 42218 664867 42224 664879
rect 43120 664867 43126 664879
rect 42218 664839 43126 664867
rect 42218 664827 42224 664839
rect 43120 664827 43126 664839
rect 43178 664827 43184 664879
rect 43120 664679 43126 664731
rect 43178 664719 43184 664731
rect 43600 664719 43606 664731
rect 43178 664691 43606 664719
rect 43178 664679 43184 664691
rect 43600 664679 43606 664691
rect 43658 664679 43664 664731
rect 42064 664161 42070 664213
rect 42122 664201 42128 664213
rect 42832 664201 42838 664213
rect 42122 664173 42838 664201
rect 42122 664161 42128 664173
rect 42832 664161 42838 664173
rect 42890 664161 42896 664213
rect 42160 663347 42166 663399
rect 42218 663387 42224 663399
rect 43024 663387 43030 663399
rect 42218 663359 43030 663387
rect 42218 663347 42224 663359
rect 43024 663347 43030 663359
rect 43082 663347 43088 663399
rect 43024 663199 43030 663251
rect 43082 663239 43088 663251
rect 43696 663239 43702 663251
rect 43082 663211 43702 663239
rect 43082 663199 43088 663211
rect 43696 663199 43702 663211
rect 43754 663199 43760 663251
rect 672112 662089 672118 662141
rect 672170 662129 672176 662141
rect 676048 662129 676054 662141
rect 672170 662101 676054 662129
rect 672170 662089 672176 662101
rect 676048 662089 676054 662101
rect 676106 662089 676112 662141
rect 672784 661645 672790 661697
rect 672842 661685 672848 661697
rect 676048 661685 676054 661697
rect 672842 661657 676054 661685
rect 672842 661645 672848 661657
rect 676048 661645 676054 661657
rect 676106 661645 676112 661697
rect 672304 661349 672310 661401
rect 672362 661389 672368 661401
rect 676240 661389 676246 661401
rect 672362 661361 676246 661389
rect 672362 661349 672368 661361
rect 676240 661349 676246 661361
rect 676298 661349 676304 661401
rect 42064 660905 42070 660957
rect 42122 660945 42128 660957
rect 42928 660945 42934 660957
rect 42122 660917 42934 660945
rect 42122 660905 42128 660917
rect 42928 660905 42934 660917
rect 42986 660905 42992 660957
rect 673168 660609 673174 660661
rect 673226 660649 673232 660661
rect 676048 660649 676054 660661
rect 673226 660621 676054 660649
rect 673226 660609 673232 660621
rect 676048 660609 676054 660621
rect 676106 660609 676112 660661
rect 42064 660387 42070 660439
rect 42122 660427 42128 660439
rect 43120 660427 43126 660439
rect 42122 660399 43126 660427
rect 42122 660387 42128 660399
rect 43120 660387 43126 660399
rect 43178 660387 43184 660439
rect 672880 660165 672886 660217
rect 672938 660205 672944 660217
rect 676048 660205 676054 660217
rect 672938 660177 676054 660205
rect 672938 660165 672944 660177
rect 676048 660165 676054 660177
rect 676106 660165 676112 660217
rect 672400 659869 672406 659921
rect 672458 659909 672464 659921
rect 676240 659909 676246 659921
rect 672458 659881 676246 659909
rect 672458 659869 672464 659881
rect 676240 659869 676246 659881
rect 676298 659869 676304 659921
rect 42160 659647 42166 659699
rect 42218 659687 42224 659699
rect 43024 659687 43030 659699
rect 42218 659659 43030 659687
rect 42218 659647 42224 659659
rect 43024 659647 43030 659659
rect 43082 659647 43088 659699
rect 43216 659425 43222 659477
rect 43274 659465 43280 659477
rect 58768 659465 58774 659477
rect 43274 659437 58774 659465
rect 43274 659425 43280 659437
rect 58768 659425 58774 659437
rect 58826 659425 58832 659477
rect 45040 659351 45046 659403
rect 45098 659391 45104 659403
rect 58672 659391 58678 659403
rect 45098 659363 58678 659391
rect 45098 659351 45104 659363
rect 58672 659351 58678 659363
rect 58730 659351 58736 659403
rect 42160 659203 42166 659255
rect 42218 659243 42224 659255
rect 43792 659243 43798 659255
rect 42218 659215 43798 659243
rect 42218 659203 42224 659215
rect 43792 659203 43798 659215
rect 43850 659203 43856 659255
rect 42064 657353 42070 657405
rect 42122 657393 42128 657405
rect 42736 657393 42742 657405
rect 42122 657365 42742 657393
rect 42122 657353 42128 657365
rect 42736 657353 42742 657365
rect 42794 657353 42800 657405
rect 654160 656761 654166 656813
rect 654218 656801 654224 656813
rect 675376 656801 675382 656813
rect 654218 656773 675382 656801
rect 654218 656761 654224 656773
rect 675376 656761 675382 656773
rect 675434 656761 675440 656813
rect 42160 656687 42166 656739
rect 42218 656727 42224 656739
rect 42832 656727 42838 656739
rect 42218 656699 42838 656727
rect 42218 656687 42224 656699
rect 42832 656687 42838 656699
rect 42890 656687 42896 656739
rect 649552 656687 649558 656739
rect 649610 656727 649616 656739
rect 679792 656727 679798 656739
rect 649610 656699 679798 656727
rect 649610 656687 649616 656699
rect 679792 656687 679798 656699
rect 679850 656687 679856 656739
rect 50320 656613 50326 656665
rect 50378 656653 50384 656665
rect 58192 656653 58198 656665
rect 50378 656625 58198 656653
rect 50378 656613 50384 656625
rect 58192 656613 58198 656625
rect 58250 656613 58256 656665
rect 47728 656539 47734 656591
rect 47786 656579 47792 656591
rect 58384 656579 58390 656591
rect 47786 656551 58390 656579
rect 47786 656539 47792 656551
rect 58384 656539 58390 656551
rect 58442 656539 58448 656591
rect 42160 656169 42166 656221
rect 42218 656209 42224 656221
rect 42928 656209 42934 656221
rect 42218 656181 42934 656209
rect 42218 656169 42224 656181
rect 42928 656169 42934 656181
rect 42986 656169 42992 656221
rect 42160 655503 42166 655555
rect 42218 655543 42224 655555
rect 43024 655543 43030 655555
rect 42218 655515 43030 655543
rect 42218 655503 42224 655515
rect 43024 655503 43030 655515
rect 43082 655503 43088 655555
rect 670864 648917 670870 648969
rect 670922 648957 670928 648969
rect 675184 648957 675190 648969
rect 670922 648929 675190 648957
rect 670922 648917 670928 648929
rect 675184 648917 675190 648929
rect 675242 648917 675248 648969
rect 672400 648251 672406 648303
rect 672458 648291 672464 648303
rect 675184 648291 675190 648303
rect 672458 648263 675190 648291
rect 672458 648251 672464 648263
rect 675184 648251 675190 648263
rect 675242 648251 675248 648303
rect 655792 648177 655798 648229
rect 655850 648217 655856 648229
rect 674992 648217 674998 648229
rect 655850 648189 674998 648217
rect 655850 648177 655856 648189
rect 674992 648177 674998 648189
rect 675050 648177 675056 648229
rect 673360 648029 673366 648081
rect 673418 648069 673424 648081
rect 675184 648069 675190 648081
rect 673418 648041 675190 648069
rect 673418 648029 673424 648041
rect 675184 648029 675190 648041
rect 675242 648029 675248 648081
rect 655984 645143 655990 645195
rect 656042 645183 656048 645195
rect 675280 645183 675286 645195
rect 656042 645155 675286 645183
rect 656042 645143 656048 645155
rect 675280 645143 675286 645155
rect 675338 645143 675344 645195
rect 41584 644847 41590 644899
rect 41642 644887 41648 644899
rect 50320 644887 50326 644899
rect 41642 644859 50326 644887
rect 41642 644847 41648 644859
rect 50320 644847 50326 644859
rect 50378 644847 50384 644899
rect 672880 644773 672886 644825
rect 672938 644813 672944 644825
rect 675376 644813 675382 644825
rect 672938 644785 675382 644813
rect 672938 644773 672944 644785
rect 675376 644773 675382 644785
rect 675434 644773 675440 644825
rect 41584 644255 41590 644307
rect 41642 644295 41648 644307
rect 47824 644295 47830 644307
rect 41642 644267 47830 644295
rect 41642 644255 41648 644267
rect 47824 644255 47830 644267
rect 47882 644255 47888 644307
rect 672784 644033 672790 644085
rect 672842 644073 672848 644085
rect 675472 644073 675478 644085
rect 672842 644045 675478 644073
rect 672842 644033 672848 644045
rect 675472 644033 675478 644045
rect 675530 644033 675536 644085
rect 41776 643959 41782 644011
rect 41834 643999 41840 644011
rect 47920 643999 47926 644011
rect 41834 643971 47926 643999
rect 41834 643959 41840 643971
rect 47920 643959 47926 643971
rect 47978 643959 47984 644011
rect 41584 643737 41590 643789
rect 41642 643777 41648 643789
rect 43504 643777 43510 643789
rect 41642 643749 43510 643777
rect 41642 643737 41648 643749
rect 43504 643737 43510 643749
rect 43562 643737 43568 643789
rect 674992 643663 674998 643715
rect 675050 643703 675056 643715
rect 675376 643703 675382 643715
rect 675050 643675 675382 643703
rect 675050 643663 675056 643675
rect 675376 643663 675382 643675
rect 675434 643663 675440 643715
rect 672688 643589 672694 643641
rect 672746 643629 672752 643641
rect 675472 643629 675478 643641
rect 672746 643601 675478 643629
rect 672746 643589 672752 643601
rect 675472 643589 675478 643601
rect 675530 643589 675536 643641
rect 41584 642775 41590 642827
rect 41642 642815 41648 642827
rect 43600 642815 43606 642827
rect 41642 642787 43606 642815
rect 41642 642775 41648 642787
rect 43600 642775 43606 642787
rect 43658 642775 43664 642827
rect 41488 642479 41494 642531
rect 41546 642519 41552 642531
rect 61936 642519 61942 642531
rect 41546 642491 61942 642519
rect 41546 642479 41552 642491
rect 61936 642479 61942 642491
rect 61994 642479 62000 642531
rect 670672 642257 670678 642309
rect 670730 642297 670736 642309
rect 675472 642297 675478 642309
rect 670730 642269 675478 642297
rect 670730 642257 670736 642269
rect 675472 642257 675478 642269
rect 675530 642257 675536 642309
rect 41584 641295 41590 641347
rect 41642 641335 41648 641347
rect 43504 641335 43510 641347
rect 41642 641307 43510 641335
rect 41642 641295 41648 641307
rect 43504 641295 43510 641307
rect 43562 641295 43568 641347
rect 41584 634487 41590 634539
rect 41642 634527 41648 634539
rect 43120 634527 43126 634539
rect 41642 634499 43126 634527
rect 41642 634487 41648 634499
rect 43120 634487 43126 634499
rect 43178 634487 43184 634539
rect 41776 634191 41782 634243
rect 41834 634231 41840 634243
rect 42928 634231 42934 634243
rect 41834 634203 42934 634231
rect 41834 634191 41840 634203
rect 42928 634191 42934 634203
rect 42986 634191 42992 634243
rect 41584 634117 41590 634169
rect 41642 634157 41648 634169
rect 43024 634157 43030 634169
rect 41642 634129 43030 634157
rect 41642 634117 41648 634129
rect 43024 634117 43030 634129
rect 43082 634117 43088 634169
rect 41776 633895 41782 633947
rect 41834 633935 41840 633947
rect 42832 633935 42838 633947
rect 41834 633907 42838 633935
rect 41834 633895 41840 633907
rect 42832 633895 42838 633907
rect 42890 633895 42896 633947
rect 41584 632267 41590 632319
rect 41642 632307 41648 632319
rect 47728 632307 47734 632319
rect 41642 632279 47734 632307
rect 41642 632267 41648 632279
rect 47728 632267 47734 632279
rect 47786 632267 47792 632319
rect 41968 632045 41974 632097
rect 42026 632085 42032 632097
rect 42736 632085 42742 632097
rect 42026 632057 42742 632085
rect 42026 632045 42032 632057
rect 42736 632045 42742 632057
rect 42794 632045 42800 632097
rect 40144 630639 40150 630691
rect 40202 630679 40208 630691
rect 42064 630679 42070 630691
rect 40202 630651 42070 630679
rect 40202 630639 40208 630651
rect 42064 630639 42070 630651
rect 42122 630639 42128 630691
rect 34384 629233 34390 629285
rect 34442 629273 34448 629285
rect 40432 629273 40438 629285
rect 34442 629245 40438 629273
rect 34442 629233 34448 629245
rect 40432 629233 40438 629245
rect 40490 629233 40496 629285
rect 37360 627901 37366 627953
rect 37418 627941 37424 627953
rect 43696 627941 43702 627953
rect 37418 627913 43702 627941
rect 37418 627901 37424 627913
rect 43696 627901 43702 627913
rect 43754 627901 43760 627953
rect 40432 627827 40438 627879
rect 40490 627867 40496 627879
rect 43216 627867 43222 627879
rect 40490 627839 43222 627867
rect 40490 627827 40496 627839
rect 43216 627827 43222 627839
rect 43274 627827 43280 627879
rect 41872 627383 41878 627435
rect 41930 627383 41936 627435
rect 42256 627383 42262 627435
rect 42314 627423 42320 627435
rect 43312 627423 43318 627435
rect 42314 627395 43318 627423
rect 42314 627383 42320 627395
rect 43312 627383 43318 627395
rect 43370 627383 43376 627435
rect 41890 627213 41918 627383
rect 41872 627161 41878 627213
rect 41930 627161 41936 627213
rect 42160 625311 42166 625363
rect 42218 625351 42224 625363
rect 42736 625351 42742 625363
rect 42218 625323 42742 625351
rect 42218 625311 42224 625323
rect 42736 625311 42742 625323
rect 42794 625311 42800 625363
rect 655408 624941 655414 624993
rect 655466 624981 655472 624993
rect 676240 624981 676246 624993
rect 655466 624953 676246 624981
rect 655466 624941 655472 624953
rect 676240 624941 676246 624953
rect 676298 624941 676304 624993
rect 42160 623979 42166 624031
rect 42218 624019 42224 624031
rect 58960 624019 58966 624031
rect 42218 623991 58966 624019
rect 42218 623979 42224 623991
rect 58960 623979 58966 623991
rect 59018 623979 59024 624031
rect 673264 623979 673270 624031
rect 673322 624019 673328 624031
rect 676048 624019 676054 624031
rect 673322 623991 676054 624019
rect 673322 623979 673328 623991
rect 676048 623979 676054 623991
rect 676106 623979 676112 624031
rect 42160 623461 42166 623513
rect 42218 623501 42224 623513
rect 42928 623501 42934 623513
rect 42218 623473 42934 623501
rect 42218 623461 42224 623473
rect 42928 623461 42934 623473
rect 42986 623461 42992 623513
rect 672304 623387 672310 623439
rect 672362 623427 672368 623439
rect 676048 623427 676054 623439
rect 672362 623399 676054 623427
rect 672362 623387 672368 623399
rect 676048 623387 676054 623399
rect 676106 623387 676112 623439
rect 42928 623313 42934 623365
rect 42986 623353 42992 623365
rect 43312 623353 43318 623365
rect 42986 623325 43318 623353
rect 42986 623313 42992 623325
rect 43312 623313 43318 623325
rect 43370 623313 43376 623365
rect 669616 622943 669622 622995
rect 669674 622983 669680 622995
rect 670768 622983 670774 622995
rect 669674 622955 670774 622983
rect 669674 622943 669680 622955
rect 670768 622943 670774 622955
rect 670826 622983 670832 622995
rect 676048 622983 676054 622995
rect 670826 622955 676054 622983
rect 670826 622943 670832 622955
rect 676048 622943 676054 622955
rect 676106 622943 676112 622995
rect 670576 622425 670582 622477
rect 670634 622465 670640 622477
rect 676048 622465 676054 622477
rect 670634 622437 676054 622465
rect 670634 622425 670640 622437
rect 676048 622425 676054 622437
rect 676106 622425 676112 622477
rect 655600 622351 655606 622403
rect 655658 622391 655664 622403
rect 676240 622391 676246 622403
rect 655658 622363 676246 622391
rect 655658 622351 655664 622363
rect 676240 622351 676246 622363
rect 676298 622351 676304 622403
rect 42160 622203 42166 622255
rect 42218 622243 42224 622255
rect 42832 622243 42838 622255
rect 42218 622215 42838 622243
rect 42218 622203 42224 622215
rect 42832 622203 42838 622215
rect 42890 622203 42896 622255
rect 655216 622203 655222 622255
rect 655274 622243 655280 622255
rect 676144 622243 676150 622255
rect 655274 622215 676150 622243
rect 655274 622203 655280 622215
rect 676144 622203 676150 622215
rect 676202 622203 676208 622255
rect 42064 622055 42070 622107
rect 42122 622095 42128 622107
rect 48016 622095 48022 622107
rect 42122 622067 48022 622095
rect 42122 622055 42128 622067
rect 48016 622055 48022 622067
rect 48074 622055 48080 622107
rect 674320 621981 674326 622033
rect 674378 622021 674384 622033
rect 676240 622021 676246 622033
rect 674378 621993 676246 622021
rect 674378 621981 674384 621993
rect 676240 621981 676246 621993
rect 676298 621981 676304 622033
rect 670960 621907 670966 621959
rect 671018 621947 671024 621959
rect 676048 621947 676054 621959
rect 671018 621919 676054 621947
rect 671018 621907 671024 621919
rect 676048 621907 676054 621919
rect 676106 621907 676112 621959
rect 42160 621611 42166 621663
rect 42218 621651 42224 621663
rect 43120 621651 43126 621663
rect 42218 621623 43126 621651
rect 42218 621611 42224 621623
rect 43120 621611 43126 621623
rect 43178 621611 43184 621663
rect 670480 621315 670486 621367
rect 670538 621355 670544 621367
rect 676048 621355 676054 621367
rect 670538 621327 676054 621355
rect 670538 621315 670544 621327
rect 676048 621315 676054 621327
rect 676106 621315 676112 621367
rect 42064 620945 42070 620997
rect 42122 620985 42128 620997
rect 43024 620985 43030 620997
rect 42122 620957 43030 620985
rect 42122 620945 42128 620957
rect 43024 620945 43030 620957
rect 43082 620945 43088 620997
rect 43216 620353 43222 620405
rect 43274 620393 43280 620405
rect 43600 620393 43606 620405
rect 43274 620365 43606 620393
rect 43274 620353 43280 620365
rect 43600 620353 43606 620365
rect 43658 620353 43664 620405
rect 42160 620131 42166 620183
rect 42218 620171 42224 620183
rect 42736 620171 42742 620183
rect 42218 620143 42742 620171
rect 42218 620131 42224 620143
rect 42736 620131 42742 620143
rect 42794 620131 42800 620183
rect 669808 619835 669814 619887
rect 669866 619875 669872 619887
rect 670960 619875 670966 619887
rect 669866 619847 670966 619875
rect 669866 619835 669872 619847
rect 670960 619835 670966 619847
rect 671018 619835 671024 619887
rect 674896 619021 674902 619073
rect 674954 619061 674960 619073
rect 676048 619061 676054 619073
rect 674954 619033 676054 619061
rect 674954 619021 674960 619033
rect 676048 619021 676054 619033
rect 676106 619021 676112 619073
rect 674512 618873 674518 618925
rect 674570 618913 674576 618925
rect 676240 618913 676246 618925
rect 674570 618885 676246 618913
rect 674570 618873 674576 618885
rect 676240 618873 676246 618885
rect 676298 618873 676304 618925
rect 42064 617837 42070 617889
rect 42122 617877 42128 617889
rect 43024 617877 43030 617889
rect 42122 617849 43030 617877
rect 42122 617837 42128 617849
rect 43024 617837 43030 617849
rect 43082 617837 43088 617889
rect 43024 617689 43030 617741
rect 43082 617729 43088 617741
rect 43600 617729 43606 617741
rect 43082 617701 43606 617729
rect 43082 617689 43088 617701
rect 43600 617689 43606 617701
rect 43658 617689 43664 617741
rect 42160 617171 42166 617223
rect 42218 617211 42224 617223
rect 42928 617211 42934 617223
rect 42218 617183 42934 617211
rect 42218 617171 42224 617183
rect 42928 617171 42934 617183
rect 42986 617171 42992 617223
rect 672592 617097 672598 617149
rect 672650 617137 672656 617149
rect 676240 617137 676246 617149
rect 672650 617109 676246 617137
rect 672650 617097 672656 617109
rect 676240 617097 676246 617109
rect 676298 617097 676304 617149
rect 42160 616653 42166 616705
rect 42218 616693 42224 616705
rect 43120 616693 43126 616705
rect 42218 616665 43126 616693
rect 42218 616653 42224 616665
rect 43120 616653 43126 616665
rect 43178 616653 43184 616705
rect 672496 616505 672502 616557
rect 672554 616545 672560 616557
rect 676048 616545 676054 616557
rect 672554 616517 676054 616545
rect 672554 616505 672560 616517
rect 676048 616505 676054 616517
rect 676106 616505 676112 616557
rect 42928 616357 42934 616409
rect 42986 616397 42992 616409
rect 58192 616397 58198 616409
rect 42986 616369 58198 616397
rect 42986 616357 42992 616369
rect 58192 616357 58198 616369
rect 58250 616357 58256 616409
rect 47920 616283 47926 616335
rect 47978 616323 47984 616335
rect 58960 616323 58966 616335
rect 47978 616295 58966 616323
rect 47978 616283 47984 616295
rect 58960 616283 58966 616295
rect 59018 616283 59024 616335
rect 48016 616209 48022 616261
rect 48074 616249 48080 616261
rect 59632 616249 59638 616261
rect 48074 616221 59638 616249
rect 48074 616209 48080 616221
rect 59632 616209 59638 616221
rect 59690 616209 59696 616261
rect 672016 615913 672022 615965
rect 672074 615953 672080 615965
rect 676048 615953 676054 615965
rect 672074 615925 676054 615953
rect 672074 615913 672080 615925
rect 676048 615913 676054 615925
rect 676106 615913 676112 615965
rect 42160 615839 42166 615891
rect 42218 615879 42224 615891
rect 42832 615879 42838 615891
rect 42218 615851 42838 615879
rect 42218 615839 42224 615851
rect 42832 615839 42838 615851
rect 42890 615839 42896 615891
rect 673072 615617 673078 615669
rect 673130 615657 673136 615669
rect 676240 615657 676246 615669
rect 673130 615629 676246 615657
rect 673130 615617 673136 615629
rect 676240 615617 676246 615629
rect 676298 615617 676304 615669
rect 672976 615173 672982 615225
rect 673034 615213 673040 615225
rect 676240 615213 676246 615225
rect 673034 615185 676246 615213
rect 673034 615173 673040 615185
rect 676240 615173 676246 615185
rect 676298 615173 676304 615225
rect 672208 614433 672214 614485
rect 672266 614473 672272 614485
rect 676048 614473 676054 614485
rect 672266 614445 676054 614473
rect 672266 614433 672272 614445
rect 676048 614433 676054 614445
rect 676106 614433 676112 614485
rect 42160 614137 42166 614189
rect 42218 614177 42224 614189
rect 43024 614177 43030 614189
rect 42218 614149 43030 614177
rect 42218 614137 42224 614149
rect 43024 614137 43030 614149
rect 43082 614137 43088 614189
rect 42160 613619 42166 613671
rect 42218 613659 42224 613671
rect 42736 613659 42742 613671
rect 42218 613631 42742 613659
rect 42218 613619 42224 613631
rect 42736 613619 42742 613631
rect 42794 613619 42800 613671
rect 655792 613471 655798 613523
rect 655850 613511 655856 613523
rect 675376 613511 675382 613523
rect 655850 613483 675382 613511
rect 655850 613471 655856 613483
rect 675376 613471 675382 613483
rect 675434 613471 675440 613523
rect 50320 613397 50326 613449
rect 50378 613437 50384 613449
rect 59632 613437 59638 613449
rect 50378 613409 59638 613437
rect 50378 613397 50384 613409
rect 59632 613397 59638 613409
rect 59690 613397 59696 613449
rect 47824 613323 47830 613375
rect 47882 613363 47888 613375
rect 59536 613363 59542 613375
rect 47882 613335 59542 613363
rect 47882 613323 47888 613335
rect 59536 613323 59542 613335
rect 59594 613323 59600 613375
rect 42064 612805 42070 612857
rect 42122 612845 42128 612857
rect 42352 612845 42358 612857
rect 42122 612817 42358 612845
rect 42122 612805 42128 612817
rect 42352 612805 42358 612817
rect 42410 612805 42416 612857
rect 42160 612139 42166 612191
rect 42218 612179 42224 612191
rect 42928 612179 42934 612191
rect 42218 612151 42934 612179
rect 42218 612139 42224 612151
rect 42928 612139 42934 612151
rect 42986 612139 42992 612191
rect 649648 610585 649654 610637
rect 649706 610625 649712 610637
rect 679984 610625 679990 610637
rect 649706 610597 679990 610625
rect 649706 610585 649712 610597
rect 679984 610585 679990 610597
rect 680042 610585 680048 610637
rect 670960 606885 670966 606937
rect 671018 606925 671024 606937
rect 675184 606925 675190 606937
rect 671018 606897 675190 606925
rect 671018 606885 671024 606897
rect 675184 606885 675190 606897
rect 675242 606885 675248 606937
rect 670768 603851 670774 603903
rect 670826 603891 670832 603903
rect 675280 603891 675286 603903
rect 670826 603863 675286 603891
rect 670826 603851 670832 603863
rect 675280 603851 675286 603863
rect 675338 603851 675344 603903
rect 673264 603037 673270 603089
rect 673322 603077 673328 603089
rect 675376 603077 675382 603089
rect 673322 603049 675382 603077
rect 673322 603037 673328 603049
rect 675376 603037 675382 603049
rect 675434 603037 675440 603089
rect 656560 602149 656566 602201
rect 656618 602189 656624 602201
rect 674896 602189 674902 602201
rect 656618 602161 674902 602189
rect 656618 602149 656624 602161
rect 674896 602149 674902 602161
rect 674954 602149 674960 602201
rect 653968 602001 653974 602053
rect 654026 602041 654032 602053
rect 674992 602041 674998 602053
rect 654026 602013 674998 602041
rect 654026 602001 654032 602013
rect 674992 602001 674998 602013
rect 675050 602001 675056 602053
rect 673168 601927 673174 601979
rect 673226 601967 673232 601979
rect 675280 601967 675286 601979
rect 673226 601939 675286 601967
rect 673226 601927 673232 601939
rect 675280 601927 675286 601939
rect 675338 601927 675344 601979
rect 41584 601631 41590 601683
rect 41642 601671 41648 601683
rect 50320 601671 50326 601683
rect 41642 601643 50326 601671
rect 41642 601631 41648 601643
rect 50320 601631 50326 601643
rect 50378 601631 50384 601683
rect 41776 601335 41782 601387
rect 41834 601375 41840 601387
rect 47824 601375 47830 601387
rect 41834 601347 47830 601375
rect 41834 601335 41840 601347
rect 47824 601335 47830 601347
rect 47882 601335 47888 601387
rect 41776 600743 41782 600795
rect 41834 600783 41840 600795
rect 47920 600783 47926 600795
rect 41834 600755 47926 600783
rect 41834 600743 41840 600755
rect 47920 600743 47926 600755
rect 47978 600743 47984 600795
rect 41776 600373 41782 600425
rect 41834 600413 41840 600425
rect 43216 600413 43222 600425
rect 41834 600385 43222 600413
rect 41834 600373 41840 600385
rect 43216 600373 43222 600385
rect 43274 600373 43280 600425
rect 41776 599781 41782 599833
rect 41834 599821 41840 599833
rect 43216 599821 43222 599833
rect 41834 599793 43222 599821
rect 41834 599781 41840 599793
rect 43216 599781 43222 599793
rect 43274 599781 43280 599833
rect 672976 599781 672982 599833
rect 673034 599821 673040 599833
rect 675376 599821 675382 599833
rect 673034 599793 675382 599821
rect 673034 599781 673040 599793
rect 675376 599781 675382 599793
rect 675434 599781 675440 599833
rect 41776 599263 41782 599315
rect 41834 599303 41840 599315
rect 43408 599303 43414 599315
rect 41834 599275 43414 599303
rect 41834 599263 41840 599275
rect 43408 599263 43414 599275
rect 43466 599263 43472 599315
rect 673072 599263 673078 599315
rect 673130 599303 673136 599315
rect 675376 599303 675382 599315
rect 673130 599275 675382 599303
rect 673130 599263 673136 599275
rect 675376 599263 675382 599275
rect 675434 599263 675440 599315
rect 672592 598893 672598 598945
rect 672650 598933 672656 598945
rect 675376 598933 675382 598945
rect 672650 598905 675382 598933
rect 672650 598893 672656 598905
rect 675376 598893 675382 598905
rect 675434 598893 675440 598945
rect 674992 598671 674998 598723
rect 675050 598711 675056 598723
rect 675472 598711 675478 598723
rect 675050 598683 675478 598711
rect 675050 598671 675056 598683
rect 675472 598671 675478 598683
rect 675530 598671 675536 598723
rect 41776 598301 41782 598353
rect 41834 598341 41840 598353
rect 43888 598341 43894 598353
rect 41834 598313 43894 598341
rect 41834 598301 41840 598313
rect 43888 598301 43894 598313
rect 43946 598301 43952 598353
rect 41776 597857 41782 597909
rect 41834 597897 41840 597909
rect 43312 597897 43318 597909
rect 41834 597869 43318 597897
rect 41834 597857 41840 597869
rect 43312 597857 43318 597869
rect 43370 597857 43376 597909
rect 672496 597117 672502 597169
rect 672554 597157 672560 597169
rect 675472 597157 675478 597169
rect 672554 597129 675478 597157
rect 672554 597117 672560 597129
rect 675472 597117 675478 597129
rect 675530 597117 675536 597169
rect 674896 596821 674902 596873
rect 674954 596861 674960 596873
rect 675376 596861 675382 596873
rect 674954 596833 675382 596861
rect 674954 596821 674960 596833
rect 675376 596821 675382 596833
rect 675434 596821 675440 596873
rect 41584 596599 41590 596651
rect 41642 596639 41648 596651
rect 43120 596639 43126 596651
rect 41642 596611 43126 596639
rect 41642 596599 41648 596611
rect 43120 596599 43126 596611
rect 43178 596599 43184 596651
rect 43312 596155 43318 596207
rect 43370 596195 43376 596207
rect 45040 596195 45046 596207
rect 43370 596167 45046 596195
rect 43370 596155 43376 596167
rect 45040 596155 45046 596167
rect 45098 596155 45104 596207
rect 41584 590975 41590 591027
rect 41642 591015 41648 591027
rect 43024 591015 43030 591027
rect 41642 590987 43030 591015
rect 41642 590975 41648 590987
rect 43024 590975 43030 590987
rect 43082 590975 43088 591027
rect 41872 590383 41878 590435
rect 41930 590423 41936 590435
rect 42928 590423 42934 590435
rect 41930 590395 42934 590423
rect 41930 590383 41936 590395
rect 42928 590383 42934 590395
rect 42986 590383 42992 590435
rect 41584 587497 41590 587549
rect 41642 587537 41648 587549
rect 56080 587537 56086 587549
rect 41642 587509 56086 587537
rect 41642 587497 41648 587509
rect 56080 587497 56086 587509
rect 56138 587497 56144 587549
rect 37360 584981 37366 585033
rect 37418 585021 37424 585033
rect 43792 585021 43798 585033
rect 37418 584993 43798 585021
rect 37418 584981 37424 584993
rect 43792 584981 43798 584993
rect 43850 584981 43856 585033
rect 40144 584833 40150 584885
rect 40202 584873 40208 584885
rect 41872 584873 41878 584885
rect 40202 584845 41878 584873
rect 40202 584833 40208 584845
rect 41872 584833 41878 584845
rect 41930 584833 41936 584885
rect 42064 584833 42070 584885
rect 42122 584873 42128 584885
rect 42544 584873 42550 584885
rect 42122 584845 42550 584873
rect 42122 584833 42128 584845
rect 42544 584833 42550 584845
rect 42602 584833 42608 584885
rect 34480 584759 34486 584811
rect 34538 584799 34544 584811
rect 43600 584799 43606 584811
rect 34538 584771 43606 584799
rect 34538 584759 34544 584771
rect 43600 584759 43606 584771
rect 43658 584759 43664 584811
rect 40240 584685 40246 584737
rect 40298 584725 40304 584737
rect 42256 584725 42262 584737
rect 40298 584697 42262 584725
rect 40298 584685 40304 584697
rect 42256 584685 42262 584697
rect 42314 584685 42320 584737
rect 42544 584685 42550 584737
rect 42602 584725 42608 584737
rect 58960 584725 58966 584737
rect 42602 584697 58966 584725
rect 42602 584685 42608 584697
rect 58960 584685 58966 584697
rect 59018 584685 59024 584737
rect 43024 584463 43030 584515
rect 43082 584503 43088 584515
rect 43504 584503 43510 584515
rect 43082 584475 43510 584503
rect 43082 584463 43088 584475
rect 43504 584463 43510 584475
rect 43562 584463 43568 584515
rect 43120 584389 43126 584441
rect 43178 584429 43184 584441
rect 43312 584429 43318 584441
rect 43178 584401 43318 584429
rect 43178 584389 43184 584401
rect 43312 584389 43318 584401
rect 43370 584389 43376 584441
rect 42160 584241 42166 584293
rect 42218 584281 42224 584293
rect 43120 584281 43126 584293
rect 42218 584253 43126 584281
rect 42218 584241 42224 584253
rect 43120 584241 43126 584253
rect 43178 584241 43184 584293
rect 41776 584167 41782 584219
rect 41834 584167 41840 584219
rect 41968 584167 41974 584219
rect 42026 584207 42032 584219
rect 42928 584207 42934 584219
rect 42026 584179 42934 584207
rect 42026 584167 42032 584179
rect 42928 584167 42934 584179
rect 42986 584167 42992 584219
rect 41794 583997 41822 584167
rect 41776 583945 41782 583997
rect 41834 583945 41840 583997
rect 42160 582095 42166 582147
rect 42218 582135 42224 582147
rect 43312 582135 43318 582147
rect 42218 582107 43318 582135
rect 42218 582095 42224 582107
rect 43312 582095 43318 582107
rect 43370 582095 43376 582147
rect 42064 581429 42070 581481
rect 42122 581469 42128 581481
rect 42544 581469 42550 581481
rect 42122 581441 42550 581469
rect 42122 581429 42128 581441
rect 42544 581429 42550 581441
rect 42602 581429 42608 581481
rect 42064 580245 42070 580297
rect 42122 580285 42128 580297
rect 43024 580285 43030 580297
rect 42122 580257 43030 580285
rect 42122 580245 42128 580257
rect 43024 580245 43030 580257
rect 43082 580245 43088 580297
rect 43024 580097 43030 580149
rect 43082 580137 43088 580149
rect 43504 580137 43510 580149
rect 43082 580109 43510 580137
rect 43082 580097 43088 580109
rect 43504 580097 43510 580109
rect 43562 580097 43568 580149
rect 42160 579283 42166 579335
rect 42218 579323 42224 579335
rect 48016 579323 48022 579335
rect 42218 579295 48022 579323
rect 42218 579283 42224 579295
rect 48016 579283 48022 579295
rect 48074 579283 48080 579335
rect 42160 578839 42166 578891
rect 42218 578879 42224 578891
rect 43024 578879 43030 578891
rect 42218 578851 43030 578879
rect 42218 578839 42224 578851
rect 43024 578839 43030 578851
rect 43082 578839 43088 578891
rect 42064 578395 42070 578447
rect 42122 578435 42128 578447
rect 42544 578435 42550 578447
rect 42122 578407 42550 578435
rect 42122 578395 42128 578407
rect 42544 578395 42550 578407
rect 42602 578395 42608 578447
rect 42160 577655 42166 577707
rect 42218 577695 42224 577707
rect 43120 577695 43126 577707
rect 42218 577667 43126 577695
rect 42218 577655 42224 577667
rect 43120 577655 43126 577667
rect 43178 577655 43184 577707
rect 43120 577507 43126 577559
rect 43178 577547 43184 577559
rect 43600 577547 43606 577559
rect 43178 577519 43606 577547
rect 43178 577507 43184 577519
rect 43600 577507 43606 577519
rect 43658 577507 43664 577559
rect 42064 577137 42070 577189
rect 42122 577177 42128 577189
rect 42928 577177 42934 577189
rect 42122 577149 42934 577177
rect 42122 577137 42128 577149
rect 42928 577137 42934 577149
rect 42986 577137 42992 577189
rect 42928 576989 42934 577041
rect 42986 577029 42992 577041
rect 43792 577029 43798 577041
rect 42986 577001 43798 577029
rect 42986 576989 42992 577001
rect 43792 576989 43798 577001
rect 43850 576989 43856 577041
rect 672304 576989 672310 577041
rect 672362 577029 672368 577041
rect 676048 577029 676054 577041
rect 672362 577001 676054 577029
rect 672362 576989 672368 577001
rect 676048 576989 676054 577001
rect 676106 576989 676112 577041
rect 655504 576471 655510 576523
rect 655562 576511 655568 576523
rect 676240 576511 676246 576523
rect 655562 576483 676246 576511
rect 655562 576471 655568 576483
rect 676240 576471 676246 576483
rect 676298 576471 676304 576523
rect 655312 576323 655318 576375
rect 655370 576363 655376 576375
rect 676144 576363 676150 576375
rect 655370 576335 676150 576363
rect 655370 576323 655376 576335
rect 676144 576323 676150 576335
rect 676202 576323 676208 576375
rect 655120 576175 655126 576227
rect 655178 576215 655184 576227
rect 676336 576215 676342 576227
rect 655178 576187 676342 576215
rect 655178 576175 655184 576187
rect 676336 576175 676342 576187
rect 676394 576175 676400 576227
rect 673840 576101 673846 576153
rect 673898 576141 673904 576153
rect 676240 576141 676246 576153
rect 673898 576113 676246 576141
rect 673898 576101 673904 576113
rect 676240 576101 676246 576113
rect 676298 576101 676304 576153
rect 670576 575879 670582 575931
rect 670634 575919 670640 575931
rect 676048 575919 676054 575931
rect 670634 575891 676054 575919
rect 670634 575879 670640 575891
rect 676048 575879 676054 575891
rect 676106 575879 676112 575931
rect 672208 575435 672214 575487
rect 672266 575475 672272 575487
rect 676048 575475 676054 575487
rect 672266 575447 676054 575475
rect 672266 575435 672272 575447
rect 676048 575435 676054 575447
rect 676106 575435 676112 575487
rect 670480 574917 670486 574969
rect 670538 574957 670544 574969
rect 676048 574957 676054 574969
rect 670538 574929 676054 574957
rect 670538 574917 670544 574929
rect 676048 574917 676054 574929
rect 676106 574917 676112 574969
rect 42160 574621 42166 574673
rect 42218 574661 42224 574673
rect 43024 574661 43030 574673
rect 42218 574633 43030 574661
rect 42218 574621 42224 574633
rect 43024 574621 43030 574633
rect 43082 574621 43088 574673
rect 672304 574325 672310 574377
rect 672362 574365 672368 574377
rect 676048 574365 676054 574377
rect 672362 574337 676054 574365
rect 672362 574325 672368 574337
rect 676048 574325 676054 574337
rect 676106 574325 676112 574377
rect 42160 574103 42166 574155
rect 42218 574143 42224 574155
rect 43120 574143 43126 574155
rect 42218 574115 43126 574143
rect 42218 574103 42224 574115
rect 43120 574103 43126 574115
rect 43178 574103 43184 574155
rect 42064 573437 42070 573489
rect 42122 573477 42128 573489
rect 42544 573477 42550 573489
rect 42122 573449 42550 573477
rect 42122 573437 42128 573449
rect 42544 573437 42550 573449
rect 42602 573437 42608 573489
rect 669904 573215 669910 573267
rect 669962 573255 669968 573267
rect 670480 573255 670486 573267
rect 669962 573227 670486 573255
rect 669962 573215 669968 573227
rect 670480 573215 670486 573227
rect 670538 573215 670544 573267
rect 42928 573141 42934 573193
rect 42986 573181 42992 573193
rect 58192 573181 58198 573193
rect 42986 573153 58198 573181
rect 42986 573141 42992 573153
rect 58192 573141 58198 573153
rect 58250 573141 58256 573193
rect 670096 573141 670102 573193
rect 670154 573181 670160 573193
rect 670576 573181 670582 573193
rect 670154 573153 670582 573181
rect 670154 573141 670160 573153
rect 670576 573141 670582 573153
rect 670634 573141 670640 573193
rect 47920 573067 47926 573119
rect 47978 573107 47984 573119
rect 58960 573107 58966 573119
rect 47978 573079 58966 573107
rect 47978 573067 47984 573079
rect 58960 573067 58966 573079
rect 59018 573067 59024 573119
rect 48016 572993 48022 573045
rect 48074 573033 48080 573045
rect 59632 573033 59638 573045
rect 48074 573005 59638 573033
rect 48074 572993 48080 573005
rect 59632 572993 59638 573005
rect 59690 572993 59696 573045
rect 42352 572105 42358 572157
rect 42410 572145 42416 572157
rect 42832 572145 42838 572157
rect 42410 572117 42838 572145
rect 42410 572105 42416 572117
rect 42832 572105 42838 572117
rect 42890 572105 42896 572157
rect 42160 570995 42166 571047
rect 42218 571035 42224 571047
rect 43024 571035 43030 571047
rect 42218 571007 43030 571035
rect 42218 570995 42224 571007
rect 43024 570995 43030 571007
rect 43082 570995 43088 571047
rect 42832 570847 42838 570899
rect 42890 570887 42896 570899
rect 43024 570887 43030 570899
rect 42890 570859 43030 570887
rect 42890 570847 42896 570859
rect 43024 570847 43030 570859
rect 43082 570847 43088 570899
rect 670864 570625 670870 570677
rect 670922 570665 670928 570677
rect 676240 570665 676246 570677
rect 670922 570637 676246 570665
rect 670922 570625 670928 570637
rect 676240 570625 676246 570637
rect 676298 570625 676304 570677
rect 42160 570403 42166 570455
rect 42218 570443 42224 570455
rect 43120 570443 43126 570455
rect 42218 570415 43126 570443
rect 42218 570403 42224 570415
rect 43120 570403 43126 570415
rect 43178 570403 43184 570455
rect 50320 570181 50326 570233
rect 50378 570221 50384 570233
rect 59344 570221 59350 570233
rect 50378 570193 59350 570221
rect 50378 570181 50384 570193
rect 59344 570181 59350 570193
rect 59402 570181 59408 570233
rect 47824 570107 47830 570159
rect 47882 570147 47888 570159
rect 59536 570147 59542 570159
rect 47882 570119 59542 570147
rect 47882 570107 47888 570119
rect 59536 570107 59542 570119
rect 59594 570107 59600 570159
rect 672400 569885 672406 569937
rect 672458 569925 672464 569937
rect 676048 569925 676054 569937
rect 672458 569897 676054 569925
rect 672458 569885 672464 569897
rect 676048 569885 676054 569897
rect 676106 569885 676112 569937
rect 42064 569737 42070 569789
rect 42122 569777 42128 569789
rect 43024 569777 43030 569789
rect 42122 569749 43030 569777
rect 42122 569737 42128 569749
rect 43024 569737 43030 569749
rect 43082 569737 43088 569789
rect 670672 569515 670678 569567
rect 670730 569555 670736 569567
rect 676048 569555 676054 569567
rect 670730 569527 676054 569555
rect 670730 569515 670736 569527
rect 676048 569515 676054 569527
rect 676106 569515 676112 569567
rect 42160 569145 42166 569197
rect 42218 569185 42224 569197
rect 42928 569185 42934 569197
rect 42218 569157 42934 569185
rect 42218 569145 42224 569157
rect 42928 569145 42934 569157
rect 42986 569145 42992 569197
rect 672784 569145 672790 569197
rect 672842 569185 672848 569197
rect 676240 569185 676246 569197
rect 672842 569157 676246 569185
rect 672842 569145 672848 569157
rect 676240 569145 676246 569157
rect 676298 569145 676304 569197
rect 673360 568405 673366 568457
rect 673418 568445 673424 568457
rect 676048 568445 676054 568457
rect 673418 568417 676054 568445
rect 673418 568405 673424 568417
rect 676048 568405 676054 568417
rect 676106 568405 676112 568457
rect 672880 567961 672886 568013
rect 672938 568001 672944 568013
rect 676048 568001 676054 568013
rect 672938 567973 676054 568001
rect 672938 567961 672944 567973
rect 676048 567961 676054 567973
rect 676106 567961 676112 568013
rect 672688 567665 672694 567717
rect 672746 567705 672752 567717
rect 676240 567705 676246 567717
rect 672746 567677 676246 567705
rect 672746 567665 672752 567677
rect 676240 567665 676246 567677
rect 676298 567665 676304 567717
rect 655696 567443 655702 567495
rect 655754 567483 655760 567495
rect 675376 567483 675382 567495
rect 655754 567455 675382 567483
rect 655754 567443 655760 567455
rect 675376 567443 675382 567455
rect 675434 567443 675440 567495
rect 649840 564483 649846 564535
rect 649898 564523 649904 564535
rect 679792 564523 679798 564535
rect 649898 564495 679798 564523
rect 649898 564483 649904 564495
rect 679792 564483 679798 564495
rect 679850 564483 679856 564535
rect 674416 559525 674422 559577
rect 674474 559565 674480 559577
rect 675376 559565 675382 559577
rect 674474 559537 675382 559565
rect 674474 559525 674480 559537
rect 675376 559525 675382 559537
rect 675434 559525 675440 559577
rect 656560 558785 656566 558837
rect 656618 558825 656624 558837
rect 674992 558825 674998 558837
rect 656618 558797 674998 558825
rect 656618 558785 656624 558797
rect 674992 558785 674998 558797
rect 675050 558785 675056 558837
rect 674512 558045 674518 558097
rect 674570 558085 674576 558097
rect 675376 558085 675382 558097
rect 674570 558057 675382 558085
rect 674570 558045 674576 558057
rect 675376 558045 675382 558057
rect 675434 558045 675440 558097
rect 672784 556047 672790 556099
rect 672842 556087 672848 556099
rect 675280 556087 675286 556099
rect 672842 556059 675286 556087
rect 672842 556047 672848 556059
rect 675280 556047 675286 556059
rect 675338 556047 675344 556099
rect 654160 555899 654166 555951
rect 654218 555939 654224 555951
rect 675280 555939 675286 555951
rect 654218 555911 675286 555939
rect 654218 555899 654224 555911
rect 675280 555899 675286 555911
rect 675338 555899 675344 555951
rect 674128 555011 674134 555063
rect 674186 555051 674192 555063
rect 675472 555051 675478 555063
rect 674186 555023 675478 555051
rect 674186 555011 674192 555023
rect 675472 555011 675478 555023
rect 675530 555011 675536 555063
rect 673360 554345 673366 554397
rect 673418 554385 673424 554397
rect 675376 554385 675382 554397
rect 673418 554357 675382 554385
rect 673418 554345 673424 554357
rect 675376 554345 675382 554357
rect 675434 554345 675440 554397
rect 672688 553901 672694 553953
rect 672746 553941 672752 553953
rect 675472 553941 675478 553953
rect 672746 553913 675478 553941
rect 672746 553901 672752 553913
rect 675472 553901 675478 553913
rect 675530 553901 675536 553953
rect 674992 553457 674998 553509
rect 675050 553497 675056 553509
rect 675376 553497 675382 553509
rect 675050 553469 675382 553497
rect 675050 553457 675056 553469
rect 675376 553457 675382 553469
rect 675434 553457 675440 553509
rect 673744 553309 673750 553361
rect 673802 553349 673808 553361
rect 675472 553349 675478 553361
rect 673802 553321 675478 553349
rect 673802 553309 673808 553321
rect 675472 553309 675478 553321
rect 675530 553309 675536 553361
rect 672880 551903 672886 551955
rect 672938 551943 672944 551955
rect 675472 551943 675478 551955
rect 672938 551915 675478 551943
rect 672938 551903 672944 551915
rect 675472 551903 675478 551915
rect 675530 551903 675536 551955
rect 674320 548869 674326 548921
rect 674378 548909 674384 548921
rect 675280 548909 675286 548921
rect 674378 548881 675286 548909
rect 674378 548869 674384 548881
rect 675280 548869 675286 548881
rect 675338 548869 675344 548921
rect 674224 548203 674230 548255
rect 674282 548243 674288 548255
rect 675280 548243 675286 548255
rect 674282 548215 675286 548243
rect 674282 548203 674288 548215
rect 675280 548203 675286 548215
rect 675338 548203 675344 548255
rect 43024 541543 43030 541595
rect 43082 541583 43088 541595
rect 57712 541583 57718 541595
rect 43082 541555 57718 541583
rect 43082 541543 43088 541555
rect 57712 541543 57718 541555
rect 57770 541543 57776 541595
rect 42928 541469 42934 541521
rect 42986 541509 42992 541521
rect 57616 541509 57622 541521
rect 42986 541481 57622 541509
rect 42986 541469 42992 541481
rect 57616 541469 57622 541481
rect 57674 541469 57680 541521
rect 42160 538139 42166 538191
rect 42218 538179 42224 538191
rect 43024 538179 43030 538191
rect 42218 538151 43030 538179
rect 42218 538139 42224 538151
rect 43024 538139 43030 538151
rect 43082 538139 43088 538191
rect 42160 536437 42166 536489
rect 42218 536477 42224 536489
rect 42928 536477 42934 536489
rect 42218 536449 42934 536477
rect 42218 536437 42224 536449
rect 42928 536437 42934 536449
rect 42986 536437 42992 536489
rect 673840 533773 673846 533825
rect 673898 533813 673904 533825
rect 675952 533813 675958 533825
rect 673898 533785 675958 533813
rect 673898 533773 673904 533785
rect 675952 533773 675958 533785
rect 676010 533773 676016 533825
rect 655600 533255 655606 533307
rect 655658 533295 655664 533307
rect 676048 533295 676054 533307
rect 655658 533267 676054 533295
rect 655658 533255 655664 533267
rect 676048 533255 676054 533267
rect 676106 533255 676112 533307
rect 655408 533107 655414 533159
rect 655466 533147 655472 533159
rect 676144 533147 676150 533159
rect 655466 533119 676150 533147
rect 655466 533107 655472 533119
rect 676144 533107 676150 533119
rect 676202 533107 676208 533159
rect 655216 532959 655222 533011
rect 655274 532999 655280 533011
rect 676240 532999 676246 533011
rect 655274 532971 676246 532999
rect 655274 532959 655280 532971
rect 676240 532959 676246 532971
rect 676298 532959 676304 533011
rect 672208 532663 672214 532715
rect 672266 532703 672272 532715
rect 672400 532703 672406 532715
rect 672266 532675 672406 532703
rect 672266 532663 672272 532675
rect 672400 532663 672406 532675
rect 672458 532703 672464 532715
rect 676048 532703 676054 532715
rect 672458 532675 676054 532703
rect 672458 532663 672464 532675
rect 676048 532663 676054 532675
rect 676106 532663 676112 532715
rect 672304 531479 672310 531531
rect 672362 531519 672368 531531
rect 676240 531519 676246 531531
rect 672362 531491 676246 531519
rect 672362 531479 672368 531491
rect 676240 531479 676246 531491
rect 676298 531479 676304 531531
rect 42928 529925 42934 529977
rect 42986 529965 42992 529977
rect 58192 529965 58198 529977
rect 42986 529937 58198 529965
rect 42986 529925 42992 529937
rect 58192 529925 58198 529937
rect 58250 529925 58256 529977
rect 670960 528001 670966 528053
rect 671018 528041 671024 528053
rect 676240 528041 676246 528053
rect 671018 528013 676246 528041
rect 671018 528001 671024 528013
rect 676240 528001 676246 528013
rect 676298 528001 676304 528053
rect 670768 527409 670774 527461
rect 670826 527449 670832 527461
rect 676240 527449 676246 527461
rect 670826 527421 676246 527449
rect 670826 527409 670832 527421
rect 676240 527409 676246 527421
rect 676298 527409 676304 527461
rect 673168 526669 673174 526721
rect 673226 526709 673232 526721
rect 676048 526709 676054 526721
rect 673226 526681 676054 526709
rect 673226 526669 673232 526681
rect 676048 526669 676054 526681
rect 676106 526669 676112 526721
rect 42160 526373 42166 526425
rect 42218 526413 42224 526425
rect 42544 526413 42550 526425
rect 42218 526385 42550 526413
rect 42218 526373 42224 526385
rect 42544 526373 42550 526385
rect 42602 526373 42608 526425
rect 672496 526299 672502 526351
rect 672554 526339 672560 526351
rect 676048 526339 676054 526351
rect 672554 526311 676054 526339
rect 672554 526299 672560 526311
rect 676048 526299 676054 526311
rect 676106 526299 676112 526351
rect 673072 525929 673078 525981
rect 673130 525969 673136 525981
rect 676240 525969 676246 525981
rect 673130 525941 676246 525969
rect 673130 525929 673136 525941
rect 676240 525929 676246 525941
rect 676298 525929 676304 525981
rect 42064 525633 42070 525685
rect 42122 525673 42128 525685
rect 42352 525673 42358 525685
rect 42122 525645 42358 525673
rect 42122 525633 42128 525645
rect 42352 525633 42358 525645
rect 42410 525633 42416 525685
rect 42160 525411 42166 525463
rect 42218 525451 42224 525463
rect 42928 525451 42934 525463
rect 42218 525423 42934 525451
rect 42218 525411 42224 525423
rect 42928 525411 42934 525423
rect 42986 525411 42992 525463
rect 673264 525189 673270 525241
rect 673322 525229 673328 525241
rect 676048 525229 676054 525241
rect 673322 525201 676054 525229
rect 673322 525189 673328 525201
rect 676048 525189 676054 525201
rect 676106 525189 676112 525241
rect 672976 524819 672982 524871
rect 673034 524859 673040 524871
rect 676048 524859 676054 524871
rect 673034 524831 676054 524859
rect 673034 524819 673040 524831
rect 676048 524819 676054 524831
rect 676106 524819 676112 524871
rect 672592 524449 672598 524501
rect 672650 524489 672656 524501
rect 676240 524489 676246 524501
rect 672650 524461 676246 524489
rect 672650 524449 672656 524461
rect 676240 524449 676246 524461
rect 676298 524449 676304 524501
rect 50320 524301 50326 524353
rect 50378 524341 50384 524353
rect 58576 524341 58582 524353
rect 50378 524313 58582 524341
rect 50378 524301 50384 524313
rect 58576 524301 58582 524313
rect 58634 524301 58640 524353
rect 47824 524227 47830 524279
rect 47882 524267 47888 524279
rect 59344 524267 59350 524279
rect 47882 524239 59350 524267
rect 47882 524227 47888 524239
rect 59344 524227 59350 524239
rect 59402 524227 59408 524279
rect 649936 521267 649942 521319
rect 649994 521307 650000 521319
rect 679792 521307 679798 521319
rect 649994 521279 679798 521307
rect 649994 521267 650000 521279
rect 679792 521267 679798 521279
rect 679850 521267 679856 521319
rect 676528 498253 676534 498305
rect 676586 498293 676592 498305
rect 679696 498293 679702 498305
rect 676586 498265 679702 498293
rect 676586 498253 676592 498265
rect 679696 498253 679702 498265
rect 679754 498253 679760 498305
rect 655504 490039 655510 490091
rect 655562 490079 655568 490091
rect 676240 490079 676246 490091
rect 655562 490051 676246 490079
rect 655562 490039 655568 490051
rect 676240 490039 676246 490051
rect 676298 490039 676304 490091
rect 655312 489891 655318 489943
rect 655370 489931 655376 489943
rect 676240 489931 676246 489943
rect 655370 489903 676246 489931
rect 655370 489891 655376 489903
rect 676240 489891 676246 489903
rect 676298 489891 676304 489943
rect 655120 489743 655126 489795
rect 655178 489783 655184 489795
rect 676144 489783 676150 489795
rect 655178 489755 676150 489783
rect 655178 489743 655184 489755
rect 676144 489743 676150 489755
rect 676202 489743 676208 489795
rect 676240 489225 676246 489277
rect 676298 489265 676304 489277
rect 676720 489265 676726 489277
rect 676298 489237 676726 489265
rect 676298 489225 676304 489237
rect 676720 489225 676726 489237
rect 676778 489225 676784 489277
rect 670288 488115 670294 488167
rect 670346 488155 670352 488167
rect 676048 488155 676054 488167
rect 670346 488127 676054 488155
rect 670346 488115 670352 488127
rect 676048 488115 676054 488127
rect 676106 488155 676112 488167
rect 676624 488155 676630 488167
rect 676106 488127 676630 488155
rect 676106 488115 676112 488127
rect 676624 488115 676630 488127
rect 676682 488115 676688 488167
rect 670000 487079 670006 487131
rect 670058 487119 670064 487131
rect 676240 487119 676246 487131
rect 670058 487091 676246 487119
rect 670058 487079 670064 487091
rect 676240 487079 676246 487091
rect 676298 487079 676304 487131
rect 674320 486635 674326 486687
rect 674378 486675 674384 486687
rect 676048 486675 676054 486687
rect 674378 486647 676054 486675
rect 674378 486635 674384 486647
rect 676048 486635 676054 486647
rect 676106 486635 676112 486687
rect 674416 486561 674422 486613
rect 674474 486601 674480 486613
rect 676240 486601 676246 486613
rect 674474 486573 676246 486601
rect 674474 486561 674480 486573
rect 676240 486561 676246 486573
rect 676298 486561 676304 486613
rect 674128 485673 674134 485725
rect 674186 485713 674192 485725
rect 676048 485713 676054 485725
rect 674186 485685 676054 485713
rect 674186 485673 674192 485685
rect 676048 485673 676054 485685
rect 676106 485673 676112 485725
rect 674512 483749 674518 483801
rect 674570 483789 674576 483801
rect 676048 483789 676054 483801
rect 674570 483761 676054 483789
rect 674570 483749 674576 483761
rect 676048 483749 676054 483761
rect 676106 483749 676112 483801
rect 674224 483675 674230 483727
rect 674282 483715 674288 483727
rect 675952 483715 675958 483727
rect 674282 483687 675958 483715
rect 674282 483675 674288 483687
rect 675952 483675 675958 483687
rect 676010 483675 676016 483727
rect 672880 481899 672886 481951
rect 672938 481939 672944 481951
rect 676048 481939 676054 481951
rect 672938 481911 676054 481939
rect 672938 481899 672944 481911
rect 676048 481899 676054 481911
rect 676106 481899 676112 481951
rect 672688 481529 672694 481581
rect 672746 481569 672752 481581
rect 676240 481569 676246 481581
rect 672746 481541 676246 481569
rect 672746 481529 672752 481541
rect 676240 481529 676246 481541
rect 676298 481529 676304 481581
rect 672784 480789 672790 480841
rect 672842 480829 672848 480841
rect 676048 480829 676054 480841
rect 672842 480801 676054 480829
rect 672842 480789 672848 480801
rect 676048 480789 676054 480801
rect 676106 480789 676112 480841
rect 673360 480419 673366 480471
rect 673418 480459 673424 480471
rect 676048 480459 676054 480471
rect 673418 480431 676054 480459
rect 673418 480419 673424 480431
rect 676048 480419 676054 480431
rect 676106 480419 676112 480471
rect 673744 480049 673750 480101
rect 673802 480089 673808 480101
rect 676240 480089 676246 480101
rect 673802 480061 676246 480089
rect 673802 480049 673808 480061
rect 676240 480049 676246 480061
rect 676298 480049 676304 480101
rect 650032 478125 650038 478177
rect 650090 478165 650096 478177
rect 679888 478165 679894 478177
rect 650090 478137 679894 478165
rect 650090 478125 650096 478137
rect 679888 478125 679894 478137
rect 679946 478125 679952 478177
rect 41776 476053 41782 476105
rect 41834 476093 41840 476105
rect 50320 476093 50326 476105
rect 41834 476065 50326 476093
rect 41834 476053 41840 476065
rect 50320 476053 50326 476065
rect 50378 476053 50384 476105
rect 41776 475535 41782 475587
rect 41834 475575 41840 475587
rect 47824 475575 47830 475587
rect 41834 475547 47830 475575
rect 41834 475535 41840 475547
rect 47824 475535 47830 475547
rect 47882 475535 47888 475587
rect 37360 475239 37366 475291
rect 37418 475279 37424 475291
rect 42352 475279 42358 475291
rect 37418 475251 42358 475279
rect 37418 475239 37424 475251
rect 42352 475239 42358 475251
rect 42410 475239 42416 475291
rect 677776 475239 677782 475291
rect 677834 475279 677840 475291
rect 679792 475279 679798 475291
rect 677834 475251 679798 475279
rect 677834 475239 677840 475251
rect 679792 475239 679798 475251
rect 679850 475239 679856 475291
rect 41872 474573 41878 474625
rect 41930 474613 41936 474625
rect 43216 474613 43222 474625
rect 41930 474585 43222 474613
rect 41930 474573 41936 474585
rect 43216 474573 43222 474585
rect 43274 474573 43280 474625
rect 41584 472427 41590 472479
rect 41642 472467 41648 472479
rect 43504 472467 43510 472479
rect 41642 472439 43510 472467
rect 41642 472427 41648 472439
rect 43504 472427 43510 472439
rect 43562 472467 43568 472479
rect 45136 472467 45142 472479
rect 43562 472439 45142 472467
rect 43562 472427 43568 472439
rect 45136 472427 45142 472439
rect 45194 472427 45200 472479
rect 41776 472353 41782 472405
rect 41834 472393 41840 472405
rect 58960 472393 58966 472405
rect 41834 472365 58966 472393
rect 41834 472353 41840 472365
rect 58960 472353 58966 472365
rect 59018 472353 59024 472405
rect 41584 469319 41590 469371
rect 41642 469359 41648 469371
rect 42544 469359 42550 469371
rect 41642 469331 42550 469359
rect 41642 469319 41648 469331
rect 42544 469319 42550 469331
rect 42602 469319 42608 469371
rect 34480 463547 34486 463599
rect 34538 463587 34544 463599
rect 41776 463587 41782 463599
rect 34538 463559 41782 463587
rect 34538 463547 34544 463559
rect 41776 463547 41782 463559
rect 41834 463587 41840 463599
rect 47824 463587 47830 463599
rect 41834 463559 47830 463587
rect 41834 463547 41840 463559
rect 47824 463547 47830 463559
rect 47882 463547 47888 463599
rect 676624 440607 676630 440659
rect 676682 440647 676688 440659
rect 677776 440647 677782 440659
rect 676682 440619 677782 440647
rect 676682 440607 676688 440619
rect 677776 440607 677782 440619
rect 677834 440607 677840 440659
rect 23056 437795 23062 437847
rect 23114 437835 23120 437847
rect 39760 437835 39766 437847
rect 23114 437807 39766 437835
rect 23114 437795 23120 437807
rect 39760 437795 39766 437807
rect 39818 437795 39824 437847
rect 39856 437795 39862 437847
rect 39914 437835 39920 437847
rect 62320 437835 62326 437847
rect 39914 437807 62326 437835
rect 39914 437795 39920 437807
rect 62320 437795 62326 437807
rect 62378 437795 62384 437847
rect 676528 434909 676534 434961
rect 676586 434949 676592 434961
rect 677872 434949 677878 434961
rect 676586 434921 677878 434949
rect 676586 434909 676592 434921
rect 677872 434909 677878 434921
rect 677930 434909 677936 434961
rect 41584 426843 41590 426895
rect 41642 426883 41648 426895
rect 53200 426883 53206 426895
rect 41642 426855 53206 426883
rect 41642 426843 41648 426855
rect 53200 426843 53206 426855
rect 53258 426843 53264 426895
rect 41776 426473 41782 426525
rect 41834 426513 41840 426525
rect 50320 426513 50326 426525
rect 41834 426485 50326 426513
rect 41834 426473 41840 426485
rect 50320 426473 50326 426485
rect 50378 426473 50384 426525
rect 41776 425955 41782 426007
rect 41834 425995 41840 426007
rect 48016 425995 48022 426007
rect 41834 425967 48022 425995
rect 41834 425955 41840 425967
rect 48016 425955 48022 425967
rect 48074 425955 48080 426007
rect 41584 424771 41590 424823
rect 41642 424811 41648 424823
rect 43312 424811 43318 424823
rect 41642 424783 43318 424811
rect 41642 424771 41648 424783
rect 43312 424771 43318 424783
rect 43370 424771 43376 424823
rect 41776 423439 41782 423491
rect 41834 423479 41840 423491
rect 43216 423479 43222 423491
rect 41834 423451 43222 423479
rect 41834 423439 41840 423451
rect 43216 423439 43222 423451
rect 43274 423439 43280 423491
rect 23056 422699 23062 422751
rect 23114 422739 23120 422751
rect 41584 422739 41590 422751
rect 23114 422711 41590 422739
rect 23114 422699 23120 422711
rect 41584 422699 41590 422711
rect 41642 422699 41648 422751
rect 41584 420479 41590 420531
rect 41642 420519 41648 420531
rect 62512 420519 62518 420531
rect 41642 420491 62518 420519
rect 41642 420479 41648 420491
rect 62512 420479 62518 420491
rect 62570 420479 62576 420531
rect 39856 417519 39862 417571
rect 39914 417559 39920 417571
rect 41776 417559 41782 417571
rect 39914 417531 41782 417559
rect 39914 417519 39920 417531
rect 41776 417519 41782 417531
rect 41834 417519 41840 417571
rect 40144 417445 40150 417497
rect 40202 417485 40208 417497
rect 42928 417485 42934 417497
rect 40202 417457 42934 417485
rect 40202 417445 40208 417457
rect 42928 417445 42934 417457
rect 42986 417445 42992 417497
rect 41584 415151 41590 415203
rect 41642 415191 41648 415203
rect 43120 415191 43126 415203
rect 41642 415163 43126 415191
rect 41642 415151 41648 415163
rect 43120 415151 43126 415163
rect 43178 415151 43184 415203
rect 41872 414707 41878 414759
rect 41930 414747 41936 414759
rect 43024 414747 43030 414759
rect 41930 414719 43030 414747
rect 41930 414707 41936 414719
rect 43024 414707 43030 414719
rect 43082 414707 43088 414759
rect 41584 414263 41590 414315
rect 41642 414303 41648 414315
rect 47920 414303 47926 414315
rect 41642 414275 47926 414303
rect 41642 414263 41648 414275
rect 47920 414263 47926 414275
rect 47978 414263 47984 414315
rect 41776 413375 41782 413427
rect 41834 413375 41840 413427
rect 41794 413205 41822 413375
rect 41776 413153 41782 413205
rect 41834 413153 41840 413205
rect 42160 409675 42166 409727
rect 42218 409715 42224 409727
rect 42832 409715 42838 409727
rect 42218 409687 42838 409715
rect 42218 409675 42224 409687
rect 42832 409675 42838 409687
rect 42890 409675 42896 409727
rect 42160 409453 42166 409505
rect 42218 409493 42224 409505
rect 42928 409493 42934 409505
rect 42218 409465 42934 409493
rect 42218 409453 42224 409465
rect 42928 409453 42934 409465
rect 42986 409453 42992 409505
rect 42160 408195 42166 408247
rect 42218 408235 42224 408247
rect 43024 408235 43030 408247
rect 42218 408207 43030 408235
rect 42218 408195 42224 408207
rect 43024 408195 43030 408207
rect 43082 408195 43088 408247
rect 42064 407973 42070 408025
rect 42122 408013 42128 408025
rect 42832 408013 42838 408025
rect 42122 407985 42838 408013
rect 42122 407973 42128 407985
rect 42832 407973 42838 407985
rect 42890 407973 42896 408025
rect 42160 406863 42166 406915
rect 42218 406903 42224 406915
rect 43120 406903 43126 406915
rect 42218 406875 43126 406903
rect 42218 406863 42224 406875
rect 43120 406863 43126 406875
rect 43178 406863 43184 406915
rect 42928 406049 42934 406101
rect 42986 406089 42992 406101
rect 58480 406089 58486 406101
rect 42986 406061 58486 406089
rect 42986 406049 42992 406061
rect 58480 406049 58486 406061
rect 58538 406049 58544 406101
rect 42832 402571 42838 402623
rect 42890 402611 42896 402623
rect 59344 402611 59350 402623
rect 42890 402583 59350 402611
rect 42890 402571 42896 402583
rect 59344 402571 59350 402583
rect 59402 402571 59408 402623
rect 655120 400573 655126 400625
rect 655178 400613 655184 400625
rect 676144 400613 676150 400625
rect 655178 400585 676150 400613
rect 655178 400573 655184 400585
rect 676144 400573 676150 400585
rect 676202 400573 676208 400625
rect 655504 400499 655510 400551
rect 655562 400539 655568 400551
rect 676240 400539 676246 400551
rect 655562 400511 676246 400539
rect 655562 400499 655568 400511
rect 676240 400499 676246 400511
rect 676298 400499 676304 400551
rect 655312 400425 655318 400477
rect 655370 400465 655376 400477
rect 676048 400465 676054 400477
rect 655370 400437 676054 400465
rect 655370 400425 655376 400437
rect 676048 400425 676054 400437
rect 676106 400425 676112 400477
rect 673840 400351 673846 400403
rect 673898 400391 673904 400403
rect 676240 400391 676246 400403
rect 673898 400363 676246 400391
rect 673898 400351 673904 400363
rect 676240 400351 676246 400363
rect 676298 400351 676304 400403
rect 53200 400277 53206 400329
rect 53258 400317 53264 400329
rect 59728 400317 59734 400329
rect 53258 400289 59734 400317
rect 53258 400277 53264 400289
rect 59728 400277 59734 400289
rect 59786 400277 59792 400329
rect 50320 400203 50326 400255
rect 50378 400243 50384 400255
rect 59536 400243 59542 400255
rect 50378 400215 59542 400243
rect 50378 400203 50384 400215
rect 59536 400203 59542 400215
rect 59594 400203 59600 400255
rect 48016 400129 48022 400181
rect 48074 400169 48080 400181
rect 59632 400169 59638 400181
rect 48074 400141 59638 400169
rect 48074 400129 48080 400141
rect 59632 400129 59638 400141
rect 59690 400129 59696 400181
rect 670192 398871 670198 398923
rect 670250 398911 670256 398923
rect 676624 398911 676630 398923
rect 670250 398883 676630 398911
rect 670250 398871 670256 398883
rect 676624 398871 676630 398883
rect 676682 398871 676688 398923
rect 674416 398723 674422 398775
rect 674474 398763 674480 398775
rect 676048 398763 676054 398775
rect 674474 398735 676054 398763
rect 674474 398723 674480 398735
rect 676048 398723 676054 398735
rect 676106 398723 676112 398775
rect 670480 398427 670486 398479
rect 670538 398467 670544 398479
rect 676528 398467 676534 398479
rect 670538 398439 676534 398467
rect 670538 398427 670544 398439
rect 676528 398427 676534 398439
rect 676586 398427 676592 398479
rect 674512 397835 674518 397887
rect 674570 397875 674576 397887
rect 676048 397875 676054 397887
rect 674570 397847 676054 397875
rect 674570 397835 674576 397847
rect 676048 397835 676054 397847
rect 676106 397835 676112 397887
rect 673168 395541 673174 395593
rect 673226 395581 673232 395593
rect 676048 395581 676054 395593
rect 673226 395553 676054 395581
rect 673226 395541 673232 395553
rect 676048 395541 676054 395553
rect 676106 395541 676112 395593
rect 42064 394505 42070 394557
rect 42122 394545 42128 394557
rect 57712 394545 57718 394557
rect 42122 394517 57718 394545
rect 42122 394505 42128 394517
rect 57712 394505 57718 394517
rect 57770 394505 57776 394557
rect 650128 388807 650134 388859
rect 650186 388847 650192 388859
rect 679792 388847 679798 388859
rect 650186 388819 679798 388847
rect 650186 388807 650192 388819
rect 679792 388807 679798 388819
rect 679850 388807 679856 388859
rect 41584 385921 41590 385973
rect 41642 385961 41648 385973
rect 53200 385961 53206 385973
rect 41642 385933 53206 385961
rect 41642 385921 41648 385933
rect 53200 385921 53206 385933
rect 53258 385921 53264 385973
rect 673360 385847 673366 385899
rect 673418 385887 673424 385899
rect 674416 385887 674422 385899
rect 673418 385859 674422 385887
rect 673418 385847 673424 385859
rect 674416 385847 674422 385859
rect 674474 385847 674480 385899
rect 673264 385773 673270 385825
rect 673322 385813 673328 385825
rect 674512 385813 674518 385825
rect 673322 385785 674518 385813
rect 673322 385773 673328 385785
rect 674512 385773 674518 385785
rect 674570 385773 674576 385825
rect 41584 385255 41590 385307
rect 41642 385295 41648 385307
rect 50320 385295 50326 385307
rect 41642 385267 50326 385295
rect 41642 385255 41648 385267
rect 50320 385255 50326 385267
rect 50378 385255 50384 385307
rect 41872 384959 41878 385011
rect 41930 384999 41936 385011
rect 48112 384999 48118 385011
rect 41930 384971 48118 384999
rect 41930 384959 41936 384971
rect 48112 384959 48118 384971
rect 48170 384959 48176 385011
rect 41584 384737 41590 384789
rect 41642 384777 41648 384789
rect 43312 384777 43318 384789
rect 41642 384749 43318 384777
rect 41642 384737 41648 384749
rect 43312 384737 43318 384749
rect 43370 384737 43376 384789
rect 41584 383775 41590 383827
rect 41642 383815 41648 383827
rect 43408 383815 43414 383827
rect 41642 383787 43414 383815
rect 41642 383775 41648 383787
rect 43408 383775 43414 383787
rect 43466 383775 43472 383827
rect 41584 382295 41590 382347
rect 41642 382335 41648 382347
rect 43504 382335 43510 382347
rect 41642 382307 43510 382335
rect 41642 382295 41648 382307
rect 43504 382295 43510 382307
rect 43562 382295 43568 382347
rect 41776 381999 41782 382051
rect 41834 382039 41840 382051
rect 43216 382039 43222 382051
rect 41834 382011 43222 382039
rect 41834 381999 41840 382011
rect 43216 381999 43222 382011
rect 43274 382039 43280 382051
rect 45328 382039 45334 382051
rect 43274 382011 45334 382039
rect 43274 381999 43280 382011
rect 45328 381999 45334 382011
rect 45386 381999 45392 382051
rect 656560 381555 656566 381607
rect 656618 381595 656624 381607
rect 675088 381595 675094 381607
rect 656618 381567 675094 381595
rect 656618 381555 656624 381567
rect 675088 381555 675094 381567
rect 675146 381555 675152 381607
rect 39472 374303 39478 374355
rect 39530 374343 39536 374355
rect 41872 374343 41878 374355
rect 39530 374315 41878 374343
rect 39530 374303 39536 374315
rect 41872 374303 41878 374315
rect 41930 374303 41936 374355
rect 41488 374229 41494 374281
rect 41546 374269 41552 374281
rect 43024 374269 43030 374281
rect 41546 374241 43030 374269
rect 41546 374229 41552 374241
rect 43024 374229 43030 374241
rect 43082 374229 43088 374281
rect 41776 373489 41782 373541
rect 41834 373529 41840 373541
rect 48016 373529 48022 373541
rect 41834 373501 48022 373529
rect 41834 373489 41840 373501
rect 48016 373489 48022 373501
rect 48074 373489 48080 373541
rect 673168 372083 673174 372135
rect 673226 372123 673232 372135
rect 675376 372123 675382 372135
rect 673226 372095 675382 372123
rect 673226 372083 673232 372095
rect 675376 372083 675382 372095
rect 675434 372083 675440 372135
rect 41584 371935 41590 371987
rect 41642 371975 41648 371987
rect 42832 371975 42838 371987
rect 41642 371947 42838 371975
rect 41642 371935 41648 371947
rect 42832 371935 42838 371947
rect 42890 371935 42896 371987
rect 41680 371787 41686 371839
rect 41738 371827 41744 371839
rect 42928 371827 42934 371839
rect 41738 371799 42934 371827
rect 41738 371787 41744 371799
rect 42928 371787 42934 371799
rect 42986 371787 42992 371839
rect 41872 370159 41878 370211
rect 41930 370159 41936 370211
rect 41890 369989 41918 370159
rect 41872 369937 41878 369989
rect 41930 369937 41936 369989
rect 42448 366681 42454 366733
rect 42506 366681 42512 366733
rect 42466 366647 42494 366681
rect 42082 366619 42494 366647
rect 42082 366289 42110 366619
rect 42160 366533 42166 366585
rect 42218 366573 42224 366585
rect 42448 366573 42454 366585
rect 42218 366545 42454 366573
rect 42218 366533 42224 366545
rect 42448 366533 42454 366545
rect 42506 366533 42512 366585
rect 42064 366237 42070 366289
rect 42122 366237 42128 366289
rect 42160 364979 42166 365031
rect 42218 365019 42224 365031
rect 42832 365019 42838 365031
rect 42218 364991 42838 365019
rect 42218 364979 42224 364991
rect 42832 364979 42838 364991
rect 42890 364979 42896 365031
rect 42064 364683 42070 364735
rect 42122 364723 42128 364735
rect 42832 364723 42838 364735
rect 42122 364695 42838 364723
rect 42122 364683 42128 364695
rect 42832 364683 42838 364695
rect 42890 364683 42896 364735
rect 42064 364239 42070 364291
rect 42122 364279 42128 364291
rect 43024 364279 43030 364291
rect 42122 364251 43030 364279
rect 42122 364239 42128 364251
rect 43024 364239 43030 364251
rect 43082 364239 43088 364291
rect 42160 363795 42166 363847
rect 42218 363835 42224 363847
rect 42928 363835 42934 363847
rect 42218 363807 42934 363835
rect 42218 363795 42224 363807
rect 42928 363795 42934 363807
rect 42986 363795 42992 363847
rect 42448 361945 42454 361997
rect 42506 361985 42512 361997
rect 59248 361985 59254 361997
rect 42506 361957 59254 361985
rect 42506 361945 42512 361957
rect 59248 361945 59254 361957
rect 59306 361945 59312 361997
rect 42832 359947 42838 359999
rect 42890 359987 42896 359999
rect 59152 359987 59158 359999
rect 42890 359959 59158 359987
rect 42890 359947 42896 359959
rect 59152 359947 59158 359959
rect 59210 359947 59216 359999
rect 655312 357283 655318 357335
rect 655370 357323 655376 357335
rect 676240 357323 676246 357335
rect 655370 357295 676246 357323
rect 655370 357283 655376 357295
rect 676240 357283 676246 357295
rect 676298 357283 676304 357335
rect 655216 357209 655222 357261
rect 655274 357249 655280 357261
rect 676144 357249 676150 357261
rect 655274 357221 676150 357249
rect 655274 357209 655280 357221
rect 676144 357209 676150 357221
rect 676202 357209 676208 357261
rect 655120 357135 655126 357187
rect 655178 357175 655184 357187
rect 676336 357175 676342 357187
rect 655178 357147 676342 357175
rect 655178 357135 655184 357147
rect 676336 357135 676342 357147
rect 676394 357135 676400 357187
rect 53200 357061 53206 357113
rect 53258 357101 53264 357113
rect 58192 357101 58198 357113
rect 53258 357073 58198 357101
rect 53258 357061 53264 357073
rect 58192 357061 58198 357073
rect 58250 357061 58256 357113
rect 48112 356987 48118 357039
rect 48170 357027 48176 357039
rect 59632 357027 59638 357039
rect 48170 356999 59638 357027
rect 48170 356987 48176 356999
rect 59632 356987 59638 356999
rect 59690 356987 59696 357039
rect 50320 356913 50326 356965
rect 50378 356953 50384 356965
rect 58576 356953 58582 356965
rect 50378 356925 58582 356953
rect 50378 356913 50384 356925
rect 58576 356913 58582 356925
rect 58634 356913 58640 356965
rect 673840 356765 673846 356817
rect 673898 356805 673904 356817
rect 676048 356805 676054 356817
rect 673898 356777 676054 356805
rect 673898 356765 673904 356777
rect 676048 356765 676054 356777
rect 676106 356765 676112 356817
rect 673360 355655 673366 355707
rect 673418 355695 673424 355707
rect 676048 355695 676054 355707
rect 673418 355667 676054 355695
rect 673418 355655 673424 355667
rect 676048 355655 676054 355667
rect 676106 355655 676112 355707
rect 673264 354619 673270 354671
rect 673322 354659 673328 354671
rect 676048 354659 676054 354671
rect 673322 354631 676054 354659
rect 673322 354619 673328 354631
rect 676048 354619 676054 354631
rect 676106 354619 676112 354671
rect 672496 354323 672502 354375
rect 672554 354363 672560 354375
rect 673360 354363 673366 354375
rect 672554 354335 673366 354363
rect 672554 354323 672560 354335
rect 673360 354323 673366 354335
rect 673418 354323 673424 354375
rect 672784 354249 672790 354301
rect 672842 354289 672848 354301
rect 673264 354289 673270 354301
rect 672842 354261 673270 354289
rect 672842 354249 672848 354261
rect 673264 354249 673270 354261
rect 673322 354249 673328 354301
rect 674992 351363 674998 351415
rect 675050 351403 675056 351415
rect 676048 351403 676054 351415
rect 675050 351375 676054 351403
rect 675050 351363 675056 351375
rect 676048 351363 676054 351375
rect 676106 351363 676112 351415
rect 42160 351289 42166 351341
rect 42218 351329 42224 351341
rect 57616 351329 57622 351341
rect 42218 351301 57622 351329
rect 42218 351289 42224 351301
rect 57616 351289 57622 351301
rect 57674 351289 57680 351341
rect 675088 350327 675094 350379
rect 675146 350367 675152 350379
rect 676048 350367 676054 350379
rect 675146 350339 676054 350367
rect 675146 350327 675152 350339
rect 676048 350327 676054 350339
rect 676106 350327 676112 350379
rect 674224 348551 674230 348603
rect 674282 348591 674288 348603
rect 676240 348591 676246 348603
rect 674282 348563 676246 348591
rect 674282 348551 674288 348563
rect 676240 348551 676246 348563
rect 676298 348551 676304 348603
rect 675184 348477 675190 348529
rect 675242 348517 675248 348529
rect 676048 348517 676054 348529
rect 675242 348489 676054 348517
rect 675242 348477 675248 348489
rect 676048 348477 676054 348489
rect 676106 348477 676112 348529
rect 650224 345813 650230 345865
rect 650282 345853 650288 345865
rect 679888 345853 679894 345865
rect 650282 345825 679894 345853
rect 650282 345813 650288 345825
rect 679888 345813 679894 345825
rect 679946 345813 679952 345865
rect 674704 345739 674710 345791
rect 674762 345779 674768 345791
rect 675952 345779 675958 345791
rect 674762 345751 675958 345779
rect 674762 345739 674768 345751
rect 675952 345739 675958 345751
rect 676010 345739 676016 345791
rect 674800 345665 674806 345717
rect 674858 345705 674864 345717
rect 676048 345705 676054 345717
rect 674858 345677 676054 345705
rect 674858 345665 674864 345677
rect 676048 345665 676054 345677
rect 676106 345665 676112 345717
rect 674896 345591 674902 345643
rect 674954 345631 674960 345643
rect 676240 345631 676246 345643
rect 674954 345603 676246 345631
rect 674954 345591 674960 345603
rect 676240 345591 676246 345603
rect 676298 345591 676304 345643
rect 41776 342779 41782 342831
rect 41834 342819 41840 342831
rect 53200 342819 53206 342831
rect 41834 342791 53206 342819
rect 41834 342779 41840 342791
rect 53200 342779 53206 342791
rect 53258 342779 53264 342831
rect 41776 342261 41782 342313
rect 41834 342301 41840 342313
rect 50320 342301 50326 342313
rect 41834 342273 50326 342301
rect 41834 342261 41840 342273
rect 50320 342261 50326 342273
rect 50378 342261 50384 342313
rect 41776 341743 41782 341795
rect 41834 341783 41840 341795
rect 48112 341783 48118 341795
rect 41834 341755 48118 341783
rect 41834 341743 41840 341755
rect 48112 341743 48118 341755
rect 48170 341743 48176 341795
rect 41776 341373 41782 341425
rect 41834 341413 41840 341425
rect 43408 341413 43414 341425
rect 41834 341385 43414 341413
rect 41834 341373 41840 341385
rect 43408 341373 43414 341385
rect 43466 341373 43472 341425
rect 675472 341413 675478 341425
rect 675394 341385 675478 341413
rect 675394 340981 675422 341385
rect 675472 341373 675478 341385
rect 675530 341373 675536 341425
rect 675376 340929 675382 340981
rect 675434 340929 675440 340981
rect 41584 340559 41590 340611
rect 41642 340599 41648 340611
rect 43216 340599 43222 340611
rect 41642 340571 43222 340599
rect 41642 340559 41648 340571
rect 43216 340559 43222 340571
rect 43274 340559 43280 340611
rect 41776 340263 41782 340315
rect 41834 340303 41840 340315
rect 43312 340303 43318 340315
rect 41834 340275 43318 340303
rect 41834 340263 41840 340275
rect 43312 340263 43318 340275
rect 43370 340263 43376 340315
rect 666736 339967 666742 340019
rect 666794 340007 666800 340019
rect 675280 340007 675286 340019
rect 666794 339979 675286 340007
rect 666794 339967 666800 339979
rect 675280 339967 675286 339979
rect 675338 339967 675344 340019
rect 675088 339819 675094 339871
rect 675146 339859 675152 339871
rect 675280 339859 675286 339871
rect 675146 339831 675286 339859
rect 675146 339819 675152 339831
rect 675280 339819 675286 339831
rect 675338 339819 675344 339871
rect 41776 339449 41782 339501
rect 41834 339489 41840 339501
rect 43504 339489 43510 339501
rect 41834 339461 43510 339489
rect 41834 339449 41840 339461
rect 43504 339449 43510 339461
rect 43562 339449 43568 339501
rect 41584 339079 41590 339131
rect 41642 339119 41648 339131
rect 43408 339119 43414 339131
rect 41642 339091 43414 339119
rect 41642 339079 41648 339091
rect 43408 339079 43414 339091
rect 43466 339079 43472 339131
rect 674992 337895 674998 337947
rect 675050 337935 675056 337947
rect 675472 337935 675478 337947
rect 675050 337907 675478 337935
rect 675050 337895 675056 337907
rect 675472 337895 675478 337907
rect 675530 337895 675536 337947
rect 675184 337229 675190 337281
rect 675242 337269 675248 337281
rect 675472 337269 675478 337281
rect 675242 337241 675478 337269
rect 675242 337229 675248 337241
rect 675472 337229 675478 337241
rect 675530 337229 675536 337281
rect 674224 336563 674230 336615
rect 674282 336603 674288 336615
rect 675376 336603 675382 336615
rect 674282 336575 675382 336603
rect 674282 336563 674288 336575
rect 675376 336563 675382 336575
rect 675434 336563 675440 336615
rect 674896 336045 674902 336097
rect 674954 336085 674960 336097
rect 675376 336085 675382 336097
rect 674954 336057 675382 336085
rect 674954 336045 674960 336057
rect 675376 336045 675382 336057
rect 675434 336045 675440 336097
rect 674800 332715 674806 332767
rect 674858 332755 674864 332767
rect 675376 332755 675382 332767
rect 674858 332727 675382 332755
rect 674858 332715 674864 332727
rect 675376 332715 675382 332727
rect 675434 332715 675440 332767
rect 674704 331531 674710 331583
rect 674762 331571 674768 331583
rect 675376 331571 675382 331583
rect 674762 331543 675382 331571
rect 674762 331531 674768 331543
rect 675376 331531 675382 331543
rect 675434 331531 675440 331583
rect 41392 331161 41398 331213
rect 41450 331201 41456 331213
rect 42736 331201 42742 331213
rect 41450 331173 42742 331201
rect 41450 331161 41456 331173
rect 42736 331161 42742 331173
rect 42794 331161 42800 331213
rect 41488 331087 41494 331139
rect 41546 331127 41552 331139
rect 43024 331127 43030 331139
rect 41546 331099 43030 331127
rect 41546 331087 41552 331099
rect 43024 331087 43030 331099
rect 43082 331087 43088 331139
rect 41872 330347 41878 330399
rect 41930 330387 41936 330399
rect 45424 330387 45430 330399
rect 41930 330359 45430 330387
rect 41930 330347 41936 330359
rect 45424 330347 45430 330359
rect 45482 330347 45488 330399
rect 41584 328793 41590 328845
rect 41642 328833 41648 328845
rect 42928 328833 42934 328845
rect 41642 328805 42934 328833
rect 41642 328793 41648 328805
rect 42928 328793 42934 328805
rect 42986 328793 42992 328845
rect 654160 328275 654166 328327
rect 654218 328315 654224 328327
rect 666736 328315 666742 328327
rect 654218 328287 666742 328315
rect 654218 328275 654224 328287
rect 666736 328275 666742 328287
rect 666794 328275 666800 328327
rect 41776 327017 41782 327069
rect 41834 327017 41840 327069
rect 41794 326773 41822 327017
rect 41776 326721 41782 326773
rect 41834 326721 41840 326773
rect 42928 325759 42934 325811
rect 42986 325799 42992 325811
rect 43120 325799 43126 325811
rect 42986 325771 43126 325799
rect 42986 325759 42992 325771
rect 43120 325759 43126 325771
rect 43178 325759 43184 325811
rect 42064 323317 42070 323369
rect 42122 323357 42128 323369
rect 42448 323357 42454 323369
rect 42122 323329 42454 323357
rect 42122 323317 42128 323329
rect 42448 323317 42454 323329
rect 42506 323317 42512 323369
rect 42160 323095 42166 323147
rect 42218 323135 42224 323147
rect 43024 323135 43030 323147
rect 42218 323107 43030 323135
rect 42218 323095 42224 323107
rect 43024 323095 43030 323107
rect 43082 323095 43088 323147
rect 41968 321615 41974 321667
rect 42026 321655 42032 321667
rect 43120 321655 43126 321667
rect 42026 321627 43126 321655
rect 42026 321615 42032 321627
rect 43120 321615 43126 321627
rect 43178 321615 43184 321667
rect 42160 321467 42166 321519
rect 42218 321507 42224 321519
rect 43120 321507 43126 321519
rect 42218 321479 43126 321507
rect 42218 321467 42224 321479
rect 43120 321467 43126 321479
rect 43178 321467 43184 321519
rect 42160 321245 42166 321297
rect 42218 321285 42224 321297
rect 43024 321285 43030 321297
rect 42218 321257 43030 321285
rect 42218 321245 42224 321257
rect 43024 321245 43030 321257
rect 43082 321245 43088 321297
rect 42448 319617 42454 319669
rect 42506 319657 42512 319669
rect 58480 319657 58486 319669
rect 42506 319629 58486 319657
rect 42506 319617 42512 319629
rect 58480 319617 58486 319629
rect 58538 319617 58544 319669
rect 43120 316731 43126 316783
rect 43178 316771 43184 316783
rect 59152 316771 59158 316783
rect 43178 316743 59158 316771
rect 43178 316731 43184 316743
rect 59152 316731 59158 316743
rect 59210 316731 59216 316783
rect 53200 313845 53206 313897
rect 53258 313885 53264 313897
rect 58192 313885 58198 313897
rect 53258 313857 58198 313885
rect 53258 313845 53264 313857
rect 58192 313845 58198 313857
rect 58250 313845 58256 313897
rect 48112 313771 48118 313823
rect 48170 313811 48176 313823
rect 59632 313811 59638 313823
rect 48170 313783 59638 313811
rect 48170 313771 48176 313783
rect 59632 313771 59638 313783
rect 59690 313771 59696 313823
rect 50320 313697 50326 313749
rect 50378 313737 50384 313749
rect 59728 313737 59734 313749
rect 50378 313709 59734 313737
rect 50378 313697 50384 313709
rect 59728 313697 59734 313709
rect 59786 313697 59792 313749
rect 654256 311181 654262 311233
rect 654314 311221 654320 311233
rect 676240 311221 676246 311233
rect 654314 311193 676246 311221
rect 654314 311181 654320 311193
rect 676240 311181 676246 311193
rect 676298 311181 676304 311233
rect 654160 311107 654166 311159
rect 654218 311147 654224 311159
rect 676144 311147 676150 311159
rect 654218 311119 676150 311147
rect 654218 311107 654224 311119
rect 676144 311107 676150 311119
rect 676202 311107 676208 311159
rect 654064 311033 654070 311085
rect 654122 311073 654128 311085
rect 676336 311073 676342 311085
rect 654122 311045 676342 311073
rect 654122 311033 654128 311045
rect 676336 311033 676342 311045
rect 676394 311033 676400 311085
rect 42160 308073 42166 308125
rect 42218 308113 42224 308125
rect 59344 308113 59350 308125
rect 42218 308085 59350 308113
rect 42218 308073 42224 308085
rect 59344 308073 59350 308085
rect 59402 308073 59408 308125
rect 674512 305335 674518 305387
rect 674570 305375 674576 305387
rect 676048 305375 676054 305387
rect 674570 305347 676054 305375
rect 674570 305335 674576 305347
rect 676048 305335 676054 305347
rect 676106 305335 676112 305387
rect 675088 305261 675094 305313
rect 675146 305301 675152 305313
rect 676240 305301 676246 305313
rect 675146 305273 676246 305301
rect 675146 305261 675152 305273
rect 676240 305261 676246 305273
rect 676298 305261 676304 305313
rect 674320 302523 674326 302575
rect 674378 302563 674384 302575
rect 675952 302563 675958 302575
rect 674378 302535 675958 302563
rect 674378 302523 674384 302535
rect 675952 302523 675958 302535
rect 676010 302523 676016 302575
rect 674416 302449 674422 302501
rect 674474 302489 674480 302501
rect 676048 302489 676054 302501
rect 674474 302461 676054 302489
rect 674474 302449 674480 302461
rect 676048 302449 676054 302461
rect 676106 302449 676112 302501
rect 674704 302375 674710 302427
rect 674762 302415 674768 302427
rect 676240 302415 676246 302427
rect 674762 302387 676246 302415
rect 674762 302375 674768 302387
rect 676240 302375 676246 302387
rect 676298 302375 676304 302427
rect 43312 300895 43318 300947
rect 43370 300935 43376 300947
rect 62800 300935 62806 300947
rect 43370 300907 62806 300935
rect 43370 300895 43376 300907
rect 62800 300895 62806 300907
rect 62858 300895 62864 300947
rect 650320 299711 650326 299763
rect 650378 299751 650384 299763
rect 679984 299751 679990 299763
rect 650378 299723 679990 299751
rect 650378 299711 650384 299723
rect 679984 299711 679990 299723
rect 680042 299711 680048 299763
rect 39760 299637 39766 299689
rect 39818 299677 39824 299689
rect 43312 299677 43318 299689
rect 39818 299649 43318 299677
rect 39818 299637 39824 299649
rect 43312 299637 43318 299649
rect 43370 299637 43376 299689
rect 674896 299637 674902 299689
rect 674954 299677 674960 299689
rect 676240 299677 676246 299689
rect 674954 299649 676246 299677
rect 674954 299637 674960 299649
rect 676240 299637 676246 299649
rect 676298 299637 676304 299689
rect 41776 299563 41782 299615
rect 41834 299603 41840 299615
rect 60208 299603 60214 299615
rect 41834 299575 60214 299603
rect 41834 299563 41840 299575
rect 60208 299563 60214 299575
rect 60266 299563 60272 299615
rect 674992 299563 674998 299615
rect 675050 299603 675056 299615
rect 676048 299603 676054 299615
rect 675050 299575 676054 299603
rect 675050 299563 675056 299575
rect 676048 299563 676054 299575
rect 676106 299563 676112 299615
rect 41776 299119 41782 299171
rect 41834 299159 41840 299171
rect 51760 299159 51766 299171
rect 41834 299131 51766 299159
rect 41834 299119 41840 299131
rect 51760 299119 51766 299131
rect 51818 299119 51824 299171
rect 41776 298157 41782 298209
rect 41834 298197 41840 298209
rect 43216 298197 43222 298209
rect 41834 298169 43222 298197
rect 41834 298157 41840 298169
rect 43216 298157 43222 298169
rect 43274 298157 43280 298209
rect 43504 298083 43510 298135
rect 43562 298123 43568 298135
rect 62992 298123 62998 298135
rect 43562 298095 62998 298123
rect 43562 298083 43568 298095
rect 62992 298083 62998 298095
rect 63050 298083 63056 298135
rect 41776 297565 41782 297617
rect 41834 297605 41840 297617
rect 43408 297605 43414 297617
rect 41834 297577 43414 297605
rect 41834 297565 41840 297577
rect 43408 297565 43414 297577
rect 43466 297565 43472 297617
rect 41776 297047 41782 297099
rect 41834 297087 41840 297099
rect 43312 297087 43318 297099
rect 41834 297059 43318 297087
rect 41834 297047 41840 297059
rect 43312 297047 43318 297059
rect 43370 297047 43376 297099
rect 39952 296677 39958 296729
rect 40010 296717 40016 296729
rect 43504 296717 43510 296729
rect 40010 296689 43510 296717
rect 40010 296677 40016 296689
rect 43504 296677 43510 296689
rect 43562 296677 43568 296729
rect 41584 295863 41590 295915
rect 41642 295903 41648 295915
rect 43216 295903 43222 295915
rect 41642 295875 43222 295903
rect 41642 295863 41648 295875
rect 43216 295863 43222 295875
rect 43274 295863 43280 295915
rect 674800 295641 674806 295693
rect 674858 295681 674864 295693
rect 675184 295681 675190 295693
rect 674858 295653 675190 295681
rect 674858 295641 674864 295653
rect 675184 295641 675190 295653
rect 675242 295641 675248 295693
rect 674704 295419 674710 295471
rect 674762 295459 674768 295471
rect 675280 295459 675286 295471
rect 674762 295431 675286 295459
rect 674762 295419 674768 295431
rect 675280 295419 675286 295431
rect 675338 295419 675344 295471
rect 674512 294531 674518 294583
rect 674570 294571 674576 294583
rect 675376 294571 675382 294583
rect 674570 294543 675382 294571
rect 674570 294531 674576 294543
rect 675376 294531 675382 294543
rect 675434 294531 675440 294583
rect 53296 293865 53302 293917
rect 53354 293905 53360 293917
rect 59632 293905 59638 293917
rect 53354 293877 59638 293905
rect 53354 293865 53360 293877
rect 59632 293865 59638 293877
rect 59690 293865 59696 293917
rect 56272 293791 56278 293843
rect 56330 293831 56336 293843
rect 60304 293831 60310 293843
rect 56330 293803 60310 293831
rect 56330 293791 56336 293803
rect 60304 293791 60310 293803
rect 60362 293791 60368 293843
rect 39664 293717 39670 293769
rect 39722 293757 39728 293769
rect 58768 293757 58774 293769
rect 39722 293729 58774 293757
rect 39722 293717 39728 293729
rect 58768 293717 58774 293729
rect 58826 293717 58832 293769
rect 674416 292015 674422 292067
rect 674474 292055 674480 292067
rect 675472 292055 675478 292067
rect 674474 292027 675478 292055
rect 674474 292015 674480 292027
rect 675472 292015 675478 292027
rect 675530 292015 675536 292067
rect 674320 291571 674326 291623
rect 674378 291611 674384 291623
rect 675376 291611 675382 291623
rect 674378 291583 675382 291611
rect 674378 291571 674384 291583
rect 675376 291571 675382 291583
rect 675434 291571 675440 291623
rect 48208 290905 48214 290957
rect 48266 290945 48272 290957
rect 58384 290945 58390 290957
rect 48266 290917 58390 290945
rect 48266 290905 48272 290917
rect 58384 290905 58390 290917
rect 58442 290905 58448 290957
rect 656560 290831 656566 290883
rect 656618 290871 656624 290883
rect 674800 290871 674806 290883
rect 656618 290843 674806 290871
rect 656618 290831 656624 290843
rect 674800 290831 674806 290843
rect 674858 290831 674864 290883
rect 51760 289499 51766 289551
rect 51818 289539 51824 289551
rect 58000 289539 58006 289551
rect 51818 289511 58006 289539
rect 51818 289499 51824 289511
rect 58000 289499 58006 289511
rect 58058 289499 58064 289551
rect 50320 288019 50326 288071
rect 50378 288059 50384 288071
rect 59632 288059 59638 288071
rect 50378 288031 59638 288059
rect 50378 288019 50384 288031
rect 59632 288019 59638 288031
rect 59690 288019 59696 288071
rect 674992 287723 674998 287775
rect 675050 287763 675056 287775
rect 675376 287763 675382 287775
rect 675050 287735 675382 287763
rect 675050 287723 675056 287735
rect 675376 287723 675382 287735
rect 675434 287723 675440 287775
rect 41872 287131 41878 287183
rect 41930 287171 41936 287183
rect 45808 287171 45814 287183
rect 41930 287143 45814 287171
rect 41930 287131 41936 287143
rect 45808 287131 45814 287143
rect 45866 287131 45872 287183
rect 674896 286761 674902 286813
rect 674954 286801 674960 286813
rect 675376 286801 675382 286813
rect 674954 286773 675382 286801
rect 674954 286761 674960 286773
rect 675376 286761 675382 286773
rect 675434 286761 675440 286813
rect 41488 285281 41494 285333
rect 41546 285321 41552 285333
rect 43120 285321 43126 285333
rect 41546 285293 43126 285321
rect 41546 285281 41552 285293
rect 43120 285281 43126 285293
rect 43178 285281 43184 285333
rect 41680 285207 41686 285259
rect 41738 285247 41744 285259
rect 43024 285247 43030 285259
rect 41738 285219 43030 285247
rect 41738 285207 41744 285219
rect 43024 285207 43030 285219
rect 43082 285207 43088 285259
rect 41584 285133 41590 285185
rect 41642 285173 41648 285185
rect 42928 285173 42934 285185
rect 41642 285145 42934 285173
rect 41642 285133 41648 285145
rect 42928 285133 42934 285145
rect 42986 285133 42992 285185
rect 53200 285133 53206 285185
rect 53258 285173 53264 285185
rect 58960 285173 58966 285185
rect 53258 285145 58966 285173
rect 53258 285133 53264 285145
rect 58960 285133 58966 285145
rect 59018 285133 59024 285185
rect 653776 284245 653782 284297
rect 653834 284285 653840 284297
rect 658000 284285 658006 284297
rect 653834 284257 658006 284285
rect 653834 284245 653840 284257
rect 658000 284245 658006 284257
rect 658058 284245 658064 284297
rect 41776 283801 41782 283853
rect 41834 283801 41840 283853
rect 41794 283557 41822 283801
rect 41776 283505 41782 283557
rect 41834 283505 41840 283557
rect 48112 282543 48118 282595
rect 48170 282583 48176 282595
rect 59632 282583 59638 282595
rect 48170 282555 59638 282583
rect 48170 282543 48176 282555
rect 59632 282543 59638 282555
rect 59690 282543 59696 282595
rect 45520 282321 45526 282373
rect 45578 282361 45584 282373
rect 58960 282361 58966 282373
rect 45578 282333 58966 282361
rect 45578 282321 45584 282333
rect 58960 282321 58966 282333
rect 59018 282321 59024 282373
rect 56176 282247 56182 282299
rect 56234 282287 56240 282299
rect 57616 282287 57622 282299
rect 56234 282259 57622 282287
rect 56234 282247 56240 282259
rect 57616 282247 57622 282259
rect 57674 282247 57680 282299
rect 42064 280101 42070 280153
rect 42122 280141 42128 280153
rect 42832 280141 42838 280153
rect 42122 280113 42838 280141
rect 42122 280101 42128 280113
rect 42832 280101 42838 280113
rect 42890 280101 42896 280153
rect 42160 279879 42166 279931
rect 42218 279919 42224 279931
rect 43120 279919 43126 279931
rect 42218 279891 43126 279919
rect 42218 279879 42224 279891
rect 43120 279879 43126 279891
rect 43178 279879 43184 279931
rect 45712 279435 45718 279487
rect 45770 279475 45776 279487
rect 59536 279475 59542 279487
rect 45770 279447 59542 279475
rect 45770 279435 45776 279447
rect 59536 279435 59542 279447
rect 59594 279435 59600 279487
rect 654160 279435 654166 279487
rect 654218 279475 654224 279487
rect 663760 279475 663766 279487
rect 654218 279447 663766 279475
rect 654218 279435 654224 279447
rect 663760 279435 663766 279447
rect 663818 279435 663824 279487
rect 45616 279361 45622 279413
rect 45674 279401 45680 279413
rect 59344 279401 59350 279413
rect 45674 279373 59350 279401
rect 45674 279361 45680 279373
rect 59344 279361 59350 279373
rect 59402 279361 59408 279413
rect 42160 278547 42166 278599
rect 42218 278587 42224 278599
rect 42928 278587 42934 278599
rect 42218 278559 42934 278587
rect 42218 278547 42224 278559
rect 42928 278547 42934 278559
rect 42986 278547 42992 278599
rect 42064 278473 42070 278525
rect 42122 278513 42128 278525
rect 43120 278513 43126 278525
rect 42122 278485 43126 278513
rect 42122 278473 42128 278485
rect 43120 278473 43126 278485
rect 43178 278473 43184 278525
rect 314896 278251 314902 278303
rect 314954 278291 314960 278303
rect 408304 278291 408310 278303
rect 314954 278263 408310 278291
rect 314954 278251 314960 278263
rect 408304 278251 408310 278263
rect 408362 278251 408368 278303
rect 319504 278177 319510 278229
rect 319562 278217 319568 278229
rect 418960 278217 418966 278229
rect 319562 278189 418966 278217
rect 319562 278177 319568 278189
rect 418960 278177 418966 278189
rect 419018 278177 419024 278229
rect 316624 278103 316630 278155
rect 316682 278143 316688 278155
rect 411856 278143 411862 278155
rect 316682 278115 411862 278143
rect 316682 278103 316688 278115
rect 411856 278103 411862 278115
rect 411914 278103 411920 278155
rect 317872 278029 317878 278081
rect 317930 278069 317936 278081
rect 415408 278069 415414 278081
rect 317930 278041 415414 278069
rect 317930 278029 317936 278041
rect 415408 278029 415414 278041
rect 415466 278029 415472 278081
rect 322096 277955 322102 278007
rect 322154 277995 322160 278007
rect 426256 277995 426262 278007
rect 322154 277967 426262 277995
rect 322154 277955 322160 277967
rect 426256 277955 426262 277967
rect 426314 277955 426320 278007
rect 382288 277881 382294 277933
rect 382346 277921 382352 277933
rect 574960 277921 574966 277933
rect 382346 277893 574966 277921
rect 382346 277881 382352 277893
rect 574960 277881 574966 277893
rect 575018 277881 575024 277933
rect 326416 277807 326422 277859
rect 326474 277847 326480 277859
rect 437008 277847 437014 277859
rect 326474 277819 437014 277847
rect 326474 277807 326480 277819
rect 437008 277807 437014 277819
rect 437066 277807 437072 277859
rect 323824 277733 323830 277785
rect 323882 277773 323888 277785
rect 429904 277773 429910 277785
rect 323882 277745 429910 277773
rect 323882 277733 323888 277745
rect 429904 277733 429910 277745
rect 429962 277733 429968 277785
rect 329296 277659 329302 277711
rect 329354 277699 329360 277711
rect 444112 277699 444118 277711
rect 329354 277671 444118 277699
rect 329354 277659 329360 277671
rect 444112 277659 444118 277671
rect 444170 277659 444176 277711
rect 332368 277585 332374 277637
rect 332426 277625 332432 277637
rect 451216 277625 451222 277637
rect 332426 277597 451222 277625
rect 332426 277585 332432 277597
rect 451216 277585 451222 277597
rect 451274 277585 451280 277637
rect 334960 277511 334966 277563
rect 335018 277551 335024 277563
rect 458224 277551 458230 277563
rect 335018 277523 458230 277551
rect 335018 277511 335024 277523
rect 458224 277511 458230 277523
rect 458282 277511 458288 277563
rect 337840 277437 337846 277489
rect 337898 277477 337904 277489
rect 465328 277477 465334 277489
rect 337898 277449 465334 277477
rect 337898 277437 337904 277449
rect 465328 277437 465334 277449
rect 465386 277437 465392 277489
rect 42064 277363 42070 277415
rect 42122 277403 42128 277415
rect 43024 277403 43030 277415
rect 42122 277375 43030 277403
rect 42122 277363 42128 277375
rect 43024 277363 43030 277375
rect 43082 277363 43088 277415
rect 341008 277363 341014 277415
rect 341066 277403 341072 277415
rect 472432 277403 472438 277415
rect 341066 277375 472438 277403
rect 341066 277363 341072 277375
rect 472432 277363 472438 277375
rect 472490 277363 472496 277415
rect 343888 277289 343894 277341
rect 343946 277329 343952 277341
rect 479536 277329 479542 277341
rect 343946 277301 479542 277329
rect 343946 277289 343952 277301
rect 479536 277289 479542 277301
rect 479594 277289 479600 277341
rect 373840 277215 373846 277267
rect 373898 277255 373904 277267
rect 554032 277255 554038 277267
rect 373898 277227 554038 277255
rect 373898 277215 373904 277227
rect 554032 277215 554038 277227
rect 554090 277215 554096 277267
rect 375088 277141 375094 277193
rect 375146 277181 375152 277193
rect 557584 277181 557590 277193
rect 375146 277153 557590 277181
rect 375146 277141 375152 277153
rect 557584 277141 557590 277153
rect 557642 277141 557648 277193
rect 376816 277067 376822 277119
rect 376874 277107 376880 277119
rect 561136 277107 561142 277119
rect 376874 277079 561142 277107
rect 376874 277067 376880 277079
rect 561136 277067 561142 277079
rect 561194 277067 561200 277119
rect 377968 276993 377974 277045
rect 378026 277033 378032 277045
rect 564688 277033 564694 277045
rect 378026 277005 564694 277033
rect 378026 276993 378032 277005
rect 564688 276993 564694 277005
rect 564746 276993 564752 277045
rect 379408 276919 379414 276971
rect 379466 276959 379472 276971
rect 568240 276959 568246 276971
rect 379466 276931 568246 276959
rect 379466 276919 379472 276931
rect 568240 276919 568246 276931
rect 568298 276919 568304 276971
rect 381040 276845 381046 276897
rect 381098 276885 381104 276897
rect 571696 276885 571702 276897
rect 381098 276857 571702 276885
rect 381098 276845 381104 276857
rect 571696 276845 571702 276857
rect 571754 276845 571760 276897
rect 383632 276771 383638 276823
rect 383690 276811 383696 276823
rect 578800 276811 578806 276823
rect 383690 276783 578806 276811
rect 383690 276771 383696 276783
rect 578800 276771 578806 276783
rect 578858 276771 578864 276823
rect 320944 276697 320950 276749
rect 321002 276737 321008 276749
rect 422800 276737 422806 276749
rect 321002 276709 422806 276737
rect 321002 276697 321008 276709
rect 422800 276697 422806 276709
rect 422858 276697 422864 276749
rect 386512 276623 386518 276675
rect 386570 276663 386576 276675
rect 585904 276663 585910 276675
rect 386570 276635 585910 276663
rect 386570 276623 386576 276635
rect 585904 276623 585910 276635
rect 585962 276623 585968 276675
rect 676528 276623 676534 276675
rect 676586 276663 676592 276675
rect 679792 276663 679798 276675
rect 676586 276635 679798 276663
rect 676586 276623 676592 276635
rect 679792 276623 679798 276635
rect 679850 276623 679856 276675
rect 385360 276549 385366 276601
rect 385418 276589 385424 276601
rect 582352 276589 582358 276601
rect 385418 276561 582358 276589
rect 385418 276549 385424 276561
rect 582352 276549 582358 276561
rect 582410 276549 582416 276601
rect 392272 276475 392278 276527
rect 392330 276515 392336 276527
rect 600112 276515 600118 276527
rect 392330 276487 600118 276515
rect 392330 276475 392336 276487
rect 600112 276475 600118 276487
rect 600170 276475 600176 276527
rect 42832 276401 42838 276453
rect 42890 276441 42896 276453
rect 53296 276441 53302 276453
rect 42890 276413 53302 276441
rect 42890 276401 42896 276413
rect 53296 276401 53302 276413
rect 53354 276401 53360 276453
rect 286096 276401 286102 276453
rect 286154 276441 286160 276453
rect 336496 276441 336502 276453
rect 286154 276413 336502 276441
rect 286154 276401 286160 276413
rect 336496 276401 336502 276413
rect 336554 276401 336560 276453
rect 359152 276401 359158 276453
rect 359210 276441 359216 276453
rect 517360 276441 517366 276453
rect 359210 276413 517366 276441
rect 359210 276401 359216 276413
rect 517360 276401 517366 276413
rect 517418 276401 517424 276453
rect 287344 276327 287350 276379
rect 287402 276367 287408 276379
rect 340048 276367 340054 276379
rect 287402 276339 340054 276367
rect 287402 276327 287408 276339
rect 340048 276327 340054 276339
rect 340106 276327 340112 276379
rect 361744 276327 361750 276379
rect 361802 276367 361808 276379
rect 524464 276367 524470 276379
rect 361802 276339 524470 276367
rect 361802 276327 361808 276339
rect 524464 276327 524470 276339
rect 524522 276327 524528 276379
rect 288688 276253 288694 276305
rect 288746 276293 288752 276305
rect 343600 276293 343606 276305
rect 288746 276265 343606 276293
rect 288746 276253 288752 276265
rect 343600 276253 343606 276265
rect 343658 276253 343664 276305
rect 364624 276253 364630 276305
rect 364682 276293 364688 276305
rect 531568 276293 531574 276305
rect 364682 276265 531574 276293
rect 364682 276253 364688 276265
rect 531568 276253 531574 276265
rect 531626 276253 531632 276305
rect 290320 276179 290326 276231
rect 290378 276219 290384 276231
rect 347152 276219 347158 276231
rect 290378 276191 347158 276219
rect 290378 276179 290384 276191
rect 347152 276179 347158 276191
rect 347210 276179 347216 276231
rect 367696 276179 367702 276231
rect 367754 276219 367760 276231
rect 538672 276219 538678 276231
rect 367754 276191 538678 276219
rect 367754 276179 367760 276191
rect 538672 276179 538678 276191
rect 538730 276179 538736 276231
rect 291856 276105 291862 276157
rect 291914 276145 291920 276157
rect 350704 276145 350710 276157
rect 291914 276117 350710 276145
rect 291914 276105 291920 276117
rect 350704 276105 350710 276117
rect 350762 276105 350768 276157
rect 370288 276105 370294 276157
rect 370346 276145 370352 276157
rect 545776 276145 545782 276157
rect 370346 276117 545782 276145
rect 370346 276105 370352 276117
rect 545776 276105 545782 276117
rect 545834 276105 545840 276157
rect 293008 276031 293014 276083
rect 293066 276071 293072 276083
rect 354256 276071 354262 276083
rect 293066 276043 354262 276071
rect 293066 276031 293072 276043
rect 354256 276031 354262 276043
rect 354314 276031 354320 276083
rect 371920 276031 371926 276083
rect 371978 276071 371984 276083
rect 549328 276071 549334 276083
rect 371978 276043 549334 276071
rect 371978 276031 371984 276043
rect 549328 276031 549334 276043
rect 549386 276031 549392 276083
rect 294640 275957 294646 276009
rect 294698 275997 294704 276009
rect 357808 275997 357814 276009
rect 294698 275969 357814 275997
rect 294698 275957 294704 275969
rect 357808 275957 357814 275969
rect 357866 275957 357872 276009
rect 371056 275957 371062 276009
rect 371114 275997 371120 276009
rect 546928 275997 546934 276009
rect 371114 275969 546934 275997
rect 371114 275957 371120 275969
rect 546928 275957 546934 275969
rect 546986 275957 546992 276009
rect 295888 275883 295894 275935
rect 295946 275923 295952 275935
rect 361360 275923 361366 275935
rect 295946 275895 361366 275923
rect 295946 275883 295952 275895
rect 361360 275883 361366 275895
rect 361418 275883 361424 275935
rect 373456 275883 373462 275935
rect 373514 275923 373520 275935
rect 552784 275923 552790 275935
rect 373514 275895 552790 275923
rect 373514 275883 373520 275895
rect 552784 275883 552790 275895
rect 552842 275883 552848 275935
rect 296464 275809 296470 275861
rect 296522 275849 296528 275861
rect 362512 275849 362518 275861
rect 296522 275821 362518 275849
rect 296522 275809 296528 275821
rect 362512 275809 362518 275821
rect 362570 275809 362576 275861
rect 374608 275809 374614 275861
rect 374666 275849 374672 275861
rect 556336 275849 556342 275861
rect 374666 275821 556342 275849
rect 374666 275809 374672 275821
rect 556336 275809 556342 275821
rect 556394 275809 556400 275861
rect 297328 275735 297334 275787
rect 297386 275775 297392 275787
rect 364912 275775 364918 275787
rect 297386 275747 364918 275775
rect 297386 275735 297392 275747
rect 364912 275735 364918 275747
rect 364970 275735 364976 275787
rect 377488 275735 377494 275787
rect 377546 275775 377552 275787
rect 563440 275775 563446 275787
rect 377546 275747 563446 275775
rect 377546 275735 377552 275747
rect 563440 275735 563446 275747
rect 563498 275735 563504 275787
rect 297808 275661 297814 275713
rect 297866 275701 297872 275713
rect 366064 275701 366070 275713
rect 297866 275673 366070 275701
rect 297866 275661 297872 275673
rect 366064 275661 366070 275673
rect 366122 275661 366128 275713
rect 376240 275661 376246 275713
rect 376298 275701 376304 275713
rect 559888 275701 559894 275713
rect 376298 275673 559894 275701
rect 376298 275661 376304 275673
rect 559888 275661 559894 275673
rect 559946 275661 559952 275713
rect 298960 275587 298966 275639
rect 299018 275627 299024 275639
rect 368464 275627 368470 275639
rect 299018 275599 368470 275627
rect 299018 275587 299024 275599
rect 368464 275587 368470 275599
rect 368522 275587 368528 275639
rect 380560 275587 380566 275639
rect 380618 275627 380624 275639
rect 570544 275627 570550 275639
rect 380618 275599 570550 275627
rect 380618 275587 380624 275599
rect 570544 275587 570550 275599
rect 570602 275587 570608 275639
rect 300208 275513 300214 275565
rect 300266 275553 300272 275565
rect 372016 275553 372022 275565
rect 300266 275525 372022 275553
rect 300266 275513 300272 275525
rect 372016 275513 372022 275525
rect 372074 275513 372080 275565
rect 381808 275513 381814 275565
rect 381866 275553 381872 275565
rect 574096 275553 574102 275565
rect 381866 275525 574102 275553
rect 381866 275513 381872 275525
rect 574096 275513 574102 275525
rect 574154 275513 574160 275565
rect 299440 275439 299446 275491
rect 299498 275479 299504 275491
rect 369616 275479 369622 275491
rect 299498 275451 369622 275479
rect 299498 275439 299504 275451
rect 369616 275439 369622 275451
rect 369674 275439 369680 275491
rect 388912 275439 388918 275491
rect 388970 275479 388976 275491
rect 591856 275479 591862 275491
rect 388970 275451 591862 275479
rect 388970 275439 388976 275451
rect 591856 275439 591862 275451
rect 591914 275439 591920 275491
rect 303280 275365 303286 275417
rect 303338 275405 303344 275417
rect 379120 275405 379126 275417
rect 303338 275377 379126 275405
rect 303338 275365 303344 275377
rect 379120 275365 379126 275377
rect 379178 275365 379184 275417
rect 389584 275365 389590 275417
rect 389642 275405 389648 275417
rect 593008 275405 593014 275417
rect 389642 275377 593014 275405
rect 389642 275365 389648 275377
rect 593008 275365 593014 275377
rect 593066 275365 593072 275417
rect 304432 275291 304438 275343
rect 304490 275331 304496 275343
rect 382576 275331 382582 275343
rect 304490 275303 382582 275331
rect 304490 275291 304496 275303
rect 382576 275291 382582 275303
rect 382634 275291 382640 275343
rect 391984 275291 391990 275343
rect 392042 275331 392048 275343
rect 598960 275331 598966 275343
rect 392042 275303 598966 275331
rect 392042 275291 392048 275303
rect 598960 275291 598966 275303
rect 599018 275291 599024 275343
rect 307312 275217 307318 275269
rect 307370 275257 307376 275269
rect 389680 275257 389686 275269
rect 307370 275229 389686 275257
rect 307370 275217 307376 275229
rect 389680 275217 389686 275229
rect 389738 275217 389744 275269
rect 396304 275217 396310 275269
rect 396362 275257 396368 275269
rect 609520 275257 609526 275269
rect 396362 275229 609526 275257
rect 396362 275217 396368 275229
rect 609520 275217 609526 275229
rect 609578 275217 609584 275269
rect 310384 275143 310390 275195
rect 310442 275183 310448 275195
rect 396784 275183 396790 275195
rect 310442 275155 396790 275183
rect 310442 275143 310448 275155
rect 396784 275143 396790 275155
rect 396842 275143 396848 275195
rect 404944 275143 404950 275195
rect 405002 275183 405008 275195
rect 405002 275155 407678 275183
rect 405002 275143 405008 275155
rect 314704 275069 314710 275121
rect 314762 275109 314768 275121
rect 407440 275109 407446 275121
rect 314762 275081 407446 275109
rect 314762 275069 314768 275081
rect 407440 275069 407446 275081
rect 407498 275069 407504 275121
rect 311632 274995 311638 275047
rect 311690 275035 311696 275047
rect 400336 275035 400342 275047
rect 311690 275007 400342 275035
rect 311690 274995 311696 275007
rect 400336 274995 400342 275007
rect 400394 274995 400400 275047
rect 407650 275035 407678 275155
rect 407728 275143 407734 275195
rect 407786 275183 407792 275195
rect 623728 275183 623734 275195
rect 407786 275155 623734 275183
rect 407786 275143 407792 275155
rect 623728 275143 623734 275155
rect 623786 275143 623792 275195
rect 408592 275069 408598 275121
rect 408650 275109 408656 275121
rect 635536 275109 635542 275121
rect 408650 275081 635542 275109
rect 408650 275069 408656 275081
rect 635536 275069 635542 275081
rect 635594 275069 635600 275121
rect 630832 275035 630838 275047
rect 407650 275007 630838 275035
rect 630832 274995 630838 275007
rect 630890 274995 630896 275047
rect 284752 274921 284758 274973
rect 284810 274961 284816 274973
rect 332944 274961 332950 274973
rect 284810 274933 332950 274961
rect 284810 274921 284816 274933
rect 332944 274921 332950 274933
rect 333002 274921 333008 274973
rect 356176 274921 356182 274973
rect 356234 274961 356240 274973
rect 510256 274961 510262 274973
rect 356234 274933 510262 274961
rect 356234 274921 356240 274933
rect 510256 274921 510262 274933
rect 510314 274921 510320 274973
rect 283024 274847 283030 274899
rect 283082 274887 283088 274899
rect 329392 274887 329398 274899
rect 283082 274859 329398 274887
rect 283082 274847 283088 274859
rect 329392 274847 329398 274859
rect 329450 274847 329456 274899
rect 344560 274847 344566 274899
rect 344618 274887 344624 274899
rect 481936 274887 481942 274899
rect 344618 274859 481942 274887
rect 344618 274847 344624 274859
rect 481936 274847 481942 274859
rect 481994 274847 482000 274899
rect 281776 274773 281782 274825
rect 281834 274813 281840 274825
rect 325840 274813 325846 274825
rect 281834 274785 325846 274813
rect 281834 274773 281840 274785
rect 325840 274773 325846 274785
rect 325898 274773 325904 274825
rect 339088 274773 339094 274825
rect 339146 274813 339152 274825
rect 467728 274813 467734 274825
rect 339146 274785 467734 274813
rect 339146 274773 339152 274785
rect 467728 274773 467734 274785
rect 467786 274773 467792 274825
rect 336016 274699 336022 274751
rect 336074 274739 336080 274751
rect 460624 274739 460630 274751
rect 336074 274711 460630 274739
rect 336074 274699 336080 274711
rect 460624 274699 460630 274711
rect 460682 274699 460688 274751
rect 333136 274625 333142 274677
rect 333194 274665 333200 274677
rect 453520 274665 453526 274677
rect 333194 274637 453526 274665
rect 333194 274625 333200 274637
rect 453520 274625 453526 274637
rect 453578 274625 453584 274677
rect 330448 274551 330454 274603
rect 330506 274591 330512 274603
rect 446416 274591 446422 274603
rect 330506 274563 446422 274591
rect 330506 274551 330512 274563
rect 446416 274551 446422 274563
rect 446474 274551 446480 274603
rect 328816 274477 328822 274529
rect 328874 274517 328880 274529
rect 442864 274517 442870 274529
rect 328874 274489 442870 274517
rect 328874 274477 328880 274489
rect 442864 274477 442870 274489
rect 442922 274477 442928 274529
rect 325936 274403 325942 274455
rect 325994 274443 326000 274455
rect 435856 274443 435862 274455
rect 325994 274415 435862 274443
rect 325994 274403 326000 274415
rect 435856 274403 435862 274415
rect 435914 274403 435920 274455
rect 323344 274329 323350 274381
rect 323402 274369 323408 274381
rect 428752 274369 428758 274381
rect 323402 274341 428758 274369
rect 323402 274329 323408 274341
rect 428752 274329 428758 274341
rect 428810 274329 428816 274381
rect 320176 274255 320182 274307
rect 320234 274295 320240 274307
rect 421648 274295 421654 274307
rect 320234 274267 421654 274295
rect 320234 274255 320240 274267
rect 421648 274255 421654 274267
rect 421706 274255 421712 274307
rect 315952 274181 315958 274233
rect 316010 274221 316016 274233
rect 410992 274221 410998 274233
rect 316010 274193 410998 274221
rect 316010 274181 316016 274193
rect 410992 274181 410998 274193
rect 411050 274181 411056 274233
rect 317296 274107 317302 274159
rect 317354 274147 317360 274159
rect 414544 274147 414550 274159
rect 317354 274119 414550 274147
rect 317354 274107 317360 274119
rect 414544 274107 414550 274119
rect 414602 274107 414608 274159
rect 348496 274033 348502 274085
rect 348554 274073 348560 274085
rect 401488 274073 401494 274085
rect 348554 274045 401494 274073
rect 348554 274033 348560 274045
rect 401488 274033 401494 274045
rect 401546 274033 401552 274085
rect 401776 274033 401782 274085
rect 401834 274073 401840 274085
rect 407728 274073 407734 274085
rect 401834 274045 407734 274073
rect 401834 274033 401840 274045
rect 407728 274033 407734 274045
rect 407786 274033 407792 274085
rect 334288 273959 334294 274011
rect 334346 273999 334352 274011
rect 380272 273999 380278 274011
rect 334346 273971 380278 273999
rect 334346 273959 334352 273971
rect 380272 273959 380278 273971
rect 380330 273959 380336 274011
rect 347056 273885 347062 273937
rect 347114 273925 347120 273937
rect 394480 273925 394486 273937
rect 347114 273897 394486 273925
rect 347114 273885 347120 273897
rect 394480 273885 394486 273897
rect 394538 273885 394544 273937
rect 326128 273811 326134 273863
rect 326186 273851 326192 273863
rect 373168 273851 373174 273863
rect 326186 273823 373174 273851
rect 326186 273811 326192 273823
rect 373168 273811 373174 273823
rect 373226 273811 373232 273863
rect 341968 273737 341974 273789
rect 342026 273777 342032 273789
rect 387376 273777 387382 273789
rect 342026 273749 387382 273777
rect 342026 273737 342032 273749
rect 387376 273737 387382 273749
rect 387434 273737 387440 273789
rect 331216 273663 331222 273715
rect 331274 273703 331280 273715
rect 376720 273703 376726 273715
rect 331274 273675 376726 273703
rect 331274 273663 331280 273675
rect 376720 273663 376726 273675
rect 376778 273663 376784 273715
rect 43120 273515 43126 273567
rect 43178 273555 43184 273567
rect 56272 273555 56278 273567
rect 43178 273527 56278 273555
rect 43178 273515 43184 273527
rect 56272 273515 56278 273527
rect 56330 273515 56336 273567
rect 160432 273515 160438 273567
rect 160490 273555 160496 273567
rect 209392 273555 209398 273567
rect 160490 273527 209398 273555
rect 160490 273515 160496 273527
rect 209392 273515 209398 273527
rect 209450 273515 209456 273567
rect 230128 273515 230134 273567
rect 230186 273555 230192 273567
rect 242896 273555 242902 273567
rect 230186 273527 242902 273555
rect 230186 273515 230192 273527
rect 242896 273515 242902 273527
rect 242954 273515 242960 273567
rect 275152 273515 275158 273567
rect 275210 273555 275216 273567
rect 309328 273555 309334 273567
rect 275210 273527 309334 273555
rect 275210 273515 275216 273527
rect 309328 273515 309334 273527
rect 309386 273515 309392 273567
rect 350032 273515 350038 273567
rect 350090 273555 350096 273567
rect 494896 273555 494902 273567
rect 350090 273527 494902 273555
rect 350090 273515 350096 273527
rect 494896 273515 494902 273527
rect 494954 273515 494960 273567
rect 522544 273515 522550 273567
rect 522602 273555 522608 273567
rect 631984 273555 631990 273567
rect 522602 273527 631990 273555
rect 522602 273515 522608 273527
rect 631984 273515 631990 273527
rect 632042 273515 632048 273567
rect 130864 273441 130870 273493
rect 130922 273481 130928 273493
rect 190096 273481 190102 273493
rect 130922 273453 190102 273481
rect 130922 273441 130928 273453
rect 190096 273441 190102 273453
rect 190154 273441 190160 273493
rect 193552 273441 193558 273493
rect 193610 273481 193616 273493
rect 219088 273481 219094 273493
rect 193610 273453 219094 273481
rect 193610 273441 193616 273453
rect 219088 273441 219094 273453
rect 219146 273441 219152 273493
rect 227824 273441 227830 273493
rect 227882 273481 227888 273493
rect 242128 273481 242134 273493
rect 227882 273453 242134 273481
rect 227882 273441 227888 273453
rect 242128 273441 242134 273453
rect 242186 273441 242192 273493
rect 277744 273441 277750 273493
rect 277802 273481 277808 273493
rect 316432 273481 316438 273493
rect 277802 273453 316438 273481
rect 277802 273441 277808 273453
rect 316432 273441 316438 273453
rect 316490 273441 316496 273493
rect 349456 273441 349462 273493
rect 349514 273481 349520 273493
rect 493744 273481 493750 273493
rect 349514 273453 493750 273481
rect 349514 273441 349520 273453
rect 493744 273441 493750 273453
rect 493802 273441 493808 273493
rect 529840 273441 529846 273493
rect 529898 273481 529904 273493
rect 624976 273481 624982 273493
rect 529898 273453 624982 273481
rect 529898 273441 529904 273453
rect 624976 273441 624982 273453
rect 625034 273441 625040 273493
rect 108400 273367 108406 273419
rect 108458 273407 108464 273419
rect 109360 273407 109366 273419
rect 108458 273379 109366 273407
rect 108458 273367 108464 273379
rect 109360 273367 109366 273379
rect 109418 273367 109424 273419
rect 122608 273367 122614 273419
rect 122666 273407 122672 273419
rect 123760 273407 123766 273419
rect 122666 273379 123766 273407
rect 122666 273367 122672 273379
rect 123760 273367 123766 273379
rect 123818 273367 123824 273419
rect 142672 273367 142678 273419
rect 142730 273407 142736 273419
rect 209680 273407 209686 273419
rect 142730 273379 209686 273407
rect 142730 273367 142736 273379
rect 209680 273367 209686 273379
rect 209738 273367 209744 273419
rect 275344 273367 275350 273419
rect 275402 273407 275408 273419
rect 310480 273407 310486 273419
rect 275402 273379 310486 273407
rect 275402 273367 275408 273379
rect 310480 273367 310486 273379
rect 310538 273367 310544 273419
rect 310576 273367 310582 273419
rect 310634 273407 310640 273419
rect 344752 273407 344758 273419
rect 310634 273379 344758 273407
rect 310634 273367 310640 273379
rect 344752 273367 344758 273379
rect 344810 273367 344816 273419
rect 352432 273367 352438 273419
rect 352490 273407 352496 273419
rect 500848 273407 500854 273419
rect 352490 273379 500854 273407
rect 352490 273367 352496 273379
rect 500848 273367 500854 273379
rect 500906 273367 500912 273419
rect 135568 273293 135574 273345
rect 135626 273333 135632 273345
rect 209872 273333 209878 273345
rect 135626 273305 209878 273333
rect 135626 273293 135632 273305
rect 209872 273293 209878 273305
rect 209930 273293 209936 273345
rect 219568 273293 219574 273345
rect 219626 273333 219632 273345
rect 238672 273333 238678 273345
rect 219626 273305 238678 273333
rect 219626 273293 219632 273305
rect 238672 273293 238678 273305
rect 238730 273293 238736 273345
rect 278224 273293 278230 273345
rect 278282 273333 278288 273345
rect 317584 273333 317590 273345
rect 278282 273305 317590 273333
rect 278282 273293 278288 273305
rect 317584 273293 317590 273305
rect 317642 273293 317648 273345
rect 352624 273293 352630 273345
rect 352682 273333 352688 273345
rect 502000 273333 502006 273345
rect 352682 273305 502006 273333
rect 352682 273293 352688 273305
rect 502000 273293 502006 273305
rect 502058 273293 502064 273345
rect 68272 273219 68278 273271
rect 68330 273259 68336 273271
rect 142480 273259 142486 273271
rect 68330 273231 142486 273259
rect 68330 273219 68336 273231
rect 142480 273219 142486 273231
rect 142538 273219 142544 273271
rect 153328 273219 153334 273271
rect 153386 273259 153392 273271
rect 209584 273259 209590 273271
rect 153386 273231 209590 273259
rect 153386 273219 153392 273231
rect 209584 273219 209590 273231
rect 209642 273219 209648 273271
rect 279664 273219 279670 273271
rect 279722 273259 279728 273271
rect 321136 273259 321142 273271
rect 279722 273231 321142 273259
rect 279722 273219 279728 273231
rect 321136 273219 321142 273231
rect 321194 273219 321200 273271
rect 355504 273219 355510 273271
rect 355562 273259 355568 273271
rect 509104 273259 509110 273271
rect 355562 273231 509110 273259
rect 355562 273219 355568 273231
rect 509104 273219 509110 273231
rect 509162 273219 509168 273271
rect 132016 273145 132022 273197
rect 132074 273185 132080 273197
rect 209776 273185 209782 273197
rect 132074 273157 209782 273185
rect 132074 273145 132080 273157
rect 209776 273145 209782 273157
rect 209834 273145 209840 273197
rect 285616 273145 285622 273197
rect 285674 273185 285680 273197
rect 335344 273185 335350 273197
rect 285674 273157 335350 273185
rect 285674 273145 285680 273157
rect 335344 273145 335350 273157
rect 335402 273145 335408 273197
rect 355024 273145 355030 273197
rect 355082 273185 355088 273197
rect 507952 273185 507958 273197
rect 355082 273157 507958 273185
rect 355082 273145 355088 273157
rect 507952 273145 507958 273157
rect 508010 273145 508016 273197
rect 508240 273145 508246 273197
rect 508298 273185 508304 273197
rect 639088 273185 639094 273197
rect 508298 273157 639094 273185
rect 508298 273145 508304 273157
rect 639088 273145 639094 273157
rect 639146 273145 639152 273197
rect 127312 273071 127318 273123
rect 127370 273111 127376 273123
rect 209968 273111 209974 273123
rect 127370 273083 209974 273111
rect 127370 273071 127376 273083
rect 209968 273071 209974 273083
rect 210026 273071 210032 273123
rect 217168 273071 217174 273123
rect 217226 273111 217232 273123
rect 237616 273111 237622 273123
rect 217226 273083 237622 273111
rect 217226 273071 217232 273083
rect 237616 273071 237622 273083
rect 237674 273071 237680 273123
rect 284944 273071 284950 273123
rect 285002 273111 285008 273123
rect 334192 273111 334198 273123
rect 285002 273083 334198 273111
rect 285002 273071 285008 273083
rect 334192 273071 334198 273083
rect 334250 273071 334256 273123
rect 358576 273071 358582 273123
rect 358634 273111 358640 273123
rect 358634 273083 375134 273111
rect 358634 273071 358640 273083
rect 128464 272997 128470 273049
rect 128522 273037 128528 273049
rect 210160 273037 210166 273049
rect 128522 273009 210166 273037
rect 128522 272997 128528 273009
rect 210160 272997 210166 273009
rect 210218 272997 210224 273049
rect 218320 272997 218326 273049
rect 218378 273037 218384 273049
rect 238096 273037 238102 273049
rect 218378 273009 238102 273037
rect 218378 272997 218384 273009
rect 238096 272997 238102 273009
rect 238154 272997 238160 273049
rect 286768 272997 286774 273049
rect 286826 273037 286832 273049
rect 338896 273037 338902 273049
rect 286826 273009 338902 273037
rect 286826 272997 286832 273009
rect 338896 272997 338902 273009
rect 338954 272997 338960 273049
rect 360976 272997 360982 273049
rect 361034 273037 361040 273049
rect 375106 273037 375134 273083
rect 375184 273071 375190 273123
rect 375242 273111 375248 273123
rect 514960 273111 514966 273123
rect 375242 273083 514966 273111
rect 375242 273071 375248 273083
rect 514960 273071 514966 273083
rect 515018 273071 515024 273123
rect 516208 273037 516214 273049
rect 361034 273009 375038 273037
rect 375106 273009 516214 273037
rect 361034 272997 361040 273009
rect 125008 272923 125014 272975
rect 125066 272963 125072 272975
rect 207280 272963 207286 272975
rect 125066 272935 207286 272963
rect 125066 272923 125072 272935
rect 207280 272923 207286 272935
rect 207338 272923 207344 272975
rect 216016 272923 216022 272975
rect 216074 272963 216080 272975
rect 236944 272963 236950 272975
rect 216074 272935 236950 272963
rect 216074 272923 216080 272935
rect 236944 272923 236950 272935
rect 237002 272923 237008 272975
rect 274192 272923 274198 272975
rect 274250 272963 274256 272975
rect 306928 272963 306934 272975
rect 274250 272935 306934 272963
rect 274250 272923 274256 272935
rect 306928 272923 306934 272935
rect 306986 272923 306992 272975
rect 307024 272923 307030 272975
rect 307082 272963 307088 272975
rect 358960 272963 358966 272975
rect 307082 272935 358966 272963
rect 307082 272923 307088 272935
rect 358960 272923 358966 272935
rect 359018 272923 359024 272975
rect 361264 272923 361270 272975
rect 361322 272963 361328 272975
rect 375010 272963 375038 273009
rect 516208 272997 516214 273009
rect 516266 272997 516272 273049
rect 516304 272997 516310 273049
rect 516362 273037 516368 273049
rect 580048 273037 580054 273049
rect 516362 273009 580054 273037
rect 516362 272997 516368 273009
rect 580048 272997 580054 273009
rect 580106 272997 580112 273049
rect 522064 272963 522070 272975
rect 361322 272935 374942 272963
rect 375010 272935 522070 272963
rect 361322 272923 361328 272935
rect 123664 272849 123670 272901
rect 123722 272889 123728 272901
rect 209008 272889 209014 272901
rect 123722 272861 209014 272889
rect 123722 272849 123728 272861
rect 209008 272849 209014 272861
rect 209066 272849 209072 272901
rect 220720 272849 220726 272901
rect 220778 272889 220784 272901
rect 239152 272889 239158 272901
rect 220778 272861 239158 272889
rect 220778 272849 220784 272861
rect 239152 272849 239158 272861
rect 239210 272849 239216 272901
rect 289936 272849 289942 272901
rect 289994 272889 290000 272901
rect 346000 272889 346006 272901
rect 289994 272861 346006 272889
rect 289994 272849 290000 272861
rect 346000 272849 346006 272861
rect 346058 272849 346064 272901
rect 363568 272849 363574 272901
rect 363626 272889 363632 272901
rect 374914 272889 374942 272935
rect 522064 272923 522070 272935
rect 522122 272923 522128 272975
rect 523312 272889 523318 272901
rect 363626 272861 374846 272889
rect 374914 272861 523318 272889
rect 363626 272849 363632 272861
rect 120208 272775 120214 272827
rect 120266 272815 120272 272827
rect 207856 272815 207862 272827
rect 120266 272787 207862 272815
rect 120266 272775 120272 272787
rect 207856 272775 207862 272787
rect 207914 272775 207920 272827
rect 211216 272775 211222 272827
rect 211274 272815 211280 272827
rect 235024 272815 235030 272827
rect 211274 272787 235030 272815
rect 211274 272775 211280 272787
rect 235024 272775 235030 272787
rect 235082 272775 235088 272827
rect 292240 272775 292246 272827
rect 292298 272815 292304 272827
rect 351856 272815 351862 272827
rect 292298 272787 351862 272815
rect 292298 272775 292304 272787
rect 351856 272775 351862 272787
rect 351914 272775 351920 272827
rect 364144 272775 364150 272827
rect 364202 272815 364208 272827
rect 374818 272815 374846 272861
rect 523312 272849 523318 272861
rect 523370 272849 523376 272901
rect 523792 272849 523798 272901
rect 523850 272889 523856 272901
rect 611920 272889 611926 272901
rect 523850 272861 611926 272889
rect 523850 272849 523856 272861
rect 611920 272849 611926 272861
rect 611978 272849 611984 272901
rect 529168 272815 529174 272827
rect 364202 272787 374750 272815
rect 374818 272787 529174 272815
rect 364202 272775 364208 272787
rect 116656 272701 116662 272753
rect 116714 272741 116720 272753
rect 207088 272741 207094 272753
rect 116714 272713 207094 272741
rect 116714 272701 116720 272713
rect 207088 272701 207094 272713
rect 207146 272701 207152 272753
rect 233680 272701 233686 272753
rect 233738 272741 233744 272753
rect 244048 272741 244054 272753
rect 233738 272713 244054 272741
rect 233738 272701 233744 272713
rect 244048 272701 244054 272713
rect 244106 272701 244112 272753
rect 292720 272701 292726 272753
rect 292778 272741 292784 272753
rect 353104 272741 353110 272753
rect 292778 272713 353110 272741
rect 292778 272701 292784 272713
rect 353104 272701 353110 272713
rect 353162 272701 353168 272753
rect 366544 272701 366550 272753
rect 366602 272741 366608 272753
rect 374722 272741 374750 272787
rect 529168 272775 529174 272787
rect 529226 272775 529232 272827
rect 530416 272741 530422 272753
rect 366602 272713 374654 272741
rect 374722 272713 530422 272741
rect 366602 272701 366608 272713
rect 113104 272627 113110 272679
rect 113162 272667 113168 272679
rect 206032 272667 206038 272679
rect 113162 272639 206038 272667
rect 113162 272627 113168 272639
rect 206032 272627 206038 272639
rect 206090 272627 206096 272679
rect 213616 272627 213622 272679
rect 213674 272667 213680 272679
rect 236272 272667 236278 272679
rect 213674 272639 236278 272667
rect 213674 272627 213680 272639
rect 236272 272627 236278 272639
rect 236330 272627 236336 272679
rect 295408 272627 295414 272679
rect 295466 272667 295472 272679
rect 360208 272667 360214 272679
rect 295466 272639 360214 272667
rect 295466 272627 295472 272639
rect 360208 272627 360214 272639
rect 360266 272627 360272 272679
rect 367120 272627 367126 272679
rect 367178 272667 367184 272679
rect 374626 272667 374654 272713
rect 530416 272701 530422 272713
rect 530474 272701 530480 272753
rect 536272 272667 536278 272679
rect 367178 272639 374558 272667
rect 374626 272639 536278 272667
rect 367178 272627 367184 272639
rect 96592 272553 96598 272605
rect 96650 272593 96656 272605
rect 106672 272593 106678 272605
rect 96650 272565 106678 272593
rect 96650 272553 96656 272565
rect 106672 272553 106678 272565
rect 106730 272553 106736 272605
rect 110800 272553 110806 272605
rect 110858 272593 110864 272605
rect 205456 272593 205462 272605
rect 110858 272565 205462 272593
rect 110858 272553 110864 272565
rect 205456 272553 205462 272565
rect 205514 272553 205520 272605
rect 214768 272553 214774 272605
rect 214826 272593 214832 272605
rect 236464 272593 236470 272605
rect 214826 272565 236470 272593
rect 214826 272553 214832 272565
rect 236464 272553 236470 272565
rect 236522 272553 236528 272605
rect 270256 272553 270262 272605
rect 270314 272593 270320 272605
rect 297520 272593 297526 272605
rect 270314 272565 297526 272593
rect 270314 272553 270320 272565
rect 297520 272553 297526 272565
rect 297578 272553 297584 272605
rect 298480 272553 298486 272605
rect 298538 272593 298544 272605
rect 367216 272593 367222 272605
rect 298538 272565 367222 272593
rect 298538 272553 298544 272565
rect 367216 272553 367222 272565
rect 367274 272553 367280 272605
rect 372688 272553 372694 272605
rect 372746 272593 372752 272605
rect 374530 272593 374558 272639
rect 536272 272627 536278 272639
rect 536330 272627 536336 272679
rect 537424 272593 537430 272605
rect 372746 272565 374462 272593
rect 374530 272565 537430 272593
rect 372746 272553 372752 272565
rect 103696 272479 103702 272531
rect 103754 272519 103760 272531
rect 203536 272519 203542 272531
rect 103754 272491 203542 272519
rect 103754 272479 103760 272491
rect 203536 272479 203542 272491
rect 203594 272479 203600 272531
rect 210064 272479 210070 272531
rect 210122 272519 210128 272531
rect 234544 272519 234550 272531
rect 210122 272491 234550 272519
rect 210122 272479 210128 272491
rect 234544 272479 234550 272491
rect 234602 272479 234608 272531
rect 236080 272479 236086 272531
rect 236138 272519 236144 272531
rect 245296 272519 245302 272531
rect 236138 272491 245302 272519
rect 236138 272479 236144 272491
rect 245296 272479 245302 272491
rect 245354 272479 245360 272531
rect 272272 272479 272278 272531
rect 272330 272519 272336 272531
rect 302224 272519 302230 272531
rect 272330 272491 302230 272519
rect 272330 272479 272336 272491
rect 302224 272479 302230 272491
rect 302282 272479 302288 272531
rect 374320 272519 374326 272531
rect 302338 272491 374326 272519
rect 106096 272405 106102 272457
rect 106154 272445 106160 272457
rect 204016 272445 204022 272457
rect 106154 272417 204022 272445
rect 106154 272405 106160 272417
rect 204016 272405 204022 272417
rect 204074 272405 204080 272457
rect 205360 272405 205366 272457
rect 205418 272445 205424 272457
rect 232624 272445 232630 272457
rect 205418 272417 232630 272445
rect 205418 272405 205424 272417
rect 232624 272405 232630 272417
rect 232682 272405 232688 272457
rect 270544 272405 270550 272457
rect 270602 272445 270608 272457
rect 298672 272445 298678 272457
rect 270602 272417 298678 272445
rect 270602 272405 270608 272417
rect 298672 272405 298678 272417
rect 298730 272405 298736 272457
rect 301360 272405 301366 272457
rect 301418 272445 301424 272457
rect 302338 272445 302366 272491
rect 374320 272479 374326 272491
rect 374378 272479 374384 272531
rect 374434 272519 374462 272565
rect 537424 272553 537430 272565
rect 537482 272553 537488 272605
rect 551632 272519 551638 272531
rect 374434 272491 551638 272519
rect 551632 272479 551638 272491
rect 551690 272479 551696 272531
rect 301418 272417 302366 272445
rect 301418 272405 301424 272417
rect 303952 272405 303958 272457
rect 304010 272445 304016 272457
rect 381424 272445 381430 272457
rect 304010 272417 381430 272445
rect 304010 272405 304016 272417
rect 381424 272405 381430 272417
rect 381482 272405 381488 272457
rect 381520 272405 381526 272457
rect 381578 272445 381584 272457
rect 572944 272445 572950 272457
rect 381578 272417 572950 272445
rect 381578 272405 381584 272417
rect 572944 272405 572950 272417
rect 573002 272405 573008 272457
rect 98992 272331 98998 272383
rect 99050 272371 99056 272383
rect 199120 272371 199126 272383
rect 99050 272343 199126 272371
rect 99050 272331 99056 272343
rect 199120 272331 199126 272343
rect 199178 272331 199184 272383
rect 207664 272331 207670 272383
rect 207722 272371 207728 272383
rect 233872 272371 233878 272383
rect 207722 272343 233878 272371
rect 207722 272331 207728 272343
rect 233872 272331 233878 272343
rect 233930 272331 233936 272383
rect 272752 272331 272758 272383
rect 272810 272371 272816 272383
rect 303472 272371 303478 272383
rect 272810 272343 303478 272371
rect 272810 272331 272816 272343
rect 303472 272331 303478 272343
rect 303530 272331 303536 272383
rect 307120 272331 307126 272383
rect 307178 272371 307184 272383
rect 388528 272371 388534 272383
rect 307178 272343 388534 272371
rect 307178 272331 307184 272343
rect 388528 272331 388534 272343
rect 388586 272331 388592 272383
rect 407440 272331 407446 272383
rect 407498 272371 407504 272383
rect 587152 272371 587158 272383
rect 407498 272343 587158 272371
rect 407498 272331 407504 272343
rect 587152 272331 587158 272343
rect 587210 272331 587216 272383
rect 76528 272257 76534 272309
rect 76586 272297 76592 272309
rect 76586 272269 106622 272297
rect 76586 272257 76592 272269
rect 84784 272183 84790 272235
rect 84842 272223 84848 272235
rect 86320 272223 86326 272235
rect 84842 272195 86326 272223
rect 84842 272183 84848 272195
rect 86320 272183 86326 272195
rect 86378 272183 86384 272235
rect 104848 272183 104854 272235
rect 104906 272223 104912 272235
rect 106480 272223 106486 272235
rect 104906 272195 106486 272223
rect 104906 272183 104912 272195
rect 106480 272183 106486 272195
rect 106538 272183 106544 272235
rect 106594 272223 106622 272269
rect 106672 272257 106678 272309
rect 106730 272297 106736 272309
rect 201616 272297 201622 272309
rect 106730 272269 201622 272297
rect 106730 272257 106736 272269
rect 201616 272257 201622 272269
rect 201674 272257 201680 272309
rect 208912 272257 208918 272309
rect 208970 272297 208976 272309
rect 234352 272297 234358 272309
rect 208970 272269 234358 272297
rect 208970 272257 208976 272269
rect 234352 272257 234358 272269
rect 234410 272257 234416 272309
rect 234928 272257 234934 272309
rect 234986 272297 234992 272309
rect 244816 272297 244822 272309
rect 234986 272269 244822 272297
rect 234986 272257 234992 272269
rect 244816 272257 244822 272269
rect 244874 272257 244880 272309
rect 273424 272257 273430 272309
rect 273482 272297 273488 272309
rect 305776 272297 305782 272309
rect 273482 272269 305782 272297
rect 273482 272257 273488 272269
rect 305776 272257 305782 272269
rect 305834 272257 305840 272309
rect 309904 272257 309910 272309
rect 309962 272297 309968 272309
rect 395632 272297 395638 272309
rect 309962 272269 395638 272297
rect 309962 272257 309968 272269
rect 395632 272257 395638 272269
rect 395690 272257 395696 272309
rect 395920 272257 395926 272309
rect 395978 272297 395984 272309
rect 608368 272297 608374 272309
rect 395978 272269 608374 272297
rect 395978 272257 395984 272269
rect 608368 272257 608374 272269
rect 608426 272257 608432 272309
rect 195664 272223 195670 272235
rect 106594 272195 195670 272223
rect 195664 272183 195670 272195
rect 195722 272183 195728 272235
rect 198256 272183 198262 272235
rect 198314 272223 198320 272235
rect 222064 272223 222070 272235
rect 198314 272195 222070 272223
rect 198314 272183 198320 272195
rect 222064 272183 222070 272195
rect 222122 272183 222128 272235
rect 276304 272183 276310 272235
rect 276362 272223 276368 272235
rect 312880 272223 312886 272235
rect 276362 272195 312886 272223
rect 276362 272183 276368 272195
rect 312880 272183 312886 272195
rect 312938 272183 312944 272235
rect 312976 272183 312982 272235
rect 313034 272223 313040 272235
rect 402736 272223 402742 272235
rect 313034 272195 402742 272223
rect 313034 272183 313040 272195
rect 402736 272183 402742 272195
rect 402794 272183 402800 272235
rect 402832 272183 402838 272235
rect 402890 272223 402896 272235
rect 622576 272223 622582 272235
rect 402890 272195 622582 272223
rect 402890 272183 402896 272195
rect 622576 272183 622582 272195
rect 622634 272183 622640 272235
rect 194704 272109 194710 272161
rect 194762 272149 194768 272161
rect 222256 272149 222262 272161
rect 194762 272121 222262 272149
rect 194762 272109 194768 272121
rect 222256 272109 222262 272121
rect 222314 272109 222320 272161
rect 228976 272109 228982 272161
rect 229034 272149 229040 272161
rect 242416 272149 242422 272161
rect 229034 272121 242422 272149
rect 229034 272109 229040 272121
rect 242416 272109 242422 272121
rect 242474 272109 242480 272161
rect 277072 272109 277078 272161
rect 277130 272149 277136 272161
rect 314032 272149 314038 272161
rect 277130 272121 314038 272149
rect 277130 272109 277136 272121
rect 314032 272109 314038 272121
rect 314090 272109 314096 272161
rect 315472 272109 315478 272161
rect 315530 272149 315536 272161
rect 409840 272149 409846 272161
rect 315530 272121 409846 272149
rect 315530 272109 315536 272121
rect 409840 272109 409846 272121
rect 409898 272109 409904 272161
rect 413680 272109 413686 272161
rect 413738 272149 413744 272161
rect 643888 272149 643894 272161
rect 413738 272121 643894 272149
rect 413738 272109 413744 272121
rect 643888 272109 643894 272121
rect 643946 272109 643952 272161
rect 119056 272035 119062 272087
rect 119114 272075 119120 272087
rect 120880 272075 120886 272087
rect 119114 272047 120886 272075
rect 119114 272035 119120 272047
rect 120880 272035 120886 272047
rect 120938 272035 120944 272087
rect 165136 272035 165142 272087
rect 165194 272075 165200 272087
rect 166960 272075 166966 272087
rect 165194 272047 166966 272075
rect 165194 272035 165200 272047
rect 166960 272035 166966 272047
rect 167018 272035 167024 272087
rect 167536 272035 167542 272087
rect 167594 272075 167600 272087
rect 213040 272075 213046 272087
rect 167594 272047 213046 272075
rect 167594 272035 167600 272047
rect 213040 272035 213046 272047
rect 213098 272035 213104 272087
rect 298096 272035 298102 272087
rect 298154 272075 298160 272087
rect 327088 272075 327094 272087
rect 298154 272047 327094 272075
rect 298154 272035 298160 272047
rect 327088 272035 327094 272047
rect 327146 272035 327152 272087
rect 346960 272035 346966 272087
rect 347018 272075 347024 272087
rect 487792 272075 487798 272087
rect 347018 272047 487798 272075
rect 347018 272035 347024 272047
rect 487792 272035 487798 272047
rect 487850 272035 487856 272087
rect 174640 271961 174646 272013
rect 174698 272001 174704 272013
rect 212848 272001 212854 272013
rect 174698 271973 212854 272001
rect 174698 271961 174704 271973
rect 212848 271961 212854 271973
rect 212906 271961 212912 272013
rect 232528 271961 232534 272013
rect 232586 272001 232592 272013
rect 243664 272001 243670 272013
rect 232586 271973 243670 272001
rect 232586 271961 232592 271973
rect 243664 271961 243670 271973
rect 243722 271961 243728 272013
rect 271024 271961 271030 272013
rect 271082 272001 271088 272013
rect 299920 272001 299926 272013
rect 271082 271973 299926 272001
rect 271082 271961 271088 271973
rect 299920 271961 299926 271973
rect 299978 271961 299984 272013
rect 328240 272001 328246 272013
rect 300034 271973 328246 272001
rect 159280 271887 159286 271939
rect 159338 271927 159344 271939
rect 195280 271927 195286 271939
rect 159338 271899 195286 271927
rect 159338 271887 159344 271899
rect 195280 271887 195286 271899
rect 195338 271887 195344 271939
rect 195856 271887 195862 271939
rect 195914 271927 195920 271939
rect 218992 271927 218998 271939
rect 195914 271899 218998 271927
rect 195914 271887 195920 271899
rect 218992 271887 218998 271899
rect 219050 271887 219056 271939
rect 231376 271887 231382 271939
rect 231434 271927 231440 271939
rect 243088 271927 243094 271939
rect 231434 271899 243094 271927
rect 231434 271887 231440 271899
rect 243088 271887 243094 271899
rect 243146 271887 243152 271939
rect 191152 271813 191158 271865
rect 191210 271853 191216 271865
rect 227152 271853 227158 271865
rect 191210 271825 227158 271853
rect 191210 271813 191216 271825
rect 227152 271813 227158 271825
rect 227210 271813 227216 271865
rect 298000 271813 298006 271865
rect 298058 271853 298064 271865
rect 300034 271853 300062 271973
rect 328240 271961 328246 271973
rect 328298 271961 328304 272013
rect 346480 271961 346486 272013
rect 346538 272001 346544 272013
rect 486640 272001 486646 272013
rect 346538 271973 486646 272001
rect 346538 271961 346544 271973
rect 486640 271961 486646 271973
rect 486698 271961 486704 272013
rect 324688 271927 324694 271939
rect 308146 271899 324694 271927
rect 298058 271825 300062 271853
rect 298058 271813 298064 271825
rect 300112 271813 300118 271865
rect 300170 271853 300176 271865
rect 308146 271853 308174 271899
rect 324688 271887 324694 271899
rect 324746 271887 324752 271939
rect 342736 271887 342742 271939
rect 342794 271927 342800 271939
rect 348304 271927 348310 271939
rect 342794 271899 348310 271927
rect 342794 271887 342800 271899
rect 348304 271887 348310 271899
rect 348362 271887 348368 271939
rect 480688 271927 480694 271939
rect 348418 271899 480694 271927
rect 300170 271825 308174 271853
rect 300170 271813 300176 271825
rect 344080 271813 344086 271865
rect 344138 271853 344144 271865
rect 348418 271853 348446 271899
rect 480688 271887 480694 271899
rect 480746 271887 480752 271939
rect 473680 271853 473686 271865
rect 344138 271825 348446 271853
rect 348514 271825 473686 271853
rect 344138 271813 344144 271825
rect 147376 271739 147382 271791
rect 147434 271779 147440 271791
rect 149680 271779 149686 271791
rect 147434 271751 149686 271779
rect 147434 271739 147440 271751
rect 149680 271739 149686 271751
rect 149738 271739 149744 271791
rect 192304 271739 192310 271791
rect 192362 271779 192368 271791
rect 222160 271779 222166 271791
rect 192362 271751 222166 271779
rect 192362 271739 192368 271751
rect 222160 271739 222166 271751
rect 222218 271739 222224 271791
rect 341488 271739 341494 271791
rect 341546 271779 341552 271791
rect 348514 271779 348542 271825
rect 473680 271813 473686 271825
rect 473738 271813 473744 271865
rect 341546 271751 348542 271779
rect 341546 271739 341552 271751
rect 348592 271739 348598 271791
rect 348650 271779 348656 271791
rect 466576 271779 466582 271791
rect 348650 271751 466582 271779
rect 348650 271739 348656 271751
rect 466576 271739 466582 271751
rect 466634 271739 466640 271791
rect 166288 271665 166294 271717
rect 166346 271705 166352 271717
rect 196336 271705 196342 271717
rect 166346 271677 196342 271705
rect 166346 271665 166352 271677
rect 196336 271665 196342 271677
rect 196394 271665 196400 271717
rect 199408 271665 199414 271717
rect 199466 271705 199472 271717
rect 218896 271705 218902 271717
rect 199466 271677 218902 271705
rect 199466 271665 199472 271677
rect 218896 271665 218902 271677
rect 218954 271665 218960 271717
rect 335440 271665 335446 271717
rect 335498 271705 335504 271717
rect 459472 271705 459478 271717
rect 335498 271677 459478 271705
rect 335498 271665 335504 271677
rect 459472 271665 459478 271677
rect 459530 271665 459536 271717
rect 75280 271591 75286 271643
rect 75338 271631 75344 271643
rect 77680 271631 77686 271643
rect 75338 271603 77686 271631
rect 75338 271591 75344 271603
rect 77680 271591 77686 271603
rect 77738 271591 77744 271643
rect 129712 271591 129718 271643
rect 129770 271631 129776 271643
rect 132400 271631 132406 271643
rect 129770 271603 132406 271631
rect 129770 271591 129776 271603
rect 132400 271591 132406 271603
rect 132458 271591 132464 271643
rect 181744 271591 181750 271643
rect 181802 271631 181808 271643
rect 212944 271631 212950 271643
rect 181802 271603 212950 271631
rect 181802 271591 181808 271603
rect 212944 271591 212950 271603
rect 213002 271591 213008 271643
rect 332560 271591 332566 271643
rect 332618 271631 332624 271643
rect 452368 271631 452374 271643
rect 332618 271603 452374 271631
rect 332618 271591 332624 271603
rect 452368 271591 452374 271603
rect 452426 271591 452432 271643
rect 89488 271517 89494 271569
rect 89546 271557 89552 271569
rect 92080 271557 92086 271569
rect 89546 271529 92086 271557
rect 89546 271517 89552 271529
rect 92080 271517 92086 271529
rect 92138 271517 92144 271569
rect 150928 271517 150934 271569
rect 150986 271557 150992 271569
rect 152368 271557 152374 271569
rect 150986 271529 152374 271557
rect 150986 271517 150992 271529
rect 152368 271517 152374 271529
rect 152426 271517 152432 271569
rect 185200 271517 185206 271569
rect 185258 271557 185264 271569
rect 212560 271557 212566 271569
rect 185258 271529 212566 271557
rect 185258 271517 185264 271529
rect 212560 271517 212566 271529
rect 212618 271517 212624 271569
rect 329968 271517 329974 271569
rect 330026 271557 330032 271569
rect 445264 271557 445270 271569
rect 330026 271529 445270 271557
rect 330026 271517 330032 271529
rect 445264 271517 445270 271529
rect 445322 271517 445328 271569
rect 173392 271443 173398 271495
rect 173450 271483 173456 271495
rect 201520 271483 201526 271495
rect 173450 271455 201526 271483
rect 173450 271443 173456 271455
rect 201520 271443 201526 271455
rect 201578 271443 201584 271495
rect 201808 271443 201814 271495
rect 201866 271483 201872 271495
rect 221968 271483 221974 271495
rect 201866 271455 221974 271483
rect 201866 271443 201872 271455
rect 221968 271443 221974 271455
rect 222026 271443 222032 271495
rect 326896 271443 326902 271495
rect 326954 271483 326960 271495
rect 438160 271483 438166 271495
rect 326954 271455 438166 271483
rect 326954 271443 326960 271455
rect 438160 271443 438166 271455
rect 438218 271443 438224 271495
rect 180496 271369 180502 271421
rect 180554 271409 180560 271421
rect 205936 271409 205942 271421
rect 180554 271381 205942 271409
rect 180554 271369 180560 271381
rect 205936 271369 205942 271381
rect 205994 271369 206000 271421
rect 212464 271369 212470 271421
rect 212522 271409 212528 271421
rect 235696 271409 235702 271421
rect 212522 271381 235702 271409
rect 212522 271369 212528 271381
rect 235696 271369 235702 271381
rect 235754 271369 235760 271421
rect 324016 271369 324022 271421
rect 324074 271409 324080 271421
rect 431056 271409 431062 271421
rect 324074 271381 431062 271409
rect 324074 271369 324080 271381
rect 431056 271369 431062 271381
rect 431114 271369 431120 271421
rect 188752 271295 188758 271347
rect 188810 271335 188816 271347
rect 212752 271335 212758 271347
rect 188810 271307 212758 271335
rect 188810 271295 188816 271307
rect 212752 271295 212758 271307
rect 212810 271295 212816 271347
rect 321424 271295 321430 271347
rect 321482 271335 321488 271347
rect 423952 271335 423958 271347
rect 321482 271307 423958 271335
rect 321482 271295 321488 271307
rect 423952 271295 423958 271307
rect 424010 271295 424016 271347
rect 161584 271221 161590 271273
rect 161642 271261 161648 271273
rect 163888 271261 163894 271273
rect 161642 271233 163894 271261
rect 161642 271221 161648 271233
rect 163888 271221 163894 271233
rect 163946 271221 163952 271273
rect 184048 271221 184054 271273
rect 184106 271261 184112 271273
rect 205744 271261 205750 271273
rect 184106 271233 205750 271261
rect 184106 271221 184112 271233
rect 205744 271221 205750 271233
rect 205802 271221 205808 271273
rect 237232 271221 237238 271273
rect 237290 271261 237296 271273
rect 245584 271261 245590 271273
rect 237290 271233 245590 271261
rect 237290 271221 237296 271233
rect 245584 271221 245590 271233
rect 245642 271221 245648 271273
rect 318352 271221 318358 271273
rect 318410 271261 318416 271273
rect 416944 271261 416950 271273
rect 318410 271233 416950 271261
rect 318410 271221 318416 271233
rect 416944 271221 416950 271233
rect 417002 271221 417008 271273
rect 175792 271147 175798 271199
rect 175850 271187 175856 271199
rect 178288 271187 178294 271199
rect 175850 271159 178294 271187
rect 175850 271147 175856 271159
rect 178288 271147 178294 271159
rect 178346 271147 178352 271199
rect 187600 271147 187606 271199
rect 187658 271187 187664 271199
rect 205840 271187 205846 271199
rect 187658 271159 205846 271187
rect 187658 271147 187664 271159
rect 205840 271147 205846 271159
rect 205898 271147 205904 271199
rect 238480 271147 238486 271199
rect 238538 271187 238544 271199
rect 246064 271187 246070 271199
rect 238538 271159 246070 271187
rect 238538 271147 238544 271159
rect 246064 271147 246070 271159
rect 246122 271147 246128 271199
rect 338608 271147 338614 271199
rect 338666 271187 338672 271199
rect 348592 271187 348598 271199
rect 338666 271159 348598 271187
rect 338666 271147 338672 271159
rect 348592 271147 348598 271159
rect 348650 271147 348656 271199
rect 357904 271147 357910 271199
rect 357962 271187 357968 271199
rect 375184 271187 375190 271199
rect 357962 271159 375190 271187
rect 357962 271147 357968 271159
rect 375184 271147 375190 271159
rect 375242 271147 375248 271199
rect 387280 271147 387286 271199
rect 387338 271187 387344 271199
rect 407440 271187 407446 271199
rect 387338 271159 407446 271187
rect 387338 271147 387344 271159
rect 407440 271147 407446 271159
rect 407498 271147 407504 271199
rect 85936 271073 85942 271125
rect 85994 271113 86000 271125
rect 198544 271113 198550 271125
rect 85994 271085 198550 271113
rect 85994 271073 86000 271085
rect 198544 271073 198550 271085
rect 198602 271073 198608 271125
rect 240784 271073 240790 271125
rect 240842 271113 240848 271125
rect 247216 271113 247222 271125
rect 240842 271085 247222 271113
rect 240842 271073 240848 271085
rect 247216 271073 247222 271085
rect 247274 271073 247280 271125
rect 221872 270999 221878 271051
rect 221930 271039 221936 271051
rect 239344 271039 239350 271051
rect 221930 271011 239350 271039
rect 221930 270999 221936 271011
rect 239344 270999 239350 271011
rect 239402 270999 239408 271051
rect 239536 270999 239542 271051
rect 239594 271039 239600 271051
rect 241264 271039 241270 271051
rect 239594 271011 241270 271039
rect 239594 270999 239600 271011
rect 241264 270999 241270 271011
rect 241322 270999 241328 271051
rect 241936 270999 241942 271051
rect 241994 271039 242000 271051
rect 247696 271039 247702 271051
rect 241994 271011 247702 271039
rect 241994 270999 242000 271011
rect 247696 270999 247702 271011
rect 247754 270999 247760 271051
rect 223024 270925 223030 270977
rect 223082 270965 223088 270977
rect 240016 270965 240022 270977
rect 223082 270937 240022 270965
rect 223082 270925 223088 270937
rect 240016 270925 240022 270937
rect 240074 270925 240080 270977
rect 243184 270925 243190 270977
rect 243242 270965 243248 270977
rect 247984 270965 247990 270977
rect 243242 270937 247990 270965
rect 243242 270925 243248 270937
rect 247984 270925 247990 270937
rect 248042 270925 248048 270977
rect 224272 270851 224278 270903
rect 224330 270891 224336 270903
rect 240496 270891 240502 270903
rect 224330 270863 240502 270891
rect 224330 270851 224336 270863
rect 240496 270851 240502 270863
rect 240554 270851 240560 270903
rect 244336 270851 244342 270903
rect 244394 270891 244400 270903
rect 248656 270891 248662 270903
rect 244394 270863 248662 270891
rect 244394 270851 244400 270863
rect 248656 270851 248662 270863
rect 248714 270851 248720 270903
rect 351376 270851 351382 270903
rect 351434 270891 351440 270903
rect 355408 270891 355414 270903
rect 351434 270863 355414 270891
rect 351434 270851 351440 270863
rect 355408 270851 355414 270863
rect 355466 270851 355472 270903
rect 225424 270777 225430 270829
rect 225482 270817 225488 270829
rect 241072 270817 241078 270829
rect 225482 270789 241078 270817
rect 225482 270777 225488 270789
rect 241072 270777 241078 270789
rect 241130 270777 241136 270829
rect 245488 270777 245494 270829
rect 245546 270817 245552 270829
rect 249136 270817 249142 270829
rect 245546 270789 249142 270817
rect 245546 270777 245552 270789
rect 249136 270777 249142 270789
rect 249194 270777 249200 270829
rect 94192 270703 94198 270755
rect 94250 270743 94256 270755
rect 94960 270743 94966 270755
rect 94250 270715 94966 270743
rect 94250 270703 94256 270715
rect 94960 270703 94966 270715
rect 95018 270703 95024 270755
rect 101296 270703 101302 270755
rect 101354 270743 101360 270755
rect 103600 270743 103606 270755
rect 101354 270715 103606 270743
rect 101354 270703 101360 270715
rect 103600 270703 103606 270715
rect 103658 270703 103664 270755
rect 115504 270703 115510 270755
rect 115562 270743 115568 270755
rect 118000 270743 118006 270755
rect 115562 270715 118006 270743
rect 115562 270703 115568 270715
rect 118000 270703 118006 270715
rect 118058 270703 118064 270755
rect 133264 270703 133270 270755
rect 133322 270743 133328 270755
rect 135280 270743 135286 270755
rect 133322 270715 135286 270743
rect 133322 270703 133328 270715
rect 135280 270703 135286 270715
rect 135338 270703 135344 270755
rect 136816 270703 136822 270755
rect 136874 270743 136880 270755
rect 138160 270743 138166 270755
rect 136874 270715 138166 270743
rect 136874 270703 136880 270715
rect 138160 270703 138166 270715
rect 138218 270703 138224 270755
rect 154480 270703 154486 270755
rect 154538 270743 154544 270755
rect 155440 270743 155446 270755
rect 154538 270715 155446 270743
rect 154538 270703 154544 270715
rect 155440 270703 155446 270715
rect 155498 270703 155504 270755
rect 168688 270703 168694 270755
rect 168746 270743 168752 270755
rect 169840 270743 169846 270755
rect 168746 270715 169846 270743
rect 168746 270703 168752 270715
rect 169840 270703 169846 270715
rect 169898 270703 169904 270755
rect 179344 270703 179350 270755
rect 179402 270743 179408 270755
rect 181360 270743 181366 270755
rect 179402 270715 181366 270743
rect 179402 270703 179408 270715
rect 181360 270703 181366 270715
rect 181418 270703 181424 270755
rect 182896 270703 182902 270755
rect 182954 270743 182960 270755
rect 184240 270743 184246 270755
rect 182954 270715 184246 270743
rect 182954 270703 182960 270715
rect 184240 270703 184246 270715
rect 184298 270703 184304 270755
rect 185488 270703 185494 270755
rect 185546 270743 185552 270755
rect 186448 270743 186454 270755
rect 185546 270715 186454 270743
rect 185546 270703 185552 270715
rect 186448 270703 186454 270715
rect 186506 270703 186512 270755
rect 226576 270703 226582 270755
rect 226634 270743 226640 270755
rect 239536 270743 239542 270755
rect 226634 270715 239542 270743
rect 226634 270703 226640 270715
rect 239536 270703 239542 270715
rect 239594 270703 239600 270755
rect 239632 270703 239638 270755
rect 239690 270743 239696 270755
rect 246448 270743 246454 270755
rect 239690 270715 246454 270743
rect 239690 270703 239696 270715
rect 246448 270703 246454 270715
rect 246506 270703 246512 270755
rect 246736 270703 246742 270755
rect 246794 270743 246800 270755
rect 249616 270743 249622 270755
rect 246794 270715 249622 270743
rect 246794 270703 246800 270715
rect 249616 270703 249622 270715
rect 249674 270703 249680 270755
rect 334096 270703 334102 270755
rect 334154 270743 334160 270755
rect 337744 270743 337750 270755
rect 334154 270715 337750 270743
rect 334154 270703 334160 270715
rect 337744 270703 337750 270715
rect 337802 270703 337808 270755
rect 338128 270703 338134 270755
rect 338186 270743 338192 270755
rect 341296 270743 341302 270755
rect 338186 270715 341302 270743
rect 338186 270703 338192 270715
rect 341296 270703 341302 270715
rect 341354 270703 341360 270755
rect 408976 270703 408982 270755
rect 409034 270743 409040 270755
rect 413392 270743 413398 270755
rect 409034 270715 413398 270743
rect 409034 270703 409040 270715
rect 413392 270703 413398 270715
rect 413450 270703 413456 270755
rect 146224 270629 146230 270681
rect 146282 270669 146288 270681
rect 214960 270669 214966 270681
rect 146282 270641 214966 270669
rect 146282 270629 146288 270641
rect 214960 270629 214966 270641
rect 215018 270629 215024 270681
rect 269200 270629 269206 270681
rect 269258 270669 269264 270681
rect 295120 270669 295126 270681
rect 269258 270641 295126 270669
rect 269258 270629 269264 270641
rect 295120 270629 295126 270641
rect 295178 270629 295184 270681
rect 295216 270629 295222 270681
rect 295274 270669 295280 270681
rect 301072 270669 301078 270681
rect 295274 270641 301078 270669
rect 295274 270629 295280 270641
rect 301072 270629 301078 270641
rect 301130 270629 301136 270681
rect 302416 270629 302422 270681
rect 302474 270669 302480 270681
rect 304624 270669 304630 270681
rect 302474 270641 304630 270669
rect 302474 270629 302480 270641
rect 304624 270629 304630 270641
rect 304682 270629 304688 270681
rect 306352 270629 306358 270681
rect 306410 270669 306416 270681
rect 341968 270669 341974 270681
rect 306410 270641 341974 270669
rect 306410 270629 306416 270641
rect 341968 270629 341974 270641
rect 342026 270629 342032 270681
rect 345424 270629 345430 270681
rect 345482 270669 345488 270681
rect 484240 270669 484246 270681
rect 345482 270641 484246 270669
rect 345482 270629 345488 270641
rect 484240 270629 484246 270641
rect 484298 270629 484304 270681
rect 141520 270555 141526 270607
rect 141578 270595 141584 270607
rect 213808 270595 213814 270607
rect 141578 270567 213814 270595
rect 141578 270555 141584 270567
rect 213808 270555 213814 270567
rect 213866 270555 213872 270607
rect 279280 270555 279286 270607
rect 279338 270595 279344 270607
rect 298192 270595 298198 270607
rect 279338 270567 298198 270595
rect 279338 270555 279344 270567
rect 298192 270555 298198 270567
rect 298250 270555 298256 270607
rect 298384 270555 298390 270607
rect 298442 270595 298448 270607
rect 318832 270595 318838 270607
rect 298442 270567 318838 270595
rect 298442 270555 298448 270567
rect 318832 270555 318838 270567
rect 318890 270555 318896 270607
rect 348112 270555 348118 270607
rect 348170 270595 348176 270607
rect 490192 270595 490198 270607
rect 348170 270567 490198 270595
rect 348170 270555 348176 270567
rect 490192 270555 490198 270567
rect 490250 270555 490256 270607
rect 137968 270481 137974 270533
rect 138026 270521 138032 270533
rect 212656 270521 212662 270533
rect 138026 270493 212662 270521
rect 138026 270481 138032 270493
rect 212656 270481 212662 270493
rect 212714 270481 212720 270533
rect 280144 270481 280150 270533
rect 280202 270521 280208 270533
rect 322384 270521 322390 270533
rect 280202 270493 322390 270521
rect 280202 270481 280208 270493
rect 322384 270481 322390 270493
rect 322442 270481 322448 270533
rect 348400 270481 348406 270533
rect 348458 270521 348464 270533
rect 491344 270521 491350 270533
rect 348458 270493 491350 270521
rect 348458 270481 348464 270493
rect 491344 270481 491350 270493
rect 491402 270481 491408 270533
rect 134416 270407 134422 270459
rect 134474 270447 134480 270459
rect 211888 270447 211894 270459
rect 134474 270419 211894 270447
rect 134474 270407 134480 270419
rect 211888 270407 211894 270419
rect 211946 270407 211952 270459
rect 253936 270407 253942 270459
rect 253994 270447 254000 270459
rect 257296 270447 257302 270459
rect 253994 270419 257302 270447
rect 253994 270407 254000 270419
rect 257296 270407 257302 270419
rect 257354 270407 257360 270459
rect 262960 270407 262966 270459
rect 263018 270447 263024 270459
rect 279760 270447 279766 270459
rect 263018 270419 279766 270447
rect 263018 270407 263024 270419
rect 279760 270407 279766 270419
rect 279818 270407 279824 270459
rect 280624 270407 280630 270459
rect 280682 270447 280688 270459
rect 323536 270447 323542 270459
rect 280682 270419 323542 270447
rect 280682 270407 280688 270419
rect 323536 270407 323542 270419
rect 323594 270407 323600 270459
rect 350704 270407 350710 270459
rect 350762 270447 350768 270459
rect 497296 270447 497302 270459
rect 350762 270419 497302 270447
rect 350762 270407 350768 270419
rect 497296 270407 497302 270419
rect 497354 270407 497360 270459
rect 121456 270333 121462 270385
rect 121514 270373 121520 270385
rect 208336 270373 208342 270385
rect 121514 270345 208342 270373
rect 121514 270333 121520 270345
rect 208336 270333 208342 270345
rect 208394 270333 208400 270385
rect 209584 270333 209590 270385
rect 209642 270373 209648 270385
rect 216880 270373 216886 270385
rect 209642 270345 216886 270373
rect 209642 270333 209648 270345
rect 216880 270333 216886 270345
rect 216938 270333 216944 270385
rect 262480 270333 262486 270385
rect 262538 270373 262544 270385
rect 278608 270373 278614 270385
rect 262538 270345 278614 270373
rect 262538 270333 262544 270345
rect 278608 270333 278614 270345
rect 278666 270333 278672 270385
rect 284176 270333 284182 270385
rect 284234 270373 284240 270385
rect 284234 270345 298142 270373
rect 284234 270333 284240 270345
rect 117904 270259 117910 270311
rect 117962 270299 117968 270311
rect 207568 270299 207574 270311
rect 117962 270271 207574 270299
rect 117962 270259 117968 270271
rect 207568 270259 207574 270271
rect 207626 270259 207632 270311
rect 212560 270259 212566 270311
rect 212618 270299 212624 270311
rect 225520 270299 225526 270311
rect 212618 270271 225526 270299
rect 212618 270259 212624 270271
rect 225520 270259 225526 270271
rect 225578 270259 225584 270311
rect 255280 270259 255286 270311
rect 255338 270299 255344 270311
rect 260848 270299 260854 270311
rect 255338 270271 260854 270299
rect 255338 270259 255344 270271
rect 260848 270259 260854 270271
rect 260906 270259 260912 270311
rect 286288 270259 286294 270311
rect 286346 270299 286352 270311
rect 286346 270271 298046 270299
rect 286346 270259 286352 270271
rect 114352 270185 114358 270237
rect 114410 270225 114416 270237
rect 206416 270225 206422 270237
rect 114410 270197 206422 270225
rect 114410 270185 114416 270197
rect 206416 270185 206422 270197
rect 206474 270185 206480 270237
rect 209776 270185 209782 270237
rect 209834 270225 209840 270237
rect 211408 270225 211414 270237
rect 209834 270197 211414 270225
rect 209834 270185 209840 270197
rect 211408 270185 211414 270197
rect 211466 270185 211472 270237
rect 212752 270185 212758 270237
rect 212810 270225 212816 270237
rect 226672 270225 226678 270237
rect 212810 270197 226678 270225
rect 212810 270185 212816 270197
rect 226672 270185 226678 270197
rect 226730 270185 226736 270237
rect 261232 270185 261238 270237
rect 261290 270225 261296 270237
rect 275056 270225 275062 270237
rect 261290 270197 275062 270225
rect 261290 270185 261296 270197
rect 275056 270185 275062 270197
rect 275114 270185 275120 270237
rect 284464 270185 284470 270237
rect 284522 270225 284528 270237
rect 293968 270225 293974 270237
rect 284522 270197 293974 270225
rect 284522 270185 284528 270197
rect 293968 270185 293974 270197
rect 294026 270185 294032 270237
rect 109552 270111 109558 270163
rect 109610 270151 109616 270163
rect 205264 270151 205270 270163
rect 109610 270123 205270 270151
rect 109610 270111 109616 270123
rect 205264 270111 205270 270123
rect 205322 270111 205328 270163
rect 209872 270111 209878 270163
rect 209930 270151 209936 270163
rect 212368 270151 212374 270163
rect 209930 270123 212374 270151
rect 209930 270111 209936 270123
rect 212368 270111 212374 270123
rect 212426 270111 212432 270163
rect 212848 270111 212854 270163
rect 212906 270151 212912 270163
rect 222832 270151 222838 270163
rect 212906 270123 222838 270151
rect 212906 270111 212912 270123
rect 222832 270111 222838 270123
rect 222890 270111 222896 270163
rect 265360 270111 265366 270163
rect 265418 270151 265424 270163
rect 285712 270151 285718 270163
rect 265418 270123 285718 270151
rect 265418 270111 265424 270123
rect 285712 270111 285718 270123
rect 285770 270111 285776 270163
rect 287920 270111 287926 270163
rect 287978 270151 287984 270163
rect 298018 270151 298046 270271
rect 298114 270225 298142 270345
rect 298192 270333 298198 270385
rect 298250 270373 298256 270385
rect 319984 270373 319990 270385
rect 298250 270345 319990 270373
rect 298250 270333 298256 270345
rect 319984 270333 319990 270345
rect 320042 270333 320048 270385
rect 351280 270333 351286 270385
rect 351338 270373 351344 270385
rect 498448 270373 498454 270385
rect 351338 270345 498454 270373
rect 351338 270333 351344 270345
rect 498448 270333 498454 270345
rect 498506 270333 498512 270385
rect 298288 270259 298294 270311
rect 298346 270299 298352 270311
rect 330640 270299 330646 270311
rect 298346 270271 330646 270299
rect 298346 270259 298352 270271
rect 330640 270259 330646 270271
rect 330698 270259 330704 270311
rect 354064 270259 354070 270311
rect 354122 270299 354128 270311
rect 505552 270299 505558 270311
rect 354122 270271 505558 270299
rect 354122 270259 354128 270271
rect 505552 270259 505558 270271
rect 505610 270259 505616 270311
rect 331792 270225 331798 270237
rect 298114 270197 331798 270225
rect 331792 270185 331798 270197
rect 331850 270185 331856 270237
rect 353680 270185 353686 270237
rect 353738 270225 353744 270237
rect 504400 270225 504406 270237
rect 353738 270197 504406 270225
rect 353738 270185 353744 270197
rect 504400 270185 504406 270197
rect 504458 270185 504464 270237
rect 334096 270151 334102 270163
rect 287978 270123 297854 270151
rect 298018 270123 334102 270151
rect 287978 270111 287984 270123
rect 102544 270037 102550 270089
rect 102602 270077 102608 270089
rect 203344 270077 203350 270089
rect 102602 270049 203350 270077
rect 102602 270037 102608 270049
rect 203344 270037 203350 270049
rect 203402 270037 203408 270089
rect 212944 270037 212950 270089
rect 213002 270077 213008 270089
rect 224752 270077 224758 270089
rect 213002 270049 224758 270077
rect 213002 270037 213008 270049
rect 224752 270037 224758 270049
rect 224810 270037 224816 270089
rect 264688 270037 264694 270089
rect 264746 270077 264752 270089
rect 288016 270077 288022 270089
rect 264746 270049 276494 270077
rect 264746 270037 264752 270049
rect 107248 269963 107254 270015
rect 107306 270003 107312 270015
rect 204688 270003 204694 270015
rect 107306 269975 204694 270003
rect 107306 269963 107312 269975
rect 204688 269963 204694 269975
rect 204746 269963 204752 270015
rect 213040 269963 213046 270015
rect 213098 270003 213104 270015
rect 221008 270003 221014 270015
rect 213098 269975 221014 270003
rect 213098 269963 213104 269975
rect 221008 269963 221014 269975
rect 221066 269963 221072 270015
rect 261808 269963 261814 270015
rect 261866 270003 261872 270015
rect 276208 270003 276214 270015
rect 261866 269975 276214 270003
rect 261866 269963 261872 269975
rect 276208 269963 276214 269975
rect 276266 269963 276272 270015
rect 276466 270003 276494 270049
rect 284674 270049 288022 270077
rect 283312 270003 283318 270015
rect 276466 269975 283318 270003
rect 283312 269963 283318 269975
rect 283370 269963 283376 270015
rect 100144 269889 100150 269941
rect 100202 269929 100208 269941
rect 202864 269929 202870 269941
rect 100202 269901 202870 269929
rect 100202 269889 100208 269901
rect 202864 269889 202870 269901
rect 202922 269889 202928 269941
rect 205936 269889 205942 269941
rect 205994 269929 206000 269941
rect 224080 269929 224086 269941
rect 205994 269901 224086 269929
rect 205994 269889 206000 269901
rect 224080 269889 224086 269901
rect 224138 269889 224144 269941
rect 256240 269889 256246 269941
rect 256298 269929 256304 269941
rect 263248 269929 263254 269941
rect 256298 269901 263254 269929
rect 256298 269889 256304 269901
rect 263248 269889 263254 269901
rect 263306 269889 263312 269941
rect 264880 269889 264886 269941
rect 264938 269929 264944 269941
rect 284560 269929 284566 269941
rect 264938 269901 284566 269929
rect 264938 269889 264944 269901
rect 284560 269889 284566 269901
rect 284618 269889 284624 269941
rect 95440 269815 95446 269867
rect 95498 269855 95504 269867
rect 195184 269855 195190 269867
rect 95498 269827 195190 269855
rect 95498 269815 95504 269827
rect 195184 269815 195190 269827
rect 195242 269815 195248 269867
rect 205840 269815 205846 269867
rect 205898 269855 205904 269867
rect 226000 269855 226006 269867
rect 205898 269827 226006 269855
rect 205898 269815 205904 269827
rect 226000 269815 226006 269827
rect 226058 269815 226064 269867
rect 260560 269815 260566 269867
rect 260618 269855 260624 269867
rect 273904 269855 273910 269867
rect 260618 269827 273910 269855
rect 260618 269815 260624 269827
rect 273904 269815 273910 269827
rect 273962 269815 273968 269867
rect 93040 269741 93046 269793
rect 93098 269781 93104 269793
rect 200944 269781 200950 269793
rect 93098 269753 200950 269781
rect 93098 269741 93104 269753
rect 200944 269741 200950 269753
rect 201002 269741 201008 269793
rect 205744 269741 205750 269793
rect 205802 269781 205808 269793
rect 225232 269781 225238 269793
rect 205802 269753 225238 269781
rect 205802 269741 205808 269753
rect 225232 269741 225238 269753
rect 225290 269741 225296 269793
rect 259888 269741 259894 269793
rect 259946 269781 259952 269793
rect 271504 269781 271510 269793
rect 259946 269753 271510 269781
rect 259946 269741 259952 269753
rect 271504 269741 271510 269753
rect 271562 269741 271568 269793
rect 284464 269781 284470 269793
rect 271618 269753 284470 269781
rect 90640 269667 90646 269719
rect 90698 269707 90704 269719
rect 199696 269707 199702 269719
rect 90698 269679 199702 269707
rect 90698 269667 90704 269679
rect 199696 269667 199702 269679
rect 199754 269667 199760 269719
rect 201520 269667 201526 269719
rect 201578 269707 201584 269719
rect 222352 269707 222358 269719
rect 201578 269679 222358 269707
rect 201578 269667 201584 269679
rect 222352 269667 222358 269679
rect 222410 269667 222416 269719
rect 258160 269667 258166 269719
rect 258218 269707 258224 269719
rect 267952 269707 267958 269719
rect 258218 269679 267958 269707
rect 258218 269667 258224 269679
rect 267952 269667 267958 269679
rect 268010 269667 268016 269719
rect 268624 269667 268630 269719
rect 268682 269707 268688 269719
rect 271618 269707 271646 269753
rect 284464 269741 284470 269753
rect 284522 269741 284528 269793
rect 268682 269679 271646 269707
rect 268682 269667 268688 269679
rect 271696 269667 271702 269719
rect 271754 269707 271760 269719
rect 284674 269707 284702 270049
rect 288016 270037 288022 270049
rect 288074 270037 288080 270089
rect 286480 269963 286486 270015
rect 286538 270003 286544 270015
rect 295216 270003 295222 270015
rect 286538 269975 295222 270003
rect 286538 269963 286544 269975
rect 295216 269963 295222 269975
rect 295274 269963 295280 270015
rect 297826 270003 297854 270123
rect 334096 270111 334102 270123
rect 334154 270111 334160 270163
rect 356752 270111 356758 270163
rect 356810 270151 356816 270163
rect 511504 270151 511510 270163
rect 356810 270123 511510 270151
rect 356810 270111 356816 270123
rect 511504 270111 511510 270123
rect 511562 270111 511568 270163
rect 298192 270037 298198 270089
rect 298250 270077 298256 270089
rect 342448 270077 342454 270089
rect 298250 270049 342454 270077
rect 298250 270037 298256 270049
rect 342448 270037 342454 270049
rect 342506 270037 342512 270089
rect 356944 270037 356950 270089
rect 357002 270077 357008 270089
rect 512656 270077 512662 270089
rect 357002 270049 512662 270077
rect 357002 270037 357008 270049
rect 512656 270037 512662 270049
rect 512714 270037 512720 270089
rect 338128 270003 338134 270015
rect 297826 269975 338134 270003
rect 338128 269963 338134 269975
rect 338186 269963 338192 270015
rect 359344 269963 359350 270015
rect 359402 270003 359408 270015
rect 518512 270003 518518 270015
rect 359402 269975 518518 270003
rect 359402 269963 359408 269975
rect 518512 269963 518518 269975
rect 518570 269963 518576 270015
rect 290608 269889 290614 269941
rect 290666 269929 290672 269941
rect 342736 269929 342742 269941
rect 290666 269901 342742 269929
rect 290666 269889 290672 269901
rect 342736 269889 342742 269901
rect 342794 269889 342800 269941
rect 359824 269889 359830 269941
rect 359882 269929 359888 269941
rect 519760 269929 519766 269941
rect 359882 269901 519766 269929
rect 359882 269889 359888 269901
rect 519760 269889 519766 269901
rect 519818 269889 519824 269941
rect 291088 269815 291094 269867
rect 291146 269855 291152 269867
rect 349552 269855 349558 269867
rect 291146 269827 349558 269855
rect 291146 269815 291152 269827
rect 349552 269815 349558 269827
rect 349610 269815 349616 269867
rect 362224 269815 362230 269867
rect 362282 269855 362288 269867
rect 525616 269855 525622 269867
rect 362282 269827 525622 269855
rect 362282 269815 362288 269827
rect 525616 269815 525622 269827
rect 525674 269815 525680 269867
rect 293968 269741 293974 269793
rect 294026 269781 294032 269793
rect 356656 269781 356662 269793
rect 294026 269753 356662 269781
rect 294026 269741 294032 269753
rect 356656 269741 356662 269753
rect 356714 269741 356720 269793
rect 362800 269741 362806 269793
rect 362858 269781 362864 269793
rect 526864 269781 526870 269793
rect 362858 269753 526870 269781
rect 362858 269741 362864 269753
rect 526864 269741 526870 269753
rect 526922 269741 526928 269793
rect 271754 269679 284702 269707
rect 271754 269667 271760 269679
rect 293488 269667 293494 269719
rect 293546 269707 293552 269719
rect 351376 269707 351382 269719
rect 293546 269679 351382 269707
rect 293546 269667 293552 269679
rect 351376 269667 351382 269679
rect 351434 269667 351440 269719
rect 365296 269667 365302 269719
rect 365354 269707 365360 269719
rect 532720 269707 532726 269719
rect 365354 269679 532726 269707
rect 365354 269667 365360 269679
rect 532720 269667 532726 269679
rect 532778 269667 532784 269719
rect 83632 269593 83638 269645
rect 83690 269633 83696 269645
rect 83690 269605 195854 269633
rect 83690 269593 83696 269605
rect 87184 269519 87190 269571
rect 87242 269559 87248 269571
rect 185680 269559 185686 269571
rect 87242 269531 185686 269559
rect 87242 269519 87248 269531
rect 185680 269519 185686 269531
rect 185738 269519 185744 269571
rect 195826 269559 195854 269605
rect 196336 269593 196342 269645
rect 196394 269633 196400 269645
rect 220528 269633 220534 269645
rect 196394 269605 220534 269633
rect 196394 269593 196400 269605
rect 220528 269593 220534 269605
rect 220586 269593 220592 269645
rect 249040 269593 249046 269645
rect 249098 269633 249104 269645
rect 250288 269633 250294 269645
rect 249098 269605 250294 269633
rect 249098 269593 249104 269605
rect 250288 269593 250294 269605
rect 250346 269593 250352 269645
rect 255760 269593 255766 269645
rect 255818 269633 255824 269645
rect 262096 269633 262102 269645
rect 255818 269605 262102 269633
rect 255818 269593 255824 269605
rect 262096 269593 262102 269605
rect 262154 269593 262160 269645
rect 267760 269593 267766 269645
rect 267818 269633 267824 269645
rect 291568 269633 291574 269645
rect 267818 269605 291574 269633
rect 267818 269593 267824 269605
rect 291568 269593 291574 269605
rect 291626 269593 291632 269645
rect 297040 269593 297046 269645
rect 297098 269633 297104 269645
rect 363664 269633 363670 269645
rect 297098 269605 363670 269633
rect 297098 269593 297104 269605
rect 363664 269593 363670 269605
rect 363722 269593 363728 269645
rect 198064 269559 198070 269571
rect 195826 269531 198070 269559
rect 198064 269519 198070 269531
rect 198122 269519 198128 269571
rect 206512 269519 206518 269571
rect 206570 269559 206576 269571
rect 233392 269559 233398 269571
rect 206570 269531 233398 269559
rect 206570 269519 206576 269531
rect 233392 269519 233398 269531
rect 233450 269519 233456 269571
rect 258640 269519 258646 269571
rect 258698 269559 258704 269571
rect 269104 269559 269110 269571
rect 258698 269531 269110 269559
rect 258698 269519 258704 269531
rect 269104 269519 269110 269531
rect 269162 269519 269168 269571
rect 271504 269519 271510 269571
rect 271562 269559 271568 269571
rect 286480 269559 286486 269571
rect 271562 269531 286486 269559
rect 271562 269519 271568 269531
rect 286480 269519 286486 269531
rect 286538 269519 286544 269571
rect 288496 269519 288502 269571
rect 288554 269559 288560 269571
rect 298192 269559 298198 269571
rect 288554 269531 298198 269559
rect 288554 269519 288560 269531
rect 298192 269519 298198 269531
rect 298250 269519 298256 269571
rect 299632 269519 299638 269571
rect 299690 269559 299696 269571
rect 370768 269559 370774 269571
rect 299690 269531 370774 269559
rect 299690 269519 299696 269531
rect 370768 269519 370774 269531
rect 370826 269519 370832 269571
rect 371248 269519 371254 269571
rect 371306 269559 371312 269571
rect 548080 269559 548086 269571
rect 371306 269531 548086 269559
rect 371306 269519 371312 269531
rect 548080 269519 548086 269531
rect 548138 269519 548144 269571
rect 81232 269445 81238 269497
rect 81290 269485 81296 269497
rect 196816 269485 196822 269497
rect 81290 269457 196822 269485
rect 81290 269445 81296 269457
rect 196816 269445 196822 269457
rect 196874 269445 196880 269497
rect 204112 269445 204118 269497
rect 204170 269485 204176 269497
rect 232144 269485 232150 269497
rect 204170 269457 232150 269485
rect 204170 269445 204176 269457
rect 232144 269445 232150 269457
rect 232202 269445 232208 269497
rect 260080 269445 260086 269497
rect 260138 269485 260144 269497
rect 272656 269485 272662 269497
rect 260138 269457 272662 269485
rect 260138 269445 260144 269457
rect 272656 269445 272662 269457
rect 272714 269445 272720 269497
rect 272944 269445 272950 269497
rect 273002 269485 273008 269497
rect 302416 269485 302422 269497
rect 273002 269457 302422 269485
rect 273002 269445 273008 269457
rect 302416 269445 302422 269457
rect 302474 269445 302480 269497
rect 302608 269445 302614 269497
rect 302666 269485 302672 269497
rect 377872 269485 377878 269497
rect 302666 269457 377878 269485
rect 302666 269445 302672 269457
rect 377872 269445 377878 269457
rect 377930 269445 377936 269497
rect 379888 269445 379894 269497
rect 379946 269485 379952 269497
rect 569392 269485 569398 269497
rect 379946 269457 569398 269485
rect 379946 269445 379952 269457
rect 569392 269445 569398 269457
rect 569450 269445 569456 269497
rect 82384 269371 82390 269423
rect 82442 269411 82448 269423
rect 197392 269411 197398 269423
rect 82442 269383 197398 269411
rect 82442 269371 82448 269383
rect 197392 269371 197398 269383
rect 197450 269371 197456 269423
rect 202960 269371 202966 269423
rect 203018 269411 203024 269423
rect 231952 269411 231958 269423
rect 203018 269383 231958 269411
rect 203018 269371 203024 269383
rect 231952 269371 231958 269383
rect 232010 269371 232016 269423
rect 266512 269371 266518 269423
rect 266570 269411 266576 269423
rect 271696 269411 271702 269423
rect 266570 269383 271702 269411
rect 266570 269371 266576 269383
rect 271696 269371 271702 269383
rect 271754 269371 271760 269423
rect 274672 269371 274678 269423
rect 274730 269411 274736 269423
rect 308176 269411 308182 269423
rect 274730 269383 308182 269411
rect 274730 269371 274736 269383
rect 308176 269371 308182 269383
rect 308234 269371 308240 269423
rect 308272 269371 308278 269423
rect 308330 269411 308336 269423
rect 392080 269411 392086 269423
rect 308330 269383 392086 269411
rect 308330 269371 308336 269383
rect 392080 269371 392086 269383
rect 392138 269371 392144 269423
rect 394384 269371 394390 269423
rect 394442 269411 394448 269423
rect 604816 269411 604822 269423
rect 394442 269383 604822 269411
rect 394442 269371 394448 269383
rect 604816 269371 604822 269383
rect 604874 269371 604880 269423
rect 74128 269297 74134 269349
rect 74186 269337 74192 269349
rect 185584 269337 185590 269349
rect 74186 269309 185590 269337
rect 74186 269297 74192 269309
rect 185584 269297 185590 269309
rect 185642 269297 185648 269349
rect 185680 269297 185686 269349
rect 185738 269337 185744 269349
rect 199024 269337 199030 269349
rect 185738 269309 199030 269337
rect 185738 269297 185744 269309
rect 199024 269297 199030 269309
rect 199082 269297 199088 269349
rect 200656 269297 200662 269349
rect 200714 269337 200720 269349
rect 230992 269337 230998 269349
rect 200714 269309 230998 269337
rect 200714 269297 200720 269309
rect 230992 269297 230998 269309
rect 231050 269297 231056 269349
rect 257680 269297 257686 269349
rect 257738 269337 257744 269349
rect 266800 269337 266806 269349
rect 257738 269309 266806 269337
rect 257738 269297 257744 269309
rect 266800 269297 266806 269309
rect 266858 269297 266864 269349
rect 266914 269309 275198 269337
rect 67024 269223 67030 269275
rect 67082 269263 67088 269275
rect 192592 269263 192598 269275
rect 67082 269235 192598 269263
rect 67082 269223 67088 269235
rect 192592 269223 192598 269235
rect 192650 269223 192656 269275
rect 197104 269223 197110 269275
rect 197162 269263 197168 269275
rect 229552 269263 229558 269275
rect 197162 269235 229558 269263
rect 197162 269223 197168 269235
rect 229552 269223 229558 269235
rect 229610 269223 229616 269275
rect 145072 269149 145078 269201
rect 145130 269189 145136 269201
rect 214480 269189 214486 269201
rect 145130 269161 214486 269189
rect 145130 269149 145136 269161
rect 214480 269149 214486 269161
rect 214538 269149 214544 269201
rect 262000 269149 262006 269201
rect 262058 269189 262064 269201
rect 266914 269189 266942 269309
rect 275170 269263 275198 269309
rect 275824 269297 275830 269349
rect 275882 269337 275888 269349
rect 275882 269309 308174 269337
rect 275882 269297 275888 269309
rect 277456 269263 277462 269275
rect 275170 269235 277462 269263
rect 277456 269223 277462 269235
rect 277514 269223 277520 269275
rect 283696 269223 283702 269275
rect 283754 269263 283760 269275
rect 298288 269263 298294 269275
rect 283754 269235 298294 269263
rect 283754 269223 283760 269235
rect 298288 269223 298294 269235
rect 298346 269223 298352 269275
rect 308146 269263 308174 269309
rect 311152 269297 311158 269349
rect 311210 269337 311216 269349
rect 399184 269337 399190 269349
rect 311210 269309 399190 269337
rect 311210 269297 311216 269309
rect 399184 269297 399190 269309
rect 399242 269297 399248 269349
rect 399952 269297 399958 269349
rect 400010 269337 400016 269349
rect 619024 269337 619030 269349
rect 400010 269309 619030 269337
rect 400010 269297 400016 269309
rect 619024 269297 619030 269309
rect 619082 269297 619088 269349
rect 311728 269263 311734 269275
rect 308146 269235 311734 269263
rect 311728 269223 311734 269235
rect 311786 269223 311792 269275
rect 314224 269223 314230 269275
rect 314282 269263 314288 269275
rect 406288 269263 406294 269275
rect 314282 269235 406294 269263
rect 314282 269223 314288 269235
rect 406288 269223 406294 269235
rect 406346 269223 406352 269275
rect 406576 269223 406582 269275
rect 406634 269263 406640 269275
rect 408592 269263 408598 269275
rect 406634 269235 408598 269263
rect 406634 269223 406640 269235
rect 408592 269223 408598 269235
rect 408650 269223 408656 269275
rect 262058 269161 266942 269189
rect 262058 269149 262064 269161
rect 269680 269149 269686 269201
rect 269738 269189 269744 269201
rect 296368 269189 296374 269201
rect 269738 269161 296374 269189
rect 269738 269149 269744 269161
rect 296368 269149 296374 269161
rect 296426 269149 296432 269201
rect 303760 269149 303766 269201
rect 303818 269189 303824 269201
rect 334288 269189 334294 269201
rect 303818 269161 334294 269189
rect 303818 269149 303824 269161
rect 334288 269149 334294 269161
rect 334346 269149 334352 269201
rect 345232 269149 345238 269201
rect 345290 269189 345296 269201
rect 483088 269189 483094 269201
rect 345290 269161 483094 269189
rect 345290 269149 345296 269161
rect 483088 269149 483094 269161
rect 483146 269149 483152 269201
rect 148624 269075 148630 269127
rect 148682 269115 148688 269127
rect 215728 269115 215734 269127
rect 148682 269087 215734 269115
rect 148682 269075 148688 269087
rect 215728 269075 215734 269087
rect 215786 269075 215792 269127
rect 253360 269075 253366 269127
rect 253418 269115 253424 269127
rect 256144 269115 256150 269127
rect 253418 269087 256150 269115
rect 253418 269075 253424 269087
rect 256144 269075 256150 269087
rect 256202 269075 256208 269127
rect 266032 269075 266038 269127
rect 266090 269115 266096 269127
rect 286864 269115 286870 269127
rect 266090 269087 286870 269115
rect 266090 269075 266096 269087
rect 286864 269075 286870 269087
rect 286922 269075 286928 269127
rect 302032 269075 302038 269127
rect 302090 269115 302096 269127
rect 331216 269115 331222 269127
rect 302090 269087 331222 269115
rect 302090 269075 302096 269087
rect 331216 269075 331222 269087
rect 331274 269075 331280 269127
rect 342640 269075 342646 269127
rect 342698 269115 342704 269127
rect 477136 269115 477142 269127
rect 342698 269087 477142 269115
rect 342698 269075 342704 269087
rect 477136 269075 477142 269087
rect 477194 269075 477200 269127
rect 149776 269001 149782 269053
rect 149834 269041 149840 269053
rect 216208 269041 216214 269053
rect 149834 269013 216214 269041
rect 149834 269001 149840 269013
rect 216208 269001 216214 269013
rect 216266 269001 216272 269053
rect 281296 269001 281302 269053
rect 281354 269041 281360 269053
rect 300112 269041 300118 269053
rect 281354 269013 300118 269041
rect 281354 269001 281360 269013
rect 300112 269001 300118 269013
rect 300170 269001 300176 269053
rect 384112 269001 384118 269053
rect 384170 269041 384176 269053
rect 516304 269041 516310 269053
rect 384170 269013 516310 269041
rect 384170 269001 384176 269013
rect 516304 269001 516310 269013
rect 516362 269001 516368 269053
rect 152176 268927 152182 268979
rect 152234 268967 152240 268979
rect 216688 268967 216694 268979
rect 152234 268939 216694 268967
rect 152234 268927 152240 268939
rect 216688 268927 216694 268939
rect 216746 268927 216752 268979
rect 259408 268927 259414 268979
rect 259466 268967 259472 268979
rect 270352 268967 270358 268979
rect 259466 268939 270358 268967
rect 259466 268927 259472 268939
rect 270352 268927 270358 268939
rect 270410 268927 270416 268979
rect 281008 268967 281014 268979
rect 276466 268939 281014 268967
rect 155728 268853 155734 268905
rect 155786 268893 155792 268905
rect 217360 268893 217366 268905
rect 155786 268865 217366 268893
rect 155786 268853 155792 268865
rect 217360 268853 217366 268865
rect 217418 268853 217424 268905
rect 263632 268853 263638 268905
rect 263690 268893 263696 268905
rect 276466 268893 276494 268939
rect 281008 268927 281014 268939
rect 281066 268927 281072 268979
rect 282064 268927 282070 268979
rect 282122 268967 282128 268979
rect 298096 268967 298102 268979
rect 282122 268939 298102 268967
rect 282122 268927 282128 268939
rect 298096 268927 298102 268939
rect 298154 268927 298160 268979
rect 300688 268927 300694 268979
rect 300746 268967 300752 268979
rect 326128 268967 326134 268979
rect 300746 268939 326134 268967
rect 300746 268927 300752 268939
rect 326128 268927 326134 268939
rect 326186 268927 326192 268979
rect 339760 268927 339766 268979
rect 339818 268967 339824 268979
rect 470128 268967 470134 268979
rect 339818 268939 470134 268967
rect 339818 268927 339824 268939
rect 470128 268927 470134 268939
rect 470186 268927 470192 268979
rect 298384 268893 298390 268905
rect 263690 268865 276494 268893
rect 287986 268865 298390 268893
rect 263690 268853 263696 268865
rect 156880 268779 156886 268831
rect 156938 268819 156944 268831
rect 218128 268819 218134 268831
rect 156938 268791 218134 268819
rect 156938 268779 156944 268791
rect 218128 268779 218134 268791
rect 218186 268779 218192 268831
rect 257488 268779 257494 268831
rect 257546 268819 257552 268831
rect 265648 268819 265654 268831
rect 257546 268791 265654 268819
rect 257546 268779 257552 268791
rect 265648 268779 265654 268791
rect 265706 268779 265712 268831
rect 278896 268779 278902 268831
rect 278954 268819 278960 268831
rect 287986 268819 288014 268865
rect 298384 268853 298390 268865
rect 298442 268853 298448 268905
rect 336880 268853 336886 268905
rect 336938 268893 336944 268905
rect 463024 268893 463030 268905
rect 336938 268865 463030 268893
rect 336938 268853 336944 268865
rect 463024 268853 463030 268865
rect 463082 268853 463088 268905
rect 278954 268791 288014 268819
rect 278954 268779 278960 268791
rect 289168 268779 289174 268831
rect 289226 268819 289232 268831
rect 310576 268819 310582 268831
rect 289226 268791 310582 268819
rect 289226 268779 289232 268791
rect 310576 268779 310582 268791
rect 310634 268779 310640 268831
rect 334288 268779 334294 268831
rect 334346 268819 334352 268831
rect 455920 268819 455926 268831
rect 334346 268791 455926 268819
rect 334346 268779 334352 268791
rect 455920 268779 455926 268791
rect 455978 268779 455984 268831
rect 162832 268705 162838 268757
rect 162890 268745 162896 268757
rect 219280 268745 219286 268757
rect 162890 268717 219286 268745
rect 162890 268705 162896 268717
rect 219280 268705 219286 268717
rect 219338 268705 219344 268757
rect 268432 268705 268438 268757
rect 268490 268745 268496 268757
rect 292816 268745 292822 268757
rect 268490 268717 292822 268745
rect 268490 268705 268496 268717
rect 292816 268705 292822 268717
rect 292874 268705 292880 268757
rect 295216 268705 295222 268757
rect 295274 268745 295280 268757
rect 307024 268745 307030 268757
rect 295274 268717 307030 268745
rect 295274 268705 295280 268717
rect 307024 268705 307030 268717
rect 307082 268705 307088 268757
rect 331216 268705 331222 268757
rect 331274 268745 331280 268757
rect 448816 268745 448822 268757
rect 331274 268717 448822 268745
rect 331274 268705 331280 268717
rect 448816 268705 448822 268717
rect 448874 268705 448880 268757
rect 163984 268631 163990 268683
rect 164042 268671 164048 268683
rect 219952 268671 219958 268683
rect 164042 268643 219958 268671
rect 164042 268631 164048 268643
rect 219952 268631 219958 268643
rect 220010 268631 220016 268683
rect 254608 268631 254614 268683
rect 254666 268671 254672 268683
rect 258544 268671 258550 268683
rect 254666 268643 258550 268671
rect 254666 268631 254672 268643
rect 258544 268631 258550 268643
rect 258602 268631 258608 268683
rect 277552 268631 277558 268683
rect 277610 268671 277616 268683
rect 315280 268671 315286 268683
rect 277610 268643 315286 268671
rect 277610 268631 277616 268643
rect 315280 268631 315286 268643
rect 315338 268631 315344 268683
rect 328336 268631 328342 268683
rect 328394 268671 328400 268683
rect 441712 268671 441718 268683
rect 328394 268643 441718 268671
rect 328394 268631 328400 268643
rect 441712 268631 441718 268643
rect 441770 268631 441776 268683
rect 42160 268557 42166 268609
rect 42218 268597 42224 268609
rect 48208 268597 48214 268609
rect 42218 268569 48214 268597
rect 42218 268557 42224 268569
rect 48208 268557 48214 268569
rect 48266 268557 48272 268609
rect 171088 268557 171094 268609
rect 171146 268597 171152 268609
rect 221776 268597 221782 268609
rect 171146 268569 221782 268597
rect 171146 268557 171152 268569
rect 221776 268557 221782 268569
rect 221834 268557 221840 268609
rect 266800 268557 266806 268609
rect 266858 268597 266864 268609
rect 289264 268597 289270 268609
rect 266858 268569 289270 268597
rect 266858 268557 266864 268569
rect 289264 268557 289270 268569
rect 289322 268557 289328 268609
rect 325744 268557 325750 268609
rect 325802 268597 325808 268609
rect 434608 268597 434614 268609
rect 325802 268569 434614 268597
rect 325802 268557 325808 268569
rect 434608 268557 434614 268569
rect 434666 268557 434672 268609
rect 169744 268483 169750 268535
rect 169802 268523 169808 268535
rect 221200 268523 221206 268535
rect 169802 268495 221206 268523
rect 169802 268483 169808 268495
rect 221200 268483 221206 268495
rect 221258 268483 221264 268535
rect 253168 268483 253174 268535
rect 253226 268523 253232 268535
rect 254992 268523 254998 268535
rect 253226 268495 254998 268523
rect 253226 268483 253232 268495
rect 254992 268483 254998 268495
rect 255050 268483 255056 268535
rect 257008 268483 257014 268535
rect 257066 268523 257072 268535
rect 264400 268523 264406 268535
rect 257066 268495 264406 268523
rect 257066 268483 257072 268495
rect 264400 268483 264406 268495
rect 264458 268483 264464 268535
rect 267280 268483 267286 268535
rect 267338 268523 267344 268535
rect 290416 268523 290422 268535
rect 267338 268495 290422 268523
rect 267338 268483 267344 268495
rect 290416 268483 290422 268495
rect 290474 268483 290480 268535
rect 322576 268483 322582 268535
rect 322634 268523 322640 268535
rect 427504 268523 427510 268535
rect 322634 268495 427510 268523
rect 322634 268483 322640 268495
rect 427504 268483 427510 268495
rect 427562 268483 427568 268535
rect 185584 268409 185590 268461
rect 185642 268449 185648 268461
rect 194992 268449 194998 268461
rect 185642 268421 194998 268449
rect 185642 268409 185648 268421
rect 194992 268409 194998 268421
rect 195050 268409 195056 268461
rect 223408 268449 223414 268461
rect 195106 268421 223414 268449
rect 176944 268261 176950 268313
rect 177002 268301 177008 268313
rect 195106 268301 195134 268421
rect 223408 268409 223414 268421
rect 223466 268409 223472 268461
rect 319696 268409 319702 268461
rect 319754 268449 319760 268461
rect 420496 268449 420502 268461
rect 319754 268421 420502 268449
rect 319754 268409 319760 268421
rect 420496 268409 420502 268421
rect 420554 268409 420560 268461
rect 195184 268335 195190 268387
rect 195242 268375 195248 268387
rect 201136 268375 201142 268387
rect 195242 268347 201142 268375
rect 195242 268335 195248 268347
rect 201136 268335 201142 268347
rect 201194 268335 201200 268387
rect 219088 268335 219094 268387
rect 219146 268375 219152 268387
rect 219146 268347 227534 268375
rect 219146 268335 219152 268347
rect 223600 268301 223606 268313
rect 177002 268273 195134 268301
rect 195202 268273 223606 268301
rect 177002 268261 177008 268273
rect 178192 268113 178198 268165
rect 178250 268153 178256 268165
rect 195202 268153 195230 268273
rect 223600 268261 223606 268273
rect 223658 268261 223664 268313
rect 227506 268301 227534 268347
rect 247888 268335 247894 268387
rect 247946 268375 247952 268387
rect 249808 268375 249814 268387
rect 247946 268347 249814 268375
rect 247946 268335 247952 268347
rect 249808 268335 249814 268347
rect 249866 268335 249872 268387
rect 255088 268335 255094 268387
rect 255146 268375 255152 268387
rect 259696 268375 259702 268387
rect 255146 268347 259702 268375
rect 255146 268335 255152 268347
rect 259696 268335 259702 268347
rect 259754 268335 259760 268387
rect 317104 268335 317110 268387
rect 317162 268375 317168 268387
rect 408976 268375 408982 268387
rect 317162 268347 408982 268375
rect 317162 268335 317168 268347
rect 408976 268335 408982 268347
rect 409034 268335 409040 268387
rect 227824 268301 227830 268313
rect 227506 268273 227830 268301
rect 227824 268261 227830 268273
rect 227882 268261 227888 268313
rect 312304 268261 312310 268313
rect 312362 268301 312368 268313
rect 348496 268301 348502 268313
rect 312362 268273 348502 268301
rect 312362 268261 312368 268273
rect 348496 268261 348502 268273
rect 348554 268261 348560 268313
rect 195280 268187 195286 268239
rect 195338 268227 195344 268239
rect 218608 268227 218614 268239
rect 195338 268199 218614 268227
rect 195338 268187 195344 268199
rect 218608 268187 218614 268199
rect 218666 268187 218672 268239
rect 222064 268187 222070 268239
rect 222122 268227 222128 268239
rect 230032 268227 230038 268239
rect 222122 268199 230038 268227
rect 222122 268187 222128 268199
rect 230032 268187 230038 268199
rect 230090 268187 230096 268239
rect 309232 268187 309238 268239
rect 309290 268227 309296 268239
rect 347056 268227 347062 268239
rect 309290 268199 347062 268227
rect 309290 268187 309296 268199
rect 347056 268187 347062 268199
rect 347114 268187 347120 268239
rect 408496 268187 408502 268239
rect 408554 268227 408560 268239
rect 640336 268227 640342 268239
rect 408554 268199 640342 268227
rect 408554 268187 408560 268199
rect 640336 268187 640342 268199
rect 640394 268187 640400 268239
rect 210736 268153 210742 268165
rect 178250 268125 195230 268153
rect 195826 268125 210742 268153
rect 178250 268113 178256 268125
rect 190096 268039 190102 268091
rect 190154 268079 190160 268091
rect 195826 268079 195854 268125
rect 210736 268113 210742 268125
rect 210794 268113 210800 268165
rect 221968 268113 221974 268165
rect 222026 268153 222032 268165
rect 231472 268153 231478 268165
rect 222026 268125 231478 268153
rect 222026 268113 222032 268125
rect 231472 268113 231478 268125
rect 231530 268113 231536 268165
rect 305680 268113 305686 268165
rect 305738 268153 305744 268165
rect 384976 268153 384982 268165
rect 305738 268125 384982 268153
rect 305738 268113 305744 268125
rect 384976 268113 384982 268125
rect 385034 268113 385040 268165
rect 190154 268051 195854 268079
rect 190154 268039 190160 268051
rect 218896 268039 218902 268091
rect 218954 268079 218960 268091
rect 230512 268079 230518 268091
rect 218954 268051 230518 268079
rect 218954 268039 218960 268051
rect 230512 268039 230518 268051
rect 230570 268039 230576 268091
rect 252688 268039 252694 268091
rect 252746 268079 252752 268091
rect 253744 268079 253750 268091
rect 252746 268051 253750 268079
rect 252746 268039 252752 268051
rect 253744 268039 253750 268051
rect 253802 268039 253808 268091
rect 264112 268039 264118 268091
rect 264170 268079 264176 268091
rect 282160 268079 282166 268091
rect 264170 268051 282166 268079
rect 264170 268039 264176 268051
rect 282160 268039 282166 268051
rect 282218 268039 282224 268091
rect 342160 268039 342166 268091
rect 342218 268079 342224 268091
rect 359440 268079 359446 268091
rect 342218 268051 359446 268079
rect 342218 268039 342224 268051
rect 359440 268039 359446 268051
rect 359498 268039 359504 268091
rect 365680 268039 365686 268091
rect 365738 268079 365744 268091
rect 533872 268079 533878 268091
rect 365738 268051 533878 268079
rect 365738 268039 365744 268051
rect 533872 268039 533878 268051
rect 533930 268039 533936 268091
rect 218992 267965 218998 268017
rect 219050 268005 219056 268017
rect 229072 268005 229078 268017
rect 219050 267977 229078 268005
rect 219050 267965 219056 267977
rect 229072 267965 229078 267977
rect 229130 267965 229136 268017
rect 336688 267965 336694 268017
rect 336746 268005 336752 268017
rect 354256 268005 354262 268017
rect 336746 267977 354262 268005
rect 336746 267965 336752 267977
rect 354256 267965 354262 267977
rect 354314 267965 354320 268017
rect 209392 267891 209398 267943
rect 209450 267931 209456 267943
rect 218896 267931 218902 267943
rect 209450 267903 218902 267931
rect 209450 267891 209456 267903
rect 218896 267891 218902 267903
rect 218954 267891 218960 267943
rect 222256 267891 222262 267943
rect 222314 267931 222320 267943
rect 228400 267931 228406 267943
rect 222314 267903 228406 267931
rect 222314 267891 222320 267903
rect 228400 267891 228406 267903
rect 228458 267891 228464 267943
rect 333616 267891 333622 267943
rect 333674 267931 333680 267943
rect 351376 267931 351382 267943
rect 333674 267903 351382 267931
rect 333674 267891 333680 267903
rect 351376 267891 351382 267903
rect 351434 267891 351440 267943
rect 199120 267817 199126 267869
rect 199178 267857 199184 267869
rect 202288 267857 202294 267869
rect 199178 267829 202294 267857
rect 199178 267817 199184 267829
rect 202288 267817 202294 267829
rect 202346 267817 202352 267869
rect 207280 267817 207286 267869
rect 207338 267857 207344 267869
rect 209488 267857 209494 267869
rect 207338 267829 209494 267857
rect 207338 267817 207344 267829
rect 209488 267817 209494 267829
rect 209546 267817 209552 267869
rect 222160 267817 222166 267869
rect 222218 267857 222224 267869
rect 227632 267857 227638 267869
rect 222218 267829 227638 267857
rect 222218 267817 222224 267829
rect 227632 267817 227638 267829
rect 227690 267817 227696 267869
rect 282544 267817 282550 267869
rect 282602 267857 282608 267869
rect 298000 267857 298006 267869
rect 282602 267829 298006 267857
rect 282602 267817 282608 267829
rect 298000 267817 298006 267829
rect 298058 267817 298064 267869
rect 339280 267817 339286 267869
rect 339338 267857 339344 267869
rect 360400 267857 360406 267869
rect 339338 267829 360406 267857
rect 339338 267817 339344 267829
rect 360400 267817 360406 267829
rect 360458 267817 360464 267869
rect 401296 267817 401302 267869
rect 401354 267857 401360 267869
rect 402832 267857 402838 267869
rect 401354 267829 402838 267857
rect 401354 267817 401360 267829
rect 402832 267817 402838 267829
rect 402890 267817 402896 267869
rect 409936 267817 409942 267869
rect 409994 267857 410000 267869
rect 413680 267857 413686 267869
rect 409994 267829 413686 267857
rect 409994 267817 410000 267829
rect 413680 267817 413686 267829
rect 413738 267817 413744 267869
rect 351952 267743 351958 267795
rect 352010 267783 352016 267795
rect 499600 267783 499606 267795
rect 352010 267755 499606 267783
rect 352010 267743 352016 267755
rect 499600 267743 499606 267755
rect 499658 267743 499664 267795
rect 354832 267669 354838 267721
rect 354890 267709 354896 267721
rect 506704 267709 506710 267721
rect 354890 267681 506710 267709
rect 354890 267669 354896 267681
rect 506704 267669 506710 267681
rect 506762 267669 506768 267721
rect 357424 267595 357430 267647
rect 357482 267635 357488 267647
rect 513808 267635 513814 267647
rect 357482 267607 513814 267635
rect 357482 267595 357488 267607
rect 513808 267595 513814 267607
rect 513866 267595 513872 267647
rect 360304 267521 360310 267573
rect 360362 267561 360368 267573
rect 520912 267561 520918 267573
rect 360362 267533 520918 267561
rect 360362 267521 360368 267533
rect 520912 267521 520918 267533
rect 520970 267521 520976 267573
rect 363376 267447 363382 267499
rect 363434 267487 363440 267499
rect 528016 267487 528022 267499
rect 363434 267459 528022 267487
rect 363434 267447 363440 267459
rect 528016 267447 528022 267459
rect 528074 267447 528080 267499
rect 365968 267373 365974 267425
rect 366026 267413 366032 267425
rect 535120 267413 535126 267425
rect 366026 267385 535126 267413
rect 366026 267373 366032 267385
rect 535120 267373 535126 267385
rect 535178 267373 535184 267425
rect 368944 267299 368950 267351
rect 369002 267339 369008 267351
rect 542224 267339 542230 267351
rect 369002 267311 542230 267339
rect 369002 267299 369008 267311
rect 542224 267299 542230 267311
rect 542282 267299 542288 267351
rect 372496 267225 372502 267277
rect 372554 267265 372560 267277
rect 550480 267265 550486 267277
rect 372554 267237 550486 267265
rect 372554 267225 372560 267237
rect 550480 267225 550486 267237
rect 550538 267225 550544 267277
rect 384880 267151 384886 267203
rect 384938 267191 384944 267203
rect 581200 267191 581206 267203
rect 384938 267163 581206 267191
rect 384938 267151 384944 267163
rect 581200 267151 581206 267163
rect 581258 267151 581264 267203
rect 386032 267077 386038 267129
rect 386090 267117 386096 267129
rect 584752 267117 584758 267129
rect 386090 267089 584758 267117
rect 386090 267077 386096 267089
rect 584752 267077 584758 267089
rect 584810 267077 584816 267129
rect 387760 267003 387766 267055
rect 387818 267043 387824 267055
rect 588304 267043 588310 267055
rect 387818 267015 588310 267043
rect 387818 267003 387824 267015
rect 588304 267003 588310 267015
rect 588362 267003 588368 267055
rect 301840 266929 301846 266981
rect 301898 266969 301904 266981
rect 375280 266969 375286 266981
rect 301898 266941 375286 266969
rect 301898 266929 301904 266941
rect 375280 266929 375286 266941
rect 375338 266929 375344 266981
rect 394672 266929 394678 266981
rect 394730 266969 394736 266981
rect 606064 266969 606070 266981
rect 394730 266941 606070 266969
rect 394730 266929 394736 266941
rect 606064 266929 606070 266941
rect 606122 266929 606128 266981
rect 305008 266855 305014 266907
rect 305066 266895 305072 266907
rect 383824 266895 383830 266907
rect 305066 266867 383830 266895
rect 305066 266855 305072 266867
rect 383824 266855 383830 266867
rect 383882 266855 383888 266907
rect 393232 266855 393238 266907
rect 393290 266895 393296 266907
rect 602512 266895 602518 266907
rect 393290 266867 602518 266895
rect 393290 266855 393296 266867
rect 602512 266855 602518 266867
rect 602570 266855 602576 266907
rect 306160 266781 306166 266833
rect 306218 266821 306224 266833
rect 386128 266821 386134 266833
rect 306218 266793 386134 266821
rect 306218 266781 306224 266793
rect 386128 266781 386134 266793
rect 386186 266781 386192 266833
rect 397552 266781 397558 266833
rect 397610 266821 397616 266833
rect 613072 266821 613078 266833
rect 397610 266793 613078 266821
rect 397610 266781 397616 266793
rect 613072 266781 613078 266793
rect 613130 266781 613136 266833
rect 308752 266707 308758 266759
rect 308810 266747 308816 266759
rect 392944 266747 392950 266759
rect 308810 266719 392950 266747
rect 308810 266707 308816 266719
rect 392944 266707 392950 266719
rect 393002 266707 393008 266759
rect 398224 266707 398230 266759
rect 398282 266747 398288 266759
rect 614320 266747 614326 266759
rect 398282 266719 614326 266747
rect 398282 266707 398288 266719
rect 614320 266707 614326 266719
rect 614378 266707 614384 266759
rect 308080 266633 308086 266685
rect 308138 266673 308144 266685
rect 390928 266673 390934 266685
rect 308138 266645 390934 266673
rect 308138 266633 308144 266645
rect 390928 266633 390934 266645
rect 390986 266633 390992 266685
rect 400624 266633 400630 266685
rect 400682 266673 400688 266685
rect 620176 266673 620182 266685
rect 400682 266645 620182 266673
rect 400682 266633 400688 266645
rect 620176 266633 620182 266645
rect 620234 266633 620240 266685
rect 310672 266559 310678 266611
rect 310730 266599 310736 266611
rect 398032 266599 398038 266611
rect 310730 266571 398038 266599
rect 310730 266559 310736 266571
rect 398032 266559 398038 266571
rect 398090 266559 398096 266611
rect 403216 266559 403222 266611
rect 403274 266599 403280 266611
rect 627280 266599 627286 266611
rect 403274 266571 627286 266599
rect 403274 266559 403280 266571
rect 627280 266559 627286 266571
rect 627338 266559 627344 266611
rect 313552 266485 313558 266537
rect 313610 266525 313616 266537
rect 405040 266525 405046 266537
rect 313610 266497 405046 266525
rect 313610 266485 313616 266497
rect 405040 266485 405046 266497
rect 405098 266485 405104 266537
rect 406096 266485 406102 266537
rect 406154 266525 406160 266537
rect 634384 266525 634390 266537
rect 406154 266497 634390 266525
rect 406154 266485 406160 266497
rect 634384 266485 634390 266497
rect 634442 266485 634448 266537
rect 187216 266411 187222 266463
rect 187274 266451 187280 266463
rect 189712 266451 189718 266463
rect 187274 266423 189718 266451
rect 187274 266411 187280 266423
rect 189712 266411 189718 266423
rect 189770 266411 189776 266463
rect 313072 266411 313078 266463
rect 313130 266451 313136 266463
rect 403888 266451 403894 266463
rect 313130 266423 403894 266451
rect 313130 266411 313136 266423
rect 403888 266411 403894 266423
rect 403946 266411 403952 266463
rect 409168 266411 409174 266463
rect 409226 266451 409232 266463
rect 641488 266451 641494 266463
rect 409226 266423 641494 266451
rect 409226 266411 409232 266423
rect 641488 266411 641494 266423
rect 641546 266411 641552 266463
rect 44944 266337 44950 266389
rect 45002 266377 45008 266389
rect 671632 266377 671638 266389
rect 45002 266349 671638 266377
rect 45002 266337 45008 266349
rect 671632 266337 671638 266349
rect 671690 266337 671696 266389
rect 348880 266263 348886 266315
rect 348938 266303 348944 266315
rect 492592 266303 492598 266315
rect 348938 266275 492598 266303
rect 348938 266263 348944 266275
rect 492592 266263 492598 266275
rect 492650 266263 492656 266315
rect 346000 266189 346006 266241
rect 346058 266229 346064 266241
rect 485488 266229 485494 266241
rect 346058 266201 485494 266229
rect 346058 266189 346064 266201
rect 485488 266189 485494 266201
rect 485546 266189 485552 266241
rect 343312 266115 343318 266167
rect 343370 266155 343376 266167
rect 478384 266155 478390 266167
rect 343370 266127 478390 266155
rect 343370 266115 343376 266127
rect 478384 266115 478390 266127
rect 478442 266115 478448 266167
rect 340240 266041 340246 266093
rect 340298 266081 340304 266093
rect 471280 266081 471286 266093
rect 340298 266053 471286 266081
rect 340298 266041 340304 266053
rect 471280 266041 471286 266053
rect 471338 266041 471344 266093
rect 337360 265967 337366 266019
rect 337418 266007 337424 266019
rect 464176 266007 464182 266019
rect 337418 265979 464182 266007
rect 337418 265967 337424 265979
rect 464176 265967 464182 265979
rect 464234 265967 464240 266019
rect 334768 265893 334774 265945
rect 334826 265933 334832 265945
rect 457072 265933 457078 265945
rect 334826 265905 457078 265933
rect 334826 265893 334832 265905
rect 457072 265893 457078 265905
rect 457130 265893 457136 265945
rect 331888 265819 331894 265871
rect 331946 265859 331952 265871
rect 449968 265859 449974 265871
rect 331946 265831 449974 265859
rect 331946 265819 331952 265831
rect 449968 265819 449974 265831
rect 450026 265819 450032 265871
rect 327568 265745 327574 265797
rect 327626 265785 327632 265797
rect 439312 265785 439318 265797
rect 327626 265757 439318 265785
rect 327626 265745 327632 265757
rect 439312 265745 439318 265757
rect 439370 265745 439376 265797
rect 324496 265671 324502 265723
rect 324554 265711 324560 265723
rect 432304 265711 432310 265723
rect 324554 265683 432310 265711
rect 324554 265671 324560 265683
rect 432304 265671 432310 265683
rect 432362 265671 432368 265723
rect 321616 265597 321622 265649
rect 321674 265637 321680 265649
rect 425200 265637 425206 265649
rect 321674 265609 425206 265637
rect 321674 265597 321680 265609
rect 425200 265597 425206 265609
rect 425258 265597 425264 265649
rect 408016 265523 408022 265575
rect 408074 265563 408080 265575
rect 508240 265563 508246 265575
rect 408074 265535 508246 265563
rect 408074 265523 408080 265535
rect 508240 265523 508246 265535
rect 508298 265523 508304 265575
rect 319024 265449 319030 265501
rect 319082 265489 319088 265501
rect 418096 265489 418102 265501
rect 319082 265461 418102 265489
rect 319082 265449 319088 265461
rect 418096 265449 418102 265461
rect 418154 265449 418160 265501
rect 656560 265375 656566 265427
rect 656618 265415 656624 265427
rect 676048 265415 676054 265427
rect 656618 265387 676054 265415
rect 656618 265375 656624 265387
rect 676048 265375 676054 265387
rect 676106 265375 676112 265427
rect 656272 265227 656278 265279
rect 656330 265267 656336 265279
rect 676240 265267 676246 265279
rect 656330 265239 676246 265267
rect 656330 265227 656336 265239
rect 676240 265227 676246 265239
rect 676298 265227 676304 265279
rect 673264 265153 673270 265205
rect 673322 265193 673328 265205
rect 676048 265193 676054 265205
rect 673322 265165 676054 265193
rect 673322 265153 673328 265165
rect 676048 265153 676054 265165
rect 676106 265153 676112 265205
rect 656080 265079 656086 265131
rect 656138 265119 656144 265131
rect 676144 265119 676150 265131
rect 656138 265091 676150 265119
rect 656138 265079 656144 265091
rect 676144 265079 676150 265091
rect 676202 265079 676208 265131
rect 23056 265005 23062 265057
rect 23114 265045 23120 265057
rect 43504 265045 43510 265057
rect 23114 265017 43510 265045
rect 23114 265005 23120 265017
rect 43504 265005 43510 265017
rect 43562 265005 43568 265057
rect 671632 265005 671638 265057
rect 671690 265045 671696 265057
rect 673360 265045 673366 265057
rect 671690 265017 673366 265045
rect 671690 265005 671696 265017
rect 673360 265005 673366 265017
rect 673418 265045 673424 265057
rect 676048 265045 676054 265057
rect 673418 265017 676054 265045
rect 673418 265005 673424 265017
rect 676048 265005 676054 265017
rect 676106 265005 676112 265057
rect 43216 264931 43222 264983
rect 43274 264971 43280 264983
rect 44080 264971 44086 264983
rect 43274 264943 44086 264971
rect 43274 264931 43280 264943
rect 44080 264931 44086 264943
rect 44138 264971 44144 264983
rect 669808 264971 669814 264983
rect 44138 264943 669814 264971
rect 44138 264931 44144 264943
rect 669808 264931 669814 264943
rect 669866 264931 669872 264983
rect 43312 264857 43318 264909
rect 43370 264897 43376 264909
rect 44176 264897 44182 264909
rect 43370 264869 44182 264897
rect 43370 264857 43376 264869
rect 44176 264857 44182 264869
rect 44234 264897 44240 264909
rect 669616 264897 669622 264909
rect 44234 264869 669622 264897
rect 44234 264857 44240 264869
rect 669616 264857 669622 264869
rect 669674 264857 669680 264909
rect 359440 264783 359446 264835
rect 359498 264823 359504 264835
rect 475984 264823 475990 264835
rect 359498 264795 475990 264823
rect 359498 264783 359504 264795
rect 475984 264783 475990 264795
rect 476042 264783 476048 264835
rect 328048 264709 328054 264761
rect 328106 264749 328112 264761
rect 440560 264749 440566 264761
rect 328106 264721 440566 264749
rect 328106 264709 328112 264721
rect 440560 264709 440566 264721
rect 440618 264709 440624 264761
rect 331120 264635 331126 264687
rect 331178 264675 331184 264687
rect 447664 264675 447670 264687
rect 331178 264647 447670 264675
rect 331178 264635 331184 264647
rect 447664 264635 447670 264647
rect 447722 264635 447728 264687
rect 354256 264561 354262 264613
rect 354314 264601 354320 264613
rect 461776 264601 461782 264613
rect 354314 264573 461782 264601
rect 354314 264561 354320 264573
rect 461776 264561 461782 264573
rect 461834 264561 461840 264613
rect 360400 264487 360406 264539
rect 360458 264527 360464 264539
rect 468880 264527 468886 264539
rect 360458 264499 468886 264527
rect 360458 264487 360464 264499
rect 468880 264487 468886 264499
rect 468938 264487 468944 264539
rect 351376 264413 351382 264465
rect 351434 264453 351440 264465
rect 454768 264453 454774 264465
rect 351434 264425 454774 264453
rect 351434 264413 351440 264425
rect 454768 264413 454774 264425
rect 454826 264413 454832 264465
rect 399376 264117 399382 264169
rect 399434 264157 399440 264169
rect 410992 264157 410998 264169
rect 399434 264129 410998 264157
rect 399434 264117 399440 264129
rect 410992 264117 410998 264129
rect 411050 264117 411056 264169
rect 324976 264043 324982 264095
rect 325034 264083 325040 264095
rect 433456 264083 433462 264095
rect 325034 264055 433462 264083
rect 325034 264043 325040 264055
rect 433456 264043 433462 264055
rect 433514 264043 433520 264095
rect 387952 263969 387958 264021
rect 388010 264009 388016 264021
rect 589456 264009 589462 264021
rect 388010 263981 589462 264009
rect 388010 263969 388016 263981
rect 589456 263969 589462 263981
rect 589514 263969 589520 264021
rect 390832 263895 390838 263947
rect 390890 263935 390896 263947
rect 596560 263935 596566 263947
rect 390890 263907 596566 263935
rect 390890 263895 390896 263907
rect 596560 263895 596566 263907
rect 596618 263895 596624 263947
rect 393904 263821 393910 263873
rect 393962 263861 393968 263873
rect 603664 263861 603670 263873
rect 393962 263833 603670 263861
rect 393962 263821 393968 263833
rect 603664 263821 603670 263833
rect 603722 263821 603728 263873
rect 396784 263747 396790 263799
rect 396842 263787 396848 263799
rect 610768 263787 610774 263799
rect 396842 263759 610774 263787
rect 396842 263747 396848 263759
rect 610768 263747 610774 263759
rect 610826 263747 610832 263799
rect 401104 263673 401110 263725
rect 401162 263713 401168 263725
rect 401162 263685 410750 263713
rect 401162 263673 401168 263685
rect 23344 263599 23350 263651
rect 23402 263639 23408 263651
rect 44176 263639 44182 263651
rect 23402 263611 44182 263639
rect 23402 263599 23408 263611
rect 44176 263599 44182 263611
rect 44234 263599 44240 263651
rect 403984 263599 403990 263651
rect 404042 263639 404048 263651
rect 410722 263639 410750 263685
rect 410992 263673 410998 263725
rect 411050 263713 411056 263725
rect 617872 263713 617878 263725
rect 411050 263685 617878 263713
rect 411050 263673 411056 263685
rect 617872 263673 617878 263685
rect 617930 263673 617936 263725
rect 621424 263639 621430 263651
rect 404042 263611 410654 263639
rect 410722 263611 621430 263639
rect 404042 263599 404048 263611
rect 23248 263525 23254 263577
rect 23306 263565 23312 263577
rect 44080 263565 44086 263577
rect 23306 263537 44086 263565
rect 23306 263525 23312 263537
rect 44080 263525 44086 263537
rect 44138 263525 44144 263577
rect 409648 263525 409654 263577
rect 409706 263525 409712 263577
rect 410626 263565 410654 263611
rect 621424 263599 621430 263611
rect 621482 263599 621488 263651
rect 628432 263565 628438 263577
rect 410626 263537 628438 263565
rect 628432 263525 628438 263537
rect 628490 263525 628496 263577
rect 409666 263491 409694 263525
rect 642640 263491 642646 263503
rect 409666 263463 642646 263491
rect 642640 263451 642646 263463
rect 642698 263451 642704 263503
rect 23152 262119 23158 262171
rect 23210 262159 23216 262171
rect 43312 262159 43318 262171
rect 23210 262131 43318 262159
rect 23210 262119 23216 262131
rect 43312 262119 43318 262131
rect 43370 262119 43376 262171
rect 420400 262119 420406 262171
rect 420458 262159 420464 262171
rect 606160 262159 606166 262171
rect 420458 262131 606166 262159
rect 420458 262119 420464 262131
rect 606160 262119 606166 262131
rect 606218 262119 606224 262171
rect 674704 259307 674710 259359
rect 674762 259347 674768 259359
rect 675952 259347 675958 259359
rect 674762 259319 675958 259347
rect 674762 259307 674768 259319
rect 675952 259307 675958 259319
rect 676010 259307 676016 259359
rect 420400 259233 420406 259285
rect 420458 259273 420464 259285
rect 606256 259273 606262 259285
rect 420458 259245 606262 259273
rect 420458 259233 420464 259245
rect 606256 259233 606262 259245
rect 606314 259233 606320 259285
rect 675184 259233 675190 259285
rect 675242 259273 675248 259285
rect 676048 259273 676054 259285
rect 675242 259245 676054 259273
rect 675242 259233 675248 259245
rect 676048 259233 676054 259245
rect 676106 259233 676112 259285
rect 674608 256939 674614 256991
rect 674666 256979 674672 256991
rect 676048 256979 676054 256991
rect 674666 256951 676054 256979
rect 674666 256939 674672 256951
rect 676048 256939 676054 256951
rect 676106 256939 676112 256991
rect 674800 256421 674806 256473
rect 674858 256461 674864 256473
rect 676048 256461 676054 256473
rect 674858 256433 676054 256461
rect 674858 256421 674864 256433
rect 676048 256421 676054 256433
rect 676106 256421 676112 256473
rect 40240 256347 40246 256399
rect 40298 256387 40304 256399
rect 59056 256387 59062 256399
rect 40298 256359 59062 256387
rect 40298 256347 40304 256359
rect 59056 256347 59062 256359
rect 59114 256347 59120 256399
rect 420400 256347 420406 256399
rect 420458 256387 420464 256399
rect 606352 256387 606358 256399
rect 420458 256359 606358 256387
rect 420458 256347 420464 256359
rect 606352 256347 606358 256359
rect 606410 256347 606416 256399
rect 674896 256347 674902 256399
rect 674954 256387 674960 256399
rect 676240 256387 676246 256399
rect 674954 256359 676246 256387
rect 674954 256347 674960 256359
rect 676240 256347 676246 256359
rect 676298 256347 676304 256399
rect 41776 255385 41782 255437
rect 41834 255425 41840 255437
rect 53200 255425 53206 255437
rect 41834 255397 53206 255425
rect 41834 255385 41840 255397
rect 53200 255385 53206 255397
rect 53258 255385 53264 255437
rect 47824 255089 47830 255141
rect 47882 255129 47888 255141
rect 186064 255129 186070 255141
rect 47882 255101 186070 255129
rect 47882 255089 47888 255101
rect 186064 255089 186070 255101
rect 186122 255089 186128 255141
rect 47440 255015 47446 255067
rect 47498 255055 47504 255067
rect 185968 255055 185974 255067
rect 47498 255027 185974 255055
rect 47498 255015 47504 255027
rect 185968 255015 185974 255027
rect 186026 255015 186032 255067
rect 41776 254941 41782 254993
rect 41834 254981 41840 254993
rect 43408 254981 43414 254993
rect 41834 254953 43414 254981
rect 41834 254941 41840 254953
rect 43408 254941 43414 254953
rect 43466 254941 43472 254993
rect 47920 254941 47926 254993
rect 47978 254981 47984 254993
rect 186544 254981 186550 254993
rect 47978 254953 186550 254981
rect 47978 254941 47984 254953
rect 186544 254941 186550 254953
rect 186602 254941 186608 254993
rect 48016 254867 48022 254919
rect 48074 254907 48080 254919
rect 186736 254907 186742 254919
rect 48074 254879 186742 254907
rect 48074 254867 48080 254879
rect 186736 254867 186742 254879
rect 186794 254867 186800 254919
rect 41776 254423 41782 254475
rect 41834 254463 41840 254475
rect 43408 254463 43414 254475
rect 41834 254435 43414 254463
rect 41834 254423 41840 254435
rect 43408 254423 43414 254435
rect 43466 254423 43472 254475
rect 674992 253535 674998 253587
rect 675050 253575 675056 253587
rect 676048 253575 676054 253587
rect 675050 253547 676054 253575
rect 675050 253535 675056 253547
rect 676048 253535 676054 253547
rect 676106 253535 676112 253587
rect 41584 253461 41590 253513
rect 41642 253501 41648 253513
rect 56176 253501 56182 253513
rect 41642 253473 56182 253501
rect 41642 253461 41648 253473
rect 56176 253461 56182 253473
rect 56234 253461 56240 253513
rect 420400 253461 420406 253513
rect 420458 253501 420464 253513
rect 603280 253501 603286 253513
rect 420458 253473 603286 253501
rect 420458 253461 420464 253473
rect 603280 253461 603286 253473
rect 603338 253461 603344 253513
rect 646672 253461 646678 253513
rect 646730 253501 646736 253513
rect 679696 253501 679702 253513
rect 646730 253473 679702 253501
rect 646730 253461 646736 253473
rect 679696 253461 679702 253473
rect 679754 253461 679760 253513
rect 106480 252277 106486 252329
rect 106538 252317 106544 252329
rect 156880 252317 156886 252329
rect 106538 252289 156886 252317
rect 106538 252277 106544 252289
rect 156880 252277 156886 252289
rect 156938 252277 156944 252329
rect 92080 252203 92086 252255
rect 92138 252243 92144 252255
rect 145456 252243 145462 252255
rect 92138 252215 145462 252243
rect 92138 252203 92144 252215
rect 145456 252203 145462 252215
rect 145514 252203 145520 252255
rect 109360 252129 109366 252181
rect 109418 252169 109424 252181
rect 171280 252169 171286 252181
rect 109418 252141 171286 252169
rect 109418 252129 109424 252141
rect 171280 252129 171286 252141
rect 171338 252129 171344 252181
rect 97840 252055 97846 252107
rect 97898 252095 97904 252107
rect 182800 252095 182806 252107
rect 97898 252067 182806 252095
rect 97898 252055 97904 252067
rect 182800 252055 182806 252067
rect 182858 252055 182864 252107
rect 56080 251981 56086 252033
rect 56138 252021 56144 252033
rect 186352 252021 186358 252033
rect 56138 251993 186358 252021
rect 56138 251981 56144 251993
rect 186352 251981 186358 251993
rect 186410 251981 186416 252033
rect 666640 250649 666646 250701
rect 666698 250689 666704 250701
rect 675376 250689 675382 250701
rect 666698 250661 675382 250689
rect 666698 250649 666704 250661
rect 675376 250649 675382 250661
rect 675434 250649 675440 250701
rect 420400 250575 420406 250627
rect 420458 250615 420464 250627
rect 603376 250615 603382 250627
rect 420458 250587 603382 250615
rect 420458 250575 420464 250587
rect 603376 250575 603382 250587
rect 603434 250575 603440 250627
rect 120880 249909 120886 249961
rect 120938 249949 120944 249961
rect 145648 249949 145654 249961
rect 120938 249921 145654 249949
rect 120938 249909 120944 249921
rect 145648 249909 145654 249921
rect 145706 249909 145712 249961
rect 132400 249835 132406 249887
rect 132458 249875 132464 249887
rect 159856 249875 159862 249887
rect 132458 249847 159862 249875
rect 132458 249835 132464 249847
rect 159856 249835 159862 249847
rect 159914 249835 159920 249887
rect 135280 249761 135286 249813
rect 135338 249801 135344 249813
rect 168496 249801 168502 249813
rect 135338 249773 168502 249801
rect 135338 249761 135344 249773
rect 168496 249761 168502 249773
rect 168554 249761 168560 249813
rect 138160 249687 138166 249739
rect 138218 249727 138224 249739
rect 171472 249727 171478 249739
rect 138218 249699 171478 249727
rect 138218 249687 138224 249699
rect 171472 249687 171478 249699
rect 171530 249687 171536 249739
rect 141040 249613 141046 249665
rect 141098 249653 141104 249665
rect 180016 249653 180022 249665
rect 141098 249625 180022 249653
rect 141098 249613 141104 249625
rect 180016 249613 180022 249625
rect 180074 249613 180080 249665
rect 123760 249539 123766 249591
rect 123818 249579 123824 249591
rect 165712 249579 165718 249591
rect 123818 249551 165718 249579
rect 123818 249539 123824 249551
rect 165712 249539 165718 249551
rect 165770 249539 165776 249591
rect 126640 249465 126646 249517
rect 126698 249505 126704 249517
rect 177040 249505 177046 249517
rect 126698 249477 177046 249505
rect 126698 249465 126704 249477
rect 177040 249465 177046 249477
rect 177098 249465 177104 249517
rect 94960 249391 94966 249443
rect 95018 249431 95024 249443
rect 154000 249431 154006 249443
rect 95018 249403 154006 249431
rect 95018 249391 95024 249403
rect 154000 249391 154006 249403
rect 154058 249391 154064 249443
rect 118000 249317 118006 249369
rect 118058 249357 118064 249369
rect 182896 249357 182902 249369
rect 118058 249329 182902 249357
rect 118058 249317 118064 249329
rect 182896 249317 182902 249329
rect 182954 249317 182960 249369
rect 77680 249243 77686 249295
rect 77738 249283 77744 249295
rect 145360 249283 145366 249295
rect 77738 249255 145366 249283
rect 77738 249243 77744 249255
rect 145360 249243 145366 249255
rect 145418 249243 145424 249295
rect 80560 249169 80566 249221
rect 80618 249209 80624 249221
rect 162640 249209 162646 249221
rect 80618 249181 162646 249209
rect 80618 249169 80624 249181
rect 162640 249169 162646 249181
rect 162698 249169 162704 249221
rect 86320 249095 86326 249147
rect 86378 249135 86384 249147
rect 174160 249135 174166 249147
rect 86378 249107 174166 249135
rect 86378 249095 86384 249107
rect 174160 249095 174166 249107
rect 174218 249095 174224 249147
rect 675184 247911 675190 247963
rect 675242 247951 675248 247963
rect 675376 247951 675382 247963
rect 675242 247923 675382 247951
rect 675242 247911 675248 247923
rect 675376 247911 675382 247923
rect 675434 247911 675440 247963
rect 420304 247763 420310 247815
rect 420362 247803 420368 247815
rect 603472 247803 603478 247815
rect 420362 247775 603478 247803
rect 420362 247763 420368 247775
rect 603472 247763 603478 247775
rect 603530 247763 603536 247815
rect 420400 247689 420406 247741
rect 420458 247729 420464 247741
rect 629200 247729 629206 247741
rect 420458 247701 629206 247729
rect 420458 247689 420464 247701
rect 629200 247689 629206 247701
rect 629258 247689 629264 247741
rect 655888 247615 655894 247667
rect 655946 247655 655952 247667
rect 666640 247655 666646 247667
rect 655946 247627 666646 247655
rect 655946 247615 655952 247627
rect 666640 247615 666646 247627
rect 666698 247615 666704 247667
rect 674704 247245 674710 247297
rect 674762 247285 674768 247297
rect 675472 247285 675478 247297
rect 674762 247257 675478 247285
rect 674762 247245 674768 247257
rect 675472 247245 675478 247257
rect 675530 247245 675536 247297
rect 103600 246727 103606 246779
rect 103658 246767 103664 246779
rect 165520 246767 165526 246779
rect 103658 246739 165526 246767
rect 103658 246727 103664 246739
rect 165520 246727 165526 246739
rect 165578 246727 165584 246779
rect 112240 246653 112246 246705
rect 112298 246693 112304 246705
rect 185776 246693 185782 246705
rect 112298 246665 185782 246693
rect 112298 246653 112304 246665
rect 185776 246653 185782 246665
rect 185834 246653 185840 246705
rect 47632 246579 47638 246631
rect 47690 246619 47696 246631
rect 186256 246619 186262 246631
rect 47690 246591 186262 246619
rect 47690 246579 47696 246591
rect 186256 246579 186262 246591
rect 186314 246579 186320 246631
rect 674608 246579 674614 246631
rect 674666 246619 674672 246631
rect 675376 246619 675382 246631
rect 674666 246591 675382 246619
rect 674666 246579 674672 246591
rect 675376 246579 675382 246591
rect 675434 246579 675440 246631
rect 47536 246505 47542 246557
rect 47594 246545 47600 246557
rect 186448 246545 186454 246557
rect 47594 246517 186454 246545
rect 47594 246505 47600 246517
rect 186448 246505 186454 246517
rect 186506 246505 186512 246557
rect 47728 246431 47734 246483
rect 47786 246471 47792 246483
rect 186640 246471 186646 246483
rect 47786 246443 186646 246471
rect 47786 246431 47792 246443
rect 186640 246431 186646 246443
rect 186698 246431 186704 246483
rect 45808 246357 45814 246409
rect 45866 246397 45872 246409
rect 187024 246397 187030 246409
rect 45866 246369 187030 246397
rect 45866 246357 45872 246369
rect 187024 246357 187030 246369
rect 187082 246357 187088 246409
rect 45424 246283 45430 246335
rect 45482 246323 45488 246335
rect 186832 246323 186838 246335
rect 45482 246295 186838 246323
rect 45482 246283 45488 246295
rect 186832 246283 186838 246295
rect 186890 246283 186896 246335
rect 44560 246209 44566 246261
rect 44618 246249 44624 246261
rect 186160 246249 186166 246261
rect 44618 246221 186166 246249
rect 44618 246209 44624 246221
rect 186160 246209 186166 246221
rect 186218 246209 186224 246261
rect 674896 246061 674902 246113
rect 674954 246101 674960 246113
rect 675376 246101 675382 246113
rect 674954 246073 675382 246101
rect 674954 246061 674960 246073
rect 675376 246061 675382 246073
rect 675434 246061 675440 246113
rect 41584 244951 41590 245003
rect 41642 244991 41648 245003
rect 145552 244991 145558 245003
rect 41642 244963 145558 244991
rect 41642 244951 41648 244963
rect 145552 244951 145558 244963
rect 145610 244951 145616 245003
rect 44752 244877 44758 244929
rect 44810 244917 44816 244929
rect 186928 244917 186934 244929
rect 44810 244889 186934 244917
rect 44810 244877 44816 244889
rect 186928 244877 186934 244889
rect 186986 244877 186992 244929
rect 41776 244803 41782 244855
rect 41834 244843 41840 244855
rect 145744 244843 145750 244855
rect 41834 244815 145750 244843
rect 41834 244803 41840 244815
rect 145744 244803 145750 244815
rect 145802 244803 145808 244855
rect 420400 244803 420406 244855
rect 420458 244843 420464 244855
rect 629296 244843 629302 244855
rect 420458 244815 629302 244843
rect 420458 244803 420464 244815
rect 629296 244803 629302 244815
rect 629354 244803 629360 244855
rect 41488 244655 41494 244707
rect 41546 244695 41552 244707
rect 42928 244695 42934 244707
rect 41546 244667 42934 244695
rect 41546 244655 41552 244667
rect 42928 244655 42934 244667
rect 42986 244655 42992 244707
rect 41392 244581 41398 244633
rect 41450 244621 41456 244633
rect 42832 244621 42838 244633
rect 41450 244593 42838 244621
rect 41450 244581 41456 244593
rect 42832 244581 42838 244593
rect 42890 244581 42896 244633
rect 41296 244507 41302 244559
rect 41354 244547 41360 244559
rect 43024 244547 43030 244559
rect 41354 244519 43030 244547
rect 41354 244507 41360 244519
rect 43024 244507 43030 244519
rect 43082 244507 43088 244559
rect 44848 242805 44854 242857
rect 44906 242845 44912 242857
rect 185680 242845 185686 242857
rect 44906 242817 185686 242845
rect 44906 242805 44912 242817
rect 185680 242805 185686 242817
rect 185738 242805 185744 242857
rect 44656 242731 44662 242783
rect 44714 242771 44720 242783
rect 185584 242771 185590 242783
rect 44714 242743 185590 242771
rect 44714 242731 44720 242743
rect 185584 242731 185590 242743
rect 185642 242731 185648 242783
rect 674800 242731 674806 242783
rect 674858 242771 674864 242783
rect 675376 242771 675382 242783
rect 674858 242743 675382 242771
rect 674858 242731 674864 242743
rect 675376 242731 675382 242743
rect 675434 242731 675440 242783
rect 44560 242657 44566 242709
rect 44618 242697 44624 242709
rect 185872 242697 185878 242709
rect 44618 242669 185878 242697
rect 44618 242657 44624 242669
rect 185872 242657 185878 242669
rect 185930 242657 185936 242709
rect 41584 242583 41590 242635
rect 41642 242623 41648 242635
rect 142576 242623 142582 242635
rect 41642 242595 142582 242623
rect 41642 242583 41648 242595
rect 142576 242583 142582 242595
rect 142634 242583 142640 242635
rect 41680 241991 41686 242043
rect 41738 242031 41744 242043
rect 42736 242031 42742 242043
rect 41738 242003 42742 242031
rect 41738 241991 41744 242003
rect 42736 241991 42742 242003
rect 42794 241991 42800 242043
rect 420304 241917 420310 241969
rect 420362 241957 420368 241969
rect 600400 241957 600406 241969
rect 420362 241929 600406 241957
rect 420362 241917 420368 241929
rect 600400 241917 600406 241929
rect 600458 241917 600464 241969
rect 674992 241547 674998 241599
rect 675050 241587 675056 241599
rect 675472 241587 675478 241599
rect 675050 241559 675478 241587
rect 675050 241547 675056 241559
rect 675472 241547 675478 241559
rect 675530 241547 675536 241599
rect 41872 240585 41878 240637
rect 41930 240585 41936 240637
rect 41890 240415 41918 240585
rect 41872 240363 41878 240415
rect 41930 240363 41936 240415
rect 380848 239919 380854 239971
rect 380906 239959 380912 239971
rect 412048 239959 412054 239971
rect 380906 239931 412054 239959
rect 380906 239919 380912 239931
rect 412048 239919 412054 239931
rect 412106 239919 412112 239971
rect 409552 239845 409558 239897
rect 409610 239885 409616 239897
rect 412144 239885 412150 239897
rect 409610 239857 412150 239885
rect 409610 239845 409616 239857
rect 412144 239845 412150 239857
rect 412202 239845 412208 239897
rect 360016 239771 360022 239823
rect 360074 239811 360080 239823
rect 434608 239811 434614 239823
rect 360074 239783 434614 239811
rect 360074 239771 360080 239783
rect 434608 239771 434614 239783
rect 434666 239771 434672 239823
rect 371440 239697 371446 239749
rect 371498 239737 371504 239749
rect 446704 239737 446710 239749
rect 371498 239709 446710 239737
rect 371498 239697 371504 239709
rect 446704 239697 446710 239709
rect 446762 239697 446768 239749
rect 378832 239623 378838 239675
rect 378890 239663 378896 239675
rect 458800 239663 458806 239675
rect 378890 239635 458806 239663
rect 378890 239623 378896 239635
rect 458800 239623 458806 239635
rect 458858 239623 458864 239675
rect 383056 239549 383062 239601
rect 383114 239589 383120 239601
rect 470896 239589 470902 239601
rect 383114 239561 470902 239589
rect 383114 239549 383120 239561
rect 470896 239549 470902 239561
rect 470954 239549 470960 239601
rect 394768 239475 394774 239527
rect 394826 239515 394832 239527
rect 532816 239515 532822 239527
rect 394826 239487 532822 239515
rect 394826 239475 394832 239487
rect 532816 239475 532822 239487
rect 532874 239475 532880 239527
rect 408946 239413 411518 239441
rect 406192 239327 406198 239379
rect 406250 239367 406256 239379
rect 408946 239367 408974 239413
rect 406250 239339 408974 239367
rect 411490 239367 411518 239413
rect 411568 239401 411574 239453
rect 411626 239441 411632 239453
rect 541456 239441 541462 239453
rect 411626 239413 541462 239441
rect 411626 239401 411632 239413
rect 541456 239401 541462 239413
rect 541514 239401 541520 239453
rect 550864 239367 550870 239379
rect 411490 239339 550870 239367
rect 406250 239327 406256 239339
rect 550864 239327 550870 239339
rect 550922 239327 550928 239379
rect 400432 239253 400438 239305
rect 400490 239293 400496 239305
rect 411376 239293 411382 239305
rect 400490 239265 411382 239293
rect 400490 239253 400496 239265
rect 411376 239253 411382 239265
rect 411434 239253 411440 239305
rect 411472 239253 411478 239305
rect 411530 239293 411536 239305
rect 412240 239293 412246 239305
rect 411530 239265 412246 239293
rect 411530 239253 411536 239265
rect 412240 239253 412246 239265
rect 412298 239253 412304 239305
rect 420304 239253 420310 239305
rect 420362 239293 420368 239305
rect 599056 239293 599062 239305
rect 420362 239265 599062 239293
rect 420362 239253 420368 239265
rect 599056 239253 599062 239265
rect 599114 239253 599120 239305
rect 341200 239179 341206 239231
rect 341258 239219 341264 239231
rect 488272 239219 488278 239231
rect 341258 239191 488278 239219
rect 341258 239179 341264 239191
rect 488272 239179 488278 239191
rect 488330 239179 488336 239231
rect 350416 239105 350422 239157
rect 350474 239145 350480 239157
rect 508624 239145 508630 239157
rect 350474 239117 508630 239145
rect 350474 239105 350480 239117
rect 508624 239105 508630 239117
rect 508682 239105 508688 239157
rect 368560 239031 368566 239083
rect 368618 239071 368624 239083
rect 544816 239071 544822 239083
rect 368618 239043 544822 239071
rect 368618 239031 368624 239043
rect 544816 239031 544822 239043
rect 544874 239031 544880 239083
rect 382768 238957 382774 239009
rect 382826 238997 382832 239009
rect 414640 238997 414646 239009
rect 382826 238969 414646 238997
rect 382826 238957 382832 238969
rect 414640 238957 414646 238969
rect 414698 238957 414704 239009
rect 324400 238883 324406 238935
rect 324458 238923 324464 238935
rect 455152 238923 455158 238935
rect 324458 238895 455158 238923
rect 324458 238883 324464 238895
rect 455152 238883 455158 238895
rect 455210 238883 455216 238935
rect 323920 238809 323926 238861
rect 323978 238849 323984 238861
rect 455056 238849 455062 238861
rect 323978 238821 455062 238849
rect 323978 238809 323984 238821
rect 455056 238809 455062 238821
rect 455114 238809 455120 238861
rect 326704 238735 326710 238787
rect 326762 238775 326768 238787
rect 462544 238775 462550 238787
rect 326762 238747 462550 238775
rect 326762 238735 326768 238747
rect 462544 238735 462550 238747
rect 462602 238735 462608 238787
rect 328912 238661 328918 238713
rect 328970 238701 328976 238713
rect 464752 238701 464758 238713
rect 328970 238673 464758 238701
rect 328970 238661 328976 238673
rect 464752 238661 464758 238673
rect 464810 238661 464816 238713
rect 329872 238587 329878 238639
rect 329930 238627 329936 238639
rect 468592 238627 468598 238639
rect 329930 238599 468598 238627
rect 329930 238587 329936 238599
rect 468592 238587 468598 238599
rect 468650 238587 468656 238639
rect 332656 238513 332662 238565
rect 332714 238553 332720 238565
rect 474640 238553 474646 238565
rect 332714 238525 474646 238553
rect 332714 238513 332720 238525
rect 474640 238513 474646 238525
rect 474698 238513 474704 238565
rect 335728 238439 335734 238491
rect 335786 238479 335792 238491
rect 478192 238479 478198 238491
rect 335786 238451 478198 238479
rect 335786 238439 335792 238451
rect 478192 238439 478198 238451
rect 478250 238439 478256 238491
rect 336688 238365 336694 238417
rect 336746 238405 336752 238417
rect 378640 238405 378646 238417
rect 336746 238377 378646 238405
rect 336746 238365 336752 238377
rect 378640 238365 378646 238377
rect 378698 238365 378704 238417
rect 397072 238365 397078 238417
rect 397130 238405 397136 238417
rect 397744 238405 397750 238417
rect 397130 238377 397750 238405
rect 397130 238365 397136 238377
rect 397744 238365 397750 238377
rect 397802 238365 397808 238417
rect 403408 238365 403414 238417
rect 403466 238405 403472 238417
rect 478384 238405 478390 238417
rect 403466 238377 478390 238405
rect 403466 238365 403472 238377
rect 478384 238365 478390 238377
rect 478442 238365 478448 238417
rect 338992 238291 338998 238343
rect 339050 238331 339056 238343
rect 486736 238331 486742 238343
rect 339050 238303 486742 238331
rect 339050 238291 339056 238303
rect 486736 238291 486742 238303
rect 486794 238291 486800 238343
rect 341776 238217 341782 238269
rect 341834 238257 341840 238269
rect 492784 238257 492790 238269
rect 341834 238229 492790 238257
rect 341834 238217 341840 238229
rect 492784 238217 492790 238229
rect 492842 238217 492848 238269
rect 345328 238143 345334 238195
rect 345386 238183 345392 238195
rect 500272 238183 500278 238195
rect 345386 238155 500278 238183
rect 345386 238143 345392 238155
rect 500272 238143 500278 238155
rect 500330 238143 500336 238195
rect 346672 238069 346678 238121
rect 346730 238109 346736 238121
rect 503344 238109 503350 238121
rect 346730 238081 503350 238109
rect 346730 238069 346736 238081
rect 503344 238069 503350 238081
rect 503402 238069 503408 238121
rect 349936 237995 349942 238047
rect 349994 238035 350000 238047
rect 509392 238035 509398 238047
rect 349994 238007 509398 238035
rect 349994 237995 350000 238007
rect 509392 237995 509398 238007
rect 509450 237995 509456 238047
rect 353488 237921 353494 237973
rect 353546 237961 353552 237973
rect 378544 237961 378550 237973
rect 353546 237933 378550 237961
rect 353546 237921 353552 237933
rect 378544 237921 378550 237933
rect 378602 237921 378608 237973
rect 378640 237921 378646 237973
rect 378698 237961 378704 237973
rect 403408 237961 403414 237973
rect 378698 237933 403414 237961
rect 378698 237921 378704 237933
rect 403408 237921 403414 237933
rect 403466 237921 403472 237973
rect 403504 237921 403510 237973
rect 403562 237961 403568 237973
rect 403696 237961 403702 237973
rect 403562 237933 403702 237961
rect 403562 237921 403568 237933
rect 403696 237921 403702 237933
rect 403754 237921 403760 237973
rect 407440 237921 407446 237973
rect 407498 237961 407504 237973
rect 512752 237961 512758 237973
rect 407498 237933 512758 237961
rect 407498 237921 407504 237933
rect 512752 237921 512758 237933
rect 512810 237921 512816 237973
rect 352720 237847 352726 237899
rect 352778 237887 352784 237899
rect 513904 237887 513910 237899
rect 352778 237859 513910 237887
rect 352778 237847 352784 237859
rect 513904 237847 513910 237859
rect 513962 237847 513968 237899
rect 355696 237773 355702 237825
rect 355754 237813 355760 237825
rect 521488 237813 521494 237825
rect 355754 237785 521494 237813
rect 355754 237773 355760 237785
rect 521488 237773 521494 237785
rect 521546 237773 521552 237825
rect 358576 237699 358582 237751
rect 358634 237739 358640 237751
rect 526000 237739 526006 237751
rect 358634 237711 526006 237739
rect 358634 237699 358640 237711
rect 526000 237699 526006 237711
rect 526058 237699 526064 237751
rect 275344 237625 275350 237677
rect 275402 237665 275408 237677
rect 359920 237665 359926 237677
rect 275402 237637 359926 237665
rect 275402 237625 275408 237637
rect 359920 237625 359926 237637
rect 359978 237625 359984 237677
rect 363088 237625 363094 237677
rect 363146 237665 363152 237677
rect 535120 237665 535126 237677
rect 363146 237637 535126 237665
rect 363146 237625 363152 237637
rect 535120 237625 535126 237637
rect 535178 237625 535184 237677
rect 277072 237551 277078 237603
rect 277130 237591 277136 237603
rect 363664 237591 363670 237603
rect 277130 237563 363670 237591
rect 277130 237551 277136 237563
rect 363664 237551 363670 237563
rect 363722 237551 363728 237603
rect 364432 237551 364438 237603
rect 364490 237591 364496 237603
rect 535792 237591 535798 237603
rect 364490 237563 535798 237591
rect 364490 237551 364496 237563
rect 535792 237551 535798 237563
rect 535850 237551 535856 237603
rect 317584 237477 317590 237529
rect 317642 237517 317648 237529
rect 444496 237517 444502 237529
rect 317642 237489 444502 237517
rect 317642 237477 317648 237489
rect 444496 237477 444502 237489
rect 444554 237477 444560 237529
rect 317104 237403 317110 237455
rect 317162 237443 317168 237455
rect 441424 237443 441430 237455
rect 317162 237415 441430 237443
rect 317162 237403 317168 237415
rect 441424 237403 441430 237415
rect 441482 237403 441488 237455
rect 314800 237329 314806 237381
rect 314858 237369 314864 237381
rect 438352 237369 438358 237381
rect 314858 237341 438358 237369
rect 314858 237329 314864 237341
rect 438352 237329 438358 237341
rect 438410 237329 438416 237381
rect 311536 237255 311542 237307
rect 311594 237295 311600 237307
rect 432400 237295 432406 237307
rect 311594 237267 432406 237295
rect 311594 237255 311600 237267
rect 432400 237255 432406 237267
rect 432458 237255 432464 237307
rect 308560 237181 308566 237233
rect 308618 237221 308624 237233
rect 426352 237221 426358 237233
rect 308618 237193 426358 237221
rect 308618 237181 308624 237193
rect 426352 237181 426358 237193
rect 426410 237181 426416 237233
rect 310768 237107 310774 237159
rect 310826 237147 310832 237159
rect 411184 237147 411190 237159
rect 310826 237119 411190 237147
rect 310826 237107 310832 237119
rect 411184 237107 411190 237119
rect 411242 237107 411248 237159
rect 420304 237147 420310 237159
rect 411298 237119 420310 237147
rect 305776 237033 305782 237085
rect 305834 237073 305840 237085
rect 411298 237073 411326 237119
rect 420304 237107 420310 237119
rect 420362 237107 420368 237159
rect 305834 237045 411326 237073
rect 305834 237033 305840 237045
rect 411376 237033 411382 237085
rect 411434 237073 411440 237085
rect 413968 237073 413974 237085
rect 411434 237045 413974 237073
rect 411434 237033 411440 237045
rect 413968 237033 413974 237045
rect 414026 237033 414032 237085
rect 300208 236959 300214 237011
rect 300266 236999 300272 237011
rect 406768 236999 406774 237011
rect 300266 236971 406774 236999
rect 300266 236959 300272 236971
rect 406768 236959 406774 236971
rect 406826 236959 406832 237011
rect 408784 236959 408790 237011
rect 408842 236999 408848 237011
rect 414256 236999 414262 237011
rect 408842 236971 414262 236999
rect 408842 236959 408848 236971
rect 414256 236959 414262 236971
rect 414314 236959 414320 237011
rect 279856 236885 279862 236937
rect 279914 236925 279920 236937
rect 368944 236925 368950 236937
rect 279914 236897 368950 236925
rect 279914 236885 279920 236897
rect 368944 236885 368950 236897
rect 369002 236885 369008 236937
rect 388432 236885 388438 236937
rect 388490 236925 388496 236937
rect 397744 236925 397750 236937
rect 388490 236897 397750 236925
rect 388490 236885 388496 236897
rect 397744 236885 397750 236897
rect 397802 236885 397808 236937
rect 405904 236885 405910 236937
rect 405962 236925 405968 236937
rect 414448 236925 414454 236937
rect 405962 236897 414454 236925
rect 405962 236885 405968 236897
rect 414448 236885 414454 236897
rect 414506 236885 414512 236937
rect 278416 236811 278422 236863
rect 278474 236851 278480 236863
rect 366736 236851 366742 236863
rect 278474 236823 366742 236851
rect 278474 236811 278480 236823
rect 366736 236811 366742 236823
rect 366794 236811 366800 236863
rect 378544 236811 378550 236863
rect 378602 236851 378608 236863
rect 407440 236851 407446 236863
rect 378602 236823 407446 236851
rect 378602 236811 378608 236823
rect 407440 236811 407446 236823
rect 407498 236811 407504 236863
rect 407554 236823 408974 236851
rect 320848 236737 320854 236789
rect 320906 236777 320912 236789
rect 407554 236777 407582 236823
rect 320906 236749 407582 236777
rect 408946 236777 408974 236823
rect 411184 236811 411190 236863
rect 411242 236851 411248 236863
rect 428656 236851 428662 236863
rect 411242 236823 428662 236851
rect 411242 236811 411248 236823
rect 428656 236811 428662 236823
rect 428714 236811 428720 236863
rect 450448 236777 450454 236789
rect 408946 236749 450454 236777
rect 320906 236737 320912 236749
rect 450448 236737 450454 236749
rect 450506 236737 450512 236789
rect 42160 236663 42166 236715
rect 42218 236703 42224 236715
rect 42736 236703 42742 236715
rect 42218 236675 42742 236703
rect 42218 236663 42224 236675
rect 42736 236663 42742 236675
rect 42794 236663 42800 236715
rect 377776 236663 377782 236715
rect 377834 236703 377840 236715
rect 388720 236703 388726 236715
rect 377834 236675 388726 236703
rect 377834 236663 377840 236675
rect 388720 236663 388726 236675
rect 388778 236663 388784 236715
rect 397456 236663 397462 236715
rect 397514 236703 397520 236715
rect 413680 236703 413686 236715
rect 397514 236675 413686 236703
rect 397514 236663 397520 236675
rect 413680 236663 413686 236675
rect 413738 236663 413744 236715
rect 400336 236589 400342 236641
rect 400394 236629 400400 236641
rect 400394 236601 429134 236629
rect 400394 236589 400400 236601
rect 42736 236515 42742 236567
rect 42794 236555 42800 236567
rect 43024 236555 43030 236567
rect 42794 236527 43030 236555
rect 42794 236515 42800 236527
rect 43024 236515 43030 236527
rect 43082 236515 43088 236567
rect 397552 236515 397558 236567
rect 397610 236555 397616 236567
rect 413392 236555 413398 236567
rect 397610 236527 413398 236555
rect 397610 236515 397616 236527
rect 413392 236515 413398 236527
rect 413450 236515 413456 236567
rect 429106 236555 429134 236601
rect 511600 236555 511606 236567
rect 429106 236527 511606 236555
rect 511600 236515 511606 236527
rect 511658 236515 511664 236567
rect 376528 236441 376534 236493
rect 376586 236481 376592 236493
rect 397360 236481 397366 236493
rect 376586 236453 397366 236481
rect 376586 236441 376592 236453
rect 397360 236441 397366 236453
rect 397418 236441 397424 236493
rect 412048 236441 412054 236493
rect 412106 236481 412112 236493
rect 430096 236481 430102 236493
rect 412106 236453 430102 236481
rect 412106 236441 412112 236453
rect 430096 236441 430102 236453
rect 430154 236441 430160 236493
rect 412720 236367 412726 236419
rect 412778 236407 412784 236419
rect 442192 236407 442198 236419
rect 412778 236379 442198 236407
rect 412778 236367 412784 236379
rect 442192 236367 442198 236379
rect 442250 236367 442256 236419
rect 391600 236293 391606 236345
rect 391658 236333 391664 236345
rect 492016 236333 492022 236345
rect 391658 236305 492022 236333
rect 391658 236293 391664 236305
rect 492016 236293 492022 236305
rect 492074 236293 492080 236345
rect 394576 236219 394582 236271
rect 394634 236259 394640 236271
rect 505648 236259 505654 236271
rect 394634 236231 505654 236259
rect 394634 236219 394640 236231
rect 505648 236219 505654 236231
rect 505706 236219 505712 236271
rect 222352 236071 222358 236123
rect 222410 236111 222416 236123
rect 243952 236111 243958 236123
rect 222410 236083 243958 236111
rect 222410 236071 222416 236083
rect 243952 236071 243958 236083
rect 244010 236071 244016 236123
rect 251056 236071 251062 236123
rect 251114 236111 251120 236123
rect 273712 236111 273718 236123
rect 251114 236083 273718 236111
rect 251114 236071 251120 236083
rect 273712 236071 273718 236083
rect 273770 236071 273776 236123
rect 277552 236071 277558 236123
rect 277610 236111 277616 236123
rect 313936 236111 313942 236123
rect 277610 236083 313942 236111
rect 277610 236071 277616 236083
rect 313936 236071 313942 236083
rect 313994 236071 314000 236123
rect 319888 236071 319894 236123
rect 319946 236111 319952 236123
rect 371440 236111 371446 236123
rect 319946 236083 371446 236111
rect 319946 236071 319952 236083
rect 371440 236071 371446 236083
rect 371498 236071 371504 236123
rect 371824 236071 371830 236123
rect 371882 236111 371888 236123
rect 406192 236111 406198 236123
rect 371882 236083 406198 236111
rect 371882 236071 371888 236083
rect 406192 236071 406198 236083
rect 406250 236071 406256 236123
rect 406288 236071 406294 236123
rect 406346 236111 406352 236123
rect 411760 236111 411766 236123
rect 406346 236083 411766 236111
rect 406346 236071 406352 236083
rect 411760 236071 411766 236083
rect 411818 236071 411824 236123
rect 208432 235997 208438 236049
rect 208490 236037 208496 236049
rect 223216 236037 223222 236049
rect 208490 236009 223222 236037
rect 208490 235997 208496 236009
rect 223216 235997 223222 236009
rect 223274 235997 223280 236049
rect 247984 235997 247990 236049
rect 248042 236037 248048 236049
rect 273616 236037 273622 236049
rect 248042 236009 273622 236037
rect 248042 235997 248048 236009
rect 273616 235997 273622 236009
rect 273674 235997 273680 236049
rect 280624 235997 280630 236049
rect 280682 236037 280688 236049
rect 322000 236037 322006 236049
rect 280682 236009 322006 236037
rect 280682 235997 280688 236009
rect 322000 235997 322006 236009
rect 322058 235997 322064 236049
rect 386704 235997 386710 236049
rect 386762 236037 386768 236049
rect 411472 236037 411478 236049
rect 386762 236009 411478 236037
rect 386762 235997 386768 236009
rect 411472 235997 411478 236009
rect 411530 235997 411536 236049
rect 207472 235923 207478 235975
rect 207530 235963 207536 235975
rect 223984 235963 223990 235975
rect 207530 235935 223990 235963
rect 207530 235923 207536 235935
rect 223984 235923 223990 235935
rect 224042 235923 224048 235975
rect 243280 235923 243286 235975
rect 243338 235963 243344 235975
rect 271024 235963 271030 235975
rect 243338 235935 271030 235963
rect 243338 235923 243344 235935
rect 271024 235923 271030 235935
rect 271082 235923 271088 235975
rect 279280 235923 279286 235975
rect 279338 235963 279344 235975
rect 319600 235963 319606 235975
rect 279338 235935 319606 235963
rect 279338 235923 279344 235935
rect 319600 235923 319606 235935
rect 319658 235923 319664 235975
rect 332560 235923 332566 235975
rect 332618 235963 332624 235975
rect 472336 235963 472342 235975
rect 332618 235935 472342 235963
rect 332618 235923 332624 235935
rect 472336 235923 472342 235935
rect 472394 235923 472400 235975
rect 209680 235849 209686 235901
rect 209738 235889 209744 235901
rect 226192 235889 226198 235901
rect 209738 235861 226198 235889
rect 209738 235849 209744 235861
rect 226192 235849 226198 235861
rect 226250 235849 226256 235901
rect 234256 235849 234262 235901
rect 234314 235889 234320 235901
rect 264880 235889 264886 235901
rect 234314 235861 264886 235889
rect 234314 235849 234320 235861
rect 264880 235849 264886 235861
rect 264938 235849 264944 235901
rect 273040 235849 273046 235901
rect 273098 235889 273104 235901
rect 305008 235889 305014 235901
rect 273098 235861 305014 235889
rect 273098 235849 273104 235861
rect 305008 235849 305014 235861
rect 305066 235849 305072 235901
rect 343504 235849 343510 235901
rect 343562 235889 343568 235901
rect 495760 235889 495766 235901
rect 343562 235861 495766 235889
rect 343562 235849 343568 235861
rect 495760 235849 495766 235861
rect 495818 235849 495824 235901
rect 208912 235775 208918 235827
rect 208970 235815 208976 235827
rect 226960 235815 226966 235827
rect 208970 235787 226966 235815
rect 208970 235775 208976 235787
rect 226960 235775 226966 235787
rect 227018 235775 227024 235827
rect 237520 235775 237526 235827
rect 237578 235815 237584 235827
rect 268144 235815 268150 235827
rect 237578 235787 268150 235815
rect 237578 235775 237584 235787
rect 268144 235775 268150 235787
rect 268202 235775 268208 235827
rect 276112 235775 276118 235827
rect 276170 235815 276176 235827
rect 308272 235815 308278 235827
rect 276170 235787 308278 235815
rect 276170 235775 276176 235787
rect 308272 235775 308278 235787
rect 308330 235775 308336 235827
rect 348880 235775 348886 235827
rect 348938 235815 348944 235827
rect 394576 235815 394582 235827
rect 348938 235787 394582 235815
rect 348938 235775 348944 235787
rect 394576 235775 394582 235787
rect 394634 235775 394640 235827
rect 403600 235775 403606 235827
rect 403658 235815 403664 235827
rect 588880 235815 588886 235827
rect 403658 235787 588886 235815
rect 403658 235775 403664 235787
rect 588880 235775 588886 235787
rect 588938 235775 588944 235827
rect 211216 235701 211222 235753
rect 211274 235741 211280 235753
rect 229264 235741 229270 235753
rect 211274 235713 229270 235741
rect 211274 235701 211280 235713
rect 229264 235701 229270 235713
rect 229322 235701 229328 235753
rect 231184 235701 231190 235753
rect 231242 235741 231248 235753
rect 259024 235741 259030 235753
rect 231242 235713 259030 235741
rect 231242 235701 231248 235713
rect 259024 235701 259030 235713
rect 259082 235701 259088 235753
rect 262864 235701 262870 235753
rect 262922 235741 262928 235753
rect 305104 235741 305110 235753
rect 262922 235713 305110 235741
rect 262922 235701 262928 235713
rect 305104 235701 305110 235713
rect 305162 235701 305168 235753
rect 313840 235701 313846 235753
rect 313898 235741 313904 235753
rect 360016 235741 360022 235753
rect 313898 235713 360022 235741
rect 313898 235701 313904 235713
rect 360016 235701 360022 235713
rect 360074 235701 360080 235753
rect 393424 235701 393430 235753
rect 393482 235741 393488 235753
rect 587056 235741 587062 235753
rect 393482 235713 587062 235741
rect 393482 235701 393488 235713
rect 587056 235701 587062 235713
rect 587114 235701 587120 235753
rect 210640 235627 210646 235679
rect 210698 235667 210704 235679
rect 230032 235667 230038 235679
rect 210698 235639 230038 235667
rect 210698 235627 210704 235639
rect 230032 235627 230038 235639
rect 230090 235627 230096 235679
rect 236464 235627 236470 235679
rect 236522 235667 236528 235679
rect 282928 235667 282934 235679
rect 236522 235639 282934 235667
rect 236522 235627 236528 235639
rect 282928 235627 282934 235639
rect 282986 235627 282992 235679
rect 285136 235627 285142 235679
rect 285194 235667 285200 235679
rect 323824 235667 323830 235679
rect 285194 235639 323830 235667
rect 285194 235627 285200 235639
rect 323824 235627 323830 235639
rect 323882 235627 323888 235679
rect 326128 235627 326134 235679
rect 326186 235667 326192 235679
rect 378832 235667 378838 235679
rect 326186 235639 378838 235667
rect 326186 235627 326192 235639
rect 378832 235627 378838 235639
rect 378890 235627 378896 235679
rect 385840 235627 385846 235679
rect 385898 235667 385904 235679
rect 580336 235667 580342 235679
rect 385898 235639 580342 235667
rect 385898 235627 385904 235639
rect 580336 235627 580342 235639
rect 580394 235627 580400 235679
rect 210064 235553 210070 235605
rect 210122 235593 210128 235605
rect 227824 235593 227830 235605
rect 210122 235565 227830 235593
rect 210122 235553 210128 235565
rect 227824 235553 227830 235565
rect 227882 235553 227888 235605
rect 239344 235553 239350 235605
rect 239402 235593 239408 235605
rect 285328 235593 285334 235605
rect 239402 235565 285334 235593
rect 239402 235553 239408 235565
rect 285328 235553 285334 235565
rect 285386 235553 285392 235605
rect 286672 235553 286678 235605
rect 286730 235593 286736 235605
rect 326704 235593 326710 235605
rect 286730 235565 326710 235593
rect 286730 235553 286736 235565
rect 326704 235553 326710 235565
rect 326762 235553 326768 235605
rect 332176 235553 332182 235605
rect 332234 235593 332240 235605
rect 383056 235593 383062 235605
rect 332234 235565 383062 235593
rect 332234 235553 332240 235565
rect 383056 235553 383062 235565
rect 383114 235553 383120 235605
rect 392176 235553 392182 235605
rect 392234 235593 392240 235605
rect 586288 235593 586294 235605
rect 392234 235565 586294 235593
rect 392234 235553 392240 235565
rect 586288 235553 586294 235565
rect 586346 235553 586352 235605
rect 212944 235479 212950 235531
rect 213002 235519 213008 235531
rect 232336 235519 232342 235531
rect 213002 235491 232342 235519
rect 213002 235479 213008 235491
rect 232336 235479 232342 235491
rect 232394 235479 232400 235531
rect 249712 235479 249718 235531
rect 249770 235519 249776 235531
rect 302320 235519 302326 235531
rect 249770 235491 302326 235519
rect 249770 235479 249776 235491
rect 302320 235479 302326 235491
rect 302378 235479 302384 235531
rect 309328 235479 309334 235531
rect 309386 235519 309392 235531
rect 362800 235519 362806 235531
rect 309386 235491 362806 235519
rect 309386 235479 309392 235491
rect 362800 235479 362806 235491
rect 362858 235479 362864 235531
rect 387664 235479 387670 235531
rect 387722 235519 387728 235531
rect 583408 235519 583414 235531
rect 387722 235491 583414 235519
rect 387722 235479 387728 235491
rect 583408 235479 583414 235491
rect 583466 235479 583472 235531
rect 42160 235405 42166 235457
rect 42218 235445 42224 235457
rect 42928 235445 42934 235457
rect 42218 235417 42934 235445
rect 42218 235405 42224 235417
rect 42928 235405 42934 235417
rect 42986 235405 42992 235457
rect 211984 235405 211990 235457
rect 212042 235445 212048 235457
rect 233008 235445 233014 235457
rect 212042 235417 233014 235445
rect 212042 235405 212048 235417
rect 233008 235405 233014 235417
rect 233066 235405 233072 235457
rect 238000 235405 238006 235457
rect 238058 235445 238064 235457
rect 285904 235445 285910 235457
rect 238058 235417 285910 235445
rect 238058 235405 238064 235417
rect 285904 235405 285910 235417
rect 285962 235405 285968 235457
rect 295216 235405 295222 235457
rect 295274 235445 295280 235457
rect 348688 235445 348694 235457
rect 295274 235417 348694 235445
rect 295274 235405 295280 235417
rect 348688 235405 348694 235417
rect 348746 235405 348752 235457
rect 389872 235405 389878 235457
rect 389930 235445 389936 235457
rect 587920 235445 587926 235457
rect 389930 235417 587926 235445
rect 389930 235405 389936 235417
rect 587920 235405 587926 235417
rect 587978 235405 587984 235457
rect 214192 235331 214198 235383
rect 214250 235371 214256 235383
rect 235312 235371 235318 235383
rect 214250 235343 235318 235371
rect 214250 235331 214256 235343
rect 235312 235331 235318 235343
rect 235370 235331 235376 235383
rect 242128 235331 242134 235383
rect 242186 235371 242192 235383
rect 293392 235371 293398 235383
rect 242186 235343 293398 235371
rect 242186 235331 242192 235343
rect 293392 235331 293398 235343
rect 293450 235331 293456 235383
rect 299824 235331 299830 235383
rect 299882 235371 299888 235383
rect 356464 235371 356470 235383
rect 299882 235343 356470 235371
rect 299882 235331 299888 235343
rect 356464 235331 356470 235343
rect 356522 235331 356528 235383
rect 385744 235371 385750 235383
rect 368626 235343 385750 235371
rect 206992 235257 206998 235309
rect 207050 235297 207056 235309
rect 221776 235297 221782 235309
rect 207050 235269 221782 235297
rect 207050 235257 207056 235269
rect 221776 235257 221782 235269
rect 221834 235257 221840 235309
rect 223888 235257 223894 235309
rect 223946 235297 223952 235309
rect 244720 235297 244726 235309
rect 223946 235269 244726 235297
rect 223946 235257 223952 235269
rect 244720 235257 244726 235269
rect 244778 235257 244784 235309
rect 246640 235257 246646 235309
rect 246698 235297 246704 235309
rect 299248 235297 299254 235309
rect 246698 235269 299254 235297
rect 246698 235257 246704 235269
rect 299248 235257 299254 235269
rect 299306 235257 299312 235309
rect 301744 235257 301750 235309
rect 301802 235297 301808 235309
rect 358576 235297 358582 235309
rect 301802 235269 358582 235297
rect 301802 235257 301808 235269
rect 358576 235257 358582 235269
rect 358634 235257 358640 235309
rect 361360 235257 361366 235309
rect 361418 235297 361424 235309
rect 368626 235297 368654 235343
rect 385744 235331 385750 235343
rect 385802 235331 385808 235383
rect 394864 235331 394870 235383
rect 394922 235371 394928 235383
rect 597712 235371 597718 235383
rect 394922 235343 597718 235371
rect 394922 235331 394928 235343
rect 597712 235331 597718 235343
rect 597770 235331 597776 235383
rect 361418 235269 368654 235297
rect 361418 235257 361424 235269
rect 370192 235257 370198 235309
rect 370250 235297 370256 235309
rect 385936 235297 385942 235309
rect 370250 235269 385942 235297
rect 370250 235257 370256 235269
rect 385936 235257 385942 235269
rect 385994 235257 386000 235309
rect 394960 235257 394966 235309
rect 395018 235297 395024 235309
rect 598480 235297 598486 235309
rect 395018 235269 598486 235297
rect 395018 235257 395024 235269
rect 598480 235257 598486 235269
rect 598538 235257 598544 235309
rect 220624 235183 220630 235235
rect 220682 235223 220688 235235
rect 240496 235223 240502 235235
rect 220682 235195 240502 235223
rect 220682 235183 220688 235195
rect 240496 235183 240502 235195
rect 240554 235183 240560 235235
rect 240592 235183 240598 235235
rect 240650 235223 240656 235235
rect 290416 235223 290422 235235
rect 240650 235195 290422 235223
rect 240650 235183 240656 235195
rect 290416 235183 290422 235195
rect 290474 235183 290480 235235
rect 342544 235183 342550 235235
rect 342602 235223 342608 235235
rect 391600 235223 391606 235235
rect 342602 235195 391606 235223
rect 342602 235183 342608 235195
rect 391600 235183 391606 235195
rect 391658 235183 391664 235235
rect 396304 235183 396310 235235
rect 396362 235223 396368 235235
rect 600784 235223 600790 235235
rect 396362 235195 600790 235223
rect 396362 235183 396368 235195
rect 600784 235183 600790 235195
rect 600842 235183 600848 235235
rect 211600 235109 211606 235161
rect 211658 235149 211664 235161
rect 230704 235149 230710 235161
rect 211658 235121 230710 235149
rect 211658 235109 211664 235121
rect 230704 235109 230710 235121
rect 230762 235109 230768 235161
rect 232912 235109 232918 235161
rect 232970 235149 232976 235161
rect 262000 235149 262006 235161
rect 232970 235121 262006 235149
rect 232970 235109 232976 235121
rect 262000 235109 262006 235121
rect 262058 235109 262064 235161
rect 266128 235109 266134 235161
rect 266186 235149 266192 235161
rect 324112 235149 324118 235161
rect 266186 235121 324118 235149
rect 266186 235109 266192 235121
rect 324112 235109 324118 235121
rect 324170 235109 324176 235161
rect 334960 235109 334966 235161
rect 335018 235149 335024 235161
rect 391696 235149 391702 235161
rect 335018 235121 391702 235149
rect 335018 235109 335024 235121
rect 391696 235109 391702 235121
rect 391754 235109 391760 235161
rect 398992 235109 398998 235161
rect 399050 235149 399056 235161
rect 605968 235149 605974 235161
rect 399050 235121 605974 235149
rect 399050 235109 399056 235121
rect 605968 235109 605974 235121
rect 606026 235109 606032 235161
rect 213424 235035 213430 235087
rect 213482 235075 213488 235087
rect 213482 235047 235646 235075
rect 213482 235035 213488 235047
rect 211024 234961 211030 235013
rect 211082 235001 211088 235013
rect 231568 235001 231574 235013
rect 211082 234973 231574 235001
rect 211082 234961 211088 234973
rect 231568 234961 231574 234973
rect 231626 234961 231632 235013
rect 235618 235001 235646 235047
rect 235696 235035 235702 235087
rect 235754 235075 235760 235087
rect 266416 235075 266422 235087
rect 235754 235047 266422 235075
rect 235754 235035 235760 235047
rect 266416 235035 266422 235047
rect 266474 235035 266480 235087
rect 268912 235035 268918 235087
rect 268970 235075 268976 235087
rect 331408 235075 331414 235087
rect 268970 235047 331414 235075
rect 268970 235035 268976 235047
rect 331408 235035 331414 235047
rect 331466 235035 331472 235087
rect 333424 235035 333430 235087
rect 333482 235075 333488 235087
rect 394672 235075 394678 235087
rect 333482 235047 394678 235075
rect 333482 235035 333488 235047
rect 394672 235035 394678 235047
rect 394730 235035 394736 235087
rect 398608 235035 398614 235087
rect 398666 235075 398672 235087
rect 605296 235075 605302 235087
rect 398666 235047 605302 235075
rect 398666 235035 398672 235047
rect 605296 235035 605302 235047
rect 605354 235035 605360 235087
rect 235984 235001 235990 235013
rect 235618 234973 235990 235001
rect 235984 234961 235990 234973
rect 236042 234961 236048 235013
rect 243856 234961 243862 235013
rect 243914 235001 243920 235013
rect 296464 235001 296470 235013
rect 243914 234973 296470 235001
rect 243914 234961 243920 234973
rect 296464 234961 296470 234973
rect 296522 234961 296528 235013
rect 296560 234961 296566 235013
rect 296618 235001 296624 235013
rect 360208 235001 360214 235013
rect 296618 234973 360214 235001
rect 296618 234961 296624 234973
rect 360208 234961 360214 234973
rect 360266 234961 360272 235013
rect 378448 234961 378454 235013
rect 378506 235001 378512 235013
rect 399568 235001 399574 235013
rect 378506 234973 399574 235001
rect 378506 234961 378512 234973
rect 399568 234961 399574 234973
rect 399626 234961 399632 235013
rect 406672 234961 406678 235013
rect 406730 235001 406736 235013
rect 621808 235001 621814 235013
rect 406730 234973 621814 235001
rect 406730 234961 406736 234973
rect 621808 234961 621814 234973
rect 621866 234961 621872 235013
rect 208816 234887 208822 234939
rect 208874 234927 208880 234939
rect 224752 234927 224758 234939
rect 208874 234899 224758 234927
rect 208874 234887 208880 234899
rect 224752 234887 224758 234899
rect 224810 234887 224816 234939
rect 225520 234887 225526 234939
rect 225578 234927 225584 234939
rect 260176 234927 260182 234939
rect 225578 234899 260182 234927
rect 225578 234887 225584 234899
rect 260176 234887 260182 234899
rect 260234 234887 260240 234939
rect 260272 234887 260278 234939
rect 260330 234927 260336 234939
rect 325264 234927 325270 234939
rect 260330 234899 325270 234927
rect 260330 234887 260336 234899
rect 325264 234887 325270 234899
rect 325322 234887 325328 234939
rect 327664 234887 327670 234939
rect 327722 234927 327728 234939
rect 392464 234927 392470 234939
rect 327722 234899 392470 234927
rect 327722 234887 327728 234899
rect 392464 234887 392470 234899
rect 392522 234887 392528 234939
rect 409168 234887 409174 234939
rect 409226 234927 409232 234939
rect 626416 234927 626422 234939
rect 409226 234899 626422 234927
rect 409226 234887 409232 234899
rect 626416 234887 626422 234899
rect 626474 234887 626480 234939
rect 42160 234813 42166 234865
rect 42218 234853 42224 234865
rect 42736 234853 42742 234865
rect 42218 234825 42742 234853
rect 42218 234813 42224 234825
rect 42736 234813 42742 234825
rect 42794 234813 42800 234865
rect 206512 234813 206518 234865
rect 206570 234853 206576 234865
rect 222448 234853 222454 234865
rect 206570 234825 222454 234853
rect 206570 234813 206576 234825
rect 222448 234813 222454 234825
rect 222506 234813 222512 234865
rect 254224 234813 254230 234865
rect 254282 234853 254288 234865
rect 306640 234853 306646 234865
rect 254282 234825 306646 234853
rect 254282 234813 254288 234825
rect 306640 234813 306646 234825
rect 306698 234813 306704 234865
rect 321616 234813 321622 234865
rect 321674 234853 321680 234865
rect 370192 234853 370198 234865
rect 321674 234825 370198 234853
rect 321674 234813 321680 234825
rect 370192 234813 370198 234825
rect 370250 234813 370256 234865
rect 370288 234813 370294 234865
rect 370346 234853 370352 234865
rect 386896 234853 386902 234865
rect 370346 234825 386902 234853
rect 370346 234813 370352 234825
rect 386896 234813 386902 234825
rect 386954 234813 386960 234865
rect 410800 234813 410806 234865
rect 410858 234853 410864 234865
rect 630160 234853 630166 234865
rect 410858 234825 630166 234853
rect 410858 234813 410864 234825
rect 630160 234813 630166 234825
rect 630218 234813 630224 234865
rect 203248 234739 203254 234791
rect 203306 234779 203312 234791
rect 203306 234751 209246 234779
rect 203306 234739 203312 234751
rect 205552 234665 205558 234717
rect 205610 234705 205616 234717
rect 207280 234705 207286 234717
rect 205610 234677 207286 234705
rect 205610 234665 205616 234677
rect 207280 234665 207286 234677
rect 207338 234665 207344 234717
rect 209218 234705 209246 234751
rect 209296 234739 209302 234791
rect 209354 234779 209360 234791
rect 228496 234779 228502 234791
rect 209354 234751 228502 234779
rect 209354 234739 209360 234751
rect 228496 234739 228502 234751
rect 228554 234739 228560 234791
rect 229744 234739 229750 234791
rect 229802 234779 229808 234791
rect 253552 234779 253558 234791
rect 229802 234751 253558 234779
rect 229802 234739 229808 234751
rect 253552 234739 253558 234751
rect 253610 234739 253616 234791
rect 257488 234739 257494 234791
rect 257546 234779 257552 234791
rect 308176 234779 308182 234791
rect 257546 234751 308182 234779
rect 257546 234739 257552 234751
rect 308176 234739 308182 234751
rect 308234 234739 308240 234791
rect 315280 234739 315286 234791
rect 315338 234779 315344 234791
rect 394864 234779 394870 234791
rect 315338 234751 394870 234779
rect 315338 234739 315344 234751
rect 394864 234739 394870 234751
rect 394922 234739 394928 234791
rect 410032 234739 410038 234791
rect 410090 234779 410096 234791
rect 628624 234779 628630 234791
rect 410090 234751 628630 234779
rect 410090 234739 410096 234751
rect 628624 234739 628630 234751
rect 628682 234739 628688 234791
rect 215824 234705 215830 234717
rect 209218 234677 215830 234705
rect 215824 234665 215830 234677
rect 215882 234665 215888 234717
rect 225136 234665 225142 234717
rect 225194 234705 225200 234717
rect 247696 234705 247702 234717
rect 225194 234677 247702 234705
rect 225194 234665 225200 234677
rect 247696 234665 247702 234677
rect 247754 234665 247760 234717
rect 251152 234665 251158 234717
rect 251210 234705 251216 234717
rect 304144 234705 304150 234717
rect 251210 234677 304150 234705
rect 251210 234665 251216 234677
rect 304144 234665 304150 234677
rect 304202 234665 304208 234717
rect 308464 234665 308470 234717
rect 308522 234705 308528 234717
rect 411568 234705 411574 234717
rect 308522 234677 411574 234705
rect 308522 234665 308528 234677
rect 411568 234665 411574 234677
rect 411626 234665 411632 234717
rect 412144 234665 412150 234717
rect 412202 234705 412208 234717
rect 632368 234705 632374 234717
rect 412202 234677 632374 234705
rect 412202 234665 412208 234677
rect 632368 234665 632374 234677
rect 632426 234665 632432 234717
rect 204784 234591 204790 234643
rect 204842 234631 204848 234643
rect 211984 234631 211990 234643
rect 204842 234603 211990 234631
rect 204842 234591 204848 234603
rect 211984 234591 211990 234603
rect 212042 234591 212048 234643
rect 240208 234591 240214 234643
rect 240266 234631 240272 234643
rect 264688 234631 264694 234643
rect 240266 234603 264694 234631
rect 240266 234591 240272 234603
rect 264688 234591 264694 234603
rect 264746 234591 264752 234643
rect 267472 234591 267478 234643
rect 267530 234631 267536 234643
rect 285040 234631 285046 234643
rect 267530 234603 285046 234631
rect 267530 234591 267536 234603
rect 285040 234591 285046 234603
rect 285098 234591 285104 234643
rect 287056 234591 287062 234643
rect 287114 234631 287120 234643
rect 318352 234631 318358 234643
rect 287114 234603 318358 234631
rect 287114 234591 287120 234603
rect 318352 234591 318358 234603
rect 318410 234591 318416 234643
rect 320272 234591 320278 234643
rect 320330 234631 320336 234643
rect 448240 234631 448246 234643
rect 320330 234603 448246 234631
rect 320330 234591 320336 234603
rect 448240 234591 448246 234603
rect 448298 234591 448304 234643
rect 202864 234517 202870 234569
rect 202922 234557 202928 234569
rect 214864 234557 214870 234569
rect 202922 234529 214870 234557
rect 202922 234517 202928 234529
rect 214864 234517 214870 234529
rect 214922 234517 214928 234569
rect 235600 234517 235606 234569
rect 235658 234557 235664 234569
rect 250576 234557 250582 234569
rect 235658 234529 250582 234557
rect 235658 234517 235664 234529
rect 250576 234517 250582 234529
rect 250634 234517 250640 234569
rect 255280 234517 255286 234569
rect 255338 234557 255344 234569
rect 278224 234557 278230 234569
rect 255338 234529 278230 234557
rect 255338 234517 255344 234529
rect 278224 234517 278230 234529
rect 278282 234517 278288 234569
rect 283888 234517 283894 234569
rect 283946 234557 283952 234569
rect 320848 234557 320854 234569
rect 283946 234529 320854 234557
rect 283946 234517 283952 234529
rect 320848 234517 320854 234529
rect 320906 234517 320912 234569
rect 329296 234517 329302 234569
rect 329354 234557 329360 234569
rect 449296 234557 449302 234569
rect 329354 234529 449302 234557
rect 329354 234517 329360 234529
rect 449296 234517 449302 234529
rect 449354 234517 449360 234569
rect 202000 234443 202006 234495
rect 202058 234483 202064 234495
rect 213424 234483 213430 234495
rect 202058 234455 213430 234483
rect 202058 234443 202064 234455
rect 213424 234443 213430 234455
rect 213482 234443 213488 234495
rect 239824 234443 239830 234495
rect 239882 234483 239888 234495
rect 260464 234483 260470 234495
rect 239882 234455 260470 234483
rect 239882 234443 239888 234455
rect 260464 234443 260470 234455
rect 260522 234443 260528 234495
rect 262480 234443 262486 234495
rect 262538 234483 262544 234495
rect 290896 234483 290902 234495
rect 262538 234455 290902 234483
rect 262538 234443 262544 234455
rect 290896 234443 290902 234455
rect 290954 234443 290960 234495
rect 297136 234443 297142 234495
rect 297194 234483 297200 234495
rect 319408 234483 319414 234495
rect 297194 234455 319414 234483
rect 297194 234443 297200 234455
rect 319408 234443 319414 234455
rect 319466 234443 319472 234495
rect 323536 234443 323542 234495
rect 323594 234483 323600 234495
rect 434896 234483 434902 234495
rect 323594 234455 434902 234483
rect 323594 234443 323600 234455
rect 434896 234443 434902 234455
rect 434954 234443 434960 234495
rect 206128 234369 206134 234421
rect 206186 234409 206192 234421
rect 221008 234409 221014 234421
rect 206186 234381 221014 234409
rect 206186 234369 206192 234381
rect 221008 234369 221014 234381
rect 221066 234369 221072 234421
rect 250480 234369 250486 234421
rect 250538 234409 250544 234421
rect 267952 234409 267958 234421
rect 250538 234381 267958 234409
rect 250538 234369 250544 234381
rect 267952 234369 267958 234381
rect 268010 234369 268016 234421
rect 271600 234369 271606 234421
rect 271658 234409 271664 234421
rect 302224 234409 302230 234421
rect 271658 234381 302230 234409
rect 271658 234369 271664 234381
rect 302224 234369 302230 234381
rect 302282 234369 302288 234421
rect 313840 234409 313846 234421
rect 306658 234381 313846 234409
rect 207856 234295 207862 234347
rect 207914 234335 207920 234347
rect 207914 234307 211934 234335
rect 207914 234295 207920 234307
rect 200272 234221 200278 234273
rect 200330 234261 200336 234273
rect 210352 234261 210358 234273
rect 200330 234233 210358 234261
rect 200330 234221 200336 234233
rect 210352 234221 210358 234233
rect 210410 234221 210416 234273
rect 200176 234147 200182 234199
rect 200234 234187 200240 234199
rect 208816 234187 208822 234199
rect 200234 234159 208822 234187
rect 200234 234147 200240 234159
rect 208816 234147 208822 234159
rect 208874 234147 208880 234199
rect 211906 234187 211934 234307
rect 237040 234295 237046 234347
rect 237098 234335 237104 234347
rect 258448 234335 258454 234347
rect 237098 234307 258454 234335
rect 237098 234295 237104 234307
rect 258448 234295 258454 234307
rect 258506 234295 258512 234347
rect 261232 234295 261238 234347
rect 261290 234335 261296 234347
rect 288016 234335 288022 234347
rect 261290 234307 288022 234335
rect 261290 234295 261296 234307
rect 288016 234295 288022 234307
rect 288074 234295 288080 234347
rect 292912 234295 292918 234347
rect 292970 234335 292976 234347
rect 306658 234335 306686 234381
rect 313840 234369 313846 234381
rect 313898 234369 313904 234421
rect 314416 234369 314422 234421
rect 314474 234409 314480 234421
rect 423376 234409 423382 234421
rect 314474 234381 423382 234409
rect 314474 234369 314480 234381
rect 423376 234369 423382 234381
rect 423434 234369 423440 234421
rect 292970 234307 306686 234335
rect 292970 234295 292976 234307
rect 312688 234295 312694 234347
rect 312746 234335 312752 234347
rect 418288 234335 418294 234347
rect 312746 234307 418294 234335
rect 312746 234295 312752 234307
rect 418288 234295 418294 234307
rect 418346 234295 418352 234347
rect 211984 234221 211990 234273
rect 212042 234261 212048 234273
rect 219376 234261 219382 234273
rect 212042 234233 219382 234261
rect 212042 234221 212048 234233
rect 219376 234221 219382 234233
rect 219434 234221 219440 234273
rect 256528 234221 256534 234273
rect 256586 234261 256592 234273
rect 278128 234261 278134 234273
rect 256586 234233 278134 234261
rect 256586 234221 256592 234233
rect 278128 234221 278134 234233
rect 278186 234221 278192 234273
rect 290320 234221 290326 234273
rect 290378 234261 290384 234273
rect 334288 234261 334294 234273
rect 290378 234233 334294 234261
rect 290378 234221 290384 234233
rect 334288 234221 334294 234233
rect 334346 234221 334352 234273
rect 339472 234221 339478 234273
rect 339530 234261 339536 234273
rect 378640 234261 378646 234273
rect 339530 234233 378646 234261
rect 339530 234221 339536 234233
rect 378640 234221 378646 234233
rect 378698 234221 378704 234273
rect 378832 234221 378838 234273
rect 378890 234261 378896 234273
rect 400048 234261 400054 234273
rect 378890 234233 400054 234261
rect 378890 234221 378896 234233
rect 400048 234221 400054 234233
rect 400106 234221 400112 234273
rect 403696 234221 403702 234273
rect 403754 234261 403760 234273
rect 501040 234261 501046 234273
rect 403754 234233 501046 234261
rect 403754 234221 403760 234233
rect 501040 234221 501046 234233
rect 501098 234221 501104 234273
rect 225520 234187 225526 234199
rect 211906 234159 225526 234187
rect 225520 234147 225526 234159
rect 225578 234147 225584 234199
rect 244336 234147 244342 234199
rect 244394 234187 244400 234199
rect 263632 234187 263638 234199
rect 244394 234159 263638 234187
rect 244394 234147 244400 234159
rect 263632 234147 263638 234159
rect 263690 234147 263696 234199
rect 268528 234147 268534 234199
rect 268586 234187 268592 234199
rect 293776 234187 293782 234199
rect 268586 234159 293782 234187
rect 268586 234147 268592 234159
rect 293776 234147 293782 234159
rect 293834 234147 293840 234199
rect 295696 234147 295702 234199
rect 295754 234187 295760 234199
rect 342352 234187 342358 234199
rect 295754 234159 342358 234187
rect 295754 234147 295760 234159
rect 342352 234147 342358 234159
rect 342410 234147 342416 234199
rect 345904 234147 345910 234199
rect 345962 234187 345968 234199
rect 400144 234187 400150 234199
rect 345962 234159 400150 234187
rect 345962 234147 345968 234159
rect 400144 234147 400150 234159
rect 400202 234147 400208 234199
rect 401776 234147 401782 234199
rect 401834 234187 401840 234199
rect 484624 234187 484630 234199
rect 401834 234159 484630 234187
rect 401834 234147 401840 234159
rect 484624 234147 484630 234159
rect 484682 234147 484688 234199
rect 198736 234073 198742 234125
rect 198794 234113 198800 234125
rect 207376 234113 207382 234125
rect 198794 234085 207382 234113
rect 198794 234073 198800 234085
rect 207376 234073 207382 234085
rect 207434 234073 207440 234125
rect 247408 234073 247414 234125
rect 247466 234113 247472 234125
rect 266320 234113 266326 234125
rect 247466 234085 266326 234113
rect 247466 234073 247472 234085
rect 266320 234073 266326 234085
rect 266378 234073 266384 234125
rect 267088 234073 267094 234125
rect 267146 234113 267152 234125
rect 290992 234113 290998 234125
rect 267146 234085 290998 234113
rect 267146 234073 267152 234085
rect 290992 234073 290998 234085
rect 291050 234073 291056 234125
rect 294448 234073 294454 234125
rect 294506 234113 294512 234125
rect 331216 234113 331222 234125
rect 294506 234085 331222 234113
rect 294506 234073 294512 234085
rect 331216 234073 331222 234085
rect 331274 234073 331280 234125
rect 338032 234073 338038 234125
rect 338090 234113 338096 234125
rect 378544 234113 378550 234125
rect 338090 234085 378550 234113
rect 338090 234073 338096 234085
rect 378544 234073 378550 234085
rect 378602 234073 378608 234125
rect 378640 234073 378646 234125
rect 378698 234113 378704 234125
rect 394576 234113 394582 234125
rect 378698 234085 394582 234113
rect 378698 234073 378704 234085
rect 394576 234073 394582 234085
rect 394634 234073 394640 234125
rect 396688 234073 396694 234125
rect 396746 234113 396752 234125
rect 475216 234113 475222 234125
rect 396746 234085 475222 234113
rect 396746 234073 396752 234085
rect 475216 234073 475222 234085
rect 475274 234073 475280 234125
rect 42064 233999 42070 234051
rect 42122 234039 42128 234051
rect 42832 234039 42838 234051
rect 42122 234011 42838 234039
rect 42122 233999 42128 234011
rect 42832 233999 42838 234011
rect 42890 233999 42896 234051
rect 198352 233999 198358 234051
rect 198410 234039 198416 234051
rect 205936 234039 205942 234051
rect 198410 234011 205942 234039
rect 198410 233999 198416 234011
rect 205936 233999 205942 234011
rect 205994 233999 206000 234051
rect 217936 234039 217942 234051
rect 206818 234011 217942 234039
rect 197488 233925 197494 233977
rect 197546 233965 197552 233977
rect 204304 233965 204310 233977
rect 197546 233937 204310 233965
rect 197546 233925 197552 233937
rect 204304 233925 204310 233937
rect 204362 233925 204368 233977
rect 204400 233925 204406 233977
rect 204458 233965 204464 233977
rect 206818 233965 206846 234011
rect 217936 233999 217942 234011
rect 217994 233999 218000 234051
rect 259792 233999 259798 234051
rect 259850 234039 259856 234051
rect 282064 234039 282070 234051
rect 259850 234011 282070 234039
rect 259850 233999 259856 234011
rect 282064 233999 282070 234011
rect 282122 233999 282128 234051
rect 305200 233999 305206 234051
rect 305258 234039 305264 234051
rect 351376 234039 351382 234051
rect 305258 234011 351382 234039
rect 305258 233999 305264 234011
rect 351376 233999 351382 234011
rect 351434 233999 351440 234051
rect 358000 233999 358006 234051
rect 358058 234039 358064 234051
rect 378832 234039 378838 234051
rect 358058 234011 378838 234039
rect 358058 233999 358064 234011
rect 378832 233999 378838 234011
rect 378890 233999 378896 234051
rect 395920 233999 395926 234051
rect 395978 234039 395984 234051
rect 398128 234039 398134 234051
rect 395978 234011 398134 234039
rect 395978 233999 395984 234011
rect 398128 233999 398134 234011
rect 398186 233999 398192 234051
rect 398224 233999 398230 234051
rect 398282 234039 398288 234051
rect 405232 234039 405238 234051
rect 398282 234011 405238 234039
rect 398282 233999 398288 234011
rect 405232 233999 405238 234011
rect 405290 233999 405296 234051
rect 204458 233937 206846 233965
rect 204458 233925 204464 233937
rect 206896 233925 206902 233977
rect 206954 233965 206960 233977
rect 220240 233965 220246 233977
rect 206954 233937 220246 233965
rect 206954 233925 206960 233937
rect 220240 233925 220246 233937
rect 220298 233925 220304 233977
rect 258352 233925 258358 233977
rect 258410 233965 258416 233977
rect 277072 233965 277078 233977
rect 258410 233937 277078 233965
rect 258410 233925 258416 233937
rect 277072 233925 277078 233937
rect 277130 233925 277136 233977
rect 294832 233925 294838 233977
rect 294890 233965 294896 233977
rect 339760 233965 339766 233977
rect 294890 233937 339766 233965
rect 294890 233925 294896 233937
rect 339760 233925 339766 233937
rect 339818 233925 339824 233977
rect 361264 233925 361270 233977
rect 361322 233965 361328 233977
rect 432016 233965 432022 233977
rect 361322 233937 432022 233965
rect 361322 233925 361328 233937
rect 432016 233925 432022 233937
rect 432074 233925 432080 233977
rect 199120 233851 199126 233903
rect 199178 233891 199184 233903
rect 205072 233891 205078 233903
rect 199178 233863 205078 233891
rect 199178 233851 199184 233863
rect 205072 233851 205078 233863
rect 205130 233851 205136 233903
rect 205168 233851 205174 233903
rect 205226 233891 205232 233903
rect 205226 233863 215678 233891
rect 205226 233851 205232 233863
rect 196912 233777 196918 233829
rect 196970 233817 196976 233829
rect 202864 233817 202870 233829
rect 196970 233789 202870 233817
rect 196970 233777 196976 233789
rect 202864 233777 202870 233789
rect 202922 233777 202928 233829
rect 204208 233777 204214 233829
rect 204266 233817 204272 233829
rect 215536 233817 215542 233829
rect 204266 233789 215542 233817
rect 204266 233777 204272 233789
rect 215536 233777 215542 233789
rect 215594 233777 215600 233829
rect 196528 233703 196534 233755
rect 196586 233743 196592 233755
rect 200560 233743 200566 233755
rect 196586 233715 200566 233743
rect 196586 233703 196592 233715
rect 200560 233703 200566 233715
rect 200618 233703 200624 233755
rect 201520 233703 201526 233755
rect 201578 233743 201584 233755
rect 211888 233743 211894 233755
rect 201578 233715 211894 233743
rect 201578 233703 201584 233715
rect 211888 233703 211894 233715
rect 211946 233703 211952 233755
rect 215650 233743 215678 233863
rect 215824 233851 215830 233903
rect 215882 233891 215888 233903
rect 216496 233891 216502 233903
rect 215882 233863 216502 233891
rect 215882 233851 215888 233863
rect 216496 233851 216502 233863
rect 216554 233851 216560 233903
rect 253456 233851 253462 233903
rect 253514 233891 253520 233903
rect 270832 233891 270838 233903
rect 253514 233863 270838 233891
rect 253514 233851 253520 233863
rect 270832 233851 270838 233863
rect 270890 233851 270896 233903
rect 296080 233851 296086 233903
rect 296138 233891 296144 233903
rect 339088 233891 339094 233903
rect 296138 233863 339094 233891
rect 296138 233851 296144 233863
rect 339088 233851 339094 233863
rect 339146 233851 339152 233903
rect 352144 233851 352150 233903
rect 352202 233891 352208 233903
rect 361072 233891 361078 233903
rect 352202 233863 361078 233891
rect 352202 233851 352208 233863
rect 361072 233851 361078 233863
rect 361130 233851 361136 233903
rect 378544 233851 378550 233903
rect 378602 233891 378608 233903
rect 386800 233891 386806 233903
rect 378602 233863 386806 233891
rect 378602 233851 378608 233863
rect 386800 233851 386806 233863
rect 386858 233851 386864 233903
rect 386896 233851 386902 233903
rect 386954 233891 386960 233903
rect 427888 233891 427894 233903
rect 386954 233863 427894 233891
rect 386954 233851 386960 233863
rect 427888 233851 427894 233863
rect 427946 233851 427952 233903
rect 306256 233777 306262 233829
rect 306314 233817 306320 233829
rect 345520 233817 345526 233829
rect 306314 233789 345526 233817
rect 306314 233777 306320 233789
rect 345520 233777 345526 233789
rect 345578 233777 345584 233829
rect 354928 233777 354934 233829
rect 354986 233817 354992 233829
rect 404656 233817 404662 233829
rect 354986 233789 404662 233817
rect 354986 233777 354992 233789
rect 404656 233777 404662 233789
rect 404714 233777 404720 233829
rect 217168 233743 217174 233755
rect 215650 233715 217174 233743
rect 217168 233703 217174 233715
rect 217226 233703 217232 233755
rect 297232 233703 297238 233755
rect 297290 233743 297296 233755
rect 328336 233743 328342 233755
rect 297290 233715 328342 233743
rect 297290 233703 297296 233715
rect 328336 233703 328342 233715
rect 328394 233703 328400 233755
rect 330736 233703 330742 233755
rect 330794 233743 330800 233755
rect 371632 233743 371638 233755
rect 330794 233715 371638 233743
rect 330794 233703 330800 233715
rect 371632 233703 371638 233715
rect 371690 233703 371696 233755
rect 383632 233703 383638 233755
rect 383690 233743 383696 233755
rect 407632 233743 407638 233755
rect 383690 233715 407638 233743
rect 383690 233703 383696 233715
rect 407632 233703 407638 233715
rect 407690 233703 407696 233755
rect 195664 233629 195670 233681
rect 195722 233669 195728 233681
rect 201328 233669 201334 233681
rect 195722 233641 201334 233669
rect 195722 233629 195728 233641
rect 201328 233629 201334 233641
rect 201386 233629 201392 233681
rect 202480 233629 202486 233681
rect 202538 233669 202544 233681
rect 212560 233669 212566 233681
rect 202538 233641 212566 233669
rect 202538 233629 202544 233641
rect 212560 233629 212566 233641
rect 212618 233629 212624 233681
rect 302896 233629 302902 233681
rect 302954 233669 302960 233681
rect 334096 233669 334102 233681
rect 302954 233641 334102 233669
rect 302954 233629 302960 233641
rect 334096 233629 334102 233641
rect 334154 233629 334160 233681
rect 360304 233629 360310 233681
rect 360362 233669 360368 233681
rect 360976 233669 360982 233681
rect 360362 233641 360982 233669
rect 360362 233629 360368 233641
rect 360976 233629 360982 233641
rect 361034 233629 361040 233681
rect 361072 233629 361078 233681
rect 361130 233669 361136 233681
rect 400336 233669 400342 233681
rect 361130 233641 400342 233669
rect 361130 233629 361136 233641
rect 400336 233629 400342 233641
rect 400394 233629 400400 233681
rect 192880 233555 192886 233607
rect 192938 233595 192944 233607
rect 195280 233595 195286 233607
rect 192938 233567 195286 233595
rect 192938 233555 192944 233567
rect 195280 233555 195286 233567
rect 195338 233555 195344 233607
rect 195568 233555 195574 233607
rect 195626 233595 195632 233607
rect 199792 233595 199798 233607
rect 195626 233567 199798 233595
rect 195626 233555 195632 233567
rect 199792 233555 199798 233567
rect 199850 233555 199856 233607
rect 201040 233555 201046 233607
rect 201098 233595 201104 233607
rect 209680 233595 209686 233607
rect 201098 233567 209686 233595
rect 201098 233555 201104 233567
rect 209680 233555 209686 233567
rect 209738 233555 209744 233607
rect 218704 233595 218710 233607
rect 210754 233567 218710 233595
rect 194224 233481 194230 233533
rect 194282 233521 194288 233533
rect 198352 233521 198358 233533
rect 194282 233493 198358 233521
rect 194282 233481 194288 233493
rect 198352 233481 198358 233493
rect 198410 233481 198416 233533
rect 200656 233481 200662 233533
rect 200714 233521 200720 233533
rect 208144 233521 208150 233533
rect 200714 233493 208150 233521
rect 200714 233481 200720 233493
rect 208144 233481 208150 233493
rect 208202 233481 208208 233533
rect 194608 233407 194614 233459
rect 194666 233447 194672 233459
rect 196048 233447 196054 233459
rect 194666 233419 196054 233447
rect 194666 233407 194672 233419
rect 196048 233407 196054 233419
rect 196106 233407 196112 233459
rect 196144 233407 196150 233459
rect 196202 233447 196208 233459
rect 199120 233447 199126 233459
rect 196202 233419 199126 233447
rect 196202 233407 196208 233419
rect 199120 233407 199126 233419
rect 199178 233407 199184 233459
rect 199696 233407 199702 233459
rect 199754 233447 199760 233459
rect 206608 233447 206614 233459
rect 199754 233419 206614 233447
rect 199754 233407 199760 233419
rect 206608 233407 206614 233419
rect 206666 233407 206672 233459
rect 207280 233407 207286 233459
rect 207338 233447 207344 233459
rect 210754 233447 210782 233567
rect 218704 233555 218710 233567
rect 218762 233555 218768 233607
rect 283984 233555 283990 233607
rect 284042 233595 284048 233607
rect 311248 233595 311254 233607
rect 284042 233567 311254 233595
rect 284042 233555 284048 233567
rect 311248 233555 311254 233567
rect 311306 233555 311312 233607
rect 319504 233555 319510 233607
rect 319562 233595 319568 233607
rect 328144 233595 328150 233607
rect 319562 233567 328150 233595
rect 319562 233555 319568 233567
rect 328144 233555 328150 233567
rect 328202 233555 328208 233607
rect 335344 233555 335350 233607
rect 335402 233595 335408 233607
rect 463600 233595 463606 233607
rect 335402 233567 463606 233595
rect 335402 233555 335408 233567
rect 463600 233555 463606 233567
rect 463658 233555 463664 233607
rect 259888 233481 259894 233533
rect 259946 233521 259952 233533
rect 267760 233521 267766 233533
rect 259946 233493 267766 233521
rect 259946 233481 259952 233493
rect 267760 233481 267766 233493
rect 267818 233481 267824 233533
rect 287440 233481 287446 233533
rect 287498 233521 287504 233533
rect 311344 233521 311350 233533
rect 287498 233493 311350 233521
rect 287498 233481 287504 233493
rect 311344 233481 311350 233493
rect 311402 233481 311408 233533
rect 324784 233481 324790 233533
rect 324842 233521 324848 233533
rect 325936 233521 325942 233533
rect 324842 233493 325942 233521
rect 324842 233481 324848 233493
rect 325936 233481 325942 233493
rect 325994 233481 326000 233533
rect 326224 233481 326230 233533
rect 326282 233521 326288 233533
rect 460240 233521 460246 233533
rect 326282 233493 460246 233521
rect 326282 233481 326288 233493
rect 460240 233481 460246 233493
rect 460298 233481 460304 233533
rect 207338 233419 210782 233447
rect 207338 233407 207344 233419
rect 226672 233407 226678 233459
rect 226730 233447 226736 233459
rect 236752 233447 236758 233459
rect 226730 233419 236758 233447
rect 226730 233407 226736 233419
rect 236752 233407 236758 233419
rect 236810 233407 236816 233459
rect 264400 233407 264406 233459
rect 264458 233447 264464 233459
rect 272368 233447 272374 233459
rect 264458 233419 272374 233447
rect 264458 233407 264464 233419
rect 272368 233407 272374 233419
rect 272426 233407 272432 233459
rect 288400 233407 288406 233459
rect 288458 233447 288464 233459
rect 311056 233447 311062 233459
rect 288458 233419 311062 233447
rect 288458 233407 288464 233419
rect 311056 233407 311062 233419
rect 311114 233407 311120 233459
rect 317200 233407 317206 233459
rect 317258 233447 317264 233459
rect 412720 233447 412726 233459
rect 317258 233419 412726 233447
rect 317258 233407 317264 233419
rect 412720 233407 412726 233419
rect 412778 233407 412784 233459
rect 192400 233333 192406 233385
rect 192458 233373 192464 233385
rect 193744 233373 193750 233385
rect 192458 233345 193750 233373
rect 192458 233333 192464 233345
rect 193744 233333 193750 233345
rect 193802 233333 193808 233385
rect 193840 233333 193846 233385
rect 193898 233373 193904 233385
rect 196816 233373 196822 233385
rect 193898 233345 196822 233373
rect 193898 233333 193904 233345
rect 196816 233333 196822 233345
rect 196874 233333 196880 233385
rect 197968 233333 197974 233385
rect 198026 233373 198032 233385
rect 203632 233373 203638 233385
rect 198026 233345 203638 233373
rect 198026 233333 198032 233345
rect 203632 233333 203638 233345
rect 203690 233333 203696 233385
rect 203920 233333 203926 233385
rect 203978 233373 203984 233385
rect 214192 233373 214198 233385
rect 203978 233345 214198 233373
rect 203978 233333 203984 233345
rect 214192 233333 214198 233345
rect 214250 233333 214256 233385
rect 228400 233333 228406 233385
rect 228458 233373 228464 233385
rect 238960 233373 238966 233385
rect 228458 233345 238966 233373
rect 228458 233333 228464 233345
rect 238960 233333 238966 233345
rect 239018 233333 239024 233385
rect 257968 233333 257974 233385
rect 258026 233373 258032 233385
rect 269872 233373 269878 233385
rect 258026 233345 269878 233373
rect 258026 233333 258032 233345
rect 269872 233333 269878 233345
rect 269930 233333 269936 233385
rect 270544 233333 270550 233385
rect 270602 233373 270608 233385
rect 274672 233373 274678 233385
rect 270602 233345 274678 233373
rect 270602 233333 270608 233345
rect 274672 233333 274678 233345
rect 274730 233333 274736 233385
rect 282544 233333 282550 233385
rect 282602 233373 282608 233385
rect 299152 233373 299158 233385
rect 282602 233345 299158 233373
rect 282602 233333 282608 233345
rect 299152 233333 299158 233345
rect 299210 233333 299216 233385
rect 311152 233333 311158 233385
rect 311210 233373 311216 233385
rect 412048 233373 412054 233385
rect 311210 233345 412054 233373
rect 311210 233333 311216 233345
rect 412048 233333 412054 233345
rect 412106 233333 412112 233385
rect 193456 233259 193462 233311
rect 193514 233299 193520 233311
rect 194608 233299 194614 233311
rect 193514 233271 194614 233299
rect 193514 233259 193520 233271
rect 194608 233259 194614 233271
rect 194666 233259 194672 233311
rect 195184 233259 195190 233311
rect 195242 233299 195248 233311
rect 197488 233299 197494 233311
rect 195242 233271 197494 233299
rect 195242 233259 195248 233271
rect 197488 233259 197494 233271
rect 197546 233259 197552 233311
rect 197872 233259 197878 233311
rect 197930 233299 197936 233311
rect 202096 233299 202102 233311
rect 197930 233271 202102 233299
rect 197930 233259 197936 233271
rect 202096 233259 202102 233271
rect 202154 233259 202160 233311
rect 202384 233259 202390 233311
rect 202442 233299 202448 233311
rect 211120 233299 211126 233311
rect 202442 233271 211126 233299
rect 202442 233259 202448 233271
rect 211120 233259 211126 233271
rect 211178 233259 211184 233311
rect 242896 233259 242902 233311
rect 242954 233299 242960 233311
rect 259504 233299 259510 233311
rect 242954 233271 259510 233299
rect 242954 233259 242960 233271
rect 259504 233259 259510 233271
rect 259562 233259 259568 233311
rect 261616 233259 261622 233311
rect 261674 233299 261680 233311
rect 269584 233299 269590 233311
rect 261674 233271 269590 233299
rect 261674 233259 261680 233271
rect 269584 233259 269590 233271
rect 269642 233259 269648 233311
rect 270256 233259 270262 233311
rect 270314 233299 270320 233311
rect 273328 233299 273334 233311
rect 270314 233271 273334 233299
rect 270314 233259 270320 233271
rect 273328 233259 273334 233271
rect 273386 233259 273392 233311
rect 285328 233259 285334 233311
rect 285386 233299 285392 233311
rect 287440 233299 287446 233311
rect 285386 233271 287446 233299
rect 285386 233259 285392 233271
rect 287440 233259 287446 233271
rect 287498 233259 287504 233311
rect 288880 233259 288886 233311
rect 288938 233299 288944 233311
rect 346960 233299 346966 233311
rect 288938 233271 346966 233299
rect 288938 233259 288944 233271
rect 346960 233259 346966 233271
rect 347018 233259 347024 233311
rect 362512 233259 362518 233311
rect 362570 233299 362576 233311
rect 394768 233299 394774 233311
rect 362570 233271 394774 233299
rect 362570 233259 362576 233271
rect 394768 233259 394774 233271
rect 394826 233259 394832 233311
rect 400240 233259 400246 233311
rect 400298 233299 400304 233311
rect 479152 233299 479158 233311
rect 400298 233271 479158 233299
rect 400298 233259 400304 233271
rect 479152 233259 479158 233271
rect 479210 233259 479216 233311
rect 258736 233185 258742 233237
rect 258794 233225 258800 233237
rect 326608 233225 326614 233237
rect 258794 233197 326614 233225
rect 258794 233185 258800 233197
rect 326608 233185 326614 233197
rect 326666 233185 326672 233237
rect 340816 233185 340822 233237
rect 340874 233225 340880 233237
rect 491248 233225 491254 233237
rect 340874 233197 491254 233225
rect 340874 233185 340880 233197
rect 491248 233185 491254 233197
rect 491306 233185 491312 233237
rect 501040 233185 501046 233237
rect 501098 233225 501104 233237
rect 614992 233225 614998 233237
rect 501098 233197 614998 233225
rect 501098 233185 501104 233197
rect 614992 233185 614998 233197
rect 615050 233185 615056 233237
rect 262096 233111 262102 233163
rect 262154 233151 262160 233163
rect 334192 233151 334198 233163
rect 262154 233123 334198 233151
rect 262154 233111 262160 233123
rect 334192 233111 334198 233123
rect 334250 233111 334256 233163
rect 347056 233111 347062 233163
rect 347114 233151 347120 233163
rect 347114 233123 501086 233151
rect 347114 233111 347120 233123
rect 501058 233089 501086 233123
rect 260656 233037 260662 233089
rect 260714 233077 260720 233089
rect 331312 233077 331318 233089
rect 260714 233049 331318 233077
rect 260714 233037 260720 233049
rect 331312 233037 331318 233049
rect 331370 233037 331376 233089
rect 350320 233037 350326 233089
rect 350378 233077 350384 233089
rect 350378 233049 500990 233077
rect 350378 233037 350384 233049
rect 265744 232963 265750 233015
rect 265802 233003 265808 233015
rect 338032 233003 338038 233015
rect 265802 232975 338038 233003
rect 265802 232963 265808 232975
rect 338032 232963 338038 232975
rect 338090 232963 338096 233015
rect 353104 232963 353110 233015
rect 353162 233003 353168 233015
rect 500848 233003 500854 233015
rect 353162 232975 500854 233003
rect 353162 232963 353168 232975
rect 500848 232963 500854 232975
rect 500906 232963 500912 233015
rect 500962 233003 500990 233049
rect 501040 233037 501046 233089
rect 501098 233037 501104 233089
rect 507088 233003 507094 233015
rect 500962 232975 507094 233003
rect 507088 232963 507094 232975
rect 507146 232963 507152 233015
rect 289936 232889 289942 232941
rect 289994 232929 290000 232941
rect 382192 232929 382198 232941
rect 289994 232901 382198 232929
rect 289994 232889 290000 232901
rect 382192 232889 382198 232901
rect 382250 232889 382256 232941
rect 411760 232889 411766 232941
rect 411818 232929 411824 232941
rect 572080 232929 572086 232941
rect 411818 232901 572086 232929
rect 411818 232889 411824 232901
rect 572080 232889 572086 232901
rect 572138 232889 572144 232941
rect 263920 232815 263926 232867
rect 263978 232855 263984 232867
rect 337264 232855 337270 232867
rect 263978 232827 337270 232855
rect 263978 232815 263984 232827
rect 337264 232815 337270 232827
rect 337322 232815 337328 232867
rect 339184 232815 339190 232867
rect 339242 232855 339248 232867
rect 356080 232855 356086 232867
rect 339242 232827 356086 232855
rect 339242 232815 339248 232827
rect 356080 232815 356086 232827
rect 356138 232815 356144 232867
rect 356272 232815 356278 232867
rect 356330 232855 356336 232867
rect 519184 232855 519190 232867
rect 356330 232827 519190 232855
rect 356330 232815 356336 232827
rect 519184 232815 519190 232827
rect 519242 232815 519248 232867
rect 237616 232741 237622 232793
rect 237674 232781 237680 232793
rect 284368 232781 284374 232793
rect 237674 232753 284374 232781
rect 237674 232741 237680 232753
rect 284368 232741 284374 232753
rect 284426 232741 284432 232793
rect 295312 232741 295318 232793
rect 295370 232781 295376 232793
rect 397360 232781 397366 232793
rect 295370 232753 397366 232781
rect 295370 232741 295376 232753
rect 397360 232741 397366 232753
rect 397418 232741 397424 232793
rect 399568 232741 399574 232793
rect 399626 232781 399632 232793
rect 566704 232781 566710 232793
rect 399626 232753 566710 232781
rect 399626 232741 399632 232753
rect 566704 232741 566710 232753
rect 566762 232741 566768 232793
rect 216592 232667 216598 232719
rect 216650 232707 216656 232719
rect 242128 232707 242134 232719
rect 216650 232679 242134 232707
rect 216650 232667 216656 232679
rect 242128 232667 242134 232679
rect 242186 232667 242192 232719
rect 265168 232667 265174 232719
rect 265226 232707 265232 232719
rect 340240 232707 340246 232719
rect 265226 232679 340246 232707
rect 265226 232667 265232 232679
rect 340240 232667 340246 232679
rect 340298 232667 340304 232719
rect 362128 232667 362134 232719
rect 362186 232707 362192 232719
rect 531280 232707 531286 232719
rect 362186 232679 531286 232707
rect 362186 232667 362192 232679
rect 531280 232667 531286 232679
rect 531338 232667 531344 232719
rect 218032 232593 218038 232645
rect 218090 232633 218096 232645
rect 245104 232633 245110 232645
rect 218090 232605 245110 232633
rect 218090 232593 218096 232605
rect 245104 232593 245110 232605
rect 245162 232593 245168 232645
rect 268432 232593 268438 232645
rect 268490 232633 268496 232645
rect 346288 232633 346294 232645
rect 268490 232605 346294 232633
rect 268490 232593 268496 232605
rect 346288 232593 346294 232605
rect 346346 232593 346352 232645
rect 365392 232593 365398 232645
rect 365450 232633 365456 232645
rect 537232 232633 537238 232645
rect 365450 232605 537238 232633
rect 365450 232593 365456 232605
rect 537232 232593 537238 232605
rect 537290 232593 537296 232645
rect 219760 232519 219766 232571
rect 219818 232559 219824 232571
rect 248080 232559 248086 232571
rect 219818 232531 248086 232559
rect 219818 232519 219824 232531
rect 248080 232519 248086 232531
rect 248138 232519 248144 232571
rect 266608 232519 266614 232571
rect 266666 232559 266672 232571
rect 266666 232531 339422 232559
rect 266666 232519 266672 232531
rect 221104 232445 221110 232497
rect 221162 232485 221168 232497
rect 251152 232485 251158 232497
rect 221162 232457 251158 232485
rect 221162 232445 221168 232457
rect 251152 232445 251158 232457
rect 251210 232445 251216 232497
rect 271216 232445 271222 232497
rect 271274 232485 271280 232497
rect 339280 232485 339286 232497
rect 271274 232457 339286 232485
rect 271274 232445 271280 232457
rect 339280 232445 339286 232457
rect 339338 232445 339344 232497
rect 339394 232485 339422 232531
rect 339472 232519 339478 232571
rect 339530 232559 339536 232571
rect 361360 232559 361366 232571
rect 339530 232531 361366 232559
rect 339530 232519 339536 232531
rect 361360 232519 361366 232531
rect 361418 232519 361424 232571
rect 368176 232519 368182 232571
rect 368234 232559 368240 232571
rect 543376 232559 543382 232571
rect 368234 232531 543382 232559
rect 368234 232519 368240 232531
rect 543376 232519 543382 232531
rect 543434 232519 543440 232571
rect 343216 232485 343222 232497
rect 339394 232457 343222 232485
rect 343216 232445 343222 232457
rect 343274 232445 343280 232497
rect 344176 232445 344182 232497
rect 344234 232485 344240 232497
rect 355312 232485 355318 232497
rect 344234 232457 355318 232485
rect 344234 232445 344240 232457
rect 355312 232445 355318 232457
rect 355370 232445 355376 232497
rect 365008 232445 365014 232497
rect 365066 232485 365072 232497
rect 539536 232485 539542 232497
rect 365066 232457 539542 232485
rect 365066 232445 365072 232457
rect 539536 232445 539542 232457
rect 539594 232445 539600 232497
rect 222544 232371 222550 232423
rect 222602 232411 222608 232423
rect 254224 232411 254230 232423
rect 222602 232383 254230 232411
rect 222602 232371 222608 232383
rect 254224 232371 254230 232383
rect 254282 232371 254288 232423
rect 269680 232371 269686 232423
rect 269738 232411 269744 232423
rect 349360 232411 349366 232423
rect 269738 232383 349366 232411
rect 269738 232371 269744 232383
rect 349360 232371 349366 232383
rect 349418 232371 349424 232423
rect 366256 232371 366262 232423
rect 366314 232411 366320 232423
rect 542608 232411 542614 232423
rect 366314 232383 542614 232411
rect 366314 232371 366320 232383
rect 542608 232371 542614 232383
rect 542666 232371 542672 232423
rect 222928 232297 222934 232349
rect 222986 232337 222992 232349
rect 255664 232337 255670 232349
rect 222986 232309 255670 232337
rect 222986 232297 222992 232309
rect 255664 232297 255670 232309
rect 255722 232297 255728 232349
rect 274864 232297 274870 232349
rect 274922 232337 274928 232349
rect 339184 232337 339190 232349
rect 274922 232309 339190 232337
rect 274922 232297 274928 232309
rect 339184 232297 339190 232309
rect 339242 232297 339248 232349
rect 339280 232297 339286 232349
rect 339338 232337 339344 232349
rect 352336 232337 352342 232349
rect 339338 232309 352342 232337
rect 339338 232297 339344 232309
rect 352336 232297 352342 232309
rect 352394 232297 352400 232349
rect 371152 232297 371158 232349
rect 371210 232337 371216 232349
rect 549424 232337 549430 232349
rect 371210 232309 549430 232337
rect 371210 232297 371216 232309
rect 549424 232297 549430 232309
rect 549482 232297 549488 232349
rect 224272 232223 224278 232275
rect 224330 232263 224336 232275
rect 257200 232263 257206 232275
rect 224330 232235 257206 232263
rect 224330 232223 224336 232235
rect 257200 232223 257206 232235
rect 257258 232223 257264 232275
rect 272944 232223 272950 232275
rect 273002 232263 273008 232275
rect 344176 232263 344182 232275
rect 273002 232235 344182 232263
rect 273002 232223 273008 232235
rect 344176 232223 344182 232235
rect 344234 232223 344240 232275
rect 344272 232223 344278 232275
rect 344330 232263 344336 232275
rect 358480 232263 358486 232275
rect 344330 232235 358486 232263
rect 344330 232223 344336 232235
rect 358480 232223 358486 232235
rect 358538 232223 358544 232275
rect 369520 232223 369526 232275
rect 369578 232263 369584 232275
rect 548560 232263 548566 232275
rect 369578 232235 548566 232263
rect 369578 232223 369584 232235
rect 548560 232223 548566 232235
rect 548618 232223 548624 232275
rect 147856 232149 147862 232201
rect 147914 232189 147920 232201
rect 154096 232189 154102 232201
rect 147914 232161 154102 232189
rect 147914 232149 147920 232161
rect 154096 232149 154102 232161
rect 154154 232149 154160 232201
rect 226288 232149 226294 232201
rect 226346 232189 226352 232201
rect 261712 232189 261718 232201
rect 226346 232161 261718 232189
rect 226346 232149 226352 232161
rect 261712 232149 261718 232161
rect 261770 232149 261776 232201
rect 274192 232149 274198 232201
rect 274250 232189 274256 232201
rect 274250 232161 347006 232189
rect 274250 232149 274256 232161
rect 227056 232075 227062 232127
rect 227114 232115 227120 232127
rect 263248 232115 263254 232127
rect 227114 232087 263254 232115
rect 227114 232075 227120 232087
rect 263248 232075 263254 232087
rect 263306 232075 263312 232127
rect 275728 232075 275734 232127
rect 275786 232115 275792 232127
rect 339472 232115 339478 232127
rect 275786 232087 339478 232115
rect 275786 232075 275792 232087
rect 339472 232075 339478 232087
rect 339530 232075 339536 232127
rect 346978 232115 347006 232161
rect 356464 232149 356470 232201
rect 356522 232189 356528 232201
rect 365200 232189 365206 232201
rect 356522 232161 365206 232189
rect 356522 232149 356528 232161
rect 365200 232149 365206 232161
rect 365258 232149 365264 232201
rect 368080 232149 368086 232201
rect 368138 232189 368144 232201
rect 545584 232189 545590 232201
rect 368138 232161 545590 232189
rect 368138 232149 368144 232161
rect 545584 232149 545590 232161
rect 545642 232149 545648 232201
rect 358192 232115 358198 232127
rect 346978 232087 358198 232115
rect 358192 232075 358198 232087
rect 358250 232075 358256 232127
rect 358576 232075 358582 232127
rect 358634 232115 358640 232127
rect 362224 232115 362230 232127
rect 358634 232087 362230 232115
rect 358634 232075 358640 232087
rect 362224 232075 362230 232087
rect 362282 232075 362288 232127
rect 370384 232115 370390 232127
rect 364546 232087 370390 232115
rect 233872 232001 233878 232053
rect 233930 232041 233936 232053
rect 274480 232041 274486 232053
rect 233930 232013 274486 232041
rect 233930 232001 233936 232013
rect 274480 232001 274486 232013
rect 274538 232001 274544 232053
rect 277456 232001 277462 232053
rect 277514 232041 277520 232053
rect 364432 232041 364438 232053
rect 277514 232013 364438 232041
rect 277514 232001 277520 232013
rect 364432 232001 364438 232013
rect 364490 232001 364496 232053
rect 233200 231927 233206 231979
rect 233258 231967 233264 231979
rect 275344 231967 275350 231979
rect 233258 231939 275350 231967
rect 233258 231927 233264 231939
rect 275344 231927 275350 231939
rect 275402 231927 275408 231979
rect 280240 231927 280246 231979
rect 280298 231967 280304 231979
rect 364546 231967 364574 232087
rect 370384 232075 370390 232087
rect 370442 232075 370448 232127
rect 372688 232075 372694 232127
rect 372746 232115 372752 232127
rect 552400 232115 552406 232127
rect 372746 232087 552406 232115
rect 372746 232075 372752 232087
rect 552400 232075 552406 232087
rect 552458 232075 552464 232127
rect 373456 232041 373462 232053
rect 280298 231939 364574 231967
rect 367618 232013 373462 232041
rect 280298 231927 280304 231939
rect 234832 231853 234838 231905
rect 234890 231893 234896 231905
rect 278320 231893 278326 231905
rect 234890 231865 278326 231893
rect 234890 231853 234896 231865
rect 278320 231853 278326 231865
rect 278378 231853 278384 231905
rect 278992 231853 278998 231905
rect 279050 231893 279056 231905
rect 367408 231893 367414 231905
rect 279050 231865 367414 231893
rect 279050 231853 279056 231865
rect 367408 231853 367414 231865
rect 367466 231853 367472 231905
rect 236080 231779 236086 231831
rect 236138 231819 236144 231831
rect 281296 231819 281302 231831
rect 236138 231791 281302 231819
rect 236138 231779 236144 231791
rect 281296 231779 281302 231791
rect 281354 231779 281360 231831
rect 281968 231779 281974 231831
rect 282026 231819 282032 231831
rect 367618 231819 367646 232013
rect 373456 232001 373462 232013
rect 373514 232001 373520 232053
rect 554704 232041 554710 232053
rect 375682 232013 554710 232041
rect 372304 231927 372310 231979
rect 372362 231967 372368 231979
rect 375682 231967 375710 232013
rect 554704 232001 554710 232013
rect 554762 232001 554768 232053
rect 372362 231939 375710 231967
rect 372362 231927 372368 231939
rect 375760 231927 375766 231979
rect 375818 231967 375824 231979
rect 558448 231967 558454 231979
rect 375818 231939 558454 231967
rect 375818 231927 375824 231939
rect 558448 231927 558454 231939
rect 558506 231927 558512 231979
rect 374512 231853 374518 231905
rect 374570 231893 374576 231905
rect 557008 231893 557014 231905
rect 374570 231865 557014 231893
rect 374570 231853 374576 231865
rect 557008 231853 557014 231865
rect 557066 231853 557072 231905
rect 282026 231791 367646 231819
rect 282026 231779 282032 231791
rect 374032 231779 374038 231831
rect 374090 231819 374096 231831
rect 557680 231819 557686 231831
rect 374090 231791 557686 231819
rect 374090 231779 374096 231791
rect 557680 231779 557686 231791
rect 557738 231779 557744 231831
rect 259120 231705 259126 231757
rect 259178 231745 259184 231757
rect 328048 231745 328054 231757
rect 259178 231717 328054 231745
rect 259178 231705 259184 231717
rect 328048 231705 328054 231717
rect 328106 231705 328112 231757
rect 358480 231705 358486 231757
rect 358538 231745 358544 231757
rect 495088 231745 495094 231757
rect 358538 231717 495094 231745
rect 358538 231705 358544 231717
rect 495088 231705 495094 231717
rect 495146 231705 495152 231757
rect 500848 231705 500854 231757
rect 500906 231745 500912 231757
rect 513136 231745 513142 231757
rect 500906 231717 513142 231745
rect 500906 231705 500912 231717
rect 513136 231705 513142 231717
rect 513194 231705 513200 231757
rect 257584 231631 257590 231683
rect 257642 231671 257648 231683
rect 325168 231671 325174 231683
rect 257642 231643 325174 231671
rect 257642 231631 257648 231643
rect 325168 231631 325174 231643
rect 325226 231631 325232 231683
rect 337552 231631 337558 231683
rect 337610 231671 337616 231683
rect 485200 231671 485206 231683
rect 337610 231643 485206 231671
rect 337610 231631 337616 231643
rect 485200 231631 485206 231643
rect 485258 231631 485264 231683
rect 256144 231557 256150 231609
rect 256202 231597 256208 231609
rect 322096 231597 322102 231609
rect 256202 231569 322102 231597
rect 256202 231557 256208 231569
rect 322096 231557 322102 231569
rect 322154 231557 322160 231609
rect 328144 231557 328150 231609
rect 328202 231597 328208 231609
rect 448912 231597 448918 231609
rect 328202 231569 448918 231597
rect 328202 231557 328208 231569
rect 448912 231557 448918 231569
rect 448970 231557 448976 231609
rect 248368 231483 248374 231535
rect 248426 231523 248432 231535
rect 305488 231523 305494 231535
rect 248426 231495 305494 231523
rect 248426 231483 248432 231495
rect 305488 231483 305494 231495
rect 305546 231483 305552 231535
rect 312208 231483 312214 231535
rect 312266 231523 312272 231535
rect 433840 231523 433846 231535
rect 312266 231495 433846 231523
rect 312266 231483 312272 231495
rect 433840 231483 433846 231495
rect 433898 231483 433904 231535
rect 281200 231409 281206 231461
rect 281258 231449 281264 231461
rect 289648 231449 289654 231461
rect 281258 231421 289654 231449
rect 281258 231409 281264 231421
rect 289648 231409 289654 231421
rect 289706 231409 289712 231461
rect 292528 231409 292534 231461
rect 292586 231449 292592 231461
rect 379984 231449 379990 231461
rect 292586 231421 379990 231449
rect 292586 231409 292592 231421
rect 379984 231409 379990 231421
rect 380042 231409 380048 231461
rect 402544 231409 402550 231461
rect 402602 231449 402608 231461
rect 520720 231449 520726 231461
rect 402602 231421 520726 231449
rect 402602 231409 402608 231421
rect 520720 231409 520726 231421
rect 520778 231409 520784 231461
rect 290800 231335 290806 231387
rect 290858 231375 290864 231387
rect 374608 231375 374614 231387
rect 290858 231347 374614 231375
rect 290858 231335 290864 231347
rect 374608 231335 374614 231347
rect 374666 231335 374672 231387
rect 400144 231335 400150 231387
rect 400202 231375 400208 231387
rect 499600 231375 499606 231387
rect 400202 231347 499606 231375
rect 400202 231335 400208 231347
rect 499600 231335 499606 231347
rect 499658 231335 499664 231387
rect 293104 231261 293110 231313
rect 293162 231301 293168 231313
rect 372784 231301 372790 231313
rect 293162 231273 372790 231301
rect 293162 231261 293168 231273
rect 372784 231261 372790 231273
rect 372842 231261 372848 231313
rect 394576 231261 394582 231313
rect 394634 231301 394640 231313
rect 485968 231301 485974 231313
rect 394634 231273 485974 231301
rect 394634 231261 394640 231273
rect 485968 231261 485974 231273
rect 486026 231261 486032 231313
rect 255760 231187 255766 231239
rect 255818 231227 255824 231239
rect 320656 231227 320662 231239
rect 255818 231199 320662 231227
rect 255818 231187 255824 231199
rect 320656 231187 320662 231199
rect 320714 231187 320720 231239
rect 334096 231187 334102 231239
rect 334154 231227 334160 231239
rect 415696 231227 415702 231239
rect 334154 231199 415702 231227
rect 334154 231187 334160 231199
rect 415696 231187 415702 231199
rect 415754 231187 415760 231239
rect 293488 231113 293494 231165
rect 293546 231153 293552 231165
rect 364048 231153 364054 231165
rect 293546 231125 364054 231153
rect 293546 231113 293552 231125
rect 364048 231113 364054 231125
rect 364106 231113 364112 231165
rect 394672 231113 394678 231165
rect 394730 231153 394736 231165
rect 473872 231153 473878 231165
rect 394730 231125 473878 231153
rect 394730 231113 394736 231125
rect 473872 231113 473878 231125
rect 473930 231113 473936 231165
rect 252976 231039 252982 231091
rect 253034 231079 253040 231091
rect 314512 231079 314518 231091
rect 253034 231051 314518 231079
rect 253034 231039 253040 231051
rect 314512 231039 314518 231051
rect 314570 231039 314576 231091
rect 345520 231039 345526 231091
rect 345578 231079 345584 231091
rect 419248 231079 419254 231091
rect 345578 231051 419254 231079
rect 345578 231039 345584 231051
rect 419248 231039 419254 231051
rect 419306 231039 419312 231091
rect 245200 230965 245206 231017
rect 245258 231005 245264 231017
rect 299440 231005 299446 231017
rect 245258 230977 299446 231005
rect 245258 230965 245264 230977
rect 299440 230965 299446 230977
rect 299498 230965 299504 231017
rect 308176 230965 308182 231017
rect 308234 231005 308240 231017
rect 323632 231005 323638 231017
rect 308234 230977 323638 231005
rect 308234 230965 308240 230977
rect 323632 230965 323638 230977
rect 323690 230965 323696 231017
rect 328336 230965 328342 231017
rect 328394 231005 328400 231017
rect 401392 231005 401398 231017
rect 328394 230977 401398 231005
rect 328394 230965 328400 230977
rect 401392 230965 401398 230977
rect 401450 230965 401456 231017
rect 411568 230965 411574 231017
rect 411626 231005 411632 231017
rect 424048 231005 424054 231017
rect 411626 230977 424054 231005
rect 411626 230965 411632 230977
rect 424048 230965 424054 230977
rect 424106 230965 424112 231017
rect 325264 230891 325270 230943
rect 325322 230931 325328 230943
rect 329584 230931 329590 230943
rect 325322 230903 329590 230931
rect 325322 230891 325328 230903
rect 329584 230891 329590 230903
rect 329642 230891 329648 230943
rect 331216 230891 331222 230943
rect 331274 230931 331280 230943
rect 395344 230931 395350 230943
rect 331274 230903 395350 230931
rect 331274 230891 331280 230903
rect 395344 230891 395350 230903
rect 395402 230891 395408 230943
rect 326704 230817 326710 230869
rect 326762 230857 326768 230869
rect 352720 230857 352726 230869
rect 326762 230829 352726 230857
rect 326762 230817 326768 230829
rect 352720 230817 352726 230829
rect 352778 230817 352784 230869
rect 358768 230817 358774 230869
rect 358826 230857 358832 230869
rect 377104 230857 377110 230869
rect 358826 230829 377110 230857
rect 358826 230817 358832 230829
rect 377104 230817 377110 230829
rect 377162 230817 377168 230869
rect 385936 230817 385942 230869
rect 385994 230857 386000 230869
rect 449680 230857 449686 230869
rect 385994 230829 449686 230857
rect 385994 230817 386000 230829
rect 449680 230817 449686 230829
rect 449738 230817 449744 230869
rect 319600 230743 319606 230795
rect 319658 230783 319664 230795
rect 358576 230783 358582 230795
rect 319658 230755 358582 230783
rect 319658 230743 319664 230755
rect 358576 230743 358582 230755
rect 358634 230743 358640 230795
rect 358864 230743 358870 230795
rect 358922 230783 358928 230795
rect 365104 230783 365110 230795
rect 358922 230755 365110 230783
rect 358922 230743 358928 230755
rect 365104 230743 365110 230755
rect 365162 230743 365168 230795
rect 365200 230743 365206 230795
rect 365258 230783 365264 230795
rect 409648 230783 409654 230795
rect 365258 230755 409654 230783
rect 365258 230743 365264 230755
rect 409648 230743 409654 230755
rect 409706 230743 409712 230795
rect 320848 230669 320854 230721
rect 320906 230709 320912 230721
rect 320906 230681 358526 230709
rect 320906 230669 320912 230681
rect 290608 230595 290614 230647
rect 290666 230635 290672 230647
rect 297328 230635 297334 230647
rect 290666 230607 297334 230635
rect 290666 230595 290672 230607
rect 297328 230595 297334 230607
rect 297386 230595 297392 230647
rect 302320 230595 302326 230647
rect 302378 230635 302384 230647
rect 308560 230635 308566 230647
rect 302378 230607 308566 230635
rect 302378 230595 302384 230607
rect 308560 230595 308566 230607
rect 308618 230595 308624 230647
rect 313936 230595 313942 230647
rect 313994 230635 314000 230647
rect 358384 230635 358390 230647
rect 313994 230607 358390 230635
rect 313994 230595 314000 230607
rect 358384 230595 358390 230607
rect 358442 230595 358448 230647
rect 306640 230521 306646 230573
rect 306698 230561 306704 230573
rect 317584 230561 317590 230573
rect 306698 230533 317590 230561
rect 306698 230521 306704 230533
rect 317584 230521 317590 230533
rect 317642 230521 317648 230573
rect 323824 230521 323830 230573
rect 323882 230561 323888 230573
rect 358498 230561 358526 230681
rect 359056 230669 359062 230721
rect 359114 230709 359120 230721
rect 380272 230709 380278 230721
rect 359114 230681 380278 230709
rect 359114 230669 359120 230681
rect 380272 230669 380278 230681
rect 380330 230669 380336 230721
rect 358576 230595 358582 230647
rect 358634 230635 358640 230647
rect 362128 230635 362134 230647
rect 358634 230607 362134 230635
rect 358634 230595 358640 230607
rect 362128 230595 362134 230607
rect 362186 230595 362192 230647
rect 362224 230595 362230 230647
rect 362282 230635 362288 230647
rect 410512 230635 410518 230647
rect 362282 230607 410518 230635
rect 362282 230595 362288 230607
rect 410512 230595 410518 230607
rect 410570 230595 410576 230647
rect 374224 230561 374230 230573
rect 323882 230533 358430 230561
rect 358498 230533 374230 230561
rect 323882 230521 323888 230533
rect 149392 230447 149398 230499
rect 149450 230487 149456 230499
rect 156976 230487 156982 230499
rect 149450 230459 156982 230487
rect 149450 230447 149456 230459
rect 156976 230447 156982 230459
rect 157034 230447 157040 230499
rect 299248 230447 299254 230499
rect 299306 230487 299312 230499
rect 302512 230487 302518 230499
rect 299306 230459 302518 230487
rect 299306 230447 299312 230459
rect 302512 230447 302518 230459
rect 302570 230447 302576 230499
rect 304144 230447 304150 230499
rect 304202 230487 304208 230499
rect 311632 230487 311638 230499
rect 304202 230459 311638 230487
rect 304202 230447 304208 230459
rect 311632 230447 311638 230459
rect 311690 230447 311696 230499
rect 322000 230447 322006 230499
rect 322058 230487 322064 230499
rect 358288 230487 358294 230499
rect 322058 230459 358294 230487
rect 322058 230447 322064 230459
rect 358288 230447 358294 230459
rect 358346 230447 358352 230499
rect 358402 230487 358430 230533
rect 374224 230521 374230 230533
rect 374282 230521 374288 230573
rect 358672 230487 358678 230499
rect 358402 230459 358678 230487
rect 358672 230447 358678 230459
rect 358730 230447 358736 230499
rect 358768 230447 358774 230499
rect 358826 230487 358832 230499
rect 368176 230487 368182 230499
rect 358826 230459 368182 230487
rect 358826 230447 358832 230459
rect 368176 230447 368182 230459
rect 368234 230447 368240 230499
rect 423376 230447 423382 230499
rect 423434 230487 423440 230499
rect 436144 230487 436150 230499
rect 423434 230459 436150 230487
rect 423434 230447 423440 230459
rect 436144 230447 436150 230459
rect 436202 230447 436208 230499
rect 241072 230373 241078 230425
rect 241130 230413 241136 230425
rect 291952 230413 291958 230425
rect 241130 230385 291958 230413
rect 241130 230373 241136 230385
rect 291952 230373 291958 230385
rect 292010 230373 292016 230425
rect 314896 230373 314902 230425
rect 314954 230413 314960 230425
rect 439984 230413 439990 230425
rect 314954 230385 439990 230413
rect 314954 230373 314960 230385
rect 439984 230373 439990 230385
rect 440042 230373 440048 230425
rect 245776 230299 245782 230351
rect 245834 230339 245840 230351
rect 300976 230339 300982 230351
rect 245834 230311 300982 230339
rect 245834 230299 245840 230311
rect 300976 230299 300982 230311
rect 301034 230299 301040 230351
rect 321232 230299 321238 230351
rect 321290 230339 321296 230351
rect 321290 230311 329150 230339
rect 321290 230299 321296 230311
rect 248944 230225 248950 230277
rect 249002 230265 249008 230277
rect 304816 230265 304822 230277
rect 249002 230237 304822 230265
rect 249002 230225 249008 230237
rect 304816 230225 304822 230237
rect 304874 230225 304880 230277
rect 305008 230225 305014 230277
rect 305066 230265 305072 230277
rect 326800 230265 326806 230277
rect 305066 230237 326806 230265
rect 305066 230225 305072 230237
rect 326800 230225 326806 230237
rect 326858 230225 326864 230277
rect 329122 230265 329150 230311
rect 329200 230299 329206 230351
rect 329258 230339 329264 230351
rect 445936 230339 445942 230351
rect 329258 230311 445942 230339
rect 329258 230299 329264 230311
rect 445936 230299 445942 230311
rect 445994 230299 446000 230351
rect 449296 230299 449302 230351
rect 449354 230339 449360 230351
rect 466384 230339 466390 230351
rect 449354 230311 466390 230339
rect 449354 230299 449360 230311
rect 466384 230299 466390 230311
rect 466442 230299 466448 230351
rect 451984 230265 451990 230277
rect 329122 230237 451990 230265
rect 451984 230225 451990 230237
rect 452042 230225 452048 230277
rect 228880 230151 228886 230203
rect 228938 230191 228944 230203
rect 267856 230191 267862 230203
rect 228938 230163 267862 230191
rect 228938 230151 228944 230163
rect 267856 230151 267862 230163
rect 267914 230151 267920 230203
rect 269872 230151 269878 230203
rect 269930 230191 269936 230203
rect 322960 230191 322966 230203
rect 269930 230163 322966 230191
rect 269930 230151 269936 230163
rect 322960 230151 322966 230163
rect 323018 230151 323024 230203
rect 325744 230151 325750 230203
rect 325802 230191 325808 230203
rect 461008 230191 461014 230203
rect 325802 230163 461014 230191
rect 325802 230151 325808 230163
rect 461008 230151 461014 230163
rect 461066 230151 461072 230203
rect 463600 230151 463606 230203
rect 463658 230191 463664 230203
rect 478288 230191 478294 230203
rect 463658 230163 478294 230191
rect 463658 230151 463664 230163
rect 478288 230151 478294 230163
rect 478346 230151 478352 230203
rect 248752 230077 248758 230129
rect 248810 230117 248816 230129
rect 307024 230117 307030 230129
rect 248810 230089 307030 230117
rect 248810 230077 248816 230089
rect 307024 230077 307030 230089
rect 307082 230077 307088 230129
rect 324016 230077 324022 230129
rect 324074 230117 324080 230129
rect 458032 230117 458038 230129
rect 324074 230089 458038 230117
rect 324074 230077 324080 230089
rect 458032 230077 458038 230089
rect 458090 230077 458096 230129
rect 466480 230077 466486 230129
rect 466538 230117 466544 230129
rect 484432 230117 484438 230129
rect 466538 230089 484438 230117
rect 466538 230077 466544 230089
rect 484432 230077 484438 230089
rect 484490 230077 484496 230129
rect 227440 230003 227446 230055
rect 227498 230043 227504 230055
rect 264784 230043 264790 230055
rect 227498 230015 264790 230043
rect 227498 230003 227504 230015
rect 264784 230003 264790 230015
rect 264842 230003 264848 230055
rect 290896 230003 290902 230055
rect 290954 230043 290960 230055
rect 331888 230043 331894 230055
rect 290954 230015 331894 230043
rect 290954 230003 290960 230015
rect 331888 230003 331894 230015
rect 331946 230003 331952 230055
rect 475216 230003 475222 230055
rect 475274 230043 475280 230055
rect 601456 230043 601462 230055
rect 475274 230015 601462 230043
rect 475274 230003 475280 230015
rect 601456 230003 601462 230015
rect 601514 230003 601520 230055
rect 251920 229929 251926 229981
rect 251978 229969 251984 229981
rect 310768 229969 310774 229981
rect 251978 229941 310774 229969
rect 251978 229929 251984 229941
rect 310768 229929 310774 229941
rect 310826 229929 310832 229981
rect 317968 229929 317974 229981
rect 318026 229969 318032 229981
rect 329200 229969 329206 229981
rect 318026 229941 329206 229969
rect 318026 229929 318032 229941
rect 329200 229929 329206 229941
rect 329258 229929 329264 229981
rect 331600 229929 331606 229981
rect 331658 229969 331664 229981
rect 473104 229969 473110 229981
rect 331658 229941 473110 229969
rect 331658 229929 331664 229941
rect 473104 229929 473110 229941
rect 473162 229929 473168 229981
rect 479152 229929 479158 229981
rect 479210 229969 479216 229981
rect 609040 229969 609046 229981
rect 479210 229941 609046 229969
rect 479210 229929 479216 229941
rect 609040 229929 609046 229941
rect 609098 229929 609104 229981
rect 250288 229855 250294 229907
rect 250346 229895 250352 229907
rect 310000 229895 310006 229907
rect 250346 229867 310006 229895
rect 250346 229855 250352 229867
rect 310000 229855 310006 229867
rect 310058 229855 310064 229907
rect 336304 229855 336310 229907
rect 336362 229895 336368 229907
rect 482128 229895 482134 229907
rect 336362 229867 482134 229895
rect 336362 229855 336368 229867
rect 482128 229855 482134 229867
rect 482186 229855 482192 229907
rect 484624 229855 484630 229907
rect 484682 229895 484688 229907
rect 612112 229895 612118 229907
rect 484682 229867 612118 229895
rect 484682 229855 484688 229867
rect 612112 229855 612118 229867
rect 612170 229855 612176 229907
rect 146896 229781 146902 229833
rect 146954 229821 146960 229833
rect 151216 229821 151222 229833
rect 146954 229793 151222 229821
rect 146954 229781 146960 229793
rect 151216 229781 151222 229793
rect 151274 229781 151280 229833
rect 251536 229781 251542 229833
rect 251594 229821 251600 229833
rect 313072 229821 313078 229833
rect 251594 229793 313078 229821
rect 251594 229781 251600 229793
rect 313072 229781 313078 229793
rect 313130 229781 313136 229833
rect 328528 229781 328534 229833
rect 328586 229821 328592 229833
rect 331120 229821 331126 229833
rect 328586 229793 331126 229821
rect 328586 229781 328592 229793
rect 331120 229781 331126 229793
rect 331178 229781 331184 229833
rect 348496 229781 348502 229833
rect 348554 229821 348560 229833
rect 504016 229821 504022 229833
rect 348554 229793 504022 229821
rect 348554 229781 348560 229793
rect 504016 229781 504022 229793
rect 504074 229781 504080 229833
rect 506800 229781 506806 229833
rect 506858 229821 506864 229833
rect 622672 229821 622678 229833
rect 506858 229793 622678 229821
rect 506858 229781 506864 229793
rect 622672 229781 622678 229793
rect 622730 229781 622736 229833
rect 244240 229707 244246 229759
rect 244298 229747 244304 229759
rect 298000 229747 298006 229759
rect 244298 229719 298006 229747
rect 244298 229707 244304 229719
rect 298000 229707 298006 229719
rect 298058 229707 298064 229759
rect 298576 229707 298582 229759
rect 298634 229747 298640 229759
rect 406768 229747 406774 229759
rect 298634 229719 406774 229747
rect 298634 229707 298640 229719
rect 406768 229707 406774 229719
rect 406826 229707 406832 229759
rect 411472 229707 411478 229759
rect 411530 229747 411536 229759
rect 565936 229747 565942 229759
rect 411530 229719 565942 229747
rect 411530 229707 411536 229719
rect 565936 229707 565942 229719
rect 565994 229707 566000 229759
rect 215248 229633 215254 229685
rect 215306 229673 215312 229685
rect 239056 229673 239062 229685
rect 215306 229645 239062 229673
rect 215306 229633 215312 229645
rect 239056 229633 239062 229645
rect 239114 229633 239120 229685
rect 253072 229633 253078 229685
rect 253130 229673 253136 229685
rect 316144 229673 316150 229685
rect 253130 229645 316150 229673
rect 253130 229633 253136 229645
rect 316144 229633 316150 229645
rect 316202 229633 316208 229685
rect 351760 229633 351766 229685
rect 351818 229673 351824 229685
rect 510160 229673 510166 229685
rect 351818 229645 510166 229673
rect 351818 229633 351824 229645
rect 510160 229633 510166 229645
rect 510218 229633 510224 229685
rect 220144 229559 220150 229611
rect 220202 229599 220208 229611
rect 249712 229599 249718 229611
rect 220202 229571 249718 229599
rect 220202 229559 220208 229571
rect 249712 229559 249718 229571
rect 249770 229559 249776 229611
rect 255184 229559 255190 229611
rect 255242 229599 255248 229611
rect 316816 229599 316822 229611
rect 255242 229571 316822 229599
rect 255242 229559 255248 229571
rect 316816 229559 316822 229571
rect 316874 229559 316880 229611
rect 354832 229559 354838 229611
rect 354890 229599 354896 229611
rect 516112 229599 516118 229611
rect 354890 229571 516118 229599
rect 354890 229559 354896 229571
rect 516112 229559 516118 229571
rect 516170 229559 516176 229611
rect 221584 229485 221590 229537
rect 221642 229525 221648 229537
rect 252592 229525 252598 229537
rect 221642 229497 252598 229525
rect 221642 229485 221648 229497
rect 252592 229485 252598 229497
rect 252650 229485 252656 229537
rect 254800 229485 254806 229537
rect 254858 229525 254864 229537
rect 319120 229525 319126 229537
rect 254858 229497 319126 229525
rect 254858 229485 254864 229497
rect 319120 229485 319126 229497
rect 319178 229485 319184 229537
rect 357616 229485 357622 229537
rect 357674 229525 357680 229537
rect 522160 229525 522166 229537
rect 357674 229497 522166 229525
rect 357674 229485 357680 229497
rect 522160 229485 522166 229497
rect 522218 229485 522224 229537
rect 264304 229411 264310 229463
rect 264362 229451 264368 229463
rect 334960 229451 334966 229463
rect 264362 229423 334966 229451
rect 264362 229411 264368 229423
rect 334960 229411 334966 229423
rect 335018 229411 335024 229463
rect 366640 229411 366646 229463
rect 366698 229451 366704 229463
rect 366698 229423 368654 229451
rect 366698 229411 366704 229423
rect 230608 229337 230614 229389
rect 230666 229377 230672 229389
rect 270736 229377 270742 229389
rect 230666 229349 270742 229377
rect 230666 229337 230672 229349
rect 270736 229337 270742 229349
rect 270794 229337 270800 229389
rect 273328 229337 273334 229389
rect 273386 229377 273392 229389
rect 347056 229377 347062 229389
rect 273386 229349 347062 229377
rect 273386 229337 273392 229349
rect 347056 229337 347062 229349
rect 347114 229337 347120 229389
rect 367024 229377 367030 229389
rect 348466 229349 367030 229377
rect 230320 229263 230326 229315
rect 230378 229303 230384 229315
rect 269296 229303 269302 229315
rect 230378 229275 269302 229303
rect 230378 229263 230384 229275
rect 269296 229263 269302 229275
rect 269354 229263 269360 229315
rect 283504 229263 283510 229315
rect 283562 229303 283568 229315
rect 348466 229303 348494 229349
rect 367024 229337 367030 229349
rect 367082 229337 367088 229389
rect 368626 229377 368654 229423
rect 369904 229411 369910 229463
rect 369962 229451 369968 229463
rect 371440 229451 371446 229463
rect 369962 229423 371446 229451
rect 369962 229411 369968 229423
rect 371440 229411 371446 229423
rect 371498 229411 371504 229463
rect 377200 229411 377206 229463
rect 377258 229451 377264 229463
rect 538864 229451 538870 229463
rect 377258 229423 538870 229451
rect 377258 229411 377264 229423
rect 538864 229411 538870 229423
rect 538922 229411 538928 229463
rect 540304 229377 540310 229389
rect 368626 229349 540310 229377
rect 540304 229337 540310 229349
rect 540362 229337 540368 229389
rect 371248 229303 371254 229315
rect 283562 229275 348494 229303
rect 354370 229275 371254 229303
rect 283562 229263 283568 229275
rect 233488 229189 233494 229241
rect 233546 229229 233552 229241
rect 276784 229229 276790 229241
rect 233546 229201 276790 229229
rect 233546 229189 233552 229201
rect 276784 229189 276790 229201
rect 276842 229189 276848 229241
rect 282160 229189 282166 229241
rect 282218 229229 282224 229241
rect 354370 229229 354398 229275
rect 371248 229263 371254 229275
rect 371306 229263 371312 229315
rect 371440 229263 371446 229315
rect 371498 229303 371504 229315
rect 546352 229303 546358 229315
rect 371498 229275 546358 229303
rect 371498 229263 371504 229275
rect 546352 229263 546358 229275
rect 546410 229263 546416 229315
rect 371536 229229 371542 229241
rect 282218 229201 354398 229229
rect 354466 229201 371542 229229
rect 282218 229189 282224 229201
rect 231952 229115 231958 229167
rect 232010 229155 232016 229167
rect 273808 229155 273814 229167
rect 232010 229127 273814 229155
rect 232010 229115 232016 229127
rect 273808 229115 273814 229127
rect 273866 229115 273872 229167
rect 284752 229115 284758 229167
rect 284810 229155 284816 229167
rect 354466 229155 354494 229201
rect 371536 229189 371542 229201
rect 371594 229189 371600 229241
rect 374320 229189 374326 229241
rect 374378 229229 374384 229241
rect 555376 229229 555382 229241
rect 374378 229201 555382 229229
rect 374378 229189 374384 229201
rect 555376 229189 555382 229201
rect 555434 229189 555440 229241
rect 374512 229155 374518 229167
rect 284810 229127 354494 229155
rect 358498 229127 374518 229155
rect 284810 229115 284816 229127
rect 235216 229041 235222 229093
rect 235274 229081 235280 229093
rect 279856 229081 279862 229093
rect 235274 229053 279862 229081
rect 235274 229041 235280 229053
rect 279856 229041 279862 229053
rect 279914 229041 279920 229093
rect 286288 229041 286294 229093
rect 286346 229081 286352 229093
rect 358498 229081 358526 229127
rect 374512 229115 374518 229127
rect 374570 229115 374576 229167
rect 377008 229115 377014 229167
rect 377066 229155 377072 229167
rect 561424 229155 561430 229167
rect 377066 229127 561430 229155
rect 377066 229115 377072 229127
rect 561424 229115 561430 229127
rect 561482 229115 561488 229167
rect 286346 229053 358526 229081
rect 286346 229041 286352 229053
rect 380464 229041 380470 229093
rect 380522 229081 380528 229093
rect 567472 229081 567478 229093
rect 380522 229053 567478 229081
rect 380522 229041 380528 229053
rect 567472 229041 567478 229053
rect 567530 229041 567536 229093
rect 238384 228967 238390 229019
rect 238442 229007 238448 229019
rect 283600 229007 283606 229019
rect 238442 228979 283606 229007
rect 238442 228967 238448 228979
rect 283600 228967 283606 228979
rect 283658 228967 283664 229019
rect 287920 228967 287926 229019
rect 287978 229007 287984 229019
rect 374416 229007 374422 229019
rect 287978 228979 374422 229007
rect 287978 228967 287984 228979
rect 374416 228967 374422 228979
rect 374474 228967 374480 229019
rect 379888 228967 379894 229019
rect 379946 229007 379952 229019
rect 569776 229007 569782 229019
rect 379946 228979 569782 229007
rect 379946 228967 379952 228979
rect 569776 228967 569782 228979
rect 569834 228967 569840 229019
rect 246160 228893 246166 228945
rect 246218 228933 246224 228945
rect 298672 228933 298678 228945
rect 246218 228905 298678 228933
rect 246218 228893 246224 228905
rect 298672 228893 298678 228905
rect 298730 228893 298736 228945
rect 308944 228893 308950 228945
rect 309002 228933 309008 228945
rect 427792 228933 427798 228945
rect 309002 228905 427798 228933
rect 309002 228893 309008 228905
rect 427792 228893 427798 228905
rect 427850 228893 427856 228945
rect 427888 228893 427894 228945
rect 427946 228933 427952 228945
rect 547888 228933 547894 228945
rect 427946 228905 547894 228933
rect 427946 228893 427952 228905
rect 547888 228893 547894 228905
rect 547946 228893 547952 228945
rect 242512 228819 242518 228871
rect 242570 228859 242576 228871
rect 294928 228859 294934 228871
rect 242570 228831 294934 228859
rect 242570 228819 242576 228831
rect 294928 228819 294934 228831
rect 294986 228819 294992 228871
rect 310672 228819 310678 228871
rect 310730 228859 310736 228871
rect 430864 228859 430870 228871
rect 310730 228831 430870 228859
rect 310730 228819 310736 228831
rect 430864 228819 430870 228831
rect 430922 228819 430928 228871
rect 432016 228819 432022 228871
rect 432074 228859 432080 228871
rect 529744 228859 529750 228871
rect 432074 228831 529750 228859
rect 432074 228819 432080 228831
rect 529744 228819 529750 228831
rect 529802 228819 529808 228871
rect 241648 228745 241654 228797
rect 241706 228785 241712 228797
rect 289744 228785 289750 228797
rect 241706 228757 289750 228785
rect 241706 228745 241712 228757
rect 289744 228745 289750 228757
rect 289802 228745 289808 228797
rect 304432 228745 304438 228797
rect 304490 228785 304496 228797
rect 418768 228785 418774 228797
rect 304490 228757 418774 228785
rect 304490 228745 304496 228757
rect 418768 228745 418774 228757
rect 418826 228745 418832 228797
rect 434896 228745 434902 228797
rect 434954 228785 434960 228797
rect 454288 228785 454294 228797
rect 434954 228757 454294 228785
rect 434954 228745 434960 228757
rect 454288 228745 454294 228757
rect 454346 228745 454352 228797
rect 239728 228671 239734 228723
rect 239786 228711 239792 228723
rect 288880 228711 288886 228723
rect 239786 228683 288886 228711
rect 239786 228671 239792 228683
rect 288880 228671 288886 228683
rect 288938 228671 288944 228723
rect 306160 228671 306166 228723
rect 306218 228711 306224 228723
rect 421840 228711 421846 228723
rect 306218 228683 421846 228711
rect 306218 228671 306224 228683
rect 421840 228671 421846 228683
rect 421898 228671 421904 228723
rect 231856 228597 231862 228649
rect 231914 228637 231920 228649
rect 272272 228637 272278 228649
rect 231914 228609 272278 228637
rect 231914 228597 231920 228609
rect 272272 228597 272278 228609
rect 272330 228597 272336 228649
rect 291184 228597 291190 228649
rect 291242 228637 291248 228649
rect 382960 228637 382966 228649
rect 291242 228609 382966 228637
rect 291242 228597 291248 228609
rect 382960 228597 382966 228609
rect 383018 228597 383024 228649
rect 404656 228597 404662 228649
rect 404714 228637 404720 228649
rect 517648 228637 517654 228649
rect 404714 228609 517654 228637
rect 404714 228597 404720 228609
rect 517648 228597 517654 228609
rect 517706 228597 517712 228649
rect 190192 228523 190198 228575
rect 190250 228563 190256 228575
rect 192304 228563 192310 228575
rect 190250 228535 192310 228563
rect 190250 228523 190256 228535
rect 192304 228523 192310 228535
rect 192362 228523 192368 228575
rect 228784 228523 228790 228575
rect 228842 228563 228848 228575
rect 266224 228563 266230 228575
rect 228842 228535 266230 228563
rect 228842 228523 228848 228535
rect 266224 228523 266230 228535
rect 266282 228523 266288 228575
rect 266320 228523 266326 228575
rect 266378 228563 266384 228575
rect 301744 228563 301750 228575
rect 266378 228535 301750 228563
rect 266378 228523 266384 228535
rect 301744 228523 301750 228535
rect 301802 228523 301808 228575
rect 303472 228523 303478 228575
rect 303530 228563 303536 228575
rect 413488 228563 413494 228575
rect 303530 228535 413494 228563
rect 303530 228523 303536 228535
rect 413488 228523 413494 228535
rect 413546 228523 413552 228575
rect 455056 228523 455062 228575
rect 455114 228563 455120 228575
rect 456496 228563 456502 228575
rect 455114 228535 456502 228563
rect 455114 228523 455120 228535
rect 456496 228523 456502 228535
rect 456554 228523 456560 228575
rect 478192 228523 478198 228575
rect 478250 228563 478256 228575
rect 480688 228563 480694 228575
rect 478250 228535 480694 228563
rect 478250 228523 478256 228535
rect 480688 228523 480694 228535
rect 480746 228523 480752 228575
rect 512752 228523 512758 228575
rect 512810 228563 512816 228575
rect 514672 228563 514678 228575
rect 512810 228535 514678 228563
rect 512810 228523 512816 228535
rect 514672 228523 514678 228535
rect 514730 228523 514736 228575
rect 535792 228523 535798 228575
rect 535850 228563 535856 228575
rect 538000 228563 538006 228575
rect 535850 228535 538006 228563
rect 535850 228523 535856 228535
rect 538000 228523 538006 228535
rect 538058 228523 538064 228575
rect 544336 228523 544342 228575
rect 544394 228563 544400 228575
rect 547120 228563 547126 228575
rect 544394 228535 547126 228563
rect 544394 228523 544400 228535
rect 547120 228523 547126 228535
rect 547178 228523 547184 228575
rect 567376 228523 567382 228575
rect 567434 228563 567440 228575
rect 569008 228563 569014 228575
rect 567434 228535 569014 228563
rect 567434 228523 567440 228535
rect 569008 228523 569014 228535
rect 569066 228523 569072 228575
rect 224368 228449 224374 228501
rect 224426 228489 224432 228501
rect 258736 228489 258742 228501
rect 224426 228461 258742 228489
rect 224426 228449 224432 228461
rect 258736 228449 258742 228461
rect 258794 228449 258800 228501
rect 260464 228449 260470 228501
rect 260522 228489 260528 228501
rect 286672 228489 286678 228501
rect 260522 228461 286678 228489
rect 260522 228449 260528 228461
rect 286672 228449 286678 228461
rect 286730 228449 286736 228501
rect 289360 228449 289366 228501
rect 289418 228489 289424 228501
rect 380080 228489 380086 228501
rect 289418 228461 380086 228489
rect 289418 228449 289424 228461
rect 380080 228449 380086 228461
rect 380138 228449 380144 228501
rect 407440 228449 407446 228501
rect 407498 228489 407504 228501
rect 502576 228489 502582 228501
rect 407498 228461 502582 228489
rect 407498 228449 407504 228461
rect 502576 228449 502582 228461
rect 502634 228449 502640 228501
rect 250576 228375 250582 228427
rect 250634 228415 250640 228427
rect 276496 228415 276502 228427
rect 250634 228387 276502 228415
rect 250634 228375 250640 228387
rect 276496 228375 276502 228387
rect 276554 228375 276560 228427
rect 288016 228375 288022 228427
rect 288074 228415 288080 228427
rect 328912 228415 328918 228427
rect 288074 228387 328918 228415
rect 288074 228375 288080 228387
rect 328912 228375 328918 228387
rect 328970 228375 328976 228427
rect 331120 228375 331126 228427
rect 331178 228415 331184 228427
rect 467056 228415 467062 228427
rect 331178 228387 467062 228415
rect 331178 228375 331184 228387
rect 467056 228375 467062 228387
rect 467114 228375 467120 228427
rect 535792 228375 535798 228427
rect 535850 228415 535856 228427
rect 537904 228415 537910 228427
rect 535850 228387 537910 228415
rect 535850 228375 535856 228387
rect 537904 228375 537910 228387
rect 537962 228375 537968 228427
rect 259504 228301 259510 228353
rect 259562 228341 259568 228353
rect 292624 228341 292630 228353
rect 259562 228313 292630 228341
rect 259562 228301 259568 228313
rect 292624 228301 292630 228313
rect 292682 228301 292688 228353
rect 293872 228301 293878 228353
rect 293930 228341 293936 228353
rect 380752 228341 380758 228353
rect 293930 228313 380758 228341
rect 293930 228301 293936 228313
rect 380752 228301 380758 228313
rect 380810 228301 380816 228353
rect 391696 228301 391702 228353
rect 391754 228341 391760 228353
rect 476944 228341 476950 228353
rect 391754 228313 476950 228341
rect 391754 228301 391760 228313
rect 476944 228301 476950 228313
rect 477002 228301 477008 228353
rect 270832 228227 270838 228279
rect 270890 228267 270896 228279
rect 313840 228267 313846 228279
rect 270890 228239 313846 228267
rect 270890 228227 270896 228239
rect 313840 228227 313846 228239
rect 313898 228227 313904 228279
rect 313936 228227 313942 228279
rect 313994 228267 314000 228279
rect 392368 228267 392374 228279
rect 313994 228239 392374 228267
rect 313994 228227 314000 228239
rect 392368 228227 392374 228239
rect 392426 228227 392432 228279
rect 392464 228227 392470 228279
rect 392522 228267 392528 228279
rect 461872 228267 461878 228279
rect 392522 228239 461878 228267
rect 392522 228227 392528 228239
rect 461872 228227 461878 228239
rect 461930 228227 461936 228279
rect 267952 228153 267958 228205
rect 268010 228193 268016 228205
rect 307696 228193 307702 228205
rect 268010 228165 307702 228193
rect 268010 228153 268016 228165
rect 307696 228153 307702 228165
rect 307754 228153 307760 228205
rect 311056 228153 311062 228205
rect 311114 228193 311120 228205
rect 383248 228193 383254 228205
rect 311114 228165 383254 228193
rect 311114 228153 311120 228165
rect 383248 228153 383254 228165
rect 383306 228153 383312 228205
rect 394864 228153 394870 228205
rect 394922 228193 394928 228205
rect 437680 228193 437686 228205
rect 394922 228165 437686 228193
rect 394922 228153 394928 228165
rect 437680 228153 437686 228165
rect 437738 228153 437744 228205
rect 293776 228079 293782 228131
rect 293834 228119 293840 228131
rect 343984 228119 343990 228131
rect 293834 228091 343990 228119
rect 293834 228079 293840 228091
rect 343984 228079 343990 228091
rect 344042 228079 344048 228131
rect 345328 228079 345334 228131
rect 345386 228119 345392 228131
rect 412720 228119 412726 228131
rect 345386 228091 412726 228119
rect 345386 228079 345392 228091
rect 412720 228079 412726 228091
rect 412778 228079 412784 228131
rect 258448 228005 258454 228057
rect 258506 228045 258512 228057
rect 280624 228045 280630 228057
rect 258506 228017 280630 228045
rect 258506 228005 258512 228017
rect 280624 228005 280630 228017
rect 280682 228005 280688 228057
rect 298096 228005 298102 228057
rect 298154 228045 298160 228057
rect 362800 228045 362806 228057
rect 298154 228017 362806 228045
rect 298154 228005 298160 228017
rect 362800 228005 362806 228017
rect 362858 228005 362864 228057
rect 362896 228005 362902 228057
rect 362954 228045 362960 228057
rect 425584 228045 425590 228057
rect 362954 228017 425590 228045
rect 362954 228005 362960 228017
rect 425584 228005 425590 228017
rect 425642 228005 425648 228057
rect 290992 227931 290998 227983
rect 291050 227971 291056 227983
rect 341008 227971 341014 227983
rect 291050 227943 341014 227971
rect 291050 227931 291056 227943
rect 341008 227931 341014 227943
rect 341066 227931 341072 227983
rect 342352 227931 342358 227983
rect 342410 227971 342416 227983
rect 398320 227971 398326 227983
rect 342410 227943 398326 227971
rect 342410 227931 342416 227943
rect 398320 227931 398326 227943
rect 398378 227931 398384 227983
rect 247024 227857 247030 227909
rect 247082 227897 247088 227909
rect 303952 227897 303958 227909
rect 247082 227869 303958 227897
rect 247082 227857 247088 227869
rect 303952 227857 303958 227869
rect 304010 227857 304016 227909
rect 308272 227857 308278 227909
rect 308330 227897 308336 227909
rect 359152 227897 359158 227909
rect 308330 227869 359158 227897
rect 308330 227857 308336 227869
rect 359152 227857 359158 227869
rect 359210 227857 359216 227909
rect 263632 227783 263638 227835
rect 263690 227823 263696 227835
rect 295696 227823 295702 227835
rect 263690 227795 295702 227823
rect 263690 227783 263696 227795
rect 295696 227783 295702 227795
rect 295754 227783 295760 227835
rect 302224 227783 302230 227835
rect 302282 227823 302288 227835
rect 350032 227823 350038 227835
rect 302282 227795 350038 227823
rect 302282 227783 302288 227795
rect 350032 227783 350038 227795
rect 350090 227783 350096 227835
rect 319408 227709 319414 227761
rect 319466 227749 319472 227761
rect 319466 227721 325982 227749
rect 319466 227709 319472 227721
rect 282064 227635 282070 227687
rect 282122 227675 282128 227687
rect 325840 227675 325846 227687
rect 282122 227647 325846 227675
rect 282122 227635 282128 227647
rect 325840 227635 325846 227647
rect 325898 227635 325904 227687
rect 149392 227561 149398 227613
rect 149450 227601 149456 227613
rect 174256 227601 174262 227613
rect 149450 227573 174262 227601
rect 149450 227561 149456 227573
rect 174256 227561 174262 227573
rect 174314 227561 174320 227613
rect 278128 227561 278134 227613
rect 278186 227601 278192 227613
rect 319888 227601 319894 227613
rect 278186 227573 319894 227601
rect 278186 227561 278192 227573
rect 319888 227561 319894 227573
rect 319946 227561 319952 227613
rect 325954 227601 325982 227721
rect 326800 227709 326806 227761
rect 326858 227749 326864 227761
rect 353104 227749 353110 227761
rect 326858 227721 353110 227749
rect 326858 227709 326864 227721
rect 353104 227709 353110 227721
rect 353162 227709 353168 227761
rect 387760 227635 387766 227687
rect 387818 227675 387824 227687
rect 396400 227675 396406 227687
rect 387818 227647 396406 227675
rect 387818 227635 387824 227647
rect 396400 227635 396406 227647
rect 396458 227635 396464 227687
rect 403696 227601 403702 227613
rect 325954 227573 403702 227601
rect 403696 227561 403702 227573
rect 403754 227561 403760 227613
rect 418288 227561 418294 227613
rect 418346 227601 418352 227613
rect 433168 227601 433174 227613
rect 418346 227573 433174 227601
rect 418346 227561 418352 227573
rect 433168 227561 433174 227573
rect 433226 227561 433232 227613
rect 187120 227487 187126 227539
rect 187178 227527 187184 227539
rect 190768 227527 190774 227539
rect 187178 227499 190774 227527
rect 187178 227487 187184 227499
rect 190768 227487 190774 227499
rect 190826 227487 190832 227539
rect 216112 227487 216118 227539
rect 216170 227527 216176 227539
rect 239824 227527 239830 227539
rect 216170 227499 239830 227527
rect 216170 227487 216176 227499
rect 239824 227487 239830 227499
rect 239882 227487 239888 227539
rect 249328 227487 249334 227539
rect 249386 227527 249392 227539
rect 306256 227527 306262 227539
rect 249386 227499 306262 227527
rect 249386 227487 249392 227499
rect 306256 227487 306262 227499
rect 306314 227487 306320 227539
rect 311248 227487 311254 227539
rect 311306 227527 311312 227539
rect 375760 227527 375766 227539
rect 311306 227499 375766 227527
rect 311306 227487 311312 227499
rect 375760 227487 375766 227499
rect 375818 227487 375824 227539
rect 389488 227487 389494 227539
rect 389546 227527 389552 227539
rect 587152 227527 587158 227539
rect 389546 227499 587158 227527
rect 389546 227487 389552 227499
rect 587152 227487 587158 227499
rect 587210 227487 587216 227539
rect 588880 227487 588886 227539
rect 588938 227527 588944 227539
rect 615856 227527 615862 227539
rect 588938 227499 615862 227527
rect 588938 227487 588944 227499
rect 615856 227487 615862 227499
rect 615914 227487 615920 227539
rect 238768 227413 238774 227465
rect 238826 227453 238832 227465
rect 252016 227453 252022 227465
rect 238826 227425 252022 227453
rect 238826 227413 238832 227425
rect 252016 227413 252022 227425
rect 252074 227413 252080 227465
rect 253840 227413 253846 227465
rect 253898 227453 253904 227465
rect 315376 227453 315382 227465
rect 253898 227425 315382 227453
rect 253898 227413 253904 227425
rect 315376 227413 315382 227425
rect 315434 227413 315440 227465
rect 318352 227413 318358 227465
rect 318410 227453 318416 227465
rect 381808 227453 381814 227465
rect 318410 227425 381814 227453
rect 318410 227413 318416 227425
rect 381808 227413 381814 227425
rect 381866 227413 381872 227465
rect 390064 227413 390070 227465
rect 390122 227453 390128 227465
rect 588592 227453 588598 227465
rect 390122 227425 588598 227453
rect 390122 227413 390128 227425
rect 588592 227413 588598 227425
rect 588650 227413 588656 227465
rect 588976 227413 588982 227465
rect 589034 227453 589040 227465
rect 618832 227453 618838 227465
rect 589034 227425 618838 227453
rect 589034 227413 589040 227425
rect 618832 227413 618838 227425
rect 618890 227413 618896 227465
rect 217072 227339 217078 227391
rect 217130 227379 217136 227391
rect 243568 227379 243574 227391
rect 217130 227351 243574 227379
rect 217130 227339 217136 227351
rect 243568 227339 243574 227351
rect 243626 227339 243632 227391
rect 311344 227339 311350 227391
rect 311402 227379 311408 227391
rect 384016 227379 384022 227391
rect 311402 227351 384022 227379
rect 311402 227339 311408 227351
rect 384016 227339 384022 227351
rect 384074 227339 384080 227391
rect 392272 227339 392278 227391
rect 392330 227379 392336 227391
rect 593104 227379 593110 227391
rect 392330 227351 593110 227379
rect 392330 227339 392336 227351
rect 593104 227339 593110 227351
rect 593162 227339 593168 227391
rect 606256 227339 606262 227391
rect 606314 227379 606320 227391
rect 639184 227379 639190 227391
rect 606314 227351 639190 227379
rect 606314 227339 606320 227351
rect 639184 227339 639190 227351
rect 639242 227339 639248 227391
rect 236752 227265 236758 227317
rect 236810 227305 236816 227317
rect 261040 227305 261046 227317
rect 236810 227277 261046 227305
rect 236810 227265 236816 227277
rect 261040 227265 261046 227277
rect 261098 227265 261104 227317
rect 274672 227265 274678 227317
rect 274730 227305 274736 227317
rect 348592 227305 348598 227317
rect 274730 227277 348598 227305
rect 274730 227265 274736 227277
rect 348592 227265 348598 227277
rect 348650 227265 348656 227317
rect 390832 227265 390838 227317
rect 390890 227305 390896 227317
rect 590128 227305 590134 227317
rect 390890 227277 590134 227305
rect 390890 227265 390896 227277
rect 590128 227265 590134 227277
rect 590186 227265 590192 227317
rect 599056 227265 599062 227317
rect 599114 227305 599120 227317
rect 633136 227305 633142 227317
rect 599114 227277 633142 227305
rect 599114 227265 599120 227277
rect 633136 227265 633142 227277
rect 633194 227265 633200 227317
rect 217840 227191 217846 227243
rect 217898 227231 217904 227243
rect 242896 227231 242902 227243
rect 217898 227203 242902 227231
rect 217898 227191 217904 227203
rect 242896 227191 242902 227203
rect 242954 227191 242960 227243
rect 253552 227191 253558 227243
rect 253610 227231 253616 227243
rect 266992 227231 266998 227243
rect 253610 227203 266998 227231
rect 253610 227191 253616 227203
rect 266992 227191 266998 227203
rect 267050 227191 267056 227243
rect 271984 227191 271990 227243
rect 272042 227231 272048 227243
rect 351568 227231 351574 227243
rect 272042 227203 351574 227231
rect 272042 227191 272048 227203
rect 351568 227191 351574 227203
rect 351626 227191 351632 227243
rect 388528 227191 388534 227243
rect 388586 227231 388592 227243
rect 585616 227231 585622 227243
rect 388586 227203 585622 227231
rect 388586 227191 388592 227203
rect 585616 227191 585622 227203
rect 585674 227191 585680 227243
rect 587344 227191 587350 227243
rect 587402 227231 587408 227243
rect 616624 227231 616630 227243
rect 587402 227203 616630 227231
rect 587402 227191 587408 227203
rect 616624 227191 616630 227203
rect 616682 227191 616688 227243
rect 215728 227117 215734 227169
rect 215786 227157 215792 227169
rect 238384 227157 238390 227169
rect 215786 227129 238390 227157
rect 215786 227117 215792 227129
rect 238384 227117 238390 227129
rect 238442 227117 238448 227169
rect 238960 227117 238966 227169
rect 239018 227157 239024 227169
rect 264016 227157 264022 227169
rect 239018 227129 264022 227157
rect 239018 227117 239024 227129
rect 264016 227117 264022 227129
rect 264074 227117 264080 227169
rect 264688 227117 264694 227169
rect 264746 227157 264752 227169
rect 288112 227157 288118 227169
rect 264746 227129 288118 227157
rect 264746 227117 264752 227129
rect 288112 227117 288118 227129
rect 288170 227117 288176 227169
rect 289648 227117 289654 227169
rect 289706 227157 289712 227169
rect 369616 227157 369622 227169
rect 289706 227129 369622 227157
rect 289706 227117 289712 227129
rect 369616 227117 369622 227129
rect 369674 227117 369680 227169
rect 385648 227117 385654 227169
rect 385706 227157 385712 227169
rect 398800 227157 398806 227169
rect 385706 227129 398806 227157
rect 385706 227117 385712 227129
rect 398800 227117 398806 227129
rect 398858 227117 398864 227169
rect 398896 227117 398902 227169
rect 398954 227157 398960 227169
rect 584848 227157 584854 227169
rect 398954 227129 584854 227157
rect 398954 227117 398960 227129
rect 584848 227117 584854 227129
rect 584906 227117 584912 227169
rect 587440 227117 587446 227169
rect 587498 227157 587504 227169
rect 619600 227157 619606 227169
rect 587498 227129 619606 227157
rect 587498 227117 587504 227129
rect 619600 227117 619606 227129
rect 619658 227117 619664 227169
rect 219472 227043 219478 227095
rect 219530 227083 219536 227095
rect 245872 227083 245878 227095
rect 219530 227055 245878 227083
rect 219530 227043 219536 227055
rect 245872 227043 245878 227055
rect 245930 227043 245936 227095
rect 276688 227043 276694 227095
rect 276746 227083 276752 227095
rect 360592 227083 360598 227095
rect 276746 227055 360598 227083
rect 276746 227043 276752 227055
rect 360592 227043 360598 227055
rect 360650 227043 360656 227095
rect 390448 227043 390454 227095
rect 390506 227083 390512 227095
rect 589360 227083 589366 227095
rect 390506 227055 589366 227083
rect 390506 227043 390512 227055
rect 589360 227043 589366 227055
rect 589418 227043 589424 227095
rect 606352 227043 606358 227095
rect 606410 227083 606416 227095
rect 638512 227083 638518 227095
rect 606410 227055 638518 227083
rect 606410 227043 606416 227055
rect 638512 227043 638518 227055
rect 638570 227043 638576 227095
rect 149392 226969 149398 227021
rect 149450 227009 149456 227021
rect 159760 227009 159766 227021
rect 149450 226981 159766 227009
rect 149450 226969 149456 226981
rect 159760 226969 159766 226981
rect 159818 226969 159824 227021
rect 213808 226969 213814 227021
rect 213866 227009 213872 227021
rect 237520 227009 237526 227021
rect 213866 226981 237526 227009
rect 213866 226969 213872 226981
rect 237520 226969 237526 226981
rect 237578 226969 237584 227021
rect 240496 226969 240502 227021
rect 240554 227009 240560 227021
rect 248848 227009 248854 227021
rect 240554 226981 248854 227009
rect 240554 226969 240560 226981
rect 248848 226969 248854 226981
rect 248906 226969 248912 227021
rect 275248 226969 275254 227021
rect 275306 227009 275312 227021
rect 357616 227009 357622 227021
rect 275306 226981 357622 227009
rect 275306 226969 275312 226981
rect 357616 226969 357622 226981
rect 357674 226969 357680 227021
rect 392656 226969 392662 227021
rect 392714 227009 392720 227021
rect 593968 227009 593974 227021
rect 392714 226981 593974 227009
rect 392714 226969 392720 226981
rect 593968 226969 593974 226981
rect 594026 226969 594032 227021
rect 603472 226969 603478 227021
rect 603530 227009 603536 227021
rect 636208 227009 636214 227021
rect 603530 226981 636214 227009
rect 603530 226969 603536 226981
rect 636208 226969 636214 226981
rect 636266 226969 636272 227021
rect 221680 226895 221686 226947
rect 221738 226935 221744 226947
rect 250384 226935 250390 226947
rect 221738 226907 250390 226935
rect 221738 226895 221744 226907
rect 250384 226895 250390 226907
rect 250442 226895 250448 226947
rect 273424 226895 273430 226947
rect 273482 226935 273488 226947
rect 354544 226935 354550 226947
rect 273482 226907 354550 226935
rect 273482 226895 273488 226907
rect 354544 226895 354550 226907
rect 354602 226895 354608 226947
rect 359824 226895 359830 226947
rect 359882 226935 359888 226947
rect 393136 226935 393142 226947
rect 359882 226907 393142 226935
rect 359882 226895 359888 226907
rect 393136 226895 393142 226907
rect 393194 226895 393200 226947
rect 395536 226895 395542 226947
rect 395594 226935 395600 226947
rect 599152 226935 599158 226947
rect 395594 226907 599158 226935
rect 395594 226895 395600 226907
rect 599152 226895 599158 226907
rect 599210 226895 599216 226947
rect 600400 226895 600406 226947
rect 600458 226935 600464 226947
rect 634672 226935 634678 226947
rect 600458 226907 634678 226935
rect 600458 226895 600464 226907
rect 634672 226895 634678 226907
rect 634730 226895 634736 226947
rect 223312 226821 223318 226873
rect 223370 226861 223376 226873
rect 253456 226861 253462 226873
rect 223370 226833 253462 226861
rect 223370 226821 223376 226833
rect 253456 226821 253462 226833
rect 253514 226821 253520 226873
rect 324112 226821 324118 226873
rect 324170 226861 324176 226873
rect 339472 226861 339478 226873
rect 324170 226833 339478 226861
rect 324170 226821 324176 226833
rect 339472 226821 339478 226833
rect 339530 226821 339536 226873
rect 364048 226821 364054 226873
rect 364106 226861 364112 226873
rect 396112 226861 396118 226873
rect 364106 226833 396118 226861
rect 364106 226821 364112 226833
rect 396112 226821 396118 226833
rect 396170 226821 396176 226873
rect 399376 226821 399382 226873
rect 399434 226861 399440 226873
rect 419344 226861 419350 226873
rect 399434 226833 419350 226861
rect 399434 226821 399440 226833
rect 419344 226821 419350 226833
rect 419402 226821 419408 226873
rect 419440 226821 419446 226873
rect 419498 226861 419504 226873
rect 603664 226861 603670 226873
rect 419498 226833 603670 226861
rect 419498 226821 419504 226833
rect 603664 226821 603670 226833
rect 603722 226821 603728 226873
rect 606160 226821 606166 226873
rect 606218 226861 606224 226873
rect 639952 226861 639958 226873
rect 606218 226833 639958 226861
rect 606218 226821 606224 226833
rect 639952 226821 639958 226833
rect 640010 226821 640016 226873
rect 224944 226747 224950 226799
rect 225002 226787 225008 226799
rect 256432 226787 256438 226799
rect 225002 226759 256438 226787
rect 225002 226747 225008 226759
rect 256432 226747 256438 226759
rect 256490 226747 256496 226799
rect 257104 226747 257110 226799
rect 257162 226787 257168 226799
rect 273232 226787 273238 226799
rect 257162 226759 273238 226787
rect 257162 226747 257168 226759
rect 273232 226747 273238 226759
rect 273290 226747 273296 226799
rect 279760 226747 279766 226799
rect 279818 226787 279824 226799
rect 298192 226787 298198 226799
rect 279818 226759 298198 226787
rect 279818 226747 279824 226759
rect 298192 226747 298198 226759
rect 298250 226747 298256 226799
rect 298384 226747 298390 226799
rect 298442 226787 298448 226799
rect 366736 226787 366742 226799
rect 298442 226759 366742 226787
rect 298442 226747 298448 226759
rect 366736 226747 366742 226759
rect 366794 226747 366800 226799
rect 374608 226747 374614 226799
rect 374666 226787 374672 226799
rect 391504 226787 391510 226799
rect 374666 226759 391510 226787
rect 374666 226747 374672 226759
rect 391504 226747 391510 226759
rect 391562 226747 391568 226799
rect 397168 226747 397174 226799
rect 397226 226787 397232 226799
rect 602992 226787 602998 226799
rect 397226 226759 419006 226787
rect 397226 226747 397232 226759
rect 227920 226673 227926 226725
rect 227978 226713 227984 226725
rect 262480 226713 262486 226725
rect 227978 226685 262486 226713
rect 227978 226673 227984 226685
rect 262480 226673 262486 226685
rect 262538 226673 262544 226725
rect 284656 226673 284662 226725
rect 284714 226713 284720 226725
rect 298096 226713 298102 226725
rect 284714 226685 298102 226713
rect 284714 226673 284720 226685
rect 298096 226673 298102 226685
rect 298154 226673 298160 226725
rect 299152 226673 299158 226725
rect 299210 226713 299216 226725
rect 372688 226713 372694 226725
rect 299210 226685 372694 226713
rect 299210 226673 299216 226685
rect 372688 226673 372694 226685
rect 372746 226673 372752 226725
rect 372784 226673 372790 226725
rect 372842 226713 372848 226725
rect 393808 226713 393814 226725
rect 372842 226685 393814 226713
rect 372842 226673 372848 226685
rect 393808 226673 393814 226685
rect 393866 226673 393872 226725
rect 400816 226673 400822 226725
rect 400874 226713 400880 226725
rect 418978 226713 419006 226759
rect 419458 226759 602998 226787
rect 419458 226713 419486 226759
rect 602992 226747 602998 226759
rect 603050 226747 603056 226799
rect 603376 226747 603382 226799
rect 603434 226787 603440 226799
rect 636880 226787 636886 226799
rect 603434 226759 636886 226787
rect 603434 226747 603440 226759
rect 636880 226747 636886 226759
rect 636938 226747 636944 226799
rect 400874 226685 418910 226713
rect 418978 226685 419486 226713
rect 400874 226673 400880 226685
rect 226576 226599 226582 226651
rect 226634 226639 226640 226651
rect 259408 226639 259414 226651
rect 226634 226611 259414 226639
rect 226634 226599 226640 226611
rect 259408 226599 259414 226611
rect 259466 226599 259472 226651
rect 268144 226599 268150 226651
rect 268202 226639 268208 226651
rect 282064 226639 282070 226651
rect 268202 226611 282070 226639
rect 268202 226599 268208 226611
rect 282064 226599 282070 226611
rect 282122 226599 282128 226651
rect 285712 226599 285718 226651
rect 285770 226639 285776 226651
rect 378736 226639 378742 226651
rect 285770 226611 378742 226639
rect 285770 226599 285776 226611
rect 378736 226599 378742 226611
rect 378794 226599 378800 226651
rect 379984 226599 379990 226651
rect 380042 226639 380048 226651
rect 394576 226639 394582 226651
rect 380042 226611 394582 226639
rect 380042 226599 380048 226611
rect 394576 226599 394582 226611
rect 394634 226599 394640 226651
rect 397648 226599 397654 226651
rect 397706 226639 397712 226651
rect 418672 226639 418678 226651
rect 397706 226611 418678 226639
rect 397706 226599 397712 226611
rect 418672 226599 418678 226611
rect 418730 226599 418736 226651
rect 418882 226639 418910 226685
rect 419632 226673 419638 226725
rect 419690 226713 419696 226725
rect 606736 226713 606742 226725
rect 419690 226685 606742 226713
rect 419690 226673 419696 226685
rect 606736 226673 606742 226685
rect 606794 226673 606800 226725
rect 609808 226639 609814 226651
rect 418882 226611 609814 226639
rect 609808 226599 609814 226611
rect 609866 226599 609872 226651
rect 629296 226599 629302 226651
rect 629354 226639 629360 226651
rect 634000 226639 634006 226651
rect 629354 226611 634006 226639
rect 629354 226599 629360 226611
rect 634000 226599 634006 226611
rect 634058 226599 634064 226651
rect 229552 226525 229558 226577
rect 229610 226565 229616 226577
rect 265552 226565 265558 226577
rect 229610 226537 265558 226565
rect 229610 226525 229616 226537
rect 265552 226525 265558 226537
rect 265610 226525 265616 226577
rect 271024 226525 271030 226577
rect 271082 226565 271088 226577
rect 294256 226565 294262 226577
rect 271082 226537 294262 226565
rect 271082 226525 271088 226537
rect 294256 226525 294262 226537
rect 294314 226525 294320 226577
rect 297328 226525 297334 226577
rect 297386 226565 297392 226577
rect 390064 226565 390070 226577
rect 297386 226537 390070 226565
rect 297386 226525 297392 226537
rect 390064 226525 390070 226537
rect 390122 226525 390128 226577
rect 401200 226525 401206 226577
rect 401258 226565 401264 226577
rect 610480 226565 610486 226577
rect 401258 226537 610486 226565
rect 401258 226525 401264 226537
rect 610480 226525 610486 226537
rect 610538 226525 610544 226577
rect 231088 226451 231094 226503
rect 231146 226491 231152 226503
rect 268528 226491 268534 226503
rect 231146 226463 268534 226491
rect 231146 226451 231152 226463
rect 268528 226451 268534 226463
rect 268586 226451 268592 226503
rect 288496 226451 288502 226503
rect 288554 226491 288560 226503
rect 288554 226463 380510 226491
rect 288554 226451 288560 226463
rect 232528 226377 232534 226429
rect 232586 226417 232592 226429
rect 271600 226417 271606 226429
rect 232586 226389 271606 226417
rect 232586 226377 232592 226389
rect 271600 226377 271606 226389
rect 271658 226377 271664 226429
rect 298096 226377 298102 226429
rect 298154 226417 298160 226429
rect 378064 226417 378070 226429
rect 298154 226389 378070 226417
rect 298154 226377 298160 226389
rect 378064 226377 378070 226389
rect 378122 226377 378128 226429
rect 380482 226417 380510 226463
rect 380560 226451 380566 226503
rect 380618 226491 380624 226503
rect 387760 226491 387766 226503
rect 380618 226463 387766 226491
rect 380618 226451 380624 226463
rect 387760 226451 387766 226463
rect 387818 226451 387824 226503
rect 388144 226451 388150 226503
rect 388202 226491 388208 226503
rect 398896 226491 398902 226503
rect 388202 226463 398902 226491
rect 388202 226451 388208 226463
rect 398896 226451 398902 226463
rect 398954 226451 398960 226503
rect 402160 226451 402166 226503
rect 402218 226491 402224 226503
rect 612784 226491 612790 226503
rect 402218 226463 612790 226491
rect 402218 226451 402224 226463
rect 612784 226451 612790 226463
rect 612842 226451 612848 226503
rect 384784 226417 384790 226429
rect 380482 226389 384790 226417
rect 384784 226377 384790 226389
rect 384842 226377 384848 226429
rect 385840 226377 385846 226429
rect 385898 226417 385904 226429
rect 388816 226417 388822 226429
rect 385898 226389 388822 226417
rect 385898 226377 385904 226389
rect 388816 226377 388822 226389
rect 388874 226377 388880 226429
rect 388912 226377 388918 226429
rect 388970 226417 388976 226429
rect 402832 226417 402838 226429
rect 388970 226389 402838 226417
rect 388970 226377 388976 226389
rect 402832 226377 402838 226389
rect 402890 226377 402896 226429
rect 404944 226377 404950 226429
rect 405002 226417 405008 226429
rect 618064 226417 618070 226429
rect 405002 226389 618070 226417
rect 405002 226377 405008 226389
rect 618064 226377 618070 226389
rect 618122 226377 618128 226429
rect 212368 226303 212374 226355
rect 212426 226343 212432 226355
rect 234544 226343 234550 226355
rect 212426 226315 234550 226343
rect 212426 226303 212432 226315
rect 234544 226303 234550 226315
rect 234602 226303 234608 226355
rect 243952 226303 243958 226355
rect 244010 226343 244016 226355
rect 251920 226343 251926 226355
rect 244010 226315 251926 226343
rect 244010 226303 244016 226315
rect 251920 226303 251926 226315
rect 251978 226303 251984 226355
rect 252016 226303 252022 226355
rect 252074 226343 252080 226355
rect 285136 226343 285142 226355
rect 252074 226315 285142 226343
rect 252074 226303 252080 226315
rect 285136 226303 285142 226315
rect 285194 226303 285200 226355
rect 291568 226303 291574 226355
rect 291626 226343 291632 226355
rect 390832 226343 390838 226355
rect 291626 226315 390838 226343
rect 291626 226303 291632 226315
rect 390832 226303 390838 226315
rect 390890 226303 390896 226355
rect 398704 226303 398710 226355
rect 398762 226343 398768 226355
rect 398762 226315 404318 226343
rect 398762 226303 398768 226315
rect 220336 226229 220342 226281
rect 220394 226269 220400 226281
rect 247408 226269 247414 226281
rect 220394 226241 247414 226269
rect 220394 226229 220400 226241
rect 247408 226229 247414 226241
rect 247466 226229 247472 226281
rect 297232 226269 297238 226281
rect 250690 226241 297238 226269
rect 215632 226155 215638 226207
rect 215690 226195 215696 226207
rect 240592 226195 240598 226207
rect 215690 226167 240598 226195
rect 215690 226155 215696 226167
rect 240592 226155 240598 226167
rect 240650 226155 240656 226207
rect 245008 226155 245014 226207
rect 245066 226195 245072 226207
rect 250690 226195 250718 226241
rect 297232 226229 297238 226241
rect 297290 226229 297296 226281
rect 297616 226229 297622 226281
rect 297674 226269 297680 226281
rect 388912 226269 388918 226281
rect 297674 226241 388918 226269
rect 297674 226229 297680 226241
rect 388912 226229 388918 226241
rect 388970 226229 388976 226281
rect 389008 226229 389014 226281
rect 389066 226269 389072 226281
rect 398992 226269 398998 226281
rect 389066 226241 398998 226269
rect 389066 226229 389072 226241
rect 398992 226229 398998 226241
rect 399050 226229 399056 226281
rect 404290 226269 404318 226315
rect 404368 226303 404374 226355
rect 404426 226343 404432 226355
rect 617296 226343 617302 226355
rect 404426 226315 617302 226343
rect 404426 226303 404432 226315
rect 617296 226303 617302 226315
rect 617354 226303 617360 226355
rect 404464 226269 404470 226281
rect 404290 226241 404470 226269
rect 404464 226229 404470 226241
rect 404522 226229 404528 226281
rect 407728 226229 407734 226281
rect 407786 226269 407792 226281
rect 624112 226269 624118 226281
rect 407786 226241 624118 226269
rect 407786 226229 407792 226241
rect 624112 226229 624118 226241
rect 624170 226229 624176 226281
rect 291184 226195 291190 226207
rect 245066 226167 250718 226195
rect 250882 226167 291190 226195
rect 245066 226155 245072 226167
rect 151120 226081 151126 226133
rect 151178 226121 151184 226133
rect 187120 226121 187126 226133
rect 151178 226093 187126 226121
rect 151178 226081 151184 226093
rect 187120 226081 187126 226093
rect 187178 226081 187184 226133
rect 214576 226007 214582 226059
rect 214634 226047 214640 226059
rect 236848 226047 236854 226059
rect 214634 226019 236854 226047
rect 214634 226007 214640 226019
rect 236848 226007 236854 226019
rect 236906 226007 236912 226059
rect 241840 226007 241846 226059
rect 241898 226047 241904 226059
rect 250882 226047 250910 226167
rect 291184 226155 291190 226167
rect 291242 226155 291248 226207
rect 300688 226155 300694 226207
rect 300746 226195 300752 226207
rect 408976 226195 408982 226207
rect 300746 226167 408982 226195
rect 300746 226155 300752 226167
rect 408976 226155 408982 226167
rect 409034 226155 409040 226207
rect 418672 226155 418678 226207
rect 418730 226195 418736 226207
rect 419440 226195 419446 226207
rect 418730 226167 419446 226195
rect 418730 226155 418736 226167
rect 419440 226155 419446 226167
rect 419498 226155 419504 226207
rect 300208 226121 300214 226133
rect 241898 226019 250910 226047
rect 256306 226093 300214 226121
rect 241898 226007 241904 226019
rect 213040 225933 213046 225985
rect 213098 225973 213104 225985
rect 233776 225973 233782 225985
rect 213098 225945 233782 225973
rect 213098 225933 213104 225945
rect 233776 225933 233782 225945
rect 233834 225933 233840 225985
rect 246544 225933 246550 225985
rect 246602 225973 246608 225985
rect 256306 225973 256334 226093
rect 300208 226081 300214 226093
rect 300266 226081 300272 226133
rect 301264 226081 301270 226133
rect 301322 226121 301328 226133
rect 411280 226121 411286 226133
rect 301322 226093 411286 226121
rect 301322 226081 301328 226093
rect 411280 226081 411286 226093
rect 411338 226081 411344 226133
rect 411664 226081 411670 226133
rect 411722 226121 411728 226133
rect 631696 226121 631702 226133
rect 411722 226093 631702 226121
rect 411722 226081 411728 226093
rect 631696 226081 631702 226093
rect 631754 226081 631760 226133
rect 264880 226007 264886 226059
rect 264938 226047 264944 226059
rect 276112 226047 276118 226059
rect 264938 226019 276118 226047
rect 264938 226007 264944 226019
rect 276112 226007 276118 226019
rect 276170 226007 276176 226059
rect 334288 226007 334294 226059
rect 334346 226047 334352 226059
rect 380560 226047 380566 226059
rect 334346 226019 380566 226047
rect 334346 226007 334352 226019
rect 380560 226007 380566 226019
rect 380618 226007 380624 226059
rect 386992 226047 386998 226059
rect 380674 226019 386998 226047
rect 246602 225945 256334 225973
rect 246602 225933 246608 225945
rect 267760 225933 267766 225985
rect 267818 225973 267824 225985
rect 267818 225945 273182 225973
rect 267818 225933 267824 225945
rect 217456 225859 217462 225911
rect 217514 225899 217520 225911
rect 241264 225899 241270 225911
rect 217514 225871 241270 225899
rect 217514 225859 217520 225871
rect 241264 225859 241270 225871
rect 241322 225859 241328 225911
rect 262000 225859 262006 225911
rect 262058 225899 262064 225911
rect 273040 225899 273046 225911
rect 262058 225871 273046 225899
rect 262058 225859 262064 225871
rect 273040 225859 273046 225871
rect 273098 225859 273104 225911
rect 273154 225899 273182 225945
rect 273232 225933 273238 225985
rect 273290 225973 273296 225985
rect 321328 225973 321334 225985
rect 273290 225945 321334 225973
rect 273290 225933 273296 225945
rect 321328 225933 321334 225945
rect 321386 225933 321392 225985
rect 380674 225973 380702 226019
rect 386992 226007 386998 226019
rect 387050 226007 387056 226059
rect 388816 226007 388822 226059
rect 388874 226047 388880 226059
rect 398704 226047 398710 226059
rect 388874 226019 398710 226047
rect 388874 226007 388880 226019
rect 398704 226007 398710 226019
rect 398762 226007 398768 226059
rect 398800 226007 398806 226059
rect 398858 226047 398864 226059
rect 398858 226019 398942 226047
rect 398858 226007 398864 226019
rect 368626 225945 380702 225973
rect 327376 225899 327382 225911
rect 273154 225871 327382 225899
rect 327376 225859 327382 225871
rect 327434 225859 327440 225911
rect 331408 225859 331414 225911
rect 331466 225899 331472 225911
rect 345520 225899 345526 225911
rect 331466 225871 345526 225899
rect 331466 225859 331472 225871
rect 345520 225859 345526 225871
rect 345578 225859 345584 225911
rect 346960 225859 346966 225911
rect 347018 225899 347024 225911
rect 368626 225899 368654 225945
rect 380752 225933 380758 225985
rect 380810 225973 380816 225985
rect 386416 225973 386422 225985
rect 380810 225945 386422 225973
rect 380810 225933 380816 225945
rect 386416 225933 386422 225945
rect 386474 225933 386480 225985
rect 386608 225933 386614 225985
rect 386666 225973 386672 225985
rect 398914 225973 398942 226019
rect 398992 226007 398998 226059
rect 399050 226047 399056 226059
rect 586384 226047 586390 226059
rect 399050 226019 586390 226047
rect 399050 226007 399056 226019
rect 586384 226007 586390 226019
rect 586442 226007 586448 226059
rect 587824 226007 587830 226059
rect 587882 226047 587888 226059
rect 594640 226047 594646 226059
rect 587882 226019 594646 226047
rect 587882 226007 587888 226019
rect 594640 226007 594646 226019
rect 594698 226007 594704 226059
rect 603280 226007 603286 226059
rect 603338 226047 603344 226059
rect 637744 226047 637750 226059
rect 603338 226019 637750 226047
rect 603338 226007 603344 226019
rect 637744 226007 637750 226019
rect 637802 226007 637808 226059
rect 579568 225973 579574 225985
rect 386666 225945 398846 225973
rect 398914 225945 579574 225973
rect 386666 225933 386672 225945
rect 347018 225871 368654 225899
rect 347018 225859 347024 225871
rect 374416 225859 374422 225911
rect 374474 225899 374480 225911
rect 385552 225899 385558 225911
rect 374474 225871 385558 225899
rect 374474 225859 374480 225871
rect 385552 225859 385558 225871
rect 385610 225859 385616 225911
rect 387280 225859 387286 225911
rect 387338 225899 387344 225911
rect 398608 225899 398614 225911
rect 387338 225871 398614 225899
rect 387338 225859 387344 225871
rect 398608 225859 398614 225871
rect 398666 225859 398672 225911
rect 218800 225785 218806 225837
rect 218858 225825 218864 225837
rect 244336 225825 244342 225837
rect 218858 225797 244342 225825
rect 218858 225785 218864 225797
rect 244336 225785 244342 225797
rect 244394 225785 244400 225837
rect 269584 225785 269590 225837
rect 269642 225825 269648 225837
rect 330448 225825 330454 225837
rect 269642 225797 330454 225825
rect 269642 225785 269648 225797
rect 330448 225785 330454 225797
rect 330506 225785 330512 225837
rect 374512 225785 374518 225837
rect 374570 225825 374576 225837
rect 382576 225825 382582 225837
rect 374570 225797 382582 225825
rect 374570 225785 374576 225797
rect 382576 225785 382582 225797
rect 382634 225785 382640 225837
rect 382960 225785 382966 225837
rect 383018 225825 383024 225837
rect 389296 225825 389302 225837
rect 383018 225797 389302 225825
rect 383018 225785 383024 225797
rect 389296 225785 389302 225797
rect 389354 225785 389360 225837
rect 398818 225825 398846 225945
rect 579568 225933 579574 225945
rect 579626 225933 579632 225985
rect 587056 225933 587062 225985
rect 587114 225973 587120 225985
rect 595408 225973 595414 225985
rect 587114 225945 595414 225973
rect 587114 225933 587120 225945
rect 595408 225933 595414 225945
rect 595466 225933 595472 225985
rect 398896 225859 398902 225911
rect 398954 225899 398960 225911
rect 582640 225899 582646 225911
rect 398954 225871 582646 225899
rect 398954 225859 398960 225871
rect 582640 225859 582646 225871
rect 582698 225859 582704 225911
rect 629200 225859 629206 225911
rect 629258 225899 629264 225911
rect 635440 225899 635446 225911
rect 629258 225871 635446 225899
rect 629258 225859 629264 225871
rect 635440 225859 635446 225871
rect 635498 225859 635504 225911
rect 581104 225825 581110 225837
rect 398818 225797 581110 225825
rect 581104 225785 581110 225797
rect 581162 225785 581168 225837
rect 218320 225711 218326 225763
rect 218378 225751 218384 225763
rect 246640 225751 246646 225763
rect 218378 225723 246646 225751
rect 218378 225711 218384 225723
rect 246640 225711 246646 225723
rect 246698 225711 246704 225763
rect 247696 225711 247702 225763
rect 247754 225751 247760 225763
rect 257968 225751 257974 225763
rect 247754 225723 257974 225751
rect 247754 225711 247760 225723
rect 257968 225711 257974 225723
rect 258026 225711 258032 225763
rect 266416 225711 266422 225763
rect 266474 225751 266480 225763
rect 279088 225751 279094 225763
rect 266474 225723 279094 225751
rect 266474 225711 266480 225723
rect 279088 225711 279094 225723
rect 279146 225711 279152 225763
rect 285040 225711 285046 225763
rect 285098 225751 285104 225763
rect 342544 225751 342550 225763
rect 285098 225723 342550 225751
rect 285098 225711 285104 225723
rect 342544 225711 342550 225723
rect 342602 225711 342608 225763
rect 371536 225711 371542 225763
rect 371594 225751 371600 225763
rect 379504 225751 379510 225763
rect 371594 225723 379510 225751
rect 371594 225711 371600 225723
rect 379504 225711 379510 225723
rect 379562 225711 379568 225763
rect 380080 225711 380086 225763
rect 380138 225751 380144 225763
rect 388624 225751 388630 225763
rect 380138 225723 388630 225751
rect 380138 225711 380144 225723
rect 388624 225711 388630 225723
rect 388682 225711 388688 225763
rect 396400 225711 396406 225763
rect 396458 225751 396464 225763
rect 584080 225751 584086 225763
rect 396458 225723 584086 225751
rect 396458 225711 396464 225723
rect 584080 225711 584086 225723
rect 584138 225711 584144 225763
rect 278224 225637 278230 225689
rect 278282 225677 278288 225689
rect 318352 225677 318358 225689
rect 278282 225649 318358 225677
rect 278282 225637 278288 225649
rect 318352 225637 318358 225649
rect 318410 225637 318416 225689
rect 321712 225637 321718 225689
rect 321770 225677 321776 225689
rect 451216 225677 451222 225689
rect 321770 225649 451222 225677
rect 321770 225637 321776 225649
rect 451216 225637 451222 225649
rect 451274 225637 451280 225689
rect 244720 225563 244726 225615
rect 244778 225603 244784 225615
rect 254896 225603 254902 225615
rect 244778 225575 254902 225603
rect 244778 225563 244784 225575
rect 254896 225563 254902 225575
rect 254954 225563 254960 225615
rect 259024 225563 259030 225615
rect 259082 225603 259088 225615
rect 269968 225603 269974 225615
rect 259082 225575 269974 225603
rect 259082 225563 259088 225575
rect 269968 225563 269974 225575
rect 270026 225563 270032 225615
rect 273712 225563 273718 225615
rect 273770 225603 273776 225615
rect 309328 225603 309334 225615
rect 273770 225575 309334 225603
rect 273770 225563 273776 225575
rect 309328 225563 309334 225575
rect 309386 225563 309392 225615
rect 315760 225563 315766 225615
rect 315818 225603 315824 225615
rect 439120 225603 439126 225615
rect 315818 225575 439126 225603
rect 315818 225563 315824 225575
rect 439120 225563 439126 225575
rect 439178 225563 439184 225615
rect 273616 225489 273622 225541
rect 273674 225529 273680 225541
rect 303184 225529 303190 225541
rect 273674 225501 303190 225529
rect 273674 225489 273680 225501
rect 303184 225489 303190 225501
rect 303242 225489 303248 225541
rect 309904 225489 309910 225541
rect 309962 225529 309968 225541
rect 427024 225529 427030 225541
rect 309962 225501 427030 225529
rect 309962 225489 309968 225501
rect 427024 225489 427030 225501
rect 427082 225489 427088 225541
rect 306736 225415 306742 225467
rect 306794 225455 306800 225467
rect 420976 225455 420982 225467
rect 306794 225427 420982 225455
rect 306794 225415 306800 225427
rect 420976 225415 420982 225427
rect 421034 225415 421040 225467
rect 303856 225341 303862 225393
rect 303914 225381 303920 225393
rect 415024 225381 415030 225393
rect 303914 225353 415030 225381
rect 303914 225341 303920 225353
rect 415024 225341 415030 225353
rect 415082 225341 415088 225393
rect 302128 225267 302134 225319
rect 302186 225307 302192 225319
rect 411952 225307 411958 225319
rect 302186 225279 411958 225307
rect 302186 225267 302192 225279
rect 411952 225267 411958 225279
rect 412010 225267 412016 225319
rect 277072 225193 277078 225245
rect 277130 225233 277136 225245
rect 324400 225233 324406 225245
rect 277130 225205 324406 225233
rect 277130 225193 277136 225205
rect 324400 225193 324406 225205
rect 324458 225193 324464 225245
rect 351376 225193 351382 225245
rect 351434 225233 351440 225245
rect 418000 225233 418006 225245
rect 351434 225205 418006 225233
rect 351434 225193 351440 225205
rect 418000 225193 418006 225205
rect 418058 225193 418064 225245
rect 305104 225119 305110 225171
rect 305162 225159 305168 225171
rect 333520 225159 333526 225171
rect 305162 225131 333526 225159
rect 305162 225119 305168 225131
rect 333520 225119 333526 225131
rect 333578 225119 333584 225171
rect 339088 225119 339094 225171
rect 339146 225159 339152 225171
rect 399952 225159 399958 225171
rect 339146 225131 399958 225159
rect 339146 225119 339152 225131
rect 399952 225119 399958 225131
rect 400010 225119 400016 225171
rect 410416 225119 410422 225171
rect 410474 225159 410480 225171
rect 629392 225159 629398 225171
rect 410474 225131 629398 225159
rect 410474 225119 410480 225131
rect 629392 225119 629398 225131
rect 629450 225119 629456 225171
rect 252688 225045 252694 225097
rect 252746 225085 252752 225097
rect 312304 225085 312310 225097
rect 252746 225057 312310 225085
rect 252746 225045 252752 225057
rect 312304 225045 312310 225057
rect 312362 225045 312368 225097
rect 339760 225045 339766 225097
rect 339818 225085 339824 225097
rect 396784 225085 396790 225097
rect 339818 225057 396790 225085
rect 339818 225045 339824 225057
rect 396784 225045 396790 225057
rect 396842 225045 396848 225097
rect 408208 225085 408214 225097
rect 396898 225057 408214 225085
rect 272368 224971 272374 225023
rect 272426 225011 272432 225023
rect 336400 225011 336406 225023
rect 272426 224983 336406 225011
rect 272426 224971 272432 224983
rect 336400 224971 336406 224983
rect 336458 224971 336464 225023
rect 354352 224971 354358 225023
rect 354410 225011 354416 225023
rect 396898 225011 396926 225057
rect 408208 225045 408214 225057
rect 408266 225045 408272 225097
rect 405136 225011 405142 225023
rect 354410 224983 396926 225011
rect 396994 224983 405142 225011
rect 354410 224971 354416 224983
rect 348688 224897 348694 224949
rect 348746 224937 348752 224949
rect 394384 224937 394390 224949
rect 348746 224909 394390 224937
rect 348746 224897 348752 224909
rect 394384 224897 394390 224909
rect 394442 224897 394448 224949
rect 362800 224823 362806 224875
rect 362858 224863 362864 224875
rect 396994 224863 397022 224983
rect 405136 224971 405142 224983
rect 405194 224971 405200 225023
rect 402160 224863 402166 224875
rect 362858 224835 397022 224863
rect 397282 224835 402166 224863
rect 362858 224823 362864 224835
rect 147088 224749 147094 224801
rect 147146 224789 147152 224801
rect 151312 224789 151318 224801
rect 147146 224761 151318 224789
rect 147146 224749 147152 224761
rect 151312 224749 151318 224761
rect 151370 224749 151376 224801
rect 360304 224749 360310 224801
rect 360362 224789 360368 224801
rect 360362 224761 363902 224789
rect 360362 224749 360368 224761
rect 149488 224675 149494 224727
rect 149546 224715 149552 224727
rect 162736 224715 162742 224727
rect 149546 224687 162742 224715
rect 149546 224675 149552 224687
rect 162736 224675 162742 224687
rect 162794 224675 162800 224727
rect 277936 224675 277942 224727
rect 277994 224715 278000 224727
rect 363760 224715 363766 224727
rect 277994 224687 363766 224715
rect 277994 224675 278000 224687
rect 363760 224675 363766 224687
rect 363818 224675 363824 224727
rect 363874 224715 363902 224761
rect 367024 224749 367030 224801
rect 367082 224789 367088 224801
rect 376432 224789 376438 224801
rect 367082 224761 376438 224789
rect 367082 224749 367088 224761
rect 376432 224749 376438 224761
rect 376490 224749 376496 224801
rect 397282 224789 397310 224835
rect 402160 224823 402166 224835
rect 402218 224823 402224 224875
rect 397648 224789 397654 224801
rect 378658 224761 397310 224789
rect 397378 224761 397654 224789
rect 378658 224715 378686 224761
rect 363874 224687 378686 224715
rect 382192 224675 382198 224727
rect 382250 224715 382256 224727
rect 386320 224715 386326 224727
rect 382250 224687 386326 224715
rect 382250 224675 382256 224687
rect 386320 224675 386326 224687
rect 386378 224675 386384 224727
rect 386416 224675 386422 224727
rect 386474 224715 386480 224727
rect 397378 224715 397406 224761
rect 397648 224749 397654 224761
rect 397706 224749 397712 224801
rect 586288 224749 586294 224801
rect 586346 224789 586352 224801
rect 592336 224789 592342 224801
rect 586346 224761 592342 224789
rect 586346 224749 586352 224761
rect 592336 224749 592342 224761
rect 592394 224749 592400 224801
rect 386474 224687 397406 224715
rect 386474 224675 386480 224687
rect 397456 224675 397462 224727
rect 397514 224715 397520 224727
rect 400624 224715 400630 224727
rect 397514 224687 400630 224715
rect 397514 224675 397520 224687
rect 400624 224675 400630 224687
rect 400682 224675 400688 224727
rect 316336 224601 316342 224653
rect 316394 224641 316400 224653
rect 441424 224641 441430 224653
rect 316394 224613 441430 224641
rect 316394 224601 316400 224613
rect 441424 224601 441430 224613
rect 441482 224601 441488 224653
rect 323152 224527 323158 224579
rect 323210 224567 323216 224579
rect 452752 224567 452758 224579
rect 323210 224539 452758 224567
rect 323210 224527 323216 224539
rect 452752 224527 452758 224539
rect 452810 224527 452816 224579
rect 319312 224453 319318 224505
rect 319370 224493 319376 224505
rect 447472 224493 447478 224505
rect 319370 224465 447478 224493
rect 319370 224453 319376 224465
rect 447472 224453 447478 224465
rect 447530 224453 447536 224505
rect 322288 224379 322294 224431
rect 322346 224419 322352 224431
rect 453424 224419 453430 224431
rect 322346 224391 453430 224419
rect 322346 224379 322352 224391
rect 453424 224379 453430 224391
rect 453482 224379 453488 224431
rect 325360 224305 325366 224357
rect 325418 224345 325424 224357
rect 459568 224345 459574 224357
rect 325418 224317 459574 224345
rect 325418 224305 325424 224317
rect 459568 224305 459574 224317
rect 459626 224305 459632 224357
rect 328240 224231 328246 224283
rect 328298 224271 328304 224283
rect 465616 224271 465622 224283
rect 328298 224243 465622 224271
rect 328298 224231 328304 224243
rect 465616 224231 465622 224243
rect 465674 224231 465680 224283
rect 331504 224157 331510 224209
rect 331562 224197 331568 224209
rect 471568 224197 471574 224209
rect 331562 224169 471574 224197
rect 331562 224157 331568 224169
rect 471568 224157 471574 224169
rect 471626 224157 471632 224209
rect 334480 224083 334486 224135
rect 334538 224123 334544 224135
rect 477616 224123 477622 224135
rect 334538 224095 477622 224123
rect 334538 224083 334544 224095
rect 477616 224083 477622 224095
rect 477674 224083 477680 224135
rect 337168 224009 337174 224061
rect 337226 224049 337232 224061
rect 483760 224049 483766 224061
rect 337226 224021 483766 224049
rect 337226 224009 337232 224021
rect 483760 224009 483766 224021
rect 483818 224009 483824 224061
rect 340432 223935 340438 223987
rect 340490 223975 340496 223987
rect 489712 223975 489718 223987
rect 340490 223947 489718 223975
rect 340490 223935 340496 223947
rect 489712 223935 489718 223947
rect 489770 223935 489776 223987
rect 343600 223861 343606 223913
rect 343658 223901 343664 223913
rect 497296 223901 497302 223913
rect 343658 223873 497302 223901
rect 343658 223861 343664 223873
rect 497296 223861 497302 223873
rect 497354 223861 497360 223913
rect 261904 223787 261910 223839
rect 261962 223827 261968 223839
rect 332656 223827 332662 223839
rect 261962 223799 332662 223827
rect 261962 223787 261968 223799
rect 332656 223787 332662 223799
rect 332714 223787 332720 223839
rect 346576 223787 346582 223839
rect 346634 223827 346640 223839
rect 501808 223827 501814 223839
rect 346634 223799 501814 223827
rect 346634 223787 346640 223799
rect 501808 223787 501814 223799
rect 501866 223787 501872 223839
rect 263536 223713 263542 223765
rect 263594 223753 263600 223765
rect 335728 223753 335734 223765
rect 263594 223725 335734 223753
rect 263594 223713 263600 223725
rect 335728 223713 335734 223725
rect 335786 223713 335792 223765
rect 348112 223713 348118 223765
rect 348170 223753 348176 223765
rect 506320 223753 506326 223765
rect 348170 223725 506326 223753
rect 348170 223713 348176 223725
rect 506320 223713 506326 223725
rect 506378 223713 506384 223765
rect 266512 223639 266518 223691
rect 266570 223679 266576 223691
rect 341776 223679 341782 223691
rect 266570 223651 341782 223679
rect 266570 223639 266576 223651
rect 341776 223639 341782 223651
rect 341834 223639 341840 223691
rect 349552 223639 349558 223691
rect 349610 223679 349616 223691
rect 507856 223679 507862 223691
rect 349610 223651 507862 223679
rect 349610 223639 349616 223651
rect 507856 223639 507862 223651
rect 507914 223639 507920 223691
rect 264592 223565 264598 223617
rect 264650 223605 264656 223617
rect 338704 223605 338710 223617
rect 264650 223577 338710 223605
rect 264650 223565 264656 223577
rect 338704 223565 338710 223577
rect 338762 223565 338768 223617
rect 351184 223565 351190 223617
rect 351242 223605 351248 223617
rect 512368 223605 512374 223617
rect 351242 223577 512374 223605
rect 351242 223565 351248 223577
rect 512368 223565 512374 223577
rect 512426 223565 512432 223617
rect 268048 223491 268054 223543
rect 268106 223531 268112 223543
rect 344848 223531 344854 223543
rect 268106 223503 344854 223531
rect 268106 223491 268112 223503
rect 344848 223491 344854 223503
rect 344906 223491 344912 223543
rect 348016 223491 348022 223543
rect 348074 223531 348080 223543
rect 504784 223531 504790 223543
rect 348074 223503 504790 223531
rect 348074 223491 348080 223503
rect 504784 223491 504790 223503
rect 504842 223491 504848 223543
rect 270928 223417 270934 223469
rect 270986 223457 270992 223469
rect 350800 223457 350806 223469
rect 270986 223429 350806 223457
rect 270986 223417 270992 223429
rect 350800 223417 350806 223429
rect 350858 223417 350864 223469
rect 351088 223417 351094 223469
rect 351146 223457 351152 223469
rect 510832 223457 510838 223469
rect 351146 223429 510838 223457
rect 351146 223417 351152 223429
rect 510832 223417 510838 223429
rect 510890 223417 510896 223469
rect 269392 223343 269398 223395
rect 269450 223383 269456 223395
rect 347728 223383 347734 223395
rect 269450 223355 347734 223383
rect 269450 223343 269456 223355
rect 347728 223343 347734 223355
rect 347786 223343 347792 223395
rect 352528 223343 352534 223395
rect 352586 223383 352592 223395
rect 514000 223383 514006 223395
rect 352586 223355 514006 223383
rect 352586 223343 352592 223355
rect 514000 223343 514006 223355
rect 514058 223343 514064 223395
rect 355600 223269 355606 223321
rect 355658 223309 355664 223321
rect 519856 223309 519862 223321
rect 355658 223281 519862 223309
rect 355658 223269 355664 223281
rect 519856 223269 519862 223281
rect 519914 223269 519920 223321
rect 354064 223195 354070 223247
rect 354122 223235 354128 223247
rect 516976 223235 516982 223247
rect 354122 223207 516982 223235
rect 354122 223195 354128 223207
rect 516976 223195 516982 223207
rect 517034 223195 517040 223247
rect 318544 223121 318550 223173
rect 318602 223161 318608 223173
rect 443728 223161 443734 223173
rect 318602 223133 443734 223161
rect 318602 223121 318608 223133
rect 443728 223121 443734 223133
rect 443786 223121 443792 223173
rect 313360 223047 313366 223099
rect 313418 223087 313424 223099
rect 435376 223087 435382 223099
rect 313418 223059 435382 223087
rect 313418 223047 313424 223059
rect 435376 223047 435382 223059
rect 435434 223047 435440 223099
rect 310288 222973 310294 223025
rect 310346 223013 310352 223025
rect 429328 223013 429334 223025
rect 310346 222985 429334 223013
rect 310346 222973 310352 222985
rect 429328 222973 429334 222985
rect 429386 222973 429392 223025
rect 307984 222899 307990 222951
rect 308042 222939 308048 222951
rect 422512 222939 422518 222951
rect 308042 222911 422518 222939
rect 308042 222899 308048 222911
rect 422512 222899 422518 222911
rect 422570 222899 422576 222951
rect 312592 222825 312598 222877
rect 312650 222865 312656 222877
rect 431536 222865 431542 222877
rect 312650 222837 431542 222865
rect 312650 222825 312656 222837
rect 431536 222825 431542 222837
rect 431594 222825 431600 222877
rect 307216 222751 307222 222803
rect 307274 222791 307280 222803
rect 423280 222791 423286 222803
rect 307274 222763 423286 222791
rect 307274 222751 307280 222763
rect 423280 222751 423286 222763
rect 423338 222751 423344 222803
rect 304240 222677 304246 222729
rect 304298 222717 304304 222729
rect 417232 222717 417238 222729
rect 304298 222689 417238 222717
rect 304298 222677 304304 222689
rect 417232 222677 417238 222689
rect 417290 222677 417296 222729
rect 302800 222603 302806 222655
rect 302858 222643 302864 222655
rect 414256 222643 414262 222655
rect 302858 222615 414262 222643
rect 302858 222603 302864 222615
rect 414256 222603 414262 222615
rect 414314 222603 414320 222655
rect 304912 222529 304918 222581
rect 304970 222569 304976 222581
rect 416464 222569 416470 222581
rect 304970 222541 416470 222569
rect 304970 222529 304976 222541
rect 416464 222529 416470 222541
rect 416522 222529 416528 222581
rect 286192 222455 286198 222507
rect 286250 222495 286256 222507
rect 381040 222495 381046 222507
rect 286250 222467 381046 222495
rect 286250 222455 286256 222467
rect 381040 222455 381046 222467
rect 381098 222455 381104 222507
rect 396976 222455 396982 222507
rect 397034 222495 397040 222507
rect 496528 222495 496534 222507
rect 397034 222467 496534 222495
rect 397034 222455 397040 222467
rect 496528 222455 496534 222467
rect 496586 222455 496592 222507
rect 272560 222381 272566 222433
rect 272618 222421 272624 222433
rect 353872 222421 353878 222433
rect 272618 222393 353878 222421
rect 272618 222381 272624 222393
rect 353872 222381 353878 222393
rect 353930 222381 353936 222433
rect 371632 222381 371638 222433
rect 371690 222421 371696 222433
rect 467824 222421 467830 222433
rect 371690 222393 467830 222421
rect 371690 222381 371696 222393
rect 467824 222381 467830 222393
rect 467882 222381 467888 222433
rect 283120 222307 283126 222359
rect 283178 222347 283184 222359
rect 374992 222347 374998 222359
rect 283178 222319 374998 222347
rect 283178 222307 283184 222319
rect 374992 222307 374998 222319
rect 375050 222307 375056 222359
rect 386800 222307 386806 222359
rect 386858 222347 386864 222359
rect 482896 222347 482902 222359
rect 386858 222319 482902 222347
rect 386858 222307 386864 222319
rect 482896 222307 482902 222319
rect 482954 222307 482960 222359
rect 281584 222233 281590 222285
rect 281642 222273 281648 222285
rect 371920 222273 371926 222285
rect 281642 222245 371926 222273
rect 281642 222233 281648 222245
rect 371920 222233 371926 222245
rect 371978 222233 371984 222285
rect 394384 222233 394390 222285
rect 394442 222273 394448 222285
rect 399088 222273 399094 222285
rect 394442 222245 399094 222273
rect 394442 222233 394448 222245
rect 399088 222233 399094 222245
rect 399146 222233 399152 222285
rect 274096 222159 274102 222211
rect 274154 222199 274160 222211
rect 356848 222199 356854 222211
rect 274154 222171 356854 222199
rect 274154 222159 274160 222171
rect 356848 222159 356854 222171
rect 356906 222159 356912 222211
rect 149392 221863 149398 221915
rect 149450 221903 149456 221915
rect 168400 221903 168406 221915
rect 149450 221875 168406 221903
rect 149450 221863 149456 221875
rect 168400 221863 168406 221875
rect 168458 221863 168464 221915
rect 149488 221789 149494 221841
rect 149546 221829 149552 221841
rect 171376 221829 171382 221841
rect 149546 221801 171382 221829
rect 149546 221789 149552 221801
rect 171376 221789 171382 221801
rect 171434 221789 171440 221841
rect 656176 221789 656182 221841
rect 656234 221829 656240 221841
rect 676240 221829 676246 221841
rect 656234 221801 676246 221829
rect 656234 221789 656240 221801
rect 676240 221789 676246 221801
rect 676298 221789 676304 221841
rect 42064 221715 42070 221767
rect 42122 221755 42128 221767
rect 50320 221755 50326 221767
rect 42122 221727 50326 221755
rect 42122 221715 42128 221727
rect 50320 221715 50326 221727
rect 50378 221715 50384 221767
rect 145744 221715 145750 221767
rect 145802 221755 145808 221767
rect 184336 221755 184342 221767
rect 145802 221727 184342 221755
rect 145802 221715 145808 221727
rect 184336 221715 184342 221727
rect 184394 221715 184400 221767
rect 276400 221715 276406 221767
rect 276458 221755 276464 221767
rect 277552 221755 277558 221767
rect 276458 221727 277558 221755
rect 276458 221715 276464 221727
rect 277552 221715 277558 221727
rect 277610 221715 277616 221767
rect 478480 221715 478486 221767
rect 478538 221755 478544 221767
rect 479968 221755 479974 221767
rect 478538 221727 479974 221755
rect 478538 221715 478544 221727
rect 479968 221715 479974 221727
rect 480026 221715 480032 221767
rect 513808 221715 513814 221767
rect 513866 221755 513872 221767
rect 515392 221755 515398 221767
rect 513866 221727 515398 221755
rect 513866 221715 513872 221727
rect 515392 221715 515398 221727
rect 515450 221715 515456 221767
rect 147280 220753 147286 220805
rect 147338 220793 147344 220805
rect 151408 220793 151414 220805
rect 147338 220765 151414 220793
rect 147338 220753 147344 220765
rect 151408 220753 151414 220765
rect 151466 220753 151472 220805
rect 673264 220605 673270 220657
rect 673322 220645 673328 220657
rect 676048 220645 676054 220657
rect 673322 220617 676054 220645
rect 673322 220605 673328 220617
rect 676048 220605 676054 220617
rect 676106 220605 676112 220657
rect 673360 219495 673366 219547
rect 673418 219535 673424 219547
rect 676048 219535 676054 219547
rect 673418 219507 676054 219535
rect 673418 219495 673424 219507
rect 676048 219495 676054 219507
rect 676106 219495 676112 219547
rect 655984 219199 655990 219251
rect 656042 219239 656048 219251
rect 676240 219239 676246 219251
rect 656042 219211 676246 219239
rect 656042 219199 656048 219211
rect 676240 219199 676246 219211
rect 676298 219199 676304 219251
rect 655792 219051 655798 219103
rect 655850 219091 655856 219103
rect 676144 219091 676150 219103
rect 655850 219063 676150 219091
rect 655850 219051 655856 219063
rect 676144 219051 676150 219063
rect 676202 219051 676208 219103
rect 149488 218977 149494 219029
rect 149546 219017 149552 219029
rect 165616 219017 165622 219029
rect 149546 218989 165622 219017
rect 149546 218977 149552 218989
rect 165616 218977 165622 218989
rect 165674 218977 165680 219029
rect 149392 218903 149398 218955
rect 149450 218943 149456 218955
rect 179920 218943 179926 218955
rect 149450 218915 179926 218943
rect 149450 218903 149456 218915
rect 179920 218903 179926 218915
rect 179978 218903 179984 218955
rect 143056 218829 143062 218881
rect 143114 218869 143120 218881
rect 184336 218869 184342 218881
rect 143114 218841 184342 218869
rect 143114 218829 143120 218841
rect 184336 218829 184342 218841
rect 184394 218829 184400 218881
rect 149488 216091 149494 216143
rect 149546 216131 149552 216143
rect 174352 216131 174358 216143
rect 149546 216103 174358 216131
rect 149546 216091 149552 216103
rect 174352 216091 174358 216103
rect 174410 216091 174416 216143
rect 149392 216017 149398 216069
rect 149450 216057 149456 216069
rect 177136 216057 177142 216069
rect 149450 216029 177142 216057
rect 149450 216017 149456 216029
rect 177136 216017 177142 216029
rect 177194 216017 177200 216069
rect 149392 214685 149398 214737
rect 149450 214725 149456 214737
rect 159952 214725 159958 214737
rect 149450 214697 159958 214725
rect 149450 214685 149456 214697
rect 159952 214685 159958 214697
rect 160010 214685 160016 214737
rect 147280 214019 147286 214071
rect 147338 214059 147344 214071
rect 151792 214059 151798 214071
rect 147338 214031 151798 214059
rect 147338 214019 147344 214031
rect 151792 214019 151798 214031
rect 151850 214019 151856 214071
rect 41776 213279 41782 213331
rect 41834 213319 41840 213331
rect 45712 213319 45718 213331
rect 41834 213291 45718 213319
rect 41834 213279 41840 213291
rect 45712 213279 45718 213291
rect 45770 213279 45776 213331
rect 675088 213205 675094 213257
rect 675146 213245 675152 213257
rect 675952 213245 675958 213257
rect 675146 213217 675958 213245
rect 675146 213205 675152 213217
rect 675952 213205 675958 213217
rect 676010 213205 676016 213257
rect 675280 213131 675286 213183
rect 675338 213171 675344 213183
rect 676048 213171 676054 213183
rect 675338 213143 676054 213171
rect 675338 213131 675344 213143
rect 676048 213131 676054 213143
rect 676106 213131 676112 213183
rect 41584 212909 41590 212961
rect 41642 212949 41648 212961
rect 45616 212949 45622 212961
rect 41642 212921 45622 212949
rect 41642 212909 41648 212921
rect 45616 212909 45622 212921
rect 45674 212909 45680 212961
rect 146896 212835 146902 212887
rect 146954 212875 146960 212887
rect 152080 212875 152086 212887
rect 146954 212847 152086 212875
rect 146954 212835 146960 212847
rect 152080 212835 152086 212847
rect 152138 212835 152144 212887
rect 41776 212169 41782 212221
rect 41834 212209 41840 212221
rect 45520 212209 45526 212221
rect 41834 212181 45526 212209
rect 41834 212169 41840 212181
rect 45520 212169 45526 212181
rect 45578 212169 45584 212221
rect 674704 212095 674710 212147
rect 674762 212135 674768 212147
rect 676048 212135 676054 212147
rect 674762 212107 676054 212135
rect 674762 212095 674768 212107
rect 676048 212095 676054 212107
rect 676106 212095 676112 212147
rect 41776 211725 41782 211777
rect 41834 211765 41840 211777
rect 43408 211765 43414 211777
rect 41834 211737 43414 211765
rect 41834 211725 41840 211737
rect 43408 211725 43414 211737
rect 43466 211725 43472 211777
rect 41584 211429 41590 211481
rect 41642 211469 41648 211481
rect 44848 211469 44854 211481
rect 41642 211441 44854 211469
rect 41642 211429 41648 211441
rect 44848 211429 44854 211441
rect 44906 211429 44912 211481
rect 147088 211281 147094 211333
rect 147146 211321 147152 211333
rect 151696 211321 151702 211333
rect 147146 211293 151702 211321
rect 147146 211281 147152 211293
rect 151696 211281 151702 211293
rect 151754 211281 151760 211333
rect 41776 210689 41782 210741
rect 41834 210729 41840 210741
rect 50608 210729 50614 210741
rect 41834 210701 50614 210729
rect 41834 210689 41840 210701
rect 50608 210689 50614 210701
rect 50666 210689 50672 210741
rect 674800 210393 674806 210445
rect 674858 210433 674864 210445
rect 675952 210433 675958 210445
rect 674858 210405 675958 210433
rect 674858 210393 674864 210405
rect 675952 210393 675958 210405
rect 676010 210393 676016 210445
rect 147472 210319 147478 210371
rect 147530 210359 147536 210371
rect 151600 210359 151606 210371
rect 147530 210331 151606 210359
rect 147530 210319 147536 210331
rect 151600 210319 151606 210331
rect 151658 210319 151664 210371
rect 674896 210319 674902 210371
rect 674954 210359 674960 210371
rect 676240 210359 676246 210371
rect 674954 210331 676246 210359
rect 674954 210319 674960 210331
rect 676240 210319 676246 210331
rect 676298 210319 676304 210371
rect 674992 210245 674998 210297
rect 675050 210285 675056 210297
rect 676048 210285 676054 210297
rect 675050 210257 676054 210285
rect 675050 210245 675056 210257
rect 676048 210245 676054 210257
rect 676106 210245 676112 210297
rect 41776 210171 41782 210223
rect 41834 210211 41840 210223
rect 43312 210211 43318 210223
rect 41834 210183 43318 210211
rect 41834 210171 41840 210183
rect 43312 210171 43318 210183
rect 43370 210171 43376 210223
rect 41584 209949 41590 210001
rect 41642 209989 41648 210001
rect 50416 209989 50422 210001
rect 41642 209961 50422 209989
rect 41642 209949 41648 209961
rect 50416 209949 50422 209961
rect 50474 209949 50480 210001
rect 41584 209357 41590 209409
rect 41642 209397 41648 209409
rect 43504 209397 43510 209409
rect 41642 209369 43510 209397
rect 41642 209357 41648 209369
rect 43504 209357 43510 209369
rect 43562 209357 43568 209409
rect 147184 207877 147190 207929
rect 147242 207917 147248 207929
rect 151504 207917 151510 207929
rect 147242 207889 151510 207917
rect 147242 207877 147248 207889
rect 151504 207877 151510 207889
rect 151562 207877 151568 207929
rect 146896 207359 146902 207411
rect 146954 207399 146960 207411
rect 151984 207399 151990 207411
rect 146954 207371 151990 207399
rect 146954 207359 146960 207371
rect 151984 207359 151990 207371
rect 152042 207359 152048 207411
rect 646768 207359 646774 207411
rect 646826 207399 646832 207411
rect 679792 207399 679798 207411
rect 646826 207371 679798 207399
rect 646826 207359 646832 207371
rect 679792 207359 679798 207371
rect 679850 207359 679856 207411
rect 675760 206101 675766 206153
rect 675818 206101 675824 206153
rect 675088 205657 675094 205709
rect 675146 205697 675152 205709
rect 675472 205697 675478 205709
rect 675146 205669 675478 205697
rect 675146 205657 675152 205669
rect 675472 205657 675478 205669
rect 675530 205657 675536 205709
rect 675778 205635 675806 206101
rect 675760 205583 675766 205635
rect 675818 205583 675824 205635
rect 147088 204547 147094 204599
rect 147146 204587 147152 204599
rect 151888 204587 151894 204599
rect 147146 204559 151894 204587
rect 147146 204547 147152 204559
rect 151888 204547 151894 204559
rect 151946 204547 151952 204599
rect 149392 204473 149398 204525
rect 149450 204513 149456 204525
rect 182992 204513 182998 204525
rect 149450 204485 182998 204513
rect 149450 204473 149456 204485
rect 182992 204473 182998 204485
rect 183050 204473 183056 204525
rect 675184 201883 675190 201935
rect 675242 201923 675248 201935
rect 675472 201923 675478 201935
rect 675242 201895 675478 201923
rect 675242 201883 675248 201895
rect 675472 201883 675478 201895
rect 675530 201883 675536 201935
rect 149392 201735 149398 201787
rect 149450 201775 149456 201787
rect 174448 201775 174454 201787
rect 149450 201747 174454 201775
rect 149450 201735 149456 201747
rect 174448 201735 174454 201747
rect 174506 201735 174512 201787
rect 41872 201661 41878 201713
rect 41930 201701 41936 201713
rect 44752 201701 44758 201713
rect 41930 201673 44758 201701
rect 41930 201661 41936 201673
rect 44752 201661 44758 201673
rect 44810 201661 44816 201713
rect 149488 201661 149494 201713
rect 149546 201701 149552 201713
rect 177232 201701 177238 201713
rect 149546 201673 177238 201701
rect 149546 201661 149552 201673
rect 177232 201661 177238 201673
rect 177290 201661 177296 201713
rect 149296 201587 149302 201639
rect 149354 201627 149360 201639
rect 180112 201627 180118 201639
rect 149354 201599 180118 201627
rect 149354 201587 149360 201599
rect 180112 201587 180118 201599
rect 180170 201587 180176 201639
rect 143056 201513 143062 201565
rect 143114 201553 143120 201565
rect 184336 201553 184342 201565
rect 143114 201525 184342 201553
rect 143114 201513 143120 201525
rect 184336 201513 184342 201525
rect 184394 201513 184400 201565
rect 655600 201513 655606 201565
rect 655658 201553 655664 201565
rect 675088 201553 675094 201565
rect 655658 201525 675094 201553
rect 655658 201513 655664 201525
rect 675088 201513 675094 201525
rect 675146 201513 675152 201565
rect 41488 201439 41494 201491
rect 41546 201479 41552 201491
rect 42928 201479 42934 201491
rect 41546 201451 42934 201479
rect 41546 201439 41552 201451
rect 42928 201439 42934 201451
rect 42986 201439 42992 201491
rect 41872 201365 41878 201417
rect 41930 201405 41936 201417
rect 44560 201405 44566 201417
rect 41930 201377 44566 201405
rect 41930 201365 41936 201377
rect 44560 201365 44566 201377
rect 44618 201365 44624 201417
rect 41488 200921 41494 200973
rect 41546 200961 41552 200973
rect 44656 200961 44662 200973
rect 41546 200933 44662 200961
rect 41546 200921 41552 200933
rect 44656 200921 44662 200933
rect 44714 200921 44720 200973
rect 674992 200847 674998 200899
rect 675050 200887 675056 200899
rect 675376 200887 675382 200899
rect 675050 200859 675382 200887
rect 675050 200847 675056 200859
rect 675376 200847 675382 200859
rect 675434 200847 675440 200899
rect 41584 198923 41590 198975
rect 41642 198963 41648 198975
rect 42736 198963 42742 198975
rect 41642 198935 42742 198963
rect 41642 198923 41648 198935
rect 42736 198923 42742 198935
rect 42794 198923 42800 198975
rect 41680 198849 41686 198901
rect 41738 198889 41744 198901
rect 42832 198889 42838 198901
rect 41738 198861 42838 198889
rect 41738 198849 41744 198861
rect 42832 198849 42838 198861
rect 42890 198849 42896 198901
rect 41776 198775 41782 198827
rect 41834 198815 41840 198827
rect 43024 198815 43030 198827
rect 41834 198787 43030 198815
rect 41834 198775 41840 198787
rect 43024 198775 43030 198787
rect 43082 198775 43088 198827
rect 147472 198775 147478 198827
rect 147530 198815 147536 198827
rect 154192 198815 154198 198827
rect 147530 198787 154198 198815
rect 147530 198775 147536 198787
rect 154192 198775 154198 198787
rect 154250 198775 154256 198827
rect 149392 198701 149398 198753
rect 149450 198741 149456 198753
rect 162832 198741 162838 198753
rect 149450 198713 162838 198741
rect 149450 198701 149456 198713
rect 162832 198701 162838 198713
rect 162890 198701 162896 198753
rect 181360 198627 181366 198679
rect 181418 198667 181424 198679
rect 184432 198667 184438 198679
rect 181418 198639 184438 198667
rect 181418 198627 181424 198639
rect 184432 198627 184438 198639
rect 184490 198627 184496 198679
rect 178288 198553 178294 198605
rect 178346 198593 178352 198605
rect 184336 198593 184342 198605
rect 178346 198565 184342 198593
rect 178346 198553 178352 198565
rect 184336 198553 184342 198565
rect 184394 198553 184400 198605
rect 674896 197739 674902 197791
rect 674954 197779 674960 197791
rect 675376 197779 675382 197791
rect 674954 197751 675382 197779
rect 674954 197739 674960 197751
rect 675376 197739 675382 197751
rect 675434 197739 675440 197791
rect 41968 197369 41974 197421
rect 42026 197369 42032 197421
rect 41986 197199 42014 197369
rect 41968 197147 41974 197199
rect 42026 197147 42032 197199
rect 674704 196999 674710 197051
rect 674762 197039 674768 197051
rect 675472 197039 675478 197051
rect 674762 197011 675478 197039
rect 674762 196999 674768 197011
rect 675472 196999 675478 197011
rect 675530 196999 675536 197051
rect 674800 196555 674806 196607
rect 674858 196595 674864 196607
rect 675376 196595 675382 196607
rect 674858 196567 675382 196595
rect 674858 196555 674864 196567
rect 675376 196555 675382 196567
rect 675434 196555 675440 196607
rect 149392 195963 149398 196015
rect 149450 196003 149456 196015
rect 168592 196003 168598 196015
rect 149450 195975 168598 196003
rect 149450 195963 149456 195975
rect 168592 195963 168598 195975
rect 168650 195963 168656 196015
rect 149488 195889 149494 195941
rect 149546 195929 149552 195941
rect 171568 195929 171574 195941
rect 149546 195901 171574 195929
rect 149546 195889 149552 195901
rect 171568 195889 171574 195901
rect 171626 195889 171632 195941
rect 149392 195815 149398 195867
rect 149450 195855 149456 195867
rect 183088 195855 183094 195867
rect 149450 195827 183094 195855
rect 149450 195815 149456 195827
rect 183088 195815 183094 195827
rect 183146 195815 183152 195867
rect 166960 195741 166966 195793
rect 167018 195781 167024 195793
rect 184528 195781 184534 195793
rect 167018 195753 184534 195781
rect 167018 195741 167024 195753
rect 184528 195741 184534 195753
rect 184586 195741 184592 195793
rect 169840 195667 169846 195719
rect 169898 195707 169904 195719
rect 184432 195707 184438 195719
rect 169898 195679 184438 195707
rect 169898 195667 169904 195679
rect 184432 195667 184438 195679
rect 184490 195667 184496 195719
rect 172720 195593 172726 195645
rect 172778 195633 172784 195645
rect 184336 195633 184342 195645
rect 172778 195605 184342 195633
rect 172778 195593 172784 195605
rect 184336 195593 184342 195605
rect 184394 195593 184400 195645
rect 42064 193447 42070 193499
rect 42122 193487 42128 193499
rect 42832 193487 42838 193499
rect 42122 193459 42838 193487
rect 42122 193447 42128 193459
rect 42832 193447 42838 193459
rect 42890 193447 42896 193499
rect 149392 193151 149398 193203
rect 149450 193191 149456 193203
rect 160048 193191 160054 193203
rect 149450 193163 160054 193191
rect 149450 193151 149456 193163
rect 160048 193151 160054 193163
rect 160106 193151 160112 193203
rect 149488 193003 149494 193055
rect 149546 193043 149552 193055
rect 165808 193043 165814 193055
rect 149546 193015 165814 193043
rect 149546 193003 149552 193015
rect 165808 193003 165814 193015
rect 165866 193003 165872 193055
rect 152368 192929 152374 192981
rect 152426 192969 152432 192981
rect 184624 192969 184630 192981
rect 152426 192941 184630 192969
rect 152426 192929 152432 192941
rect 184624 192929 184630 192941
rect 184682 192929 184688 192981
rect 155440 192855 155446 192907
rect 155498 192895 155504 192907
rect 184528 192895 184534 192907
rect 155498 192867 184534 192895
rect 155498 192855 155504 192867
rect 184528 192855 184534 192867
rect 184586 192855 184592 192907
rect 158128 192781 158134 192833
rect 158186 192821 158192 192833
rect 184336 192821 184342 192833
rect 158186 192793 184342 192821
rect 158186 192781 158192 192793
rect 184336 192781 184342 192793
rect 184394 192781 184400 192833
rect 163888 192707 163894 192759
rect 163946 192747 163952 192759
rect 184432 192747 184438 192759
rect 163946 192719 184438 192747
rect 163946 192707 163952 192719
rect 184432 192707 184438 192719
rect 184490 192707 184496 192759
rect 42160 192189 42166 192241
rect 42218 192229 42224 192241
rect 42736 192229 42742 192241
rect 42218 192201 42742 192229
rect 42218 192189 42224 192201
rect 42736 192189 42742 192201
rect 42794 192189 42800 192241
rect 42064 191449 42070 191501
rect 42122 191489 42128 191501
rect 43024 191489 43030 191501
rect 42122 191461 43030 191489
rect 42122 191449 42128 191461
rect 43024 191449 43030 191461
rect 43082 191449 43088 191501
rect 42160 191005 42166 191057
rect 42218 191045 42224 191057
rect 42928 191045 42934 191057
rect 42218 191017 42934 191045
rect 42218 191005 42224 191017
rect 42928 191005 42934 191017
rect 42986 191005 42992 191057
rect 147376 190191 147382 190243
rect 147434 190231 147440 190243
rect 154288 190231 154294 190243
rect 147434 190203 154294 190231
rect 147434 190191 147440 190203
rect 154288 190191 154294 190203
rect 154346 190191 154352 190243
rect 149392 190117 149398 190169
rect 149450 190157 149456 190169
rect 157072 190157 157078 190169
rect 149450 190129 157078 190157
rect 149450 190117 149456 190129
rect 157072 190117 157078 190129
rect 157130 190117 157136 190169
rect 143920 190043 143926 190095
rect 143978 190083 143984 190095
rect 184528 190083 184534 190095
rect 143978 190055 184534 190083
rect 143978 190043 143984 190055
rect 184528 190043 184534 190055
rect 184586 190043 184592 190095
rect 149680 189969 149686 190021
rect 149738 190009 149744 190021
rect 184336 190009 184342 190021
rect 149738 189981 184342 190009
rect 149738 189969 149744 189981
rect 184336 189969 184342 189981
rect 184394 189969 184400 190021
rect 171472 189895 171478 189947
rect 171530 189935 171536 189947
rect 184432 189935 184438 189947
rect 171530 189907 184438 189935
rect 171530 189895 171536 189907
rect 184432 189895 184438 189907
rect 184490 189895 184496 189947
rect 180016 189821 180022 189873
rect 180074 189861 180080 189873
rect 184336 189861 184342 189873
rect 180074 189833 184342 189861
rect 180074 189821 180080 189833
rect 184336 189821 184342 189833
rect 184394 189821 184400 189873
rect 159856 187157 159862 187209
rect 159914 187197 159920 187209
rect 184432 187197 184438 187209
rect 159914 187169 184438 187197
rect 159914 187157 159920 187169
rect 184432 187157 184438 187169
rect 184490 187157 184496 187209
rect 165712 187083 165718 187135
rect 165770 187123 165776 187135
rect 184528 187123 184534 187135
rect 165770 187095 184534 187123
rect 165770 187083 165776 187095
rect 184528 187083 184534 187095
rect 184586 187083 184592 187135
rect 168496 187009 168502 187061
rect 168554 187049 168560 187061
rect 184336 187049 184342 187061
rect 168554 187021 184342 187049
rect 168554 187009 168560 187021
rect 184336 187009 184342 187021
rect 184394 187009 184400 187061
rect 177040 186935 177046 186987
rect 177098 186975 177104 186987
rect 184624 186975 184630 186987
rect 177098 186947 184630 186975
rect 177098 186935 177104 186947
rect 184624 186935 184630 186947
rect 184682 186935 184688 186987
rect 149392 185751 149398 185803
rect 149450 185791 149456 185803
rect 185968 185791 185974 185803
rect 149450 185763 185974 185791
rect 149450 185751 149456 185763
rect 185968 185751 185974 185763
rect 186026 185751 186032 185803
rect 145648 184271 145654 184323
rect 145706 184311 145712 184323
rect 184336 184311 184342 184323
rect 145706 184283 184342 184311
rect 145706 184271 145712 184283
rect 184336 184271 184342 184283
rect 184394 184271 184400 184323
rect 171280 184197 171286 184249
rect 171338 184237 171344 184249
rect 184432 184237 184438 184249
rect 171338 184209 184438 184237
rect 171338 184197 171344 184209
rect 184432 184197 184438 184209
rect 184490 184197 184496 184249
rect 182896 184123 182902 184175
rect 182954 184163 182960 184175
rect 186736 184163 186742 184175
rect 182954 184135 186742 184163
rect 182954 184123 182960 184135
rect 186736 184123 186742 184135
rect 186794 184123 186800 184175
rect 645136 183087 645142 183139
rect 645194 183127 645200 183139
rect 649360 183127 649366 183139
rect 645194 183099 649366 183127
rect 645194 183087 645200 183099
rect 649360 183087 649366 183099
rect 649418 183087 649424 183139
rect 149296 182939 149302 182991
rect 149354 182979 149360 182991
rect 186256 182979 186262 182991
rect 149354 182951 186262 182979
rect 149354 182939 149360 182951
rect 186256 182939 186262 182951
rect 186314 182939 186320 182991
rect 149488 182865 149494 182917
rect 149546 182905 149552 182917
rect 186064 182905 186070 182917
rect 149546 182877 186070 182905
rect 149546 182865 149552 182877
rect 186064 182865 186070 182877
rect 186122 182865 186128 182917
rect 42160 182199 42166 182251
rect 42218 182239 42224 182251
rect 48112 182239 48118 182251
rect 42218 182211 48118 182239
rect 42218 182199 42224 182211
rect 48112 182199 48118 182211
rect 48170 182199 48176 182251
rect 149392 181459 149398 181511
rect 149450 181499 149456 181511
rect 171472 181499 171478 181511
rect 149450 181471 171478 181499
rect 149450 181459 149456 181471
rect 171472 181459 171478 181471
rect 171530 181459 171536 181511
rect 182800 181385 182806 181437
rect 182858 181425 182864 181437
rect 184624 181425 184630 181437
rect 182858 181397 184630 181425
rect 182858 181385 182864 181397
rect 184624 181385 184630 181397
rect 184682 181385 184688 181437
rect 156880 181311 156886 181363
rect 156938 181351 156944 181363
rect 184336 181351 184342 181363
rect 156938 181323 184342 181351
rect 156938 181311 156944 181323
rect 184336 181311 184342 181323
rect 184394 181311 184400 181363
rect 165520 181237 165526 181289
rect 165578 181277 165584 181289
rect 184432 181277 184438 181289
rect 165578 181249 184438 181277
rect 165578 181237 165584 181249
rect 184432 181237 184438 181249
rect 184490 181237 184496 181289
rect 154000 181163 154006 181215
rect 154058 181203 154064 181215
rect 184528 181203 184534 181215
rect 154058 181175 184534 181203
rect 154058 181163 154064 181175
rect 184528 181163 184534 181175
rect 184586 181163 184592 181215
rect 149584 180053 149590 180105
rect 149642 180093 149648 180105
rect 185488 180093 185494 180105
rect 149642 180065 185494 180093
rect 149642 180053 149648 180065
rect 185488 180053 185494 180065
rect 185546 180053 185552 180105
rect 149200 179979 149206 180031
rect 149258 180019 149264 180031
rect 186448 180019 186454 180031
rect 149258 179991 186454 180019
rect 149258 179979 149264 179991
rect 186448 179979 186454 179991
rect 186506 179979 186512 180031
rect 645136 179387 645142 179439
rect 645194 179427 645200 179439
rect 649456 179427 649462 179439
rect 645194 179399 649462 179427
rect 645194 179387 645200 179399
rect 649456 179387 649462 179399
rect 649514 179387 649520 179439
rect 149392 178721 149398 178773
rect 149450 178761 149456 178773
rect 162928 178761 162934 178773
rect 149450 178733 162934 178761
rect 149450 178721 149456 178733
rect 162928 178721 162934 178733
rect 162986 178721 162992 178773
rect 149488 178647 149494 178699
rect 149546 178687 149552 178699
rect 165712 178687 165718 178699
rect 149546 178659 165718 178687
rect 149546 178647 149552 178659
rect 165712 178647 165718 178659
rect 165770 178647 165776 178699
rect 149296 178573 149302 178625
rect 149354 178613 149360 178625
rect 168496 178613 168502 178625
rect 149354 178585 168502 178613
rect 149354 178573 149360 178585
rect 168496 178573 168502 178585
rect 168554 178573 168560 178625
rect 145456 178499 145462 178551
rect 145514 178539 145520 178551
rect 184432 178539 184438 178551
rect 145514 178511 184438 178539
rect 145514 178499 145520 178511
rect 184432 178499 184438 178511
rect 184490 178499 184496 178551
rect 162640 178425 162646 178477
rect 162698 178465 162704 178477
rect 184528 178465 184534 178477
rect 162698 178437 184534 178465
rect 162698 178425 162704 178437
rect 184528 178425 184534 178437
rect 184586 178425 184592 178477
rect 174160 178351 174166 178403
rect 174218 178391 174224 178403
rect 184336 178391 184342 178403
rect 174218 178363 184342 178391
rect 174218 178351 174224 178363
rect 184336 178351 184342 178363
rect 184394 178351 184400 178403
rect 149392 177241 149398 177293
rect 149450 177281 149456 177293
rect 156880 177281 156886 177293
rect 149450 177253 156886 177281
rect 149450 177241 149456 177253
rect 156880 177241 156886 177253
rect 156938 177241 156944 177293
rect 655696 176131 655702 176183
rect 655754 176171 655760 176183
rect 676240 176171 676246 176183
rect 655754 176143 676246 176171
rect 655754 176131 655760 176143
rect 676240 176131 676246 176143
rect 676298 176131 676304 176183
rect 147760 175983 147766 176035
rect 147818 176023 147824 176035
rect 154000 176023 154006 176035
rect 147818 175995 154006 176023
rect 147818 175983 147824 175995
rect 154000 175983 154006 175995
rect 154058 175983 154064 176035
rect 655504 175983 655510 176035
rect 655562 176023 655568 176035
rect 676336 176023 676342 176035
rect 655562 175995 676342 176023
rect 655562 175983 655568 175995
rect 676336 175983 676342 175995
rect 676394 175983 676400 176035
rect 655408 175835 655414 175887
rect 655466 175875 655472 175887
rect 676144 175875 676150 175887
rect 655466 175847 676150 175875
rect 655466 175835 655472 175847
rect 676144 175835 676150 175847
rect 676202 175835 676208 175887
rect 145360 175613 145366 175665
rect 145418 175653 145424 175665
rect 184336 175653 184342 175665
rect 145418 175625 184342 175653
rect 145418 175613 145424 175625
rect 184336 175613 184342 175625
rect 184394 175613 184400 175665
rect 145552 175539 145558 175591
rect 145610 175579 145616 175591
rect 184432 175579 184438 175591
rect 145610 175551 184438 175579
rect 145610 175539 145616 175551
rect 184432 175539 184438 175551
rect 184490 175539 184496 175591
rect 645136 174873 645142 174925
rect 645194 174913 645200 174925
rect 649552 174913 649558 174925
rect 645194 174885 649558 174913
rect 645194 174873 645200 174885
rect 649552 174873 649558 174885
rect 649610 174873 649616 174925
rect 149200 174207 149206 174259
rect 149258 174247 149264 174259
rect 186160 174247 186166 174259
rect 149258 174219 186166 174247
rect 149258 174207 149264 174219
rect 186160 174207 186166 174219
rect 186218 174207 186224 174259
rect 149392 172801 149398 172853
rect 149450 172841 149456 172853
rect 182800 172841 182806 172853
rect 149450 172813 182806 172841
rect 149450 172801 149456 172813
rect 182800 172801 182806 172813
rect 182858 172801 182864 172853
rect 148336 172727 148342 172779
rect 148394 172767 148400 172779
rect 184528 172767 184534 172779
rect 148394 172739 184534 172767
rect 148394 172727 148400 172739
rect 184528 172727 184534 172739
rect 184586 172727 184592 172779
rect 149008 172653 149014 172705
rect 149066 172693 149072 172705
rect 184624 172693 184630 172705
rect 149066 172665 184630 172693
rect 149066 172653 149072 172665
rect 184624 172653 184630 172665
rect 184682 172653 184688 172705
rect 148720 172579 148726 172631
rect 148778 172619 148784 172631
rect 184336 172619 184342 172631
rect 148778 172591 184342 172619
rect 148778 172579 148784 172591
rect 184336 172579 184342 172591
rect 184394 172579 184400 172631
rect 148528 172505 148534 172557
rect 148586 172545 148592 172557
rect 184432 172545 184438 172557
rect 148586 172517 184438 172545
rect 148586 172505 148592 172517
rect 184432 172505 184438 172517
rect 184490 172505 184496 172557
rect 645136 171025 645142 171077
rect 645194 171065 645200 171077
rect 649648 171065 649654 171077
rect 645194 171037 649654 171065
rect 645194 171025 645200 171037
rect 649648 171025 649654 171037
rect 649706 171025 649712 171077
rect 675280 169989 675286 170041
rect 675338 170029 675344 170041
rect 676240 170029 676246 170041
rect 675338 170001 676246 170029
rect 675338 169989 675344 170001
rect 676240 169989 676246 170001
rect 676298 169989 676304 170041
rect 675088 169915 675094 169967
rect 675146 169955 675152 169967
rect 676048 169955 676054 169967
rect 675146 169927 676054 169955
rect 675146 169915 675152 169927
rect 676048 169915 676054 169927
rect 676106 169915 676112 169967
rect 148432 169841 148438 169893
rect 148490 169881 148496 169893
rect 184528 169881 184534 169893
rect 148490 169853 184534 169881
rect 148490 169841 148496 169853
rect 184528 169841 184534 169853
rect 184586 169841 184592 169893
rect 148240 169767 148246 169819
rect 148298 169807 148304 169819
rect 184336 169807 184342 169819
rect 148298 169779 184342 169807
rect 148298 169767 148304 169779
rect 184336 169767 184342 169779
rect 184394 169767 184400 169819
rect 149296 169693 149302 169745
rect 149354 169733 149360 169745
rect 184624 169733 184630 169745
rect 149354 169705 184630 169733
rect 149354 169693 149360 169705
rect 184624 169693 184630 169705
rect 184682 169693 184688 169745
rect 148912 169619 148918 169671
rect 148970 169659 148976 169671
rect 184432 169659 184438 169671
rect 148970 169631 184438 169659
rect 148970 169619 148976 169631
rect 184432 169619 184438 169631
rect 184490 169619 184496 169671
rect 645136 168213 645142 168265
rect 645194 168253 645200 168265
rect 649840 168253 649846 168265
rect 645194 168225 649846 168253
rect 645194 168213 645200 168225
rect 649840 168213 649846 168225
rect 649898 168213 649904 168265
rect 674896 167103 674902 167155
rect 674954 167143 674960 167155
rect 676240 167143 676246 167155
rect 674954 167115 676246 167143
rect 674954 167103 674960 167115
rect 676240 167103 676246 167115
rect 676298 167103 676304 167155
rect 674992 167029 674998 167081
rect 675050 167069 675056 167081
rect 676048 167069 676054 167081
rect 675050 167041 676054 167069
rect 675050 167029 675056 167041
rect 676048 167029 676054 167041
rect 676106 167029 676112 167081
rect 148816 166955 148822 167007
rect 148874 166995 148880 167007
rect 184336 166995 184342 167007
rect 148874 166967 184342 166995
rect 148874 166955 148880 166967
rect 184336 166955 184342 166967
rect 184394 166955 184400 167007
rect 148624 166881 148630 166933
rect 148682 166921 148688 166933
rect 184432 166921 184438 166933
rect 148682 166893 184438 166921
rect 148682 166881 148688 166893
rect 184432 166881 184438 166893
rect 184490 166881 184496 166933
rect 154096 166807 154102 166859
rect 154154 166847 154160 166859
rect 184528 166847 184534 166859
rect 154154 166819 184534 166847
rect 154154 166807 154160 166819
rect 184528 166807 184534 166819
rect 184586 166807 184592 166859
rect 674128 166215 674134 166267
rect 674186 166255 674192 166267
rect 676048 166255 676054 166267
rect 674186 166227 676054 166255
rect 674186 166215 674192 166227
rect 676048 166215 676054 166227
rect 676106 166215 676112 166267
rect 646864 164365 646870 164417
rect 646922 164405 646928 164417
rect 676048 164405 676054 164417
rect 646922 164377 676054 164405
rect 646922 164365 646928 164377
rect 676048 164365 676054 164377
rect 676106 164365 676112 164417
rect 647056 164291 647062 164343
rect 647114 164331 647120 164343
rect 676240 164331 676246 164343
rect 647114 164303 676246 164331
rect 647114 164291 647120 164303
rect 676240 164291 676246 164303
rect 676298 164291 676304 164343
rect 646960 164217 646966 164269
rect 647018 164257 647024 164269
rect 676144 164257 676150 164269
rect 647018 164229 676150 164257
rect 647018 164217 647024 164229
rect 676144 164217 676150 164229
rect 676202 164217 676208 164269
rect 151216 164069 151222 164121
rect 151274 164109 151280 164121
rect 184528 164109 184534 164121
rect 151274 164081 184534 164109
rect 151274 164069 151280 164081
rect 184528 164069 184534 164081
rect 184586 164069 184592 164121
rect 156976 163995 156982 164047
rect 157034 164035 157040 164047
rect 184336 164035 184342 164047
rect 157034 164007 184342 164035
rect 157034 163995 157040 164007
rect 184336 163995 184342 164007
rect 184394 163995 184400 164047
rect 159760 163921 159766 163973
rect 159818 163961 159824 163973
rect 184432 163961 184438 163973
rect 159818 163933 184438 163961
rect 159818 163921 159824 163933
rect 184432 163921 184438 163933
rect 184490 163921 184496 163973
rect 174256 163847 174262 163899
rect 174314 163887 174320 163899
rect 184336 163887 184342 163899
rect 174314 163859 184342 163887
rect 174314 163847 174320 163859
rect 184336 163847 184342 163859
rect 184394 163847 184400 163899
rect 645136 163329 645142 163381
rect 645194 163369 645200 163381
rect 649936 163369 649942 163381
rect 645194 163341 649942 163369
rect 645194 163329 645200 163341
rect 649936 163329 649942 163341
rect 649994 163329 650000 163381
rect 151312 161183 151318 161235
rect 151370 161223 151376 161235
rect 184432 161223 184438 161235
rect 151370 161195 184438 161223
rect 151370 161183 151376 161195
rect 184432 161183 184438 161195
rect 184490 161183 184496 161235
rect 162736 161109 162742 161161
rect 162794 161149 162800 161161
rect 184528 161149 184534 161161
rect 162794 161121 184534 161149
rect 162794 161109 162800 161121
rect 184528 161109 184534 161121
rect 184586 161109 184592 161161
rect 168400 161035 168406 161087
rect 168458 161075 168464 161087
rect 184624 161075 184630 161087
rect 168458 161047 184630 161075
rect 168458 161035 168464 161047
rect 184624 161035 184630 161047
rect 184682 161035 184688 161087
rect 171376 160961 171382 161013
rect 171434 161001 171440 161013
rect 184336 161001 184342 161013
rect 171434 160973 184342 161001
rect 171434 160961 171440 160973
rect 184336 160961 184342 160973
rect 184394 160961 184400 161013
rect 675088 160591 675094 160643
rect 675146 160631 675152 160643
rect 675376 160631 675382 160643
rect 675146 160603 675382 160631
rect 675146 160591 675152 160603
rect 675376 160591 675382 160603
rect 675434 160591 675440 160643
rect 645136 159703 645142 159755
rect 645194 159743 645200 159755
rect 650032 159743 650038 159755
rect 645194 159715 650038 159743
rect 645194 159703 645200 159715
rect 650032 159703 650038 159715
rect 650090 159703 650096 159755
rect 147472 158889 147478 158941
rect 147530 158929 147536 158941
rect 152176 158929 152182 158941
rect 147530 158901 152182 158929
rect 147530 158889 147536 158901
rect 152176 158889 152182 158901
rect 152234 158889 152240 158941
rect 151408 158371 151414 158423
rect 151466 158411 151472 158423
rect 184336 158411 184342 158423
rect 151466 158383 184342 158411
rect 151466 158371 151472 158383
rect 184336 158371 184342 158383
rect 184394 158371 184400 158423
rect 165616 158297 165622 158349
rect 165674 158337 165680 158349
rect 184432 158337 184438 158349
rect 165674 158309 184438 158337
rect 165674 158297 165680 158309
rect 184432 158297 184438 158309
rect 184490 158297 184496 158349
rect 179920 158223 179926 158275
rect 179978 158263 179984 158275
rect 184528 158263 184534 158275
rect 179978 158235 184534 158263
rect 179978 158223 179984 158235
rect 184528 158223 184534 158235
rect 184586 158223 184592 158275
rect 177136 158149 177142 158201
rect 177194 158189 177200 158201
rect 184624 158189 184630 158201
rect 177194 158161 184630 158189
rect 177194 158149 177200 158161
rect 184624 158149 184630 158161
rect 184682 158149 184688 158201
rect 674992 157039 674998 157091
rect 675050 157079 675056 157091
rect 675472 157079 675478 157091
rect 675050 157051 675478 157079
rect 675050 157039 675056 157051
rect 675472 157039 675478 157051
rect 675530 157039 675536 157091
rect 674896 156299 674902 156351
rect 674954 156339 674960 156351
rect 675376 156339 675382 156351
rect 674954 156311 675382 156339
rect 674954 156299 674960 156311
rect 675376 156299 675382 156311
rect 675434 156299 675440 156351
rect 146896 156151 146902 156203
rect 146954 156191 146960 156203
rect 151216 156191 151222 156203
rect 146954 156163 151222 156191
rect 146954 156151 146960 156163
rect 151216 156151 151222 156163
rect 151274 156151 151280 156203
rect 645136 156003 645142 156055
rect 645194 156043 645200 156055
rect 650128 156043 650134 156055
rect 645194 156015 650134 156043
rect 645194 156003 645200 156015
rect 650128 156003 650134 156015
rect 650186 156003 650192 156055
rect 149296 155707 149302 155759
rect 149354 155747 149360 155759
rect 180016 155747 180022 155759
rect 149354 155719 180022 155747
rect 149354 155707 149360 155719
rect 180016 155707 180022 155719
rect 180074 155707 180080 155759
rect 149392 155633 149398 155685
rect 149450 155673 149456 155685
rect 177040 155673 177046 155685
rect 149450 155645 177046 155673
rect 149450 155633 149456 155645
rect 177040 155633 177046 155645
rect 177098 155633 177104 155685
rect 151792 155485 151798 155537
rect 151850 155525 151856 155537
rect 184528 155525 184534 155537
rect 151850 155497 184534 155525
rect 151850 155485 151856 155497
rect 184528 155485 184534 155497
rect 184586 155485 184592 155537
rect 658000 155485 658006 155537
rect 658058 155525 658064 155537
rect 675088 155525 675094 155537
rect 658058 155497 675094 155525
rect 658058 155485 658064 155497
rect 675088 155485 675094 155497
rect 675146 155485 675152 155537
rect 152080 155411 152086 155463
rect 152138 155451 152144 155463
rect 184624 155451 184630 155463
rect 152138 155423 184630 155451
rect 152138 155411 152144 155423
rect 184624 155411 184630 155423
rect 184682 155411 184688 155463
rect 159952 155337 159958 155389
rect 160010 155377 160016 155389
rect 184432 155377 184438 155389
rect 160010 155349 184438 155377
rect 160010 155337 160016 155349
rect 184432 155337 184438 155349
rect 184490 155337 184496 155389
rect 174352 155263 174358 155315
rect 174410 155303 174416 155315
rect 184336 155303 184342 155315
rect 174410 155275 184342 155303
rect 174410 155263 174416 155275
rect 184336 155263 184342 155275
rect 184394 155263 184400 155315
rect 149392 152747 149398 152799
rect 149450 152787 149456 152799
rect 174160 152787 174166 152799
rect 149450 152759 174166 152787
rect 149450 152747 149456 152759
rect 174160 152747 174166 152759
rect 174218 152747 174224 152799
rect 149296 152673 149302 152725
rect 149354 152713 149360 152725
rect 182896 152713 182902 152725
rect 149354 152685 182902 152713
rect 149354 152673 149360 152685
rect 182896 152673 182902 152685
rect 182954 152673 182960 152725
rect 151984 152599 151990 152651
rect 152042 152639 152048 152651
rect 184528 152639 184534 152651
rect 152042 152611 184534 152639
rect 152042 152599 152048 152611
rect 184528 152599 184534 152611
rect 184586 152599 184592 152651
rect 151600 152525 151606 152577
rect 151658 152565 151664 152577
rect 184432 152565 184438 152577
rect 151658 152537 184438 152565
rect 151658 152525 151664 152537
rect 184432 152525 184438 152537
rect 184490 152525 184496 152577
rect 645136 152525 645142 152577
rect 645194 152565 645200 152577
rect 650224 152565 650230 152577
rect 645194 152537 650230 152565
rect 645194 152525 645200 152537
rect 650224 152525 650230 152537
rect 650282 152525 650288 152577
rect 151696 152451 151702 152503
rect 151754 152491 151760 152503
rect 184336 152491 184342 152503
rect 151754 152463 184342 152491
rect 151754 152451 151760 152463
rect 184336 152451 184342 152463
rect 184394 152451 184400 152503
rect 674128 151415 674134 151467
rect 674186 151455 674192 151467
rect 675376 151455 675382 151467
rect 674186 151427 675382 151455
rect 674186 151415 674192 151427
rect 675376 151415 675382 151427
rect 675434 151415 675440 151467
rect 149296 149935 149302 149987
rect 149354 149975 149360 149987
rect 171376 149975 171382 149987
rect 149354 149947 171382 149975
rect 149354 149935 149360 149947
rect 171376 149935 171382 149947
rect 171434 149935 171440 149987
rect 149392 149861 149398 149913
rect 149450 149901 149456 149913
rect 174256 149901 174262 149913
rect 149450 149873 174262 149901
rect 149450 149861 149456 149873
rect 174256 149861 174262 149873
rect 174314 149861 174320 149913
rect 149200 149787 149206 149839
rect 149258 149827 149264 149839
rect 180208 149827 180214 149839
rect 149258 149799 180214 149827
rect 149258 149787 149264 149799
rect 180208 149787 180214 149799
rect 180266 149787 180272 149839
rect 182992 149713 182998 149765
rect 183050 149753 183056 149765
rect 184720 149753 184726 149765
rect 183050 149725 184726 149753
rect 183050 149713 183056 149725
rect 184720 149713 184726 149725
rect 184778 149713 184784 149765
rect 151888 149639 151894 149691
rect 151946 149679 151952 149691
rect 184432 149679 184438 149691
rect 151946 149651 184438 149679
rect 151946 149639 151952 149651
rect 184432 149639 184438 149651
rect 184490 149639 184496 149691
rect 180112 149565 180118 149617
rect 180170 149605 180176 149617
rect 184528 149605 184534 149617
rect 180170 149577 184534 149605
rect 180170 149565 180176 149577
rect 184528 149565 184534 149577
rect 184586 149565 184592 149617
rect 151504 149491 151510 149543
rect 151562 149531 151568 149543
rect 184336 149531 184342 149543
rect 151562 149503 184342 149531
rect 151562 149491 151568 149503
rect 184336 149491 184342 149503
rect 184394 149491 184400 149543
rect 645136 148159 645142 148211
rect 645194 148199 645200 148211
rect 650320 148199 650326 148211
rect 645194 148171 650326 148199
rect 645194 148159 645200 148171
rect 650320 148159 650326 148171
rect 650378 148159 650384 148211
rect 149392 146975 149398 147027
rect 149450 147015 149456 147027
rect 168400 147015 168406 147027
rect 149450 146987 168406 147015
rect 149450 146975 149456 146987
rect 168400 146975 168406 146987
rect 168458 146975 168464 147027
rect 149296 146901 149302 146953
rect 149354 146941 149360 146953
rect 177136 146941 177142 146953
rect 149354 146913 177142 146941
rect 149354 146901 149360 146913
rect 177136 146901 177142 146913
rect 177194 146901 177200 146953
rect 154192 146827 154198 146879
rect 154250 146867 154256 146879
rect 184528 146867 184534 146879
rect 154250 146839 184534 146867
rect 154250 146827 154256 146839
rect 184528 146827 184534 146839
rect 184586 146827 184592 146879
rect 162832 146753 162838 146805
rect 162890 146793 162896 146805
rect 184432 146793 184438 146805
rect 162890 146765 184438 146793
rect 162890 146753 162896 146765
rect 184432 146753 184438 146765
rect 184490 146753 184496 146805
rect 174448 146679 174454 146731
rect 174506 146719 174512 146731
rect 184336 146719 184342 146731
rect 174506 146691 184342 146719
rect 174506 146679 174512 146691
rect 184336 146679 184342 146691
rect 184394 146679 184400 146731
rect 177232 146605 177238 146657
rect 177290 146645 177296 146657
rect 184624 146645 184630 146657
rect 177290 146617 184630 146645
rect 177290 146605 177296 146617
rect 184624 146605 184630 146617
rect 184682 146605 184688 146657
rect 147664 145717 147670 145769
rect 147722 145757 147728 145769
rect 165520 145757 165526 145769
rect 147722 145729 165526 145757
rect 147722 145717 147728 145729
rect 165520 145717 165526 145729
rect 165578 145717 165584 145769
rect 147472 144015 147478 144067
rect 147530 144055 147536 144067
rect 162736 144055 162742 144067
rect 147530 144027 162742 144055
rect 147530 144015 147536 144027
rect 162736 144015 162742 144027
rect 162794 144015 162800 144067
rect 183088 143941 183094 143993
rect 183146 143981 183152 143993
rect 184624 143981 184630 143993
rect 183146 143953 184630 143981
rect 183146 143941 183152 143953
rect 184624 143941 184630 143953
rect 184682 143941 184688 143993
rect 168592 143867 168598 143919
rect 168650 143907 168656 143919
rect 184432 143907 184438 143919
rect 168650 143879 184438 143907
rect 168650 143867 168656 143879
rect 184432 143867 184438 143879
rect 184490 143867 184496 143919
rect 171568 143793 171574 143845
rect 171626 143833 171632 143845
rect 184336 143833 184342 143845
rect 171626 143805 184342 143833
rect 171626 143793 171632 143805
rect 184336 143793 184342 143805
rect 184394 143793 184400 143845
rect 165808 143719 165814 143771
rect 165866 143759 165872 143771
rect 184528 143759 184534 143771
rect 165866 143731 184534 143759
rect 165866 143719 165872 143731
rect 184528 143719 184534 143731
rect 184586 143719 184592 143771
rect 147472 143349 147478 143401
rect 147530 143389 147536 143401
rect 159856 143389 159862 143401
rect 147530 143361 159862 143389
rect 147530 143349 147536 143361
rect 159856 143349 159862 143361
rect 159914 143349 159920 143401
rect 147664 142387 147670 142439
rect 147722 142427 147728 142439
rect 156976 142427 156982 142439
rect 147722 142399 156982 142427
rect 147722 142387 147728 142399
rect 156976 142387 156982 142399
rect 157034 142387 157040 142439
rect 149680 141203 149686 141255
rect 149738 141243 149744 141255
rect 154096 141243 154102 141255
rect 149738 141215 154102 141243
rect 149738 141203 149744 141215
rect 154096 141203 154102 141215
rect 154154 141203 154160 141255
rect 154288 141055 154294 141107
rect 154346 141095 154352 141107
rect 184528 141095 184534 141107
rect 154346 141067 184534 141095
rect 154346 141055 154352 141067
rect 184528 141055 184534 141067
rect 184586 141055 184592 141107
rect 157072 140981 157078 141033
rect 157130 141021 157136 141033
rect 184432 141021 184438 141033
rect 157130 140993 184438 141021
rect 157130 140981 157136 140993
rect 184432 140981 184438 140993
rect 184490 140981 184496 141033
rect 160048 140907 160054 140959
rect 160106 140947 160112 140959
rect 184336 140947 184342 140959
rect 160106 140919 184342 140947
rect 160106 140907 160112 140919
rect 184336 140907 184342 140919
rect 184394 140907 184400 140959
rect 147472 140315 147478 140367
rect 147530 140355 147536 140367
rect 151120 140355 151126 140367
rect 147530 140327 151126 140355
rect 147530 140315 147536 140327
rect 151120 140315 151126 140327
rect 151178 140315 151184 140367
rect 147472 138243 147478 138295
rect 147530 138283 147536 138295
rect 159760 138283 159766 138295
rect 147530 138255 159766 138283
rect 147530 138243 147536 138255
rect 159760 138243 159766 138255
rect 159818 138243 159824 138295
rect 148048 137059 148054 137111
rect 148106 137099 148112 137111
rect 148432 137099 148438 137111
rect 148106 137071 148438 137099
rect 148106 137059 148112 137071
rect 148432 137059 148438 137071
rect 148490 137059 148496 137111
rect 148240 136985 148246 137037
rect 148298 137025 148304 137037
rect 148720 137025 148726 137037
rect 148298 136997 148726 137025
rect 148298 136985 148304 136997
rect 148720 136985 148726 136997
rect 148778 136985 148784 137037
rect 148432 136911 148438 136963
rect 148490 136951 148496 136963
rect 148624 136951 148630 136963
rect 148490 136923 148630 136951
rect 148490 136911 148496 136923
rect 148624 136911 148630 136923
rect 148682 136911 148688 136963
rect 148912 136911 148918 136963
rect 148970 136911 148976 136963
rect 148720 136689 148726 136741
rect 148778 136729 148784 136741
rect 148930 136729 148958 136911
rect 148778 136701 148958 136729
rect 148778 136689 148784 136701
rect 149680 135431 149686 135483
rect 149738 135471 149744 135483
rect 171280 135471 171286 135483
rect 149738 135443 171286 135471
rect 149738 135431 149744 135443
rect 171280 135431 171286 135443
rect 171338 135431 171344 135483
rect 149584 135357 149590 135409
rect 149642 135397 149648 135409
rect 179920 135397 179926 135409
rect 149642 135369 179926 135397
rect 149642 135357 149648 135369
rect 179920 135357 179926 135369
rect 179978 135357 179984 135409
rect 168496 135283 168502 135335
rect 168554 135323 168560 135335
rect 184432 135323 184438 135335
rect 168554 135295 184438 135323
rect 168554 135283 168560 135295
rect 184432 135283 184438 135295
rect 184490 135283 184496 135335
rect 171472 135209 171478 135261
rect 171530 135249 171536 135261
rect 184336 135249 184342 135261
rect 171530 135221 184342 135249
rect 171530 135209 171536 135221
rect 184336 135209 184342 135221
rect 184394 135209 184400 135261
rect 177136 132545 177142 132597
rect 177194 132585 177200 132597
rect 184720 132585 184726 132597
rect 177194 132557 184726 132585
rect 177194 132545 177200 132557
rect 184720 132545 184726 132557
rect 184778 132545 184784 132597
rect 149680 132471 149686 132523
rect 149738 132511 149744 132523
rect 182992 132511 182998 132523
rect 149738 132483 182998 132511
rect 149738 132471 149744 132483
rect 182992 132471 182998 132483
rect 183050 132471 183056 132523
rect 154000 132397 154006 132449
rect 154058 132437 154064 132449
rect 184624 132437 184630 132449
rect 154058 132409 184630 132437
rect 154058 132397 154064 132409
rect 184624 132397 184630 132409
rect 184682 132397 184688 132449
rect 156880 132323 156886 132375
rect 156938 132363 156944 132375
rect 184528 132363 184534 132375
rect 156938 132335 184534 132363
rect 156938 132323 156944 132335
rect 184528 132323 184534 132335
rect 184586 132323 184592 132375
rect 162928 132249 162934 132301
rect 162986 132289 162992 132301
rect 184432 132289 184438 132301
rect 162986 132261 184438 132289
rect 162986 132249 162992 132261
rect 184432 132249 184438 132261
rect 184490 132249 184496 132301
rect 165712 132175 165718 132227
rect 165770 132215 165776 132227
rect 184336 132215 184342 132227
rect 165770 132187 184342 132215
rect 165770 132175 165776 132187
rect 184336 132175 184342 132187
rect 184394 132175 184400 132227
rect 180208 132027 180214 132079
rect 180266 132067 180272 132079
rect 185584 132067 185590 132079
rect 180266 132039 185590 132067
rect 180266 132027 180272 132039
rect 185584 132027 185590 132039
rect 185642 132027 185648 132079
rect 655312 130103 655318 130155
rect 655370 130143 655376 130155
rect 676144 130143 676150 130155
rect 655370 130115 676150 130143
rect 655370 130103 655376 130115
rect 676144 130103 676150 130115
rect 676202 130103 676208 130155
rect 655216 129955 655222 130007
rect 655274 129995 655280 130007
rect 676240 129995 676246 130007
rect 655274 129967 676246 129995
rect 655274 129955 655280 129967
rect 676240 129955 676246 129967
rect 676298 129955 676304 130007
rect 655120 129807 655126 129859
rect 655178 129847 655184 129859
rect 676336 129847 676342 129859
rect 655178 129819 676342 129847
rect 655178 129807 655184 129819
rect 676336 129807 676342 129819
rect 676394 129807 676400 129859
rect 147472 129659 147478 129711
rect 147530 129699 147536 129711
rect 165616 129699 165622 129711
rect 147530 129671 165622 129699
rect 147530 129659 147536 129671
rect 165616 129659 165622 129671
rect 165674 129659 165680 129711
rect 149680 129585 149686 129637
rect 149738 129625 149744 129637
rect 168496 129625 168502 129637
rect 149738 129597 168502 129625
rect 149738 129585 149744 129597
rect 168496 129585 168502 129597
rect 168554 129585 168560 129637
rect 645712 129585 645718 129637
rect 645770 129625 645776 129637
rect 676240 129625 676246 129637
rect 645770 129597 676246 129625
rect 645770 129585 645776 129597
rect 676240 129585 676246 129597
rect 676298 129585 676304 129637
rect 182800 129511 182806 129563
rect 182858 129551 182864 129563
rect 186736 129551 186742 129563
rect 182858 129523 186742 129551
rect 182858 129511 182864 129523
rect 186736 129511 186742 129523
rect 186794 129511 186800 129563
rect 149488 129437 149494 129489
rect 149546 129477 149552 129489
rect 184432 129477 184438 129489
rect 149546 129449 184438 129477
rect 149546 129437 149552 129449
rect 184432 129437 184438 129449
rect 184490 129437 184496 129489
rect 149392 129363 149398 129415
rect 149450 129403 149456 129415
rect 184528 129403 184534 129415
rect 149450 129375 184534 129403
rect 149450 129363 149456 129375
rect 184528 129363 184534 129375
rect 184586 129363 184592 129415
rect 149104 129289 149110 129341
rect 149162 129329 149168 129341
rect 184336 129329 184342 129341
rect 149162 129301 184342 129329
rect 149162 129289 149168 129301
rect 184336 129289 184342 129301
rect 184394 129289 184400 129341
rect 147472 127809 147478 127861
rect 147530 127849 147536 127861
rect 162640 127849 162646 127861
rect 147530 127821 162646 127849
rect 147530 127809 147536 127821
rect 162640 127809 162646 127821
rect 162698 127809 162704 127861
rect 646480 126921 646486 126973
rect 646538 126961 646544 126973
rect 676240 126961 676246 126973
rect 646538 126933 676246 126961
rect 646538 126921 646544 126933
rect 676240 126921 676246 126933
rect 676298 126921 676304 126973
rect 646576 126773 646582 126825
rect 646634 126813 646640 126825
rect 676144 126813 676150 126825
rect 646634 126785 676150 126813
rect 646634 126773 646640 126785
rect 676144 126773 676150 126785
rect 676202 126773 676208 126825
rect 674320 126699 674326 126751
rect 674378 126739 674384 126751
rect 676048 126739 676054 126751
rect 674378 126711 676054 126739
rect 674378 126699 674384 126711
rect 676048 126699 676054 126711
rect 676106 126699 676112 126751
rect 148336 126625 148342 126677
rect 148394 126665 148400 126677
rect 184528 126665 184534 126677
rect 148394 126637 184534 126665
rect 148394 126625 148400 126637
rect 184528 126625 184534 126637
rect 184586 126625 184592 126677
rect 148528 126551 148534 126603
rect 148586 126591 148592 126603
rect 184432 126591 184438 126603
rect 148586 126563 184438 126591
rect 148586 126551 148592 126563
rect 184432 126551 184438 126563
rect 184490 126551 184496 126603
rect 148912 126477 148918 126529
rect 148970 126517 148976 126529
rect 184336 126517 184342 126529
rect 148970 126489 184342 126517
rect 148970 126477 148976 126489
rect 184336 126477 184342 126489
rect 184394 126477 184400 126529
rect 149392 124183 149398 124235
rect 149450 124223 149456 124235
rect 156880 124223 156886 124235
rect 149450 124195 156886 124223
rect 149450 124183 149456 124195
rect 156880 124183 156886 124195
rect 156938 124183 156944 124235
rect 674608 124183 674614 124235
rect 674666 124223 674672 124235
rect 676048 124223 676054 124235
rect 674666 124195 676054 124223
rect 674666 124183 674672 124195
rect 676048 124183 676054 124195
rect 676106 124183 676112 124235
rect 674800 123961 674806 124013
rect 674858 124001 674864 124013
rect 676048 124001 676054 124013
rect 674858 123973 676054 124001
rect 674858 123961 674864 123973
rect 676048 123961 676054 123973
rect 676106 123961 676112 124013
rect 675280 123887 675286 123939
rect 675338 123927 675344 123939
rect 676240 123927 676246 123939
rect 675338 123899 676246 123927
rect 675338 123887 675344 123899
rect 676240 123887 676246 123899
rect 676298 123887 676304 123939
rect 148144 123813 148150 123865
rect 148202 123853 148208 123865
rect 184624 123853 184630 123865
rect 148202 123825 184630 123853
rect 148202 123813 148208 123825
rect 184624 123813 184630 123825
rect 184682 123813 184688 123865
rect 148720 123739 148726 123791
rect 148778 123779 148784 123791
rect 184528 123779 184534 123791
rect 148778 123751 184534 123779
rect 148778 123739 148784 123751
rect 184528 123739 184534 123751
rect 184586 123739 184592 123791
rect 148048 123665 148054 123717
rect 148106 123705 148112 123717
rect 184432 123705 184438 123717
rect 148106 123677 184438 123705
rect 148106 123665 148112 123677
rect 184432 123665 184438 123677
rect 184490 123665 184496 123717
rect 148240 123591 148246 123643
rect 148298 123631 148304 123643
rect 184336 123631 184342 123643
rect 148298 123603 184342 123631
rect 148298 123591 148304 123603
rect 184336 123591 184342 123603
rect 184394 123591 184400 123643
rect 174256 122407 174262 122459
rect 174314 122447 174320 122459
rect 186160 122447 186166 122459
rect 174314 122419 186166 122447
rect 174314 122407 174320 122419
rect 186160 122407 186166 122419
rect 186218 122407 186224 122459
rect 675088 122111 675094 122163
rect 675146 122151 675152 122163
rect 676048 122151 676054 122163
rect 675146 122123 676054 122151
rect 675146 122111 675152 122123
rect 676048 122111 676054 122123
rect 676106 122111 676112 122163
rect 674704 121149 674710 121201
rect 674762 121189 674768 121201
rect 675952 121189 675958 121201
rect 674762 121161 675958 121189
rect 674762 121149 674768 121161
rect 675952 121149 675958 121161
rect 676010 121149 676016 121201
rect 674896 121075 674902 121127
rect 674954 121115 674960 121127
rect 676240 121115 676246 121127
rect 674954 121087 676246 121115
rect 674954 121075 674960 121087
rect 676240 121075 676246 121087
rect 676298 121075 676304 121127
rect 674992 121001 674998 121053
rect 675050 121041 675056 121053
rect 676048 121041 676054 121053
rect 675050 121013 676054 121041
rect 675050 121001 675056 121013
rect 676048 121001 676054 121013
rect 676106 121001 676112 121053
rect 148624 120927 148630 120979
rect 148682 120967 148688 120979
rect 184528 120967 184534 120979
rect 148682 120939 184534 120967
rect 148682 120927 148688 120939
rect 184528 120927 184534 120939
rect 184586 120927 184592 120979
rect 148432 120853 148438 120905
rect 148490 120893 148496 120905
rect 184336 120893 184342 120905
rect 148490 120865 184342 120893
rect 148490 120853 148496 120865
rect 184336 120853 184342 120865
rect 184394 120853 184400 120905
rect 171376 120779 171382 120831
rect 171434 120819 171440 120831
rect 184432 120819 184438 120831
rect 171434 120791 184438 120819
rect 171434 120779 171440 120791
rect 184432 120779 184438 120791
rect 184490 120779 184496 120831
rect 147856 120483 147862 120535
rect 147914 120523 147920 120535
rect 154480 120523 154486 120535
rect 147914 120495 154486 120523
rect 147914 120483 147920 120495
rect 154480 120483 154486 120495
rect 154538 120483 154544 120535
rect 647824 118337 647830 118389
rect 647882 118377 647888 118389
rect 676240 118377 676246 118389
rect 647882 118349 676246 118377
rect 647882 118337 647888 118349
rect 676240 118337 676246 118349
rect 676298 118337 676304 118389
rect 149392 118189 149398 118241
rect 149450 118229 149456 118241
rect 168592 118229 168598 118241
rect 149450 118201 168598 118229
rect 149450 118189 149456 118201
rect 168592 118189 168598 118201
rect 168650 118189 168656 118241
rect 647920 118189 647926 118241
rect 647978 118229 647984 118241
rect 676144 118229 676150 118241
rect 647978 118201 676150 118229
rect 647978 118189 647984 118201
rect 676144 118189 676150 118201
rect 676202 118189 676208 118241
rect 149488 118115 149494 118167
rect 149546 118155 149552 118167
rect 174256 118155 174262 118167
rect 149546 118127 174262 118155
rect 149546 118115 149552 118127
rect 174256 118115 174262 118127
rect 174314 118115 174320 118167
rect 645232 118115 645238 118167
rect 645290 118155 645296 118167
rect 676048 118155 676054 118167
rect 645290 118127 676054 118155
rect 645290 118115 645296 118127
rect 676048 118115 676054 118127
rect 676106 118115 676112 118167
rect 159856 118041 159862 118093
rect 159914 118081 159920 118093
rect 184624 118081 184630 118093
rect 159914 118053 184630 118081
rect 159914 118041 159920 118053
rect 184624 118041 184630 118053
rect 184682 118041 184688 118093
rect 162736 117967 162742 118019
rect 162794 118007 162800 118019
rect 184528 118007 184534 118019
rect 162794 117979 184534 118007
rect 162794 117967 162800 117979
rect 184528 117967 184534 117979
rect 184586 117967 184592 118019
rect 165520 117893 165526 117945
rect 165578 117933 165584 117945
rect 184432 117933 184438 117945
rect 165578 117905 184438 117933
rect 165578 117893 165584 117905
rect 184432 117893 184438 117905
rect 184490 117893 184496 117945
rect 168400 117819 168406 117871
rect 168458 117859 168464 117871
rect 184336 117859 184342 117871
rect 168458 117831 184342 117859
rect 168458 117819 168464 117831
rect 184336 117819 184342 117831
rect 184394 117819 184400 117871
rect 675568 115969 675574 116021
rect 675626 115969 675632 116021
rect 675586 115355 675614 115969
rect 149392 115303 149398 115355
rect 149450 115343 149456 115355
rect 162832 115343 162838 115355
rect 149450 115315 162838 115343
rect 149450 115303 149456 115315
rect 162832 115303 162838 115315
rect 162890 115303 162896 115355
rect 675568 115303 675574 115355
rect 675626 115303 675632 115355
rect 149488 115229 149494 115281
rect 149546 115269 149552 115281
rect 165712 115269 165718 115281
rect 149546 115241 165718 115269
rect 149546 115229 149552 115241
rect 165712 115229 165718 115241
rect 165770 115229 165776 115281
rect 647920 115229 647926 115281
rect 647978 115269 647984 115281
rect 665296 115269 665302 115281
rect 647978 115241 665302 115269
rect 647978 115229 647984 115241
rect 665296 115229 665302 115241
rect 665354 115229 665360 115281
rect 670384 115229 670390 115281
rect 670442 115269 670448 115281
rect 675472 115269 675478 115281
rect 670442 115241 675478 115269
rect 670442 115229 670448 115241
rect 675472 115229 675478 115241
rect 675530 115229 675536 115281
rect 152176 115155 152182 115207
rect 152234 115195 152240 115207
rect 184528 115195 184534 115207
rect 152234 115167 184534 115195
rect 152234 115155 152240 115167
rect 184528 115155 184534 115167
rect 184586 115155 184592 115207
rect 154096 115081 154102 115133
rect 154154 115121 154160 115133
rect 184432 115121 184438 115133
rect 154154 115093 184438 115121
rect 154154 115081 154160 115093
rect 184432 115081 184438 115093
rect 184490 115081 184496 115133
rect 156976 115007 156982 115059
rect 157034 115047 157040 115059
rect 184336 115047 184342 115059
rect 157034 115019 184342 115047
rect 157034 115007 157040 115019
rect 184336 115007 184342 115019
rect 184394 115007 184400 115059
rect 180016 114119 180022 114171
rect 180074 114159 180080 114171
rect 184624 114159 184630 114171
rect 180074 114131 184630 114159
rect 180074 114119 180080 114131
rect 184624 114119 184630 114131
rect 184682 114119 184688 114171
rect 674320 114119 674326 114171
rect 674378 114159 674384 114171
rect 675376 114159 675382 114171
rect 674378 114131 675382 114159
rect 674378 114119 674384 114131
rect 675376 114119 675382 114131
rect 675434 114119 675440 114171
rect 149392 114045 149398 114097
rect 149450 114085 149456 114097
rect 159856 114085 159862 114097
rect 149450 114057 159862 114085
rect 149450 114045 149456 114057
rect 159856 114045 159862 114057
rect 159914 114045 159920 114097
rect 663760 112935 663766 112987
rect 663818 112975 663824 112987
rect 665200 112975 665206 112987
rect 663818 112947 665206 112975
rect 663818 112935 663824 112947
rect 665200 112935 665206 112947
rect 665258 112935 665264 112987
rect 674608 112491 674614 112543
rect 674666 112531 674672 112543
rect 675376 112531 675382 112543
rect 674666 112503 675382 112531
rect 674666 112491 674672 112503
rect 675376 112491 675382 112503
rect 675434 112491 675440 112543
rect 149392 112343 149398 112395
rect 149450 112383 149456 112395
rect 177136 112383 177142 112395
rect 149450 112355 177142 112383
rect 149450 112343 149456 112355
rect 177136 112343 177142 112355
rect 177194 112343 177200 112395
rect 151216 112269 151222 112321
rect 151274 112309 151280 112321
rect 184336 112309 184342 112321
rect 151274 112281 184342 112309
rect 151274 112269 151280 112281
rect 184336 112269 184342 112281
rect 184394 112269 184400 112321
rect 665200 112269 665206 112321
rect 665258 112309 665264 112321
rect 670384 112309 670390 112321
rect 665258 112281 670390 112309
rect 665258 112269 665264 112281
rect 670384 112269 670390 112281
rect 670442 112269 670448 112321
rect 182896 112195 182902 112247
rect 182954 112235 182960 112247
rect 184528 112235 184534 112247
rect 182954 112207 184534 112235
rect 182954 112195 182960 112207
rect 184528 112195 184534 112207
rect 184586 112195 184592 112247
rect 177040 112121 177046 112173
rect 177098 112161 177104 112173
rect 184432 112161 184438 112173
rect 177098 112133 184438 112161
rect 177098 112121 177104 112133
rect 184432 112121 184438 112133
rect 184490 112121 184496 112173
rect 674800 111825 674806 111877
rect 674858 111865 674864 111877
rect 675376 111865 675382 111877
rect 674858 111837 675382 111865
rect 674858 111825 674864 111837
rect 675376 111825 675382 111837
rect 675434 111825 675440 111877
rect 675184 111159 675190 111211
rect 675242 111199 675248 111211
rect 675376 111199 675382 111211
rect 675242 111171 675382 111199
rect 675242 111159 675248 111171
rect 675376 111159 675382 111171
rect 675434 111159 675440 111211
rect 674992 110641 674998 110693
rect 675050 110681 675056 110693
rect 675376 110681 675382 110693
rect 675050 110653 675382 110681
rect 675050 110641 675056 110653
rect 675376 110641 675382 110653
rect 675434 110641 675440 110693
rect 148624 109531 148630 109583
rect 148682 109571 148688 109583
rect 154000 109571 154006 109583
rect 148682 109543 154006 109571
rect 148682 109531 148688 109543
rect 154000 109531 154006 109543
rect 154058 109531 154064 109583
rect 149392 109457 149398 109509
rect 149450 109497 149456 109509
rect 156976 109497 156982 109509
rect 149450 109469 156982 109497
rect 149450 109457 149456 109469
rect 156976 109457 156982 109469
rect 157034 109457 157040 109509
rect 159760 109383 159766 109435
rect 159818 109423 159824 109435
rect 184432 109423 184438 109435
rect 159818 109395 184438 109423
rect 159818 109383 159824 109395
rect 184432 109383 184438 109395
rect 184490 109383 184496 109435
rect 174160 109309 174166 109361
rect 174218 109349 174224 109361
rect 184336 109349 184342 109361
rect 174218 109321 184342 109349
rect 174218 109309 174224 109321
rect 184336 109309 184342 109321
rect 184394 109309 184400 109361
rect 147184 108273 147190 108325
rect 147242 108313 147248 108325
rect 151120 108313 151126 108325
rect 147242 108285 151126 108313
rect 147242 108273 147248 108285
rect 151120 108273 151126 108285
rect 151178 108273 151184 108325
rect 674896 107533 674902 107585
rect 674954 107573 674960 107585
rect 675376 107573 675382 107585
rect 674954 107545 675382 107573
rect 674954 107533 674960 107545
rect 675376 107533 675382 107545
rect 675434 107533 675440 107585
rect 182992 106497 182998 106549
rect 183050 106537 183056 106549
rect 184528 106537 184534 106549
rect 183050 106509 184534 106537
rect 183050 106497 183056 106509
rect 184528 106497 184534 106509
rect 184586 106497 184592 106549
rect 171280 106423 171286 106475
rect 171338 106463 171344 106475
rect 184336 106463 184342 106475
rect 171338 106435 184342 106463
rect 171338 106423 171344 106435
rect 184336 106423 184342 106435
rect 184394 106423 184400 106475
rect 179920 106349 179926 106401
rect 179978 106389 179984 106401
rect 185296 106389 185302 106401
rect 179978 106361 185302 106389
rect 179978 106349 179984 106361
rect 185296 106349 185302 106361
rect 185354 106349 185360 106401
rect 674800 106349 674806 106401
rect 674858 106389 674864 106401
rect 675376 106389 675382 106401
rect 674858 106361 675382 106389
rect 674858 106349 674864 106361
rect 675376 106349 675382 106361
rect 675434 106349 675440 106401
rect 149488 106275 149494 106327
rect 149546 106315 149552 106327
rect 184432 106315 184438 106327
rect 149546 106287 184438 106315
rect 149546 106275 149552 106287
rect 184432 106275 184438 106287
rect 184490 106275 184496 106327
rect 154480 105091 154486 105143
rect 154538 105131 154544 105143
rect 184720 105131 184726 105143
rect 154538 105103 184726 105131
rect 154538 105091 154544 105103
rect 184720 105091 184726 105103
rect 184778 105091 184784 105143
rect 647920 103907 647926 103959
rect 647978 103947 647984 103959
rect 661168 103947 661174 103959
rect 647978 103919 661174 103947
rect 647978 103907 647984 103919
rect 661168 103907 661174 103919
rect 661226 103907 661232 103959
rect 645904 103685 645910 103737
rect 645962 103725 645968 103737
rect 657520 103725 657526 103737
rect 645962 103697 657526 103725
rect 645962 103685 645968 103697
rect 657520 103685 657526 103697
rect 657578 103685 657584 103737
rect 149008 103611 149014 103663
rect 149066 103651 149072 103663
rect 184432 103651 184438 103663
rect 149066 103623 184438 103651
rect 149066 103611 149072 103623
rect 184432 103611 184438 103623
rect 184490 103611 184496 103663
rect 149104 103537 149110 103589
rect 149162 103577 149168 103589
rect 184624 103577 184630 103589
rect 149162 103549 184630 103577
rect 149162 103537 149168 103549
rect 184624 103537 184630 103549
rect 184682 103537 184688 103589
rect 165616 103463 165622 103515
rect 165674 103503 165680 103515
rect 184528 103503 184534 103515
rect 165674 103475 184534 103503
rect 165674 103463 165680 103475
rect 184528 103463 184534 103475
rect 184586 103463 184592 103515
rect 168496 103389 168502 103441
rect 168554 103429 168560 103441
rect 184336 103429 184342 103441
rect 168554 103401 184342 103429
rect 168554 103389 168560 103401
rect 184336 103389 184342 103401
rect 184394 103389 184400 103441
rect 645136 102057 645142 102109
rect 645194 102097 645200 102109
rect 652432 102097 652438 102109
rect 645194 102069 652438 102097
rect 645194 102057 645200 102069
rect 652432 102057 652438 102069
rect 652490 102057 652496 102109
rect 149392 100799 149398 100851
rect 149450 100839 149456 100851
rect 171280 100839 171286 100851
rect 149450 100811 171286 100839
rect 149450 100799 149456 100811
rect 171280 100799 171286 100811
rect 171338 100799 171344 100851
rect 149584 100725 149590 100777
rect 149642 100765 149648 100777
rect 184624 100765 184630 100777
rect 149642 100737 184630 100765
rect 149642 100725 149648 100737
rect 184624 100725 184630 100737
rect 184682 100725 184688 100777
rect 149296 100651 149302 100703
rect 149354 100691 149360 100703
rect 184432 100691 184438 100703
rect 149354 100663 184438 100691
rect 149354 100651 149360 100663
rect 184432 100651 184438 100663
rect 184490 100651 184496 100703
rect 156880 100577 156886 100629
rect 156938 100617 156944 100629
rect 184528 100617 184534 100629
rect 156938 100589 184534 100617
rect 156938 100577 156944 100589
rect 184528 100577 184534 100589
rect 184586 100577 184592 100629
rect 162640 100503 162646 100555
rect 162698 100543 162704 100555
rect 184336 100543 184342 100555
rect 162698 100515 184342 100543
rect 162698 100503 162704 100515
rect 184336 100503 184342 100515
rect 184394 100503 184400 100555
rect 149392 97987 149398 98039
rect 149450 98027 149456 98039
rect 184240 98027 184246 98039
rect 149450 97999 184246 98027
rect 149450 97987 149456 97999
rect 184240 97987 184246 97999
rect 184298 97987 184304 98039
rect 149488 97913 149494 97965
rect 149546 97953 149552 97965
rect 186160 97953 186166 97965
rect 149546 97925 186166 97953
rect 149546 97913 149552 97925
rect 186160 97913 186166 97925
rect 186218 97913 186224 97965
rect 647920 97913 647926 97965
rect 647978 97953 647984 97965
rect 662512 97953 662518 97965
rect 647978 97925 662518 97953
rect 647978 97913 647984 97925
rect 662512 97913 662518 97925
rect 662570 97913 662576 97965
rect 148336 97839 148342 97891
rect 148394 97879 148400 97891
rect 184336 97879 184342 97891
rect 148394 97851 184342 97879
rect 148394 97839 148400 97851
rect 184336 97839 184342 97851
rect 184394 97839 184400 97891
rect 148528 97765 148534 97817
rect 148586 97805 148592 97817
rect 184432 97805 184438 97817
rect 148586 97777 184438 97805
rect 148586 97765 148592 97777
rect 184432 97765 184438 97777
rect 184490 97765 184496 97817
rect 642256 96433 642262 96485
rect 642314 96473 642320 96485
rect 665200 96473 665206 96485
rect 642314 96445 665206 96473
rect 642314 96433 642320 96445
rect 665200 96433 665206 96445
rect 665258 96433 665264 96485
rect 645424 95915 645430 95967
rect 645482 95955 645488 95967
rect 653680 95955 653686 95967
rect 645482 95927 653686 95955
rect 645482 95915 645488 95927
rect 653680 95915 653686 95927
rect 653738 95915 653744 95967
rect 149488 95101 149494 95153
rect 149546 95141 149552 95153
rect 168208 95141 168214 95153
rect 149546 95113 168214 95141
rect 149546 95101 149552 95113
rect 168208 95101 168214 95113
rect 168266 95101 168272 95153
rect 149392 95027 149398 95079
rect 149450 95067 149456 95079
rect 179920 95067 179926 95079
rect 149450 95039 179926 95067
rect 149450 95027 149456 95039
rect 179920 95027 179926 95039
rect 179978 95027 179984 95079
rect 162832 94953 162838 95005
rect 162890 94993 162896 95005
rect 184624 94993 184630 95005
rect 162890 94965 184630 94993
rect 162890 94953 162896 94965
rect 184624 94953 184630 94965
rect 184682 94953 184688 95005
rect 165712 94879 165718 94931
rect 165770 94919 165776 94931
rect 184528 94919 184534 94931
rect 165770 94891 184534 94919
rect 165770 94879 165776 94891
rect 184528 94879 184534 94891
rect 184586 94879 184592 94931
rect 168592 94805 168598 94857
rect 168650 94845 168656 94857
rect 184432 94845 184438 94857
rect 168650 94817 184438 94845
rect 168650 94805 168656 94817
rect 184432 94805 184438 94817
rect 184490 94805 184496 94857
rect 174256 94731 174262 94783
rect 174314 94771 174320 94783
rect 184336 94771 184342 94783
rect 174314 94743 184342 94771
rect 174314 94731 174320 94743
rect 184336 94731 184342 94743
rect 184394 94731 184400 94783
rect 646768 92659 646774 92711
rect 646826 92699 646832 92711
rect 663088 92699 663094 92711
rect 646826 92671 663094 92699
rect 646826 92659 646832 92671
rect 663088 92659 663094 92671
rect 663146 92659 663152 92711
rect 646480 92363 646486 92415
rect 646538 92403 646544 92415
rect 660688 92403 660694 92415
rect 646538 92375 660694 92403
rect 646538 92363 646544 92375
rect 660688 92363 660694 92375
rect 660746 92363 660752 92415
rect 645520 92289 645526 92341
rect 645578 92329 645584 92341
rect 661744 92329 661750 92341
rect 645578 92301 661750 92329
rect 645578 92289 645584 92301
rect 661744 92289 661750 92301
rect 661802 92289 661808 92341
rect 149392 92215 149398 92267
rect 149450 92255 149456 92267
rect 162448 92255 162454 92267
rect 149450 92227 162454 92255
rect 149450 92215 149456 92227
rect 162448 92215 162454 92227
rect 162506 92215 162512 92267
rect 646864 92215 646870 92267
rect 646922 92255 646928 92267
rect 659824 92255 659830 92267
rect 646922 92227 659830 92255
rect 646922 92215 646928 92227
rect 659824 92215 659830 92227
rect 659882 92215 659888 92267
rect 149488 92141 149494 92193
rect 149546 92181 149552 92193
rect 165232 92181 165238 92193
rect 149546 92153 165238 92181
rect 149546 92141 149552 92153
rect 165232 92141 165238 92153
rect 165290 92141 165296 92193
rect 646960 92141 646966 92193
rect 647018 92181 647024 92193
rect 658864 92181 658870 92193
rect 647018 92153 658870 92181
rect 647018 92141 647024 92153
rect 658864 92141 658870 92153
rect 658922 92141 658928 92193
rect 148240 92067 148246 92119
rect 148298 92107 148304 92119
rect 184432 92107 184438 92119
rect 148298 92079 184438 92107
rect 148298 92067 148304 92079
rect 184432 92067 184438 92079
rect 184490 92067 184496 92119
rect 156976 91993 156982 92045
rect 157034 92033 157040 92045
rect 184528 92033 184534 92045
rect 157034 92005 184534 92033
rect 157034 91993 157040 92005
rect 184528 91993 184534 92005
rect 184586 91993 184592 92045
rect 159856 91919 159862 91971
rect 159914 91959 159920 91971
rect 184336 91959 184342 91971
rect 159914 91931 184342 91959
rect 159914 91919 159920 91931
rect 184336 91919 184342 91931
rect 184394 91919 184400 91971
rect 177136 91845 177142 91897
rect 177194 91885 177200 91897
rect 184624 91885 184630 91897
rect 177194 91857 184630 91885
rect 177194 91845 177200 91857
rect 184624 91845 184630 91857
rect 184682 91845 184688 91897
rect 149392 90069 149398 90121
rect 149450 90109 149456 90121
rect 159760 90109 159766 90121
rect 149450 90081 159766 90109
rect 149450 90069 149456 90081
rect 159760 90069 159766 90081
rect 159818 90069 159824 90121
rect 148432 89181 148438 89233
rect 148490 89221 148496 89233
rect 184528 89221 184534 89233
rect 148490 89193 184534 89221
rect 148490 89181 148496 89193
rect 184528 89181 184534 89193
rect 184586 89181 184592 89233
rect 148816 89107 148822 89159
rect 148874 89147 148880 89159
rect 184624 89147 184630 89159
rect 148874 89119 184630 89147
rect 148874 89107 148880 89119
rect 184624 89107 184630 89119
rect 184682 89107 184688 89159
rect 151120 89033 151126 89085
rect 151178 89073 151184 89085
rect 184432 89073 184438 89085
rect 151178 89045 184438 89073
rect 151178 89033 151184 89045
rect 184432 89033 184438 89045
rect 184490 89033 184496 89085
rect 154000 88959 154006 89011
rect 154058 88999 154064 89011
rect 184336 88999 184342 89011
rect 154058 88971 184342 88999
rect 154058 88959 154064 88971
rect 184336 88959 184342 88971
rect 184394 88959 184400 89011
rect 645904 87479 645910 87531
rect 645962 87519 645968 87531
rect 650896 87519 650902 87531
rect 645962 87491 650902 87519
rect 645962 87479 645968 87491
rect 650896 87479 650902 87491
rect 650954 87479 650960 87531
rect 647920 87257 647926 87309
rect 647978 87297 647984 87309
rect 658000 87297 658006 87309
rect 647978 87269 658006 87297
rect 647978 87257 647984 87269
rect 658000 87257 658006 87269
rect 658058 87257 658064 87309
rect 647056 87035 647062 87087
rect 647114 87075 647120 87087
rect 663280 87075 663286 87087
rect 647114 87047 663286 87075
rect 647114 87035 647120 87047
rect 663280 87035 663286 87047
rect 663338 87035 663344 87087
rect 149488 86739 149494 86791
rect 149546 86779 149552 86791
rect 156496 86779 156502 86791
rect 149546 86751 156502 86779
rect 149546 86739 149552 86751
rect 156496 86739 156502 86751
rect 156554 86739 156560 86791
rect 148816 86443 148822 86495
rect 148874 86483 148880 86495
rect 154096 86483 154102 86495
rect 148874 86455 154102 86483
rect 148874 86443 148880 86455
rect 154096 86443 154102 86455
rect 154154 86443 154160 86495
rect 148624 86369 148630 86421
rect 148682 86409 148688 86421
rect 184336 86409 184342 86421
rect 148682 86381 184342 86409
rect 148682 86369 148688 86381
rect 184336 86369 184342 86381
rect 184394 86369 184400 86421
rect 148720 86295 148726 86347
rect 148778 86335 148784 86347
rect 184432 86335 184438 86347
rect 148778 86307 184438 86335
rect 148778 86295 148784 86307
rect 184432 86295 184438 86307
rect 184490 86295 184496 86347
rect 148912 86221 148918 86273
rect 148970 86261 148976 86273
rect 184528 86261 184534 86273
rect 148970 86233 184534 86261
rect 148970 86221 148976 86233
rect 184528 86221 184534 86233
rect 184586 86221 184592 86273
rect 645904 84149 645910 84201
rect 645962 84189 645968 84201
rect 657040 84189 657046 84201
rect 645962 84161 657046 84189
rect 645962 84149 645968 84161
rect 657040 84149 657046 84161
rect 657098 84149 657104 84201
rect 147088 83557 147094 83609
rect 147146 83597 147152 83609
rect 151120 83597 151126 83609
rect 147146 83569 151126 83597
rect 147146 83557 147152 83569
rect 151120 83557 151126 83569
rect 151178 83557 151184 83609
rect 646768 83557 646774 83609
rect 646826 83597 646832 83609
rect 651760 83597 651766 83609
rect 646826 83569 651766 83597
rect 646826 83557 646832 83569
rect 651760 83557 651766 83569
rect 651818 83557 651824 83609
rect 168208 83483 168214 83535
rect 168266 83523 168272 83535
rect 184432 83523 184438 83535
rect 168266 83495 184438 83523
rect 168266 83483 168272 83495
rect 184432 83483 184438 83495
rect 184490 83483 184496 83535
rect 640720 83483 640726 83535
rect 640778 83523 640784 83535
rect 642256 83523 642262 83535
rect 640778 83495 642262 83523
rect 640778 83483 640784 83495
rect 642256 83483 642262 83495
rect 642314 83483 642320 83535
rect 171280 83409 171286 83461
rect 171338 83449 171344 83461
rect 184336 83449 184342 83461
rect 171338 83421 184342 83449
rect 171338 83409 171344 83421
rect 184336 83409 184342 83421
rect 184394 83409 184400 83461
rect 647920 81855 647926 81907
rect 647978 81895 647984 81907
rect 663280 81895 663286 81907
rect 647978 81867 663286 81895
rect 647978 81855 647984 81867
rect 663280 81855 663286 81867
rect 663338 81855 663344 81907
rect 647824 81781 647830 81833
rect 647882 81821 647888 81833
rect 663376 81821 663382 81833
rect 647882 81793 663382 81821
rect 647882 81781 647888 81793
rect 663376 81781 663382 81793
rect 663434 81781 663440 81833
rect 657040 81633 657046 81685
rect 657098 81673 657104 81685
rect 658576 81673 658582 81685
rect 657098 81645 658582 81673
rect 657098 81633 657104 81645
rect 658576 81633 658582 81645
rect 658634 81633 658640 81685
rect 647728 81559 647734 81611
rect 647786 81599 647792 81611
rect 662416 81599 662422 81611
rect 647786 81571 662422 81599
rect 647786 81559 647792 81571
rect 662416 81559 662422 81571
rect 662474 81559 662480 81611
rect 647920 80745 647926 80797
rect 647978 80785 647984 80797
rect 662512 80785 662518 80797
rect 647978 80757 662518 80785
rect 647978 80745 647984 80757
rect 662512 80745 662518 80757
rect 662570 80745 662576 80797
rect 659440 80671 659446 80723
rect 659498 80711 659504 80723
rect 659536 80711 659542 80723
rect 659498 80683 659542 80711
rect 659498 80671 659504 80683
rect 659536 80671 659542 80683
rect 659594 80671 659600 80723
rect 149584 80597 149590 80649
rect 149642 80637 149648 80649
rect 184432 80637 184438 80649
rect 149642 80609 184438 80637
rect 149642 80597 149648 80609
rect 184432 80597 184438 80609
rect 184490 80597 184496 80649
rect 162448 80523 162454 80575
rect 162506 80563 162512 80575
rect 184528 80563 184534 80575
rect 162506 80535 184534 80563
rect 162506 80523 162512 80535
rect 184528 80523 184534 80535
rect 184586 80523 184592 80575
rect 165232 80449 165238 80501
rect 165290 80489 165296 80501
rect 184336 80489 184342 80501
rect 165290 80461 184342 80489
rect 165290 80449 165296 80461
rect 184336 80449 184342 80461
rect 184394 80449 184400 80501
rect 179920 80375 179926 80427
rect 179978 80415 179984 80427
rect 184624 80415 184630 80427
rect 179978 80387 184630 80415
rect 179978 80375 179984 80387
rect 184624 80375 184630 80387
rect 184682 80375 184688 80427
rect 149296 77711 149302 77763
rect 149354 77751 149360 77763
rect 184432 77751 184438 77763
rect 149354 77723 184438 77751
rect 149354 77711 149360 77723
rect 184432 77711 184438 77723
rect 184490 77711 184496 77763
rect 647152 77711 647158 77763
rect 647210 77751 647216 77763
rect 658288 77751 658294 77763
rect 647210 77723 658294 77751
rect 647210 77711 647216 77723
rect 658288 77711 658294 77723
rect 658346 77711 658352 77763
rect 149392 77637 149398 77689
rect 149450 77677 149456 77689
rect 184528 77677 184534 77689
rect 149450 77649 184534 77677
rect 149450 77637 149456 77649
rect 184528 77637 184534 77649
rect 184586 77637 184592 77689
rect 646576 77637 646582 77689
rect 646634 77677 646640 77689
rect 659440 77677 659446 77689
rect 646634 77649 659446 77677
rect 646634 77637 646640 77649
rect 659440 77637 659446 77649
rect 659498 77637 659504 77689
rect 156496 77563 156502 77615
rect 156554 77603 156560 77615
rect 184624 77603 184630 77615
rect 156554 77575 184630 77603
rect 156554 77563 156560 77575
rect 184624 77563 184630 77575
rect 184682 77563 184688 77615
rect 646672 77563 646678 77615
rect 646730 77603 646736 77615
rect 661744 77603 661750 77615
rect 646730 77575 661750 77603
rect 646730 77563 646736 77575
rect 661744 77563 661750 77575
rect 661802 77563 661808 77615
rect 159760 77489 159766 77541
rect 159818 77529 159824 77541
rect 184336 77529 184342 77541
rect 159818 77501 184342 77529
rect 159818 77489 159824 77501
rect 184336 77489 184342 77501
rect 184394 77489 184400 77541
rect 647920 77489 647926 77541
rect 647978 77529 647984 77541
rect 656944 77529 656950 77541
rect 647978 77501 656950 77529
rect 647978 77489 647984 77501
rect 656944 77489 656950 77501
rect 657002 77489 657008 77541
rect 646000 76083 646006 76135
rect 646058 76123 646064 76135
rect 657520 76123 657526 76135
rect 646058 76095 657526 76123
rect 646058 76083 646064 76095
rect 657520 76083 657526 76095
rect 657578 76083 657584 76135
rect 647056 74899 647062 74951
rect 647114 74939 647120 74951
rect 660112 74939 660118 74951
rect 647114 74911 660118 74939
rect 647114 74899 647120 74911
rect 660112 74899 660118 74911
rect 660170 74899 660176 74951
rect 148816 74825 148822 74877
rect 148874 74865 148880 74877
rect 184528 74865 184534 74877
rect 148874 74837 184534 74865
rect 148874 74825 148880 74837
rect 184528 74825 184534 74837
rect 184586 74825 184592 74877
rect 149104 74751 149110 74803
rect 149162 74791 149168 74803
rect 184624 74791 184630 74803
rect 149162 74763 184630 74791
rect 149162 74751 149168 74763
rect 184624 74751 184630 74763
rect 184682 74751 184688 74803
rect 151120 74677 151126 74729
rect 151178 74717 151184 74729
rect 184432 74717 184438 74729
rect 151178 74689 184438 74717
rect 151178 74677 151184 74689
rect 184432 74677 184438 74689
rect 184490 74677 184496 74729
rect 154096 74603 154102 74655
rect 154154 74643 154160 74655
rect 184336 74643 184342 74655
rect 154154 74615 184342 74643
rect 154154 74603 154160 74615
rect 184336 74603 184342 74615
rect 184394 74603 184400 74655
rect 647920 72161 647926 72213
rect 647978 72201 647984 72213
rect 660688 72201 660694 72213
rect 647978 72173 660694 72201
rect 647978 72161 647984 72173
rect 660688 72161 660694 72173
rect 660746 72161 660752 72213
rect 148432 71939 148438 71991
rect 148490 71979 148496 71991
rect 184432 71979 184438 71991
rect 148490 71951 184438 71979
rect 148490 71939 148496 71951
rect 184432 71939 184438 71951
rect 184490 71939 184496 71991
rect 149680 71865 149686 71917
rect 149738 71905 149744 71917
rect 184528 71905 184534 71917
rect 149738 71877 184534 71905
rect 149738 71865 149744 71877
rect 184528 71865 184534 71877
rect 184586 71865 184592 71917
rect 149584 71791 149590 71843
rect 149642 71831 149648 71843
rect 184336 71831 184342 71843
rect 149642 71803 184342 71831
rect 149642 71791 149648 71803
rect 184336 71791 184342 71803
rect 184394 71791 184400 71843
rect 647920 69571 647926 69623
rect 647978 69611 647984 69623
rect 661456 69611 661462 69623
rect 647978 69583 661462 69611
rect 647978 69571 647984 69583
rect 661456 69571 661462 69583
rect 661514 69571 661520 69623
rect 149584 69053 149590 69105
rect 149642 69093 149648 69105
rect 184528 69093 184534 69105
rect 149642 69065 184534 69093
rect 149642 69053 149648 69065
rect 184528 69053 184534 69065
rect 184586 69053 184592 69105
rect 148912 68979 148918 69031
rect 148970 69019 148976 69031
rect 184336 69019 184342 69031
rect 148970 68991 184342 69019
rect 148970 68979 148976 68991
rect 184336 68979 184342 68991
rect 184394 68979 184400 69031
rect 149200 68905 149206 68957
rect 149258 68945 149264 68957
rect 184432 68945 184438 68957
rect 149258 68917 184438 68945
rect 149258 68905 149264 68917
rect 184432 68905 184438 68917
rect 184490 68905 184496 68957
rect 149296 68831 149302 68883
rect 149354 68871 149360 68883
rect 184336 68871 184342 68883
rect 149354 68843 184342 68871
rect 149354 68831 149360 68843
rect 184336 68831 184342 68843
rect 184394 68831 184400 68883
rect 149104 66167 149110 66219
rect 149162 66207 149168 66219
rect 184528 66207 184534 66219
rect 149162 66179 184534 66207
rect 149162 66167 149168 66179
rect 184528 66167 184534 66179
rect 184586 66167 184592 66219
rect 646000 66167 646006 66219
rect 646058 66207 646064 66219
rect 652336 66207 652342 66219
rect 646058 66179 652342 66207
rect 646058 66167 646064 66179
rect 652336 66167 652342 66179
rect 652394 66167 652400 66219
rect 149392 66093 149398 66145
rect 149450 66133 149456 66145
rect 184624 66133 184630 66145
rect 149450 66105 184630 66133
rect 149450 66093 149456 66105
rect 184624 66093 184630 66105
rect 184682 66093 184688 66145
rect 149488 66019 149494 66071
rect 149546 66059 149552 66071
rect 184432 66059 184438 66071
rect 149546 66031 184438 66059
rect 149546 66019 149552 66031
rect 184432 66019 184438 66031
rect 184490 66019 184496 66071
rect 149008 65945 149014 65997
rect 149066 65985 149072 65997
rect 184336 65985 184342 65997
rect 149066 65957 184342 65985
rect 149066 65945 149072 65957
rect 184336 65945 184342 65957
rect 184394 65945 184400 65997
rect 647920 63577 647926 63629
rect 647978 63617 647984 63629
rect 663184 63617 663190 63629
rect 647978 63589 663190 63617
rect 647978 63577 647984 63589
rect 663184 63577 663190 63589
rect 663242 63577 663248 63629
rect 149200 63281 149206 63333
rect 149258 63321 149264 63333
rect 184432 63321 184438 63333
rect 149258 63293 184438 63321
rect 149258 63281 149264 63293
rect 184432 63281 184438 63293
rect 184490 63281 184496 63333
rect 149488 63207 149494 63259
rect 149546 63247 149552 63259
rect 184528 63247 184534 63259
rect 149546 63219 184534 63247
rect 149546 63207 149552 63219
rect 184528 63207 184534 63219
rect 184586 63207 184592 63259
rect 149392 63133 149398 63185
rect 149450 63173 149456 63185
rect 184624 63173 184630 63185
rect 149450 63145 184630 63173
rect 149450 63133 149456 63145
rect 184624 63133 184630 63145
rect 184682 63133 184688 63185
rect 149584 63059 149590 63111
rect 149642 63099 149648 63111
rect 184336 63099 184342 63111
rect 149642 63071 184342 63099
rect 149642 63059 149648 63071
rect 184336 63059 184342 63071
rect 184394 63059 184400 63111
rect 647920 60987 647926 61039
rect 647978 61027 647984 61039
rect 663472 61027 663478 61039
rect 647978 60999 663478 61027
rect 647978 60987 647984 60999
rect 663472 60987 663478 60999
rect 663530 60987 663536 61039
rect 149296 60395 149302 60447
rect 149354 60435 149360 60447
rect 184432 60435 184438 60447
rect 149354 60407 184438 60435
rect 149354 60395 149360 60407
rect 184432 60395 184438 60407
rect 184490 60395 184496 60447
rect 149488 60321 149494 60373
rect 149546 60361 149552 60373
rect 184528 60361 184534 60373
rect 149546 60333 184534 60361
rect 149546 60321 149552 60333
rect 184528 60321 184534 60333
rect 184586 60321 184592 60373
rect 149392 60247 149398 60299
rect 149450 60287 149456 60299
rect 184336 60287 184342 60299
rect 149450 60259 184342 60287
rect 149450 60247 149456 60259
rect 184336 60247 184342 60259
rect 184394 60247 184400 60299
rect 646000 59063 646006 59115
rect 646058 59103 646064 59115
rect 652240 59103 652246 59115
rect 646058 59075 652246 59103
rect 646058 59063 646064 59075
rect 652240 59063 652246 59075
rect 652298 59063 652304 59115
rect 149392 58989 149398 59041
rect 149450 59029 149456 59041
rect 184336 59029 184342 59041
rect 149450 59001 184342 59029
rect 149450 58989 149456 59001
rect 184336 58989 184342 59001
rect 184394 58989 184400 59041
rect 149392 57509 149398 57561
rect 149450 57549 149456 57561
rect 184336 57549 184342 57561
rect 149450 57521 184342 57549
rect 149450 57509 149456 57521
rect 184336 57509 184342 57521
rect 184394 57509 184400 57561
rect 149392 56177 149398 56229
rect 149450 56217 149456 56229
rect 184432 56217 184438 56229
rect 149450 56189 184438 56217
rect 149450 56177 149456 56189
rect 184432 56177 184438 56189
rect 184490 56177 184496 56229
rect 149488 56103 149494 56155
rect 149546 56143 149552 56155
rect 184336 56143 184342 56155
rect 149546 56115 184342 56143
rect 149546 56103 149552 56115
rect 184336 56103 184342 56115
rect 184394 56103 184400 56155
rect 149680 54623 149686 54675
rect 149738 54663 149744 54675
rect 184336 54663 184342 54675
rect 149738 54635 184342 54663
rect 149738 54623 149744 54635
rect 184336 54623 184342 54635
rect 184394 54623 184400 54675
rect 149392 53217 149398 53269
rect 149450 53257 149456 53269
rect 184336 53257 184342 53269
rect 149450 53229 184342 53257
rect 149450 53217 149456 53229
rect 184336 53217 184342 53229
rect 184394 53217 184400 53269
rect 175600 53143 175606 53195
rect 175658 53183 175664 53195
rect 668272 53183 668278 53195
rect 175658 53155 668278 53183
rect 175658 53143 175664 53155
rect 668272 53143 668278 53155
rect 668330 53143 668336 53195
rect 633616 48999 633622 49051
rect 633674 49039 633680 49051
rect 640720 49039 640726 49051
rect 633674 49011 640726 49039
rect 633674 48999 633680 49011
rect 640720 48999 640726 49011
rect 640778 48999 640784 49051
rect 480976 48111 480982 48163
rect 481034 48151 481040 48163
rect 527920 48151 527926 48163
rect 481034 48123 527926 48151
rect 481034 48111 481040 48123
rect 527920 48111 527926 48123
rect 527978 48111 527984 48163
rect 460336 48037 460342 48089
rect 460394 48077 460400 48089
rect 510352 48077 510358 48089
rect 460394 48049 510358 48077
rect 460394 48037 460400 48049
rect 510352 48037 510358 48049
rect 510410 48037 510416 48089
rect 417520 47963 417526 48015
rect 417578 48003 417584 48015
rect 492976 48003 492982 48015
rect 417578 47975 492982 48003
rect 417578 47963 417584 47975
rect 492976 47963 492982 47975
rect 493034 47963 493040 48015
rect 311056 47889 311062 47941
rect 311114 47929 311120 47941
rect 371920 47929 371926 47941
rect 311114 47901 371926 47929
rect 311114 47889 311120 47901
rect 371920 47889 371926 47901
rect 371978 47889 371984 47941
rect 405520 47889 405526 47941
rect 405578 47929 405584 47941
rect 441328 47929 441334 47941
rect 405578 47901 441334 47929
rect 405578 47889 405584 47901
rect 441328 47889 441334 47901
rect 441386 47889 441392 47941
rect 472240 47889 472246 47941
rect 472298 47929 472304 47941
rect 562480 47929 562486 47941
rect 472298 47901 562486 47929
rect 472298 47889 472304 47901
rect 562480 47889 562486 47901
rect 562538 47889 562544 47941
rect 302896 47815 302902 47867
rect 302954 47855 302960 47867
rect 506800 47855 506806 47867
rect 302954 47827 506806 47855
rect 302954 47815 302960 47827
rect 506800 47815 506806 47827
rect 506858 47815 506864 47867
rect 320176 47741 320182 47793
rect 320234 47781 320240 47793
rect 529264 47781 529270 47793
rect 320234 47753 529270 47781
rect 320234 47741 320240 47753
rect 529264 47741 529270 47753
rect 529322 47741 529328 47793
rect 233680 47667 233686 47719
rect 233738 47707 233744 47719
rect 475504 47707 475510 47719
rect 233738 47679 475510 47707
rect 233738 47667 233744 47679
rect 475504 47667 475510 47679
rect 475562 47667 475568 47719
rect 268528 47593 268534 47645
rect 268586 47633 268592 47645
rect 520624 47633 520630 47645
rect 268586 47605 520630 47633
rect 268586 47593 268592 47605
rect 520624 47593 520630 47605
rect 520682 47593 520688 47645
rect 250960 47519 250966 47571
rect 251018 47559 251024 47571
rect 521200 47559 521206 47571
rect 251018 47531 521206 47559
rect 251018 47519 251024 47531
rect 521200 47519 521206 47531
rect 521258 47519 521264 47571
rect 418864 47445 418870 47497
rect 418922 47485 418928 47497
rect 424048 47485 424054 47497
rect 418922 47457 424054 47485
rect 418922 47445 418928 47457
rect 424048 47445 424054 47457
rect 424106 47445 424112 47497
rect 145360 47075 145366 47127
rect 145418 47115 145424 47127
rect 199120 47115 199126 47127
rect 145418 47087 199126 47115
rect 145418 47075 145424 47087
rect 199120 47075 199126 47087
rect 199178 47075 199184 47127
rect 331216 46557 331222 46609
rect 331274 46597 331280 46609
rect 337456 46597 337462 46609
rect 331274 46569 337462 46597
rect 331274 46557 331280 46569
rect 337456 46557 337462 46569
rect 337514 46557 337520 46609
rect 464848 46409 464854 46461
rect 464906 46449 464912 46461
rect 475696 46449 475702 46461
rect 464906 46421 475702 46449
rect 464906 46409 464912 46421
rect 475696 46409 475702 46421
rect 475754 46409 475760 46461
rect 539728 46187 539734 46239
rect 539786 46227 539792 46239
rect 545200 46227 545206 46239
rect 539786 46199 545206 46227
rect 539786 46187 539792 46199
rect 545200 46187 545206 46199
rect 545258 46187 545264 46239
rect 207376 46113 207382 46165
rect 207434 46153 207440 46165
rect 216400 46153 216406 46165
rect 207434 46125 216406 46153
rect 207434 46113 207440 46125
rect 216400 46113 216406 46125
rect 216458 46113 216464 46165
rect 402160 46113 402166 46165
rect 402218 46153 402224 46165
rect 406768 46153 406774 46165
rect 402218 46125 406774 46153
rect 402218 46113 402224 46125
rect 406768 46113 406774 46125
rect 406826 46113 406832 46165
rect 506800 44855 506806 44907
rect 506858 44895 506864 44907
rect 512176 44895 512182 44907
rect 506858 44867 512182 44895
rect 506858 44855 506864 44867
rect 512176 44855 512182 44867
rect 512234 44855 512240 44907
rect 175600 44140 175606 44192
rect 175658 44140 175664 44192
rect 285808 43227 285814 43279
rect 285866 43267 285872 43279
rect 518704 43267 518710 43279
rect 285866 43239 518710 43267
rect 285866 43227 285872 43239
rect 518704 43227 518710 43239
rect 518762 43227 518768 43279
rect 629008 43227 629014 43279
rect 629066 43267 629072 43279
rect 633616 43267 633622 43279
rect 629066 43239 633622 43267
rect 629066 43227 629072 43239
rect 633616 43227 633622 43239
rect 633674 43227 633680 43279
rect 403504 43153 403510 43205
rect 403562 43193 403568 43205
rect 418864 43193 418870 43205
rect 403562 43165 418870 43193
rect 403562 43153 403568 43165
rect 418864 43153 418870 43165
rect 418922 43153 418928 43205
rect 444880 43153 444886 43205
rect 444938 43193 444944 43205
rect 458608 43193 458614 43205
rect 444938 43165 458614 43193
rect 444938 43153 444944 43165
rect 458608 43153 458614 43165
rect 458666 43153 458672 43205
rect 302896 42117 302902 42169
rect 302954 42157 302960 42169
rect 311152 42157 311158 42169
rect 302954 42129 311158 42157
rect 302954 42117 302960 42129
rect 311152 42117 311158 42129
rect 311210 42117 311216 42169
rect 357712 42117 357718 42169
rect 357770 42157 357776 42169
rect 357770 42129 377294 42157
rect 357770 42117 357776 42129
rect 307216 42043 307222 42095
rect 307274 42083 307280 42095
rect 311056 42083 311062 42095
rect 307274 42055 311062 42083
rect 307274 42043 307280 42055
rect 311056 42043 311062 42055
rect 311114 42043 311120 42095
rect 335440 42043 335446 42095
rect 335498 42083 335504 42095
rect 354832 42083 354838 42095
rect 335498 42055 354838 42083
rect 335498 42043 335504 42055
rect 354832 42043 354838 42055
rect 354890 42043 354896 42095
rect 362032 42043 362038 42095
rect 362090 42083 362096 42095
rect 365968 42083 365974 42095
rect 362090 42055 365974 42083
rect 362090 42043 362096 42055
rect 365968 42043 365974 42055
rect 366026 42043 366032 42095
rect 377266 42083 377294 42129
rect 402160 42083 402166 42095
rect 377266 42055 402166 42083
rect 402160 42043 402166 42055
rect 402218 42043 402224 42095
rect 471664 42043 471670 42095
rect 471722 42083 471728 42095
rect 480976 42083 480982 42095
rect 471722 42055 480982 42083
rect 471722 42043 471728 42055
rect 480976 42043 480982 42055
rect 481034 42043 481040 42095
rect 186256 41969 186262 42021
rect 186314 42009 186320 42021
rect 187024 42009 187030 42021
rect 186314 41981 187030 42009
rect 186314 41969 186320 41981
rect 187024 41969 187030 41981
rect 187082 41969 187088 42021
rect 194320 41969 194326 42021
rect 194378 42009 194384 42021
rect 629008 42009 629014 42021
rect 194378 41981 629014 42009
rect 194378 41969 194384 41981
rect 629008 41969 629014 41981
rect 629066 41969 629072 42021
rect 514000 41747 514006 41799
rect 514058 41787 514064 41799
rect 514864 41787 514870 41799
rect 514058 41759 514870 41787
rect 514058 41747 514064 41759
rect 514864 41747 514870 41759
rect 514922 41747 514928 41799
rect 186256 41451 186262 41503
rect 186314 41491 186320 41503
rect 207376 41491 207382 41503
rect 186314 41463 207382 41491
rect 186314 41451 186320 41463
rect 207376 41451 207382 41463
rect 207434 41451 207440 41503
rect 403504 37495 403510 37507
rect 397426 37467 403510 37495
rect 365872 37381 365878 37433
rect 365930 37421 365936 37433
rect 397426 37421 397454 37467
rect 403504 37455 403510 37467
rect 403562 37455 403568 37507
rect 365930 37393 397454 37421
rect 365930 37381 365936 37393
rect 475504 37381 475510 37433
rect 475562 37421 475568 37433
rect 514000 37421 514006 37433
rect 475562 37393 514006 37421
rect 475562 37381 475568 37393
rect 514000 37381 514006 37393
rect 514058 37381 514064 37433
rect 365968 37307 365974 37359
rect 366026 37347 366032 37359
rect 389200 37347 389206 37359
rect 366026 37319 389206 37347
rect 366026 37307 366032 37319
rect 389200 37307 389206 37319
rect 389258 37307 389264 37359
rect 420784 34495 420790 34547
rect 420842 34535 420848 34547
rect 444880 34535 444886 34547
rect 420842 34507 444886 34535
rect 420842 34495 420848 34507
rect 444880 34495 444886 34507
rect 444938 34495 444944 34547
rect 328336 31609 328342 31661
rect 328394 31649 328400 31661
rect 335440 31649 335446 31661
rect 328394 31621 335446 31649
rect 328394 31609 328400 31621
rect 335440 31609 335446 31621
rect 335498 31609 335504 31661
<< via1 >>
rect 181462 1002267 181514 1002319
rect 184054 1002267 184106 1002319
rect 482614 1002267 482666 1002319
rect 483862 1002267 483914 1002319
rect 181366 992203 181418 992255
rect 184246 992203 184298 992255
rect 535702 992129 535754 992181
rect 538582 992129 538634 992181
rect 394582 991463 394634 991515
rect 397462 991463 397514 991515
rect 240886 982953 240938 983005
rect 241942 982953 241994 983005
rect 391606 982879 391658 982931
rect 649462 982879 649514 982931
rect 394582 982805 394634 982857
rect 656662 982953 656714 983005
rect 649462 981991 649514 982043
rect 652246 981991 652298 982043
rect 656662 979253 656714 979305
rect 679702 979253 679754 979305
rect 652246 979179 652298 979231
rect 677590 979179 677642 979231
rect 677494 967635 677546 967687
rect 679702 967635 679754 967687
rect 40150 959051 40202 959103
rect 60022 959051 60074 959103
rect 653782 950319 653834 950371
rect 676822 950319 676874 950371
rect 655414 892969 655466 893021
rect 676150 892969 676202 893021
rect 655222 892895 655274 892947
rect 676246 892895 676298 892947
rect 655126 892821 655178 892873
rect 676054 892821 676106 892873
rect 673366 892377 673418 892429
rect 676054 892377 676106 892429
rect 670966 891415 671018 891467
rect 676054 891415 676106 891467
rect 670870 890379 670922 890431
rect 676054 890379 676106 890431
rect 673942 887863 673994 887915
rect 676246 887863 676298 887915
rect 674134 887123 674186 887175
rect 676054 887123 676106 887175
rect 674230 887049 674282 887101
rect 676246 887049 676298 887101
rect 674038 885051 674090 885103
rect 676054 885051 676106 885103
rect 674518 884237 674570 884289
rect 676054 884237 676106 884289
rect 674422 883571 674474 883623
rect 676054 883571 676106 883623
rect 675286 883201 675338 883253
rect 679990 883201 680042 883253
rect 675094 883127 675146 883179
rect 680182 883127 680234 883179
rect 674998 883053 675050 883105
rect 676054 883053 676106 883105
rect 674998 882831 675050 882883
rect 679702 882831 679754 882883
rect 649462 881425 649514 881477
rect 679702 881425 679754 881477
rect 655318 881351 655370 881403
rect 675478 881351 675530 881403
rect 674326 881203 674378 881255
rect 680086 881203 680138 881255
rect 674614 880093 674666 880145
rect 679798 880093 679850 880145
rect 675190 879501 675242 879553
rect 679894 879501 679946 879553
rect 674902 878317 674954 878369
rect 675766 878317 675818 878369
rect 674998 877207 675050 877259
rect 675478 877207 675530 877259
rect 675190 876615 675242 876667
rect 675190 876171 675242 876223
rect 674230 876097 674282 876149
rect 675094 876097 675146 876149
rect 674518 875431 674570 875483
rect 674998 875431 675050 875483
rect 673942 875209 673994 875261
rect 674422 875209 674474 875261
rect 674326 874913 674378 874965
rect 675478 874913 675530 874965
rect 674614 874247 674666 874299
rect 675478 874247 675530 874299
rect 675190 873507 675242 873559
rect 675382 873507 675434 873559
rect 674902 872915 674954 872967
rect 675382 872915 675434 872967
rect 654166 872619 654218 872671
rect 674614 872619 674666 872671
rect 674518 869807 674570 869859
rect 675382 869807 675434 869859
rect 674134 868105 674186 868157
rect 674998 868105 675050 868157
rect 674614 868031 674666 868083
rect 675094 868031 675146 868083
rect 674038 867365 674090 867417
rect 675478 867365 675530 867417
rect 674422 865737 674474 865789
rect 675190 865737 675242 865789
rect 653782 863961 653834 864013
rect 675094 863961 675146 864013
rect 41782 817933 41834 817985
rect 47446 817933 47498 817985
rect 41782 817267 41834 817319
rect 44854 817267 44906 817319
rect 41590 816527 41642 816579
rect 44950 816527 45002 816579
rect 41782 815787 41834 815839
rect 43222 815787 43274 815839
rect 41782 814825 41834 814877
rect 44662 814825 44714 814877
rect 41590 813567 41642 813619
rect 44758 813567 44810 813619
rect 41590 812383 41642 812435
rect 42934 812383 42986 812435
rect 41590 809867 41642 809919
rect 42838 809867 42890 809919
rect 41782 809793 41834 809845
rect 42742 809793 42794 809845
rect 41782 808609 41834 808661
rect 43126 808609 43178 808661
rect 41782 807351 41834 807403
rect 42646 807351 42698 807403
rect 41590 806611 41642 806663
rect 43030 806611 43082 806663
rect 41590 805131 41642 805183
rect 44566 805131 44618 805183
rect 42838 800765 42890 800817
rect 43510 800765 43562 800817
rect 42742 800691 42794 800743
rect 57718 800691 57770 800743
rect 42838 800617 42890 800669
rect 57622 800617 57674 800669
rect 41878 800173 41930 800225
rect 42166 800173 42218 800225
rect 43318 800173 43370 800225
rect 41878 799951 41930 800003
rect 42166 798101 42218 798153
rect 42550 798101 42602 798153
rect 42646 797879 42698 797931
rect 42070 797287 42122 797339
rect 42742 797287 42794 797339
rect 42742 796843 42794 796895
rect 42166 796251 42218 796303
rect 43126 796251 43178 796303
rect 43222 796251 43274 796303
rect 43222 796029 43274 796081
rect 42070 795585 42122 795637
rect 42838 795585 42890 795637
rect 42166 794771 42218 794823
rect 43030 794771 43082 794823
rect 43030 794623 43082 794675
rect 43510 794623 43562 794675
rect 42166 793587 42218 793639
rect 42742 793587 42794 793639
rect 42934 792107 42986 792159
rect 43510 792107 43562 792159
rect 655126 792033 655178 792085
rect 675382 792033 675434 792085
rect 42166 790627 42218 790679
rect 43126 790627 43178 790679
rect 43126 790479 43178 790531
rect 43510 790479 43562 790531
rect 42166 789443 42218 789495
rect 42742 789443 42794 789495
rect 42934 789147 42986 789199
rect 58198 789147 58250 789199
rect 44950 789073 45002 789125
rect 58390 789073 58442 789125
rect 42166 788703 42218 788755
rect 43030 788703 43082 788755
rect 42166 786853 42218 786905
rect 43126 786853 43178 786905
rect 42166 786409 42218 786461
rect 42742 786409 42794 786461
rect 42070 785595 42122 785647
rect 42838 785595 42890 785647
rect 44854 785521 44906 785573
rect 59158 785521 59210 785573
rect 47446 785373 47498 785425
rect 59638 785373 59690 785425
rect 42166 785003 42218 785055
rect 42934 785003 42986 785055
rect 656566 783449 656618 783501
rect 674998 783449 675050 783501
rect 654358 780489 654410 780541
rect 675286 780489 675338 780541
rect 674998 778861 675050 778913
rect 675382 778861 675434 778913
rect 673078 778713 673130 778765
rect 675478 778713 675530 778765
rect 41782 774643 41834 774695
rect 47542 774643 47594 774695
rect 41590 773903 41642 773955
rect 44854 773903 44906 773955
rect 674518 773607 674570 773659
rect 675286 773607 675338 773659
rect 41590 773311 41642 773363
rect 44950 773311 45002 773363
rect 41782 773237 41834 773289
rect 43414 773237 43466 773289
rect 41782 772571 41834 772623
rect 43318 772571 43370 772623
rect 42742 771905 42794 771957
rect 62038 771905 62090 771957
rect 41590 771831 41642 771883
rect 61846 771831 61898 771883
rect 41782 768131 41834 768183
rect 42838 768131 42890 768183
rect 41782 765097 41834 765149
rect 42934 765097 42986 765149
rect 41782 764135 41834 764187
rect 43030 764135 43082 764187
rect 41590 763395 41642 763447
rect 43126 763395 43178 763447
rect 41782 762063 41834 762115
rect 47446 762063 47498 762115
rect 42934 757623 42986 757675
rect 43222 757623 43274 757675
rect 42934 757475 42986 757527
rect 58678 757475 58730 757527
rect 41398 757327 41450 757379
rect 43606 757327 43658 757379
rect 41494 757253 41546 757305
rect 43510 757253 43562 757305
rect 41878 756957 41930 757009
rect 41878 756735 41930 756787
rect 42166 754219 42218 754271
rect 42934 754219 42986 754271
rect 42070 753035 42122 753087
rect 42358 753035 42410 753087
rect 42358 752887 42410 752939
rect 43030 752887 43082 752939
rect 42070 751777 42122 751829
rect 43222 751777 43274 751829
rect 42070 751481 42122 751533
rect 42934 751481 42986 751533
rect 42070 751111 42122 751163
rect 43126 751111 43178 751163
rect 43126 750963 43178 751015
rect 43510 750963 43562 751015
rect 42166 750593 42218 750645
rect 42358 750593 42410 750645
rect 42070 749779 42122 749831
rect 42934 749779 42986 749831
rect 42934 749631 42986 749683
rect 43606 749631 43658 749683
rect 655702 748817 655754 748869
rect 675382 748817 675434 748869
rect 42070 746079 42122 746131
rect 43126 746079 43178 746131
rect 43126 745931 43178 745983
rect 54646 745931 54698 745983
rect 54742 745931 54794 745983
rect 57622 745931 57674 745983
rect 42166 745487 42218 745539
rect 42454 745487 42506 745539
rect 43222 745265 43274 745317
rect 59638 745265 59690 745317
rect 44950 745117 45002 745169
rect 58198 745117 58250 745169
rect 42166 743563 42218 743615
rect 43030 743563 43082 743615
rect 42070 743193 42122 743245
rect 42934 743193 42986 743245
rect 47542 742971 47594 743023
rect 59638 742971 59690 743023
rect 44854 742897 44906 742949
rect 59734 742897 59786 742949
rect 42166 742601 42218 742653
rect 42454 742601 42506 742653
rect 674422 742083 674474 742135
rect 675190 742083 675242 742135
rect 42166 741935 42218 741987
rect 43126 741935 43178 741987
rect 673174 738235 673226 738287
rect 675382 738235 675434 738287
rect 672118 737569 672170 737621
rect 675286 737569 675338 737621
rect 654070 737421 654122 737473
rect 675286 737421 675338 737473
rect 654166 737347 654218 737399
rect 674614 737347 674666 737399
rect 672886 734757 672938 734809
rect 675382 734757 675434 734809
rect 672310 734387 672362 734439
rect 675382 734387 675434 734439
rect 672406 734165 672458 734217
rect 675382 734165 675434 734217
rect 675190 733869 675242 733921
rect 675478 733869 675530 733921
rect 672790 732315 672842 732367
rect 675478 732315 675530 732367
rect 674614 732019 674666 732071
rect 675382 732019 675434 732071
rect 41782 731427 41834 731479
rect 47638 731427 47690 731479
rect 41590 730687 41642 730739
rect 44854 730687 44906 730739
rect 674422 730465 674474 730517
rect 675478 730465 675530 730517
rect 41782 730317 41834 730369
rect 44950 730317 45002 730369
rect 41590 730169 41642 730221
rect 43318 730169 43370 730221
rect 41590 729207 41642 729259
rect 43894 729207 43946 729259
rect 41782 728763 41834 728815
rect 43798 728763 43850 728815
rect 40438 728689 40490 728741
rect 62230 728689 62282 728741
rect 41398 728615 41450 728667
rect 62422 728615 62474 728667
rect 674230 728615 674282 728667
rect 675478 728615 675530 728667
rect 41782 727875 41834 727927
rect 43702 727875 43754 727927
rect 41878 722917 41930 722969
rect 42934 722917 42986 722969
rect 41590 720401 41642 720453
rect 43030 720401 43082 720453
rect 41590 720179 41642 720231
rect 43126 720179 43178 720231
rect 41590 718699 41642 718751
rect 47542 718699 47594 718751
rect 655606 714703 655658 714755
rect 676246 714703 676298 714755
rect 655414 714555 655466 714607
rect 676342 714555 676394 714607
rect 655222 714407 655274 714459
rect 676150 714407 676202 714459
rect 43222 714259 43274 714311
rect 59638 714259 59690 714311
rect 673366 714185 673418 714237
rect 676054 714185 676106 714237
rect 41686 714037 41738 714089
rect 43510 714037 43562 714089
rect 42166 713889 42218 713941
rect 43414 713889 43466 713941
rect 41782 713815 41834 713867
rect 41782 713519 41834 713571
rect 672694 713371 672746 713423
rect 676246 713371 676298 713423
rect 669718 713075 669770 713127
rect 670966 713075 671018 713127
rect 676054 713075 676106 713127
rect 670678 712631 670730 712683
rect 676054 712631 676106 712683
rect 42454 711965 42506 712017
rect 43222 711965 43274 712017
rect 669526 711891 669578 711943
rect 670870 711891 670922 711943
rect 676246 711891 676298 711943
rect 43222 711817 43274 711869
rect 43798 711817 43850 711869
rect 43030 711521 43082 711573
rect 43414 711521 43466 711573
rect 670774 711521 670826 711573
rect 676054 711521 676106 711573
rect 43414 711373 43466 711425
rect 43894 711373 43946 711425
rect 674902 711299 674954 711351
rect 676054 711299 676106 711351
rect 43030 711151 43082 711203
rect 43606 711077 43658 711129
rect 674518 711077 674570 711129
rect 676054 711077 676106 711129
rect 42166 710855 42218 710907
rect 42454 710855 42506 710907
rect 42166 709893 42218 709945
rect 43510 709893 43562 709945
rect 42070 708487 42122 708539
rect 43510 708487 43562 708539
rect 674998 708413 675050 708465
rect 676054 708413 676106 708465
rect 42070 708339 42122 708391
rect 43126 708339 43178 708391
rect 43126 708191 43178 708243
rect 43606 708191 43658 708243
rect 42166 708043 42218 708095
rect 42934 708043 42986 708095
rect 42166 706563 42218 706615
rect 43126 706563 43178 706615
rect 42934 706415 42986 706467
rect 43126 706415 43178 706467
rect 42454 704935 42506 704987
rect 42166 704269 42218 704321
rect 673078 704861 673130 704913
rect 676246 704861 676298 704913
rect 42070 703677 42122 703729
rect 43030 703677 43082 703729
rect 653782 702789 653834 702841
rect 675382 702789 675434 702841
rect 649462 702715 649514 702767
rect 679990 702715 680042 702767
rect 42166 702641 42218 702693
rect 42358 702641 42410 702693
rect 43510 702641 43562 702693
rect 58774 702641 58826 702693
rect 44950 702567 45002 702619
rect 58678 702567 58730 702619
rect 42166 702271 42218 702323
rect 43126 702271 43178 702323
rect 42070 700495 42122 700547
rect 43030 700495 43082 700547
rect 47638 699755 47690 699807
rect 59254 699755 59306 699807
rect 44854 699681 44906 699733
rect 58870 699681 58922 699733
rect 42166 699385 42218 699437
rect 42934 699385 42986 699437
rect 42070 698719 42122 698771
rect 45238 698719 45290 698771
rect 654166 694131 654218 694183
rect 674998 694131 675050 694183
rect 672598 693613 672650 693665
rect 675478 693613 675530 693665
rect 673078 692873 673130 692925
rect 675382 692873 675434 692925
rect 654070 691319 654122 691371
rect 675190 691319 675242 691371
rect 674902 690431 674954 690483
rect 675478 690431 675530 690483
rect 672982 689765 673034 689817
rect 675382 689765 675434 689817
rect 672022 689321 672074 689373
rect 675382 689321 675434 689373
rect 672214 689099 672266 689151
rect 675382 689099 675434 689151
rect 674998 688877 675050 688929
rect 675478 688877 675530 688929
rect 41782 688211 41834 688263
rect 50326 688211 50378 688263
rect 41590 687471 41642 687523
rect 47734 687471 47786 687523
rect 672502 687323 672554 687375
rect 675478 687323 675530 687375
rect 41782 687175 41834 687227
rect 45046 687175 45098 687227
rect 675190 687027 675242 687079
rect 675478 687027 675530 687079
rect 41590 686953 41642 687005
rect 43414 686953 43466 687005
rect 41590 685991 41642 686043
rect 43510 685991 43562 686043
rect 674326 685473 674378 685525
rect 675478 685473 675530 685525
rect 41782 685325 41834 685377
rect 43222 685325 43274 685377
rect 44950 685325 45002 685377
rect 41782 684141 41834 684193
rect 43318 684141 43370 684193
rect 44854 684141 44906 684193
rect 674518 683623 674570 683675
rect 675478 683623 675530 683675
rect 41782 683031 41834 683083
rect 42934 683031 42986 683083
rect 41590 677259 41642 677311
rect 43126 677259 43178 677311
rect 41590 676963 41642 677015
rect 43030 676963 43082 677015
rect 41590 675483 41642 675535
rect 47638 675483 47690 675535
rect 34486 672449 34538 672501
rect 40342 672449 40394 672501
rect 37366 671265 37418 671317
rect 43702 671265 43754 671317
rect 39862 671191 39914 671243
rect 43606 671191 43658 671243
rect 40342 671117 40394 671169
rect 43318 671117 43370 671169
rect 42742 671043 42794 671095
rect 59638 671043 59690 671095
rect 43510 670969 43562 671021
rect 41686 670821 41738 670873
rect 42838 670821 42890 670873
rect 43030 670821 43082 670873
rect 43318 670821 43370 670873
rect 42262 670747 42314 670799
rect 42070 670673 42122 670725
rect 43126 670673 43178 670725
rect 43414 670673 43466 670725
rect 43510 670673 43562 670725
rect 41782 670599 41834 670651
rect 41878 670599 41930 670651
rect 43030 670599 43082 670651
rect 41782 670303 41834 670355
rect 672694 669193 672746 669245
rect 676054 669193 676106 669245
rect 42166 668527 42218 668579
rect 42934 668527 42986 668579
rect 655510 668527 655562 668579
rect 676150 668527 676202 668579
rect 673270 668453 673322 668505
rect 676054 668453 676106 668505
rect 42934 668379 42986 668431
rect 43222 668379 43274 668431
rect 655318 668379 655370 668431
rect 676246 668379 676298 668431
rect 655126 668157 655178 668209
rect 676342 668157 676394 668209
rect 674422 668083 674474 668135
rect 676054 668083 676106 668135
rect 670678 668009 670730 668061
rect 675958 668009 676010 668061
rect 42166 667861 42218 667913
rect 42742 667861 42794 667913
rect 42742 667713 42794 667765
rect 43318 667713 43370 667765
rect 670774 667639 670826 667691
rect 675958 667639 676010 667691
rect 652246 666751 652298 666803
rect 670870 666751 670922 666803
rect 676246 666751 676298 666803
rect 42166 666677 42218 666729
rect 42934 666677 42986 666729
rect 649750 666677 649802 666729
rect 670678 666677 670730 666729
rect 42934 666529 42986 666581
rect 43414 666529 43466 666581
rect 670966 666307 671018 666359
rect 676246 666307 676298 666359
rect 42166 665271 42218 665323
rect 43222 665271 43274 665323
rect 674230 665197 674282 665249
rect 676054 665197 676106 665249
rect 42166 665123 42218 665175
rect 42742 665123 42794 665175
rect 42166 664827 42218 664879
rect 43126 664827 43178 664879
rect 43126 664679 43178 664731
rect 43606 664679 43658 664731
rect 42070 664161 42122 664213
rect 42838 664161 42890 664213
rect 42166 663347 42218 663399
rect 43030 663347 43082 663399
rect 43030 663199 43082 663251
rect 43702 663199 43754 663251
rect 672118 662089 672170 662141
rect 676054 662089 676106 662141
rect 672790 661645 672842 661697
rect 676054 661645 676106 661697
rect 672310 661349 672362 661401
rect 676246 661349 676298 661401
rect 42070 660905 42122 660957
rect 42934 660905 42986 660957
rect 673174 660609 673226 660661
rect 676054 660609 676106 660661
rect 42070 660387 42122 660439
rect 43126 660387 43178 660439
rect 672886 660165 672938 660217
rect 676054 660165 676106 660217
rect 672406 659869 672458 659921
rect 676246 659869 676298 659921
rect 42166 659647 42218 659699
rect 43030 659647 43082 659699
rect 43222 659425 43274 659477
rect 58774 659425 58826 659477
rect 45046 659351 45098 659403
rect 58678 659351 58730 659403
rect 42166 659203 42218 659255
rect 43798 659203 43850 659255
rect 42070 657353 42122 657405
rect 42742 657353 42794 657405
rect 654166 656761 654218 656813
rect 675382 656761 675434 656813
rect 42166 656687 42218 656739
rect 42838 656687 42890 656739
rect 649558 656687 649610 656739
rect 679798 656687 679850 656739
rect 50326 656613 50378 656665
rect 58198 656613 58250 656665
rect 47734 656539 47786 656591
rect 58390 656539 58442 656591
rect 42166 656169 42218 656221
rect 42934 656169 42986 656221
rect 42166 655503 42218 655555
rect 43030 655503 43082 655555
rect 670870 648917 670922 648969
rect 675190 648917 675242 648969
rect 672406 648251 672458 648303
rect 675190 648251 675242 648303
rect 655798 648177 655850 648229
rect 674998 648177 675050 648229
rect 673366 648029 673418 648081
rect 675190 648029 675242 648081
rect 655990 645143 656042 645195
rect 675286 645143 675338 645195
rect 41590 644847 41642 644899
rect 50326 644847 50378 644899
rect 672886 644773 672938 644825
rect 675382 644773 675434 644825
rect 41590 644255 41642 644307
rect 47830 644255 47882 644307
rect 672790 644033 672842 644085
rect 675478 644033 675530 644085
rect 41782 643959 41834 644011
rect 47926 643959 47978 644011
rect 41590 643737 41642 643789
rect 43510 643737 43562 643789
rect 674998 643663 675050 643715
rect 675382 643663 675434 643715
rect 672694 643589 672746 643641
rect 675478 643589 675530 643641
rect 41590 642775 41642 642827
rect 43606 642775 43658 642827
rect 41494 642479 41546 642531
rect 61942 642479 61994 642531
rect 670678 642257 670730 642309
rect 675478 642257 675530 642309
rect 41590 641295 41642 641347
rect 43510 641295 43562 641347
rect 41590 634487 41642 634539
rect 43126 634487 43178 634539
rect 41782 634191 41834 634243
rect 42934 634191 42986 634243
rect 41590 634117 41642 634169
rect 43030 634117 43082 634169
rect 41782 633895 41834 633947
rect 42838 633895 42890 633947
rect 41590 632267 41642 632319
rect 47734 632267 47786 632319
rect 41974 632045 42026 632097
rect 42742 632045 42794 632097
rect 40150 630639 40202 630691
rect 42070 630639 42122 630691
rect 34390 629233 34442 629285
rect 40438 629233 40490 629285
rect 37366 627901 37418 627953
rect 43702 627901 43754 627953
rect 40438 627827 40490 627879
rect 43222 627827 43274 627879
rect 41878 627383 41930 627435
rect 42262 627383 42314 627435
rect 43318 627383 43370 627435
rect 41878 627161 41930 627213
rect 42166 625311 42218 625363
rect 42742 625311 42794 625363
rect 655414 624941 655466 624993
rect 676246 624941 676298 624993
rect 42166 623979 42218 624031
rect 58966 623979 59018 624031
rect 673270 623979 673322 624031
rect 676054 623979 676106 624031
rect 42166 623461 42218 623513
rect 42934 623461 42986 623513
rect 672310 623387 672362 623439
rect 676054 623387 676106 623439
rect 42934 623313 42986 623365
rect 43318 623313 43370 623365
rect 669622 622943 669674 622995
rect 670774 622943 670826 622995
rect 676054 622943 676106 622995
rect 670582 622425 670634 622477
rect 676054 622425 676106 622477
rect 655606 622351 655658 622403
rect 676246 622351 676298 622403
rect 42166 622203 42218 622255
rect 42838 622203 42890 622255
rect 655222 622203 655274 622255
rect 676150 622203 676202 622255
rect 42070 622055 42122 622107
rect 48022 622055 48074 622107
rect 674326 621981 674378 622033
rect 676246 621981 676298 622033
rect 670966 621907 671018 621959
rect 676054 621907 676106 621959
rect 42166 621611 42218 621663
rect 43126 621611 43178 621663
rect 670486 621315 670538 621367
rect 676054 621315 676106 621367
rect 42070 620945 42122 620997
rect 43030 620945 43082 620997
rect 43222 620353 43274 620405
rect 43606 620353 43658 620405
rect 42166 620131 42218 620183
rect 42742 620131 42794 620183
rect 669814 619835 669866 619887
rect 670966 619835 671018 619887
rect 674902 619021 674954 619073
rect 676054 619021 676106 619073
rect 674518 618873 674570 618925
rect 676246 618873 676298 618925
rect 42070 617837 42122 617889
rect 43030 617837 43082 617889
rect 43030 617689 43082 617741
rect 43606 617689 43658 617741
rect 42166 617171 42218 617223
rect 42934 617171 42986 617223
rect 672598 617097 672650 617149
rect 676246 617097 676298 617149
rect 42166 616653 42218 616705
rect 43126 616653 43178 616705
rect 672502 616505 672554 616557
rect 676054 616505 676106 616557
rect 42934 616357 42986 616409
rect 58198 616357 58250 616409
rect 47926 616283 47978 616335
rect 58966 616283 59018 616335
rect 48022 616209 48074 616261
rect 59638 616209 59690 616261
rect 672022 615913 672074 615965
rect 676054 615913 676106 615965
rect 42166 615839 42218 615891
rect 42838 615839 42890 615891
rect 673078 615617 673130 615669
rect 676246 615617 676298 615669
rect 672982 615173 673034 615225
rect 676246 615173 676298 615225
rect 672214 614433 672266 614485
rect 676054 614433 676106 614485
rect 42166 614137 42218 614189
rect 43030 614137 43082 614189
rect 42166 613619 42218 613671
rect 42742 613619 42794 613671
rect 655798 613471 655850 613523
rect 675382 613471 675434 613523
rect 50326 613397 50378 613449
rect 59638 613397 59690 613449
rect 47830 613323 47882 613375
rect 59542 613323 59594 613375
rect 42070 612805 42122 612857
rect 42358 612805 42410 612857
rect 42166 612139 42218 612191
rect 42934 612139 42986 612191
rect 649654 610585 649706 610637
rect 679990 610585 680042 610637
rect 670966 606885 671018 606937
rect 675190 606885 675242 606937
rect 670774 603851 670826 603903
rect 675286 603851 675338 603903
rect 673270 603037 673322 603089
rect 675382 603037 675434 603089
rect 656566 602149 656618 602201
rect 674902 602149 674954 602201
rect 653974 602001 654026 602053
rect 674998 602001 675050 602053
rect 673174 601927 673226 601979
rect 675286 601927 675338 601979
rect 41590 601631 41642 601683
rect 50326 601631 50378 601683
rect 41782 601335 41834 601387
rect 47830 601335 47882 601387
rect 41782 600743 41834 600795
rect 47926 600743 47978 600795
rect 41782 600373 41834 600425
rect 43222 600373 43274 600425
rect 41782 599781 41834 599833
rect 43222 599781 43274 599833
rect 672982 599781 673034 599833
rect 675382 599781 675434 599833
rect 41782 599263 41834 599315
rect 43414 599263 43466 599315
rect 673078 599263 673130 599315
rect 675382 599263 675434 599315
rect 672598 598893 672650 598945
rect 675382 598893 675434 598945
rect 674998 598671 675050 598723
rect 675478 598671 675530 598723
rect 41782 598301 41834 598353
rect 43894 598301 43946 598353
rect 41782 597857 41834 597909
rect 43318 597857 43370 597909
rect 672502 597117 672554 597169
rect 675478 597117 675530 597169
rect 674902 596821 674954 596873
rect 675382 596821 675434 596873
rect 41590 596599 41642 596651
rect 43126 596599 43178 596651
rect 43318 596155 43370 596207
rect 45046 596155 45098 596207
rect 41590 590975 41642 591027
rect 43030 590975 43082 591027
rect 41878 590383 41930 590435
rect 42934 590383 42986 590435
rect 41590 587497 41642 587549
rect 56086 587497 56138 587549
rect 37366 584981 37418 585033
rect 43798 584981 43850 585033
rect 40150 584833 40202 584885
rect 41878 584833 41930 584885
rect 42070 584833 42122 584885
rect 42550 584833 42602 584885
rect 34486 584759 34538 584811
rect 43606 584759 43658 584811
rect 40246 584685 40298 584737
rect 42262 584685 42314 584737
rect 42550 584685 42602 584737
rect 58966 584685 59018 584737
rect 43030 584463 43082 584515
rect 43510 584463 43562 584515
rect 43126 584389 43178 584441
rect 43318 584389 43370 584441
rect 42166 584241 42218 584293
rect 43126 584241 43178 584293
rect 41782 584167 41834 584219
rect 41974 584167 42026 584219
rect 42934 584167 42986 584219
rect 41782 583945 41834 583997
rect 42166 582095 42218 582147
rect 43318 582095 43370 582147
rect 42070 581429 42122 581481
rect 42550 581429 42602 581481
rect 42070 580245 42122 580297
rect 43030 580245 43082 580297
rect 43030 580097 43082 580149
rect 43510 580097 43562 580149
rect 42166 579283 42218 579335
rect 48022 579283 48074 579335
rect 42166 578839 42218 578891
rect 43030 578839 43082 578891
rect 42070 578395 42122 578447
rect 42550 578395 42602 578447
rect 42166 577655 42218 577707
rect 43126 577655 43178 577707
rect 43126 577507 43178 577559
rect 43606 577507 43658 577559
rect 42070 577137 42122 577189
rect 42934 577137 42986 577189
rect 42934 576989 42986 577041
rect 43798 576989 43850 577041
rect 672310 576989 672362 577041
rect 676054 576989 676106 577041
rect 655510 576471 655562 576523
rect 676246 576471 676298 576523
rect 655318 576323 655370 576375
rect 676150 576323 676202 576375
rect 655126 576175 655178 576227
rect 676342 576175 676394 576227
rect 673846 576101 673898 576153
rect 676246 576101 676298 576153
rect 670582 575879 670634 575931
rect 676054 575879 676106 575931
rect 672214 575435 672266 575487
rect 676054 575435 676106 575487
rect 670486 574917 670538 574969
rect 676054 574917 676106 574969
rect 42166 574621 42218 574673
rect 43030 574621 43082 574673
rect 672310 574325 672362 574377
rect 676054 574325 676106 574377
rect 42166 574103 42218 574155
rect 43126 574103 43178 574155
rect 42070 573437 42122 573489
rect 42550 573437 42602 573489
rect 669910 573215 669962 573267
rect 670486 573215 670538 573267
rect 42934 573141 42986 573193
rect 58198 573141 58250 573193
rect 670102 573141 670154 573193
rect 670582 573141 670634 573193
rect 47926 573067 47978 573119
rect 58966 573067 59018 573119
rect 48022 572993 48074 573045
rect 59638 572993 59690 573045
rect 42358 572105 42410 572157
rect 42838 572105 42890 572157
rect 42166 570995 42218 571047
rect 43030 570995 43082 571047
rect 42838 570847 42890 570899
rect 43030 570847 43082 570899
rect 670870 570625 670922 570677
rect 676246 570625 676298 570677
rect 42166 570403 42218 570455
rect 43126 570403 43178 570455
rect 50326 570181 50378 570233
rect 59350 570181 59402 570233
rect 47830 570107 47882 570159
rect 59542 570107 59594 570159
rect 672406 569885 672458 569937
rect 676054 569885 676106 569937
rect 42070 569737 42122 569789
rect 43030 569737 43082 569789
rect 670678 569515 670730 569567
rect 676054 569515 676106 569567
rect 42166 569145 42218 569197
rect 42934 569145 42986 569197
rect 672790 569145 672842 569197
rect 676246 569145 676298 569197
rect 673366 568405 673418 568457
rect 676054 568405 676106 568457
rect 672886 567961 672938 568013
rect 676054 567961 676106 568013
rect 672694 567665 672746 567717
rect 676246 567665 676298 567717
rect 655702 567443 655754 567495
rect 675382 567443 675434 567495
rect 649846 564483 649898 564535
rect 679798 564483 679850 564535
rect 674422 559525 674474 559577
rect 675382 559525 675434 559577
rect 656566 558785 656618 558837
rect 674998 558785 675050 558837
rect 674518 558045 674570 558097
rect 675382 558045 675434 558097
rect 672790 556047 672842 556099
rect 675286 556047 675338 556099
rect 654166 555899 654218 555951
rect 675286 555899 675338 555951
rect 674134 555011 674186 555063
rect 675478 555011 675530 555063
rect 673366 554345 673418 554397
rect 675382 554345 675434 554397
rect 672694 553901 672746 553953
rect 675478 553901 675530 553953
rect 674998 553457 675050 553509
rect 675382 553457 675434 553509
rect 673750 553309 673802 553361
rect 675478 553309 675530 553361
rect 672886 551903 672938 551955
rect 675478 551903 675530 551955
rect 674326 548869 674378 548921
rect 675286 548869 675338 548921
rect 674230 548203 674282 548255
rect 675286 548203 675338 548255
rect 43030 541543 43082 541595
rect 57718 541543 57770 541595
rect 42934 541469 42986 541521
rect 57622 541469 57674 541521
rect 42166 538139 42218 538191
rect 43030 538139 43082 538191
rect 42166 536437 42218 536489
rect 42934 536437 42986 536489
rect 673846 533773 673898 533825
rect 675958 533773 676010 533825
rect 655606 533255 655658 533307
rect 676054 533255 676106 533307
rect 655414 533107 655466 533159
rect 676150 533107 676202 533159
rect 655222 532959 655274 533011
rect 676246 532959 676298 533011
rect 672214 532663 672266 532715
rect 672406 532663 672458 532715
rect 676054 532663 676106 532715
rect 672310 531479 672362 531531
rect 676246 531479 676298 531531
rect 42934 529925 42986 529977
rect 58198 529925 58250 529977
rect 670966 528001 671018 528053
rect 676246 528001 676298 528053
rect 670774 527409 670826 527461
rect 676246 527409 676298 527461
rect 673174 526669 673226 526721
rect 676054 526669 676106 526721
rect 42166 526373 42218 526425
rect 42550 526373 42602 526425
rect 672502 526299 672554 526351
rect 676054 526299 676106 526351
rect 673078 525929 673130 525981
rect 676246 525929 676298 525981
rect 42070 525633 42122 525685
rect 42358 525633 42410 525685
rect 42166 525411 42218 525463
rect 42934 525411 42986 525463
rect 673270 525189 673322 525241
rect 676054 525189 676106 525241
rect 672982 524819 673034 524871
rect 676054 524819 676106 524871
rect 672598 524449 672650 524501
rect 676246 524449 676298 524501
rect 50326 524301 50378 524353
rect 58582 524301 58634 524353
rect 47830 524227 47882 524279
rect 59350 524227 59402 524279
rect 649942 521267 649994 521319
rect 679798 521267 679850 521319
rect 676534 498253 676586 498305
rect 679702 498253 679754 498305
rect 655510 490039 655562 490091
rect 676246 490039 676298 490091
rect 655318 489891 655370 489943
rect 676246 489891 676298 489943
rect 655126 489743 655178 489795
rect 676150 489743 676202 489795
rect 676246 489225 676298 489277
rect 676726 489225 676778 489277
rect 670294 488115 670346 488167
rect 676054 488115 676106 488167
rect 676630 488115 676682 488167
rect 670006 487079 670058 487131
rect 676246 487079 676298 487131
rect 674326 486635 674378 486687
rect 676054 486635 676106 486687
rect 674422 486561 674474 486613
rect 676246 486561 676298 486613
rect 674134 485673 674186 485725
rect 676054 485673 676106 485725
rect 674518 483749 674570 483801
rect 676054 483749 676106 483801
rect 674230 483675 674282 483727
rect 675958 483675 676010 483727
rect 672886 481899 672938 481951
rect 676054 481899 676106 481951
rect 672694 481529 672746 481581
rect 676246 481529 676298 481581
rect 672790 480789 672842 480841
rect 676054 480789 676106 480841
rect 673366 480419 673418 480471
rect 676054 480419 676106 480471
rect 673750 480049 673802 480101
rect 676246 480049 676298 480101
rect 650038 478125 650090 478177
rect 679894 478125 679946 478177
rect 41782 476053 41834 476105
rect 50326 476053 50378 476105
rect 41782 475535 41834 475587
rect 47830 475535 47882 475587
rect 37366 475239 37418 475291
rect 42358 475239 42410 475291
rect 677782 475239 677834 475291
rect 679798 475239 679850 475291
rect 41878 474573 41930 474625
rect 43222 474573 43274 474625
rect 41590 472427 41642 472479
rect 43510 472427 43562 472479
rect 45142 472427 45194 472479
rect 41782 472353 41834 472405
rect 58966 472353 59018 472405
rect 41590 469319 41642 469371
rect 42550 469319 42602 469371
rect 34486 463547 34538 463599
rect 41782 463547 41834 463599
rect 47830 463547 47882 463599
rect 676630 440607 676682 440659
rect 677782 440607 677834 440659
rect 23062 437795 23114 437847
rect 39766 437795 39818 437847
rect 39862 437795 39914 437847
rect 62326 437795 62378 437847
rect 676534 434909 676586 434961
rect 677878 434909 677930 434961
rect 41590 426843 41642 426895
rect 53206 426843 53258 426895
rect 41782 426473 41834 426525
rect 50326 426473 50378 426525
rect 41782 425955 41834 426007
rect 48022 425955 48074 426007
rect 41590 424771 41642 424823
rect 43318 424771 43370 424823
rect 41782 423439 41834 423491
rect 43222 423439 43274 423491
rect 23062 422699 23114 422751
rect 41590 422699 41642 422751
rect 41590 420479 41642 420531
rect 62518 420479 62570 420531
rect 39862 417519 39914 417571
rect 41782 417519 41834 417571
rect 40150 417445 40202 417497
rect 42934 417445 42986 417497
rect 41590 415151 41642 415203
rect 43126 415151 43178 415203
rect 41878 414707 41930 414759
rect 43030 414707 43082 414759
rect 41590 414263 41642 414315
rect 47926 414263 47978 414315
rect 41782 413375 41834 413427
rect 41782 413153 41834 413205
rect 42166 409675 42218 409727
rect 42838 409675 42890 409727
rect 42166 409453 42218 409505
rect 42934 409453 42986 409505
rect 42166 408195 42218 408247
rect 43030 408195 43082 408247
rect 42070 407973 42122 408025
rect 42838 407973 42890 408025
rect 42166 406863 42218 406915
rect 43126 406863 43178 406915
rect 42934 406049 42986 406101
rect 58486 406049 58538 406101
rect 42838 402571 42890 402623
rect 59350 402571 59402 402623
rect 655126 400573 655178 400625
rect 676150 400573 676202 400625
rect 655510 400499 655562 400551
rect 676246 400499 676298 400551
rect 655318 400425 655370 400477
rect 676054 400425 676106 400477
rect 673846 400351 673898 400403
rect 676246 400351 676298 400403
rect 53206 400277 53258 400329
rect 59734 400277 59786 400329
rect 50326 400203 50378 400255
rect 59542 400203 59594 400255
rect 48022 400129 48074 400181
rect 59638 400129 59690 400181
rect 670198 398871 670250 398923
rect 676630 398871 676682 398923
rect 674422 398723 674474 398775
rect 676054 398723 676106 398775
rect 670486 398427 670538 398479
rect 676534 398427 676586 398479
rect 674518 397835 674570 397887
rect 676054 397835 676106 397887
rect 673174 395541 673226 395593
rect 676054 395541 676106 395593
rect 42070 394505 42122 394557
rect 57718 394505 57770 394557
rect 650134 388807 650186 388859
rect 679798 388807 679850 388859
rect 41590 385921 41642 385973
rect 53206 385921 53258 385973
rect 673366 385847 673418 385899
rect 674422 385847 674474 385899
rect 673270 385773 673322 385825
rect 674518 385773 674570 385825
rect 41590 385255 41642 385307
rect 50326 385255 50378 385307
rect 41878 384959 41930 385011
rect 48118 384959 48170 385011
rect 41590 384737 41642 384789
rect 43318 384737 43370 384789
rect 41590 383775 41642 383827
rect 43414 383775 43466 383827
rect 41590 382295 41642 382347
rect 43510 382295 43562 382347
rect 41782 381999 41834 382051
rect 43222 381999 43274 382051
rect 45334 381999 45386 382051
rect 656566 381555 656618 381607
rect 675094 381555 675146 381607
rect 39478 374303 39530 374355
rect 41878 374303 41930 374355
rect 41494 374229 41546 374281
rect 43030 374229 43082 374281
rect 41782 373489 41834 373541
rect 48022 373489 48074 373541
rect 673174 372083 673226 372135
rect 675382 372083 675434 372135
rect 41590 371935 41642 371987
rect 42838 371935 42890 371987
rect 41686 371787 41738 371839
rect 42934 371787 42986 371839
rect 41878 370159 41930 370211
rect 41878 369937 41930 369989
rect 42454 366681 42506 366733
rect 42166 366533 42218 366585
rect 42454 366533 42506 366585
rect 42070 366237 42122 366289
rect 42166 364979 42218 365031
rect 42838 364979 42890 365031
rect 42070 364683 42122 364735
rect 42838 364683 42890 364735
rect 42070 364239 42122 364291
rect 43030 364239 43082 364291
rect 42166 363795 42218 363847
rect 42934 363795 42986 363847
rect 42454 361945 42506 361997
rect 59254 361945 59306 361997
rect 42838 359947 42890 359999
rect 59158 359947 59210 359999
rect 655318 357283 655370 357335
rect 676246 357283 676298 357335
rect 655222 357209 655274 357261
rect 676150 357209 676202 357261
rect 655126 357135 655178 357187
rect 676342 357135 676394 357187
rect 53206 357061 53258 357113
rect 58198 357061 58250 357113
rect 48118 356987 48170 357039
rect 59638 356987 59690 357039
rect 50326 356913 50378 356965
rect 58582 356913 58634 356965
rect 673846 356765 673898 356817
rect 676054 356765 676106 356817
rect 673366 355655 673418 355707
rect 676054 355655 676106 355707
rect 673270 354619 673322 354671
rect 676054 354619 676106 354671
rect 672502 354323 672554 354375
rect 673366 354323 673418 354375
rect 672790 354249 672842 354301
rect 673270 354249 673322 354301
rect 674998 351363 675050 351415
rect 676054 351363 676106 351415
rect 42166 351289 42218 351341
rect 57622 351289 57674 351341
rect 675094 350327 675146 350379
rect 676054 350327 676106 350379
rect 674230 348551 674282 348603
rect 676246 348551 676298 348603
rect 675190 348477 675242 348529
rect 676054 348477 676106 348529
rect 650230 345813 650282 345865
rect 679894 345813 679946 345865
rect 674710 345739 674762 345791
rect 675958 345739 676010 345791
rect 674806 345665 674858 345717
rect 676054 345665 676106 345717
rect 674902 345591 674954 345643
rect 676246 345591 676298 345643
rect 41782 342779 41834 342831
rect 53206 342779 53258 342831
rect 41782 342261 41834 342313
rect 50326 342261 50378 342313
rect 41782 341743 41834 341795
rect 48118 341743 48170 341795
rect 41782 341373 41834 341425
rect 43414 341373 43466 341425
rect 675478 341373 675530 341425
rect 675382 340929 675434 340981
rect 41590 340559 41642 340611
rect 43222 340559 43274 340611
rect 41782 340263 41834 340315
rect 43318 340263 43370 340315
rect 666742 339967 666794 340019
rect 675286 339967 675338 340019
rect 675094 339819 675146 339871
rect 675286 339819 675338 339871
rect 41782 339449 41834 339501
rect 43510 339449 43562 339501
rect 41590 339079 41642 339131
rect 43414 339079 43466 339131
rect 674998 337895 675050 337947
rect 675478 337895 675530 337947
rect 675190 337229 675242 337281
rect 675478 337229 675530 337281
rect 674230 336563 674282 336615
rect 675382 336563 675434 336615
rect 674902 336045 674954 336097
rect 675382 336045 675434 336097
rect 674806 332715 674858 332767
rect 675382 332715 675434 332767
rect 674710 331531 674762 331583
rect 675382 331531 675434 331583
rect 41398 331161 41450 331213
rect 42742 331161 42794 331213
rect 41494 331087 41546 331139
rect 43030 331087 43082 331139
rect 41878 330347 41930 330399
rect 45430 330347 45482 330399
rect 41590 328793 41642 328845
rect 42934 328793 42986 328845
rect 654166 328275 654218 328327
rect 666742 328275 666794 328327
rect 41782 327017 41834 327069
rect 41782 326721 41834 326773
rect 42934 325759 42986 325811
rect 43126 325759 43178 325811
rect 42070 323317 42122 323369
rect 42454 323317 42506 323369
rect 42166 323095 42218 323147
rect 43030 323095 43082 323147
rect 41974 321615 42026 321667
rect 43126 321615 43178 321667
rect 42166 321467 42218 321519
rect 43126 321467 43178 321519
rect 42166 321245 42218 321297
rect 43030 321245 43082 321297
rect 42454 319617 42506 319669
rect 58486 319617 58538 319669
rect 43126 316731 43178 316783
rect 59158 316731 59210 316783
rect 53206 313845 53258 313897
rect 58198 313845 58250 313897
rect 48118 313771 48170 313823
rect 59638 313771 59690 313823
rect 50326 313697 50378 313749
rect 59734 313697 59786 313749
rect 654262 311181 654314 311233
rect 676246 311181 676298 311233
rect 654166 311107 654218 311159
rect 676150 311107 676202 311159
rect 654070 311033 654122 311085
rect 676342 311033 676394 311085
rect 42166 308073 42218 308125
rect 59350 308073 59402 308125
rect 674518 305335 674570 305387
rect 676054 305335 676106 305387
rect 675094 305261 675146 305313
rect 676246 305261 676298 305313
rect 674326 302523 674378 302575
rect 675958 302523 676010 302575
rect 674422 302449 674474 302501
rect 676054 302449 676106 302501
rect 674710 302375 674762 302427
rect 676246 302375 676298 302427
rect 43318 300895 43370 300947
rect 62806 300895 62858 300947
rect 650326 299711 650378 299763
rect 679990 299711 680042 299763
rect 39766 299637 39818 299689
rect 43318 299637 43370 299689
rect 674902 299637 674954 299689
rect 676246 299637 676298 299689
rect 41782 299563 41834 299615
rect 60214 299563 60266 299615
rect 674998 299563 675050 299615
rect 676054 299563 676106 299615
rect 41782 299119 41834 299171
rect 51766 299119 51818 299171
rect 41782 298157 41834 298209
rect 43222 298157 43274 298209
rect 43510 298083 43562 298135
rect 62998 298083 63050 298135
rect 41782 297565 41834 297617
rect 43414 297565 43466 297617
rect 41782 297047 41834 297099
rect 43318 297047 43370 297099
rect 39958 296677 40010 296729
rect 43510 296677 43562 296729
rect 41590 295863 41642 295915
rect 43222 295863 43274 295915
rect 674806 295641 674858 295693
rect 675190 295641 675242 295693
rect 674710 295419 674762 295471
rect 675286 295419 675338 295471
rect 674518 294531 674570 294583
rect 675382 294531 675434 294583
rect 53302 293865 53354 293917
rect 59638 293865 59690 293917
rect 56278 293791 56330 293843
rect 60310 293791 60362 293843
rect 39670 293717 39722 293769
rect 58774 293717 58826 293769
rect 674422 292015 674474 292067
rect 675478 292015 675530 292067
rect 674326 291571 674378 291623
rect 675382 291571 675434 291623
rect 48214 290905 48266 290957
rect 58390 290905 58442 290957
rect 656566 290831 656618 290883
rect 674806 290831 674858 290883
rect 51766 289499 51818 289551
rect 58006 289499 58058 289551
rect 50326 288019 50378 288071
rect 59638 288019 59690 288071
rect 674998 287723 675050 287775
rect 675382 287723 675434 287775
rect 41878 287131 41930 287183
rect 45814 287131 45866 287183
rect 674902 286761 674954 286813
rect 675382 286761 675434 286813
rect 41494 285281 41546 285333
rect 43126 285281 43178 285333
rect 41686 285207 41738 285259
rect 43030 285207 43082 285259
rect 41590 285133 41642 285185
rect 42934 285133 42986 285185
rect 53206 285133 53258 285185
rect 58966 285133 59018 285185
rect 653782 284245 653834 284297
rect 658006 284245 658058 284297
rect 41782 283801 41834 283853
rect 41782 283505 41834 283557
rect 48118 282543 48170 282595
rect 59638 282543 59690 282595
rect 45526 282321 45578 282373
rect 58966 282321 59018 282373
rect 56182 282247 56234 282299
rect 57622 282247 57674 282299
rect 42070 280101 42122 280153
rect 42838 280101 42890 280153
rect 42166 279879 42218 279931
rect 43126 279879 43178 279931
rect 45718 279435 45770 279487
rect 59542 279435 59594 279487
rect 654166 279435 654218 279487
rect 663766 279435 663818 279487
rect 45622 279361 45674 279413
rect 59350 279361 59402 279413
rect 42166 278547 42218 278599
rect 42934 278547 42986 278599
rect 42070 278473 42122 278525
rect 43126 278473 43178 278525
rect 314902 278251 314954 278303
rect 408310 278251 408362 278303
rect 319510 278177 319562 278229
rect 418966 278177 419018 278229
rect 316630 278103 316682 278155
rect 411862 278103 411914 278155
rect 317878 278029 317930 278081
rect 415414 278029 415466 278081
rect 322102 277955 322154 278007
rect 426262 277955 426314 278007
rect 382294 277881 382346 277933
rect 574966 277881 575018 277933
rect 326422 277807 326474 277859
rect 437014 277807 437066 277859
rect 323830 277733 323882 277785
rect 429910 277733 429962 277785
rect 329302 277659 329354 277711
rect 444118 277659 444170 277711
rect 332374 277585 332426 277637
rect 451222 277585 451274 277637
rect 334966 277511 335018 277563
rect 458230 277511 458282 277563
rect 337846 277437 337898 277489
rect 465334 277437 465386 277489
rect 42070 277363 42122 277415
rect 43030 277363 43082 277415
rect 341014 277363 341066 277415
rect 472438 277363 472490 277415
rect 343894 277289 343946 277341
rect 479542 277289 479594 277341
rect 373846 277215 373898 277267
rect 554038 277215 554090 277267
rect 375094 277141 375146 277193
rect 557590 277141 557642 277193
rect 376822 277067 376874 277119
rect 561142 277067 561194 277119
rect 377974 276993 378026 277045
rect 564694 276993 564746 277045
rect 379414 276919 379466 276971
rect 568246 276919 568298 276971
rect 381046 276845 381098 276897
rect 571702 276845 571754 276897
rect 383638 276771 383690 276823
rect 578806 276771 578858 276823
rect 320950 276697 321002 276749
rect 422806 276697 422858 276749
rect 386518 276623 386570 276675
rect 585910 276623 585962 276675
rect 676534 276623 676586 276675
rect 679798 276623 679850 276675
rect 385366 276549 385418 276601
rect 582358 276549 582410 276601
rect 392278 276475 392330 276527
rect 600118 276475 600170 276527
rect 42838 276401 42890 276453
rect 53302 276401 53354 276453
rect 286102 276401 286154 276453
rect 336502 276401 336554 276453
rect 359158 276401 359210 276453
rect 517366 276401 517418 276453
rect 287350 276327 287402 276379
rect 340054 276327 340106 276379
rect 361750 276327 361802 276379
rect 524470 276327 524522 276379
rect 288694 276253 288746 276305
rect 343606 276253 343658 276305
rect 364630 276253 364682 276305
rect 531574 276253 531626 276305
rect 290326 276179 290378 276231
rect 347158 276179 347210 276231
rect 367702 276179 367754 276231
rect 538678 276179 538730 276231
rect 291862 276105 291914 276157
rect 350710 276105 350762 276157
rect 370294 276105 370346 276157
rect 545782 276105 545834 276157
rect 293014 276031 293066 276083
rect 354262 276031 354314 276083
rect 371926 276031 371978 276083
rect 549334 276031 549386 276083
rect 294646 275957 294698 276009
rect 357814 275957 357866 276009
rect 371062 275957 371114 276009
rect 546934 275957 546986 276009
rect 295894 275883 295946 275935
rect 361366 275883 361418 275935
rect 373462 275883 373514 275935
rect 552790 275883 552842 275935
rect 296470 275809 296522 275861
rect 362518 275809 362570 275861
rect 374614 275809 374666 275861
rect 556342 275809 556394 275861
rect 297334 275735 297386 275787
rect 364918 275735 364970 275787
rect 377494 275735 377546 275787
rect 563446 275735 563498 275787
rect 297814 275661 297866 275713
rect 366070 275661 366122 275713
rect 376246 275661 376298 275713
rect 559894 275661 559946 275713
rect 298966 275587 299018 275639
rect 368470 275587 368522 275639
rect 380566 275587 380618 275639
rect 570550 275587 570602 275639
rect 300214 275513 300266 275565
rect 372022 275513 372074 275565
rect 381814 275513 381866 275565
rect 574102 275513 574154 275565
rect 299446 275439 299498 275491
rect 369622 275439 369674 275491
rect 388918 275439 388970 275491
rect 591862 275439 591914 275491
rect 303286 275365 303338 275417
rect 379126 275365 379178 275417
rect 389590 275365 389642 275417
rect 593014 275365 593066 275417
rect 304438 275291 304490 275343
rect 382582 275291 382634 275343
rect 391990 275291 392042 275343
rect 598966 275291 599018 275343
rect 307318 275217 307370 275269
rect 389686 275217 389738 275269
rect 396310 275217 396362 275269
rect 609526 275217 609578 275269
rect 310390 275143 310442 275195
rect 396790 275143 396842 275195
rect 404950 275143 405002 275195
rect 314710 275069 314762 275121
rect 407446 275069 407498 275121
rect 311638 274995 311690 275047
rect 400342 274995 400394 275047
rect 407734 275143 407786 275195
rect 623734 275143 623786 275195
rect 408598 275069 408650 275121
rect 635542 275069 635594 275121
rect 630838 274995 630890 275047
rect 284758 274921 284810 274973
rect 332950 274921 333002 274973
rect 356182 274921 356234 274973
rect 510262 274921 510314 274973
rect 283030 274847 283082 274899
rect 329398 274847 329450 274899
rect 344566 274847 344618 274899
rect 481942 274847 481994 274899
rect 281782 274773 281834 274825
rect 325846 274773 325898 274825
rect 339094 274773 339146 274825
rect 467734 274773 467786 274825
rect 336022 274699 336074 274751
rect 460630 274699 460682 274751
rect 333142 274625 333194 274677
rect 453526 274625 453578 274677
rect 330454 274551 330506 274603
rect 446422 274551 446474 274603
rect 328822 274477 328874 274529
rect 442870 274477 442922 274529
rect 325942 274403 325994 274455
rect 435862 274403 435914 274455
rect 323350 274329 323402 274381
rect 428758 274329 428810 274381
rect 320182 274255 320234 274307
rect 421654 274255 421706 274307
rect 315958 274181 316010 274233
rect 410998 274181 411050 274233
rect 317302 274107 317354 274159
rect 414550 274107 414602 274159
rect 348502 274033 348554 274085
rect 401494 274033 401546 274085
rect 401782 274033 401834 274085
rect 407734 274033 407786 274085
rect 334294 273959 334346 274011
rect 380278 273959 380330 274011
rect 347062 273885 347114 273937
rect 394486 273885 394538 273937
rect 326134 273811 326186 273863
rect 373174 273811 373226 273863
rect 341974 273737 342026 273789
rect 387382 273737 387434 273789
rect 331222 273663 331274 273715
rect 376726 273663 376778 273715
rect 43126 273515 43178 273567
rect 56278 273515 56330 273567
rect 160438 273515 160490 273567
rect 209398 273515 209450 273567
rect 230134 273515 230186 273567
rect 242902 273515 242954 273567
rect 275158 273515 275210 273567
rect 309334 273515 309386 273567
rect 350038 273515 350090 273567
rect 494902 273515 494954 273567
rect 522550 273515 522602 273567
rect 631990 273515 632042 273567
rect 130870 273441 130922 273493
rect 190102 273441 190154 273493
rect 193558 273441 193610 273493
rect 219094 273441 219146 273493
rect 227830 273441 227882 273493
rect 242134 273441 242186 273493
rect 277750 273441 277802 273493
rect 316438 273441 316490 273493
rect 349462 273441 349514 273493
rect 493750 273441 493802 273493
rect 529846 273441 529898 273493
rect 624982 273441 625034 273493
rect 108406 273367 108458 273419
rect 109366 273367 109418 273419
rect 122614 273367 122666 273419
rect 123766 273367 123818 273419
rect 142678 273367 142730 273419
rect 209686 273367 209738 273419
rect 275350 273367 275402 273419
rect 310486 273367 310538 273419
rect 310582 273367 310634 273419
rect 344758 273367 344810 273419
rect 352438 273367 352490 273419
rect 500854 273367 500906 273419
rect 135574 273293 135626 273345
rect 209878 273293 209930 273345
rect 219574 273293 219626 273345
rect 238678 273293 238730 273345
rect 278230 273293 278282 273345
rect 317590 273293 317642 273345
rect 352630 273293 352682 273345
rect 502006 273293 502058 273345
rect 68278 273219 68330 273271
rect 142486 273219 142538 273271
rect 153334 273219 153386 273271
rect 209590 273219 209642 273271
rect 279670 273219 279722 273271
rect 321142 273219 321194 273271
rect 355510 273219 355562 273271
rect 509110 273219 509162 273271
rect 132022 273145 132074 273197
rect 209782 273145 209834 273197
rect 285622 273145 285674 273197
rect 335350 273145 335402 273197
rect 355030 273145 355082 273197
rect 507958 273145 508010 273197
rect 508246 273145 508298 273197
rect 639094 273145 639146 273197
rect 127318 273071 127370 273123
rect 209974 273071 210026 273123
rect 217174 273071 217226 273123
rect 237622 273071 237674 273123
rect 284950 273071 285002 273123
rect 334198 273071 334250 273123
rect 358582 273071 358634 273123
rect 128470 272997 128522 273049
rect 210166 272997 210218 273049
rect 218326 272997 218378 273049
rect 238102 272997 238154 273049
rect 286774 272997 286826 273049
rect 338902 272997 338954 273049
rect 360982 272997 361034 273049
rect 375190 273071 375242 273123
rect 514966 273071 515018 273123
rect 125014 272923 125066 272975
rect 207286 272923 207338 272975
rect 216022 272923 216074 272975
rect 236950 272923 237002 272975
rect 274198 272923 274250 272975
rect 306934 272923 306986 272975
rect 307030 272923 307082 272975
rect 358966 272923 359018 272975
rect 361270 272923 361322 272975
rect 516214 272997 516266 273049
rect 516310 272997 516362 273049
rect 580054 272997 580106 273049
rect 123670 272849 123722 272901
rect 209014 272849 209066 272901
rect 220726 272849 220778 272901
rect 239158 272849 239210 272901
rect 289942 272849 289994 272901
rect 346006 272849 346058 272901
rect 363574 272849 363626 272901
rect 522070 272923 522122 272975
rect 120214 272775 120266 272827
rect 207862 272775 207914 272827
rect 211222 272775 211274 272827
rect 235030 272775 235082 272827
rect 292246 272775 292298 272827
rect 351862 272775 351914 272827
rect 364150 272775 364202 272827
rect 523318 272849 523370 272901
rect 523798 272849 523850 272901
rect 611926 272849 611978 272901
rect 116662 272701 116714 272753
rect 207094 272701 207146 272753
rect 233686 272701 233738 272753
rect 244054 272701 244106 272753
rect 292726 272701 292778 272753
rect 353110 272701 353162 272753
rect 366550 272701 366602 272753
rect 529174 272775 529226 272827
rect 113110 272627 113162 272679
rect 206038 272627 206090 272679
rect 213622 272627 213674 272679
rect 236278 272627 236330 272679
rect 295414 272627 295466 272679
rect 360214 272627 360266 272679
rect 367126 272627 367178 272679
rect 530422 272701 530474 272753
rect 96598 272553 96650 272605
rect 106678 272553 106730 272605
rect 110806 272553 110858 272605
rect 205462 272553 205514 272605
rect 214774 272553 214826 272605
rect 236470 272553 236522 272605
rect 270262 272553 270314 272605
rect 297526 272553 297578 272605
rect 298486 272553 298538 272605
rect 367222 272553 367274 272605
rect 372694 272553 372746 272605
rect 536278 272627 536330 272679
rect 103702 272479 103754 272531
rect 203542 272479 203594 272531
rect 210070 272479 210122 272531
rect 234550 272479 234602 272531
rect 236086 272479 236138 272531
rect 245302 272479 245354 272531
rect 272278 272479 272330 272531
rect 302230 272479 302282 272531
rect 106102 272405 106154 272457
rect 204022 272405 204074 272457
rect 205366 272405 205418 272457
rect 232630 272405 232682 272457
rect 270550 272405 270602 272457
rect 298678 272405 298730 272457
rect 301366 272405 301418 272457
rect 374326 272479 374378 272531
rect 537430 272553 537482 272605
rect 551638 272479 551690 272531
rect 303958 272405 304010 272457
rect 381430 272405 381482 272457
rect 381526 272405 381578 272457
rect 572950 272405 573002 272457
rect 98998 272331 99050 272383
rect 199126 272331 199178 272383
rect 207670 272331 207722 272383
rect 233878 272331 233930 272383
rect 272758 272331 272810 272383
rect 303478 272331 303530 272383
rect 307126 272331 307178 272383
rect 388534 272331 388586 272383
rect 407446 272331 407498 272383
rect 587158 272331 587210 272383
rect 76534 272257 76586 272309
rect 84790 272183 84842 272235
rect 86326 272183 86378 272235
rect 104854 272183 104906 272235
rect 106486 272183 106538 272235
rect 106678 272257 106730 272309
rect 201622 272257 201674 272309
rect 208918 272257 208970 272309
rect 234358 272257 234410 272309
rect 234934 272257 234986 272309
rect 244822 272257 244874 272309
rect 273430 272257 273482 272309
rect 305782 272257 305834 272309
rect 309910 272257 309962 272309
rect 395638 272257 395690 272309
rect 395926 272257 395978 272309
rect 608374 272257 608426 272309
rect 195670 272183 195722 272235
rect 198262 272183 198314 272235
rect 222070 272183 222122 272235
rect 276310 272183 276362 272235
rect 312886 272183 312938 272235
rect 312982 272183 313034 272235
rect 402742 272183 402794 272235
rect 402838 272183 402890 272235
rect 622582 272183 622634 272235
rect 194710 272109 194762 272161
rect 222262 272109 222314 272161
rect 228982 272109 229034 272161
rect 242422 272109 242474 272161
rect 277078 272109 277130 272161
rect 314038 272109 314090 272161
rect 315478 272109 315530 272161
rect 409846 272109 409898 272161
rect 413686 272109 413738 272161
rect 643894 272109 643946 272161
rect 119062 272035 119114 272087
rect 120886 272035 120938 272087
rect 165142 272035 165194 272087
rect 166966 272035 167018 272087
rect 167542 272035 167594 272087
rect 213046 272035 213098 272087
rect 298102 272035 298154 272087
rect 327094 272035 327146 272087
rect 346966 272035 347018 272087
rect 487798 272035 487850 272087
rect 174646 271961 174698 272013
rect 212854 271961 212906 272013
rect 232534 271961 232586 272013
rect 243670 271961 243722 272013
rect 271030 271961 271082 272013
rect 299926 271961 299978 272013
rect 159286 271887 159338 271939
rect 195286 271887 195338 271939
rect 195862 271887 195914 271939
rect 218998 271887 219050 271939
rect 231382 271887 231434 271939
rect 243094 271887 243146 271939
rect 191158 271813 191210 271865
rect 227158 271813 227210 271865
rect 298006 271813 298058 271865
rect 328246 271961 328298 272013
rect 346486 271961 346538 272013
rect 486646 271961 486698 272013
rect 300118 271813 300170 271865
rect 324694 271887 324746 271939
rect 342742 271887 342794 271939
rect 348310 271887 348362 271939
rect 344086 271813 344138 271865
rect 480694 271887 480746 271939
rect 147382 271739 147434 271791
rect 149686 271739 149738 271791
rect 192310 271739 192362 271791
rect 222166 271739 222218 271791
rect 341494 271739 341546 271791
rect 473686 271813 473738 271865
rect 348598 271739 348650 271791
rect 466582 271739 466634 271791
rect 166294 271665 166346 271717
rect 196342 271665 196394 271717
rect 199414 271665 199466 271717
rect 218902 271665 218954 271717
rect 335446 271665 335498 271717
rect 459478 271665 459530 271717
rect 75286 271591 75338 271643
rect 77686 271591 77738 271643
rect 129718 271591 129770 271643
rect 132406 271591 132458 271643
rect 181750 271591 181802 271643
rect 212950 271591 213002 271643
rect 332566 271591 332618 271643
rect 452374 271591 452426 271643
rect 89494 271517 89546 271569
rect 92086 271517 92138 271569
rect 150934 271517 150986 271569
rect 152374 271517 152426 271569
rect 185206 271517 185258 271569
rect 212566 271517 212618 271569
rect 329974 271517 330026 271569
rect 445270 271517 445322 271569
rect 173398 271443 173450 271495
rect 201526 271443 201578 271495
rect 201814 271443 201866 271495
rect 221974 271443 222026 271495
rect 326902 271443 326954 271495
rect 438166 271443 438218 271495
rect 180502 271369 180554 271421
rect 205942 271369 205994 271421
rect 212470 271369 212522 271421
rect 235702 271369 235754 271421
rect 324022 271369 324074 271421
rect 431062 271369 431114 271421
rect 188758 271295 188810 271347
rect 212758 271295 212810 271347
rect 321430 271295 321482 271347
rect 423958 271295 424010 271347
rect 161590 271221 161642 271273
rect 163894 271221 163946 271273
rect 184054 271221 184106 271273
rect 205750 271221 205802 271273
rect 237238 271221 237290 271273
rect 245590 271221 245642 271273
rect 318358 271221 318410 271273
rect 416950 271221 417002 271273
rect 175798 271147 175850 271199
rect 178294 271147 178346 271199
rect 187606 271147 187658 271199
rect 205846 271147 205898 271199
rect 238486 271147 238538 271199
rect 246070 271147 246122 271199
rect 338614 271147 338666 271199
rect 348598 271147 348650 271199
rect 357910 271147 357962 271199
rect 375190 271147 375242 271199
rect 387286 271147 387338 271199
rect 407446 271147 407498 271199
rect 85942 271073 85994 271125
rect 198550 271073 198602 271125
rect 240790 271073 240842 271125
rect 247222 271073 247274 271125
rect 221878 270999 221930 271051
rect 239350 270999 239402 271051
rect 239542 270999 239594 271051
rect 241270 270999 241322 271051
rect 241942 270999 241994 271051
rect 247702 270999 247754 271051
rect 223030 270925 223082 270977
rect 240022 270925 240074 270977
rect 243190 270925 243242 270977
rect 247990 270925 248042 270977
rect 224278 270851 224330 270903
rect 240502 270851 240554 270903
rect 244342 270851 244394 270903
rect 248662 270851 248714 270903
rect 351382 270851 351434 270903
rect 355414 270851 355466 270903
rect 225430 270777 225482 270829
rect 241078 270777 241130 270829
rect 245494 270777 245546 270829
rect 249142 270777 249194 270829
rect 94198 270703 94250 270755
rect 94966 270703 95018 270755
rect 101302 270703 101354 270755
rect 103606 270703 103658 270755
rect 115510 270703 115562 270755
rect 118006 270703 118058 270755
rect 133270 270703 133322 270755
rect 135286 270703 135338 270755
rect 136822 270703 136874 270755
rect 138166 270703 138218 270755
rect 154486 270703 154538 270755
rect 155446 270703 155498 270755
rect 168694 270703 168746 270755
rect 169846 270703 169898 270755
rect 179350 270703 179402 270755
rect 181366 270703 181418 270755
rect 182902 270703 182954 270755
rect 184246 270703 184298 270755
rect 185494 270703 185546 270755
rect 186454 270703 186506 270755
rect 226582 270703 226634 270755
rect 239542 270703 239594 270755
rect 239638 270703 239690 270755
rect 246454 270703 246506 270755
rect 246742 270703 246794 270755
rect 249622 270703 249674 270755
rect 334102 270703 334154 270755
rect 337750 270703 337802 270755
rect 338134 270703 338186 270755
rect 341302 270703 341354 270755
rect 408982 270703 409034 270755
rect 413398 270703 413450 270755
rect 146230 270629 146282 270681
rect 214966 270629 215018 270681
rect 269206 270629 269258 270681
rect 295126 270629 295178 270681
rect 295222 270629 295274 270681
rect 301078 270629 301130 270681
rect 302422 270629 302474 270681
rect 304630 270629 304682 270681
rect 306358 270629 306410 270681
rect 341974 270629 342026 270681
rect 345430 270629 345482 270681
rect 484246 270629 484298 270681
rect 141526 270555 141578 270607
rect 213814 270555 213866 270607
rect 279286 270555 279338 270607
rect 298198 270555 298250 270607
rect 298390 270555 298442 270607
rect 318838 270555 318890 270607
rect 348118 270555 348170 270607
rect 490198 270555 490250 270607
rect 137974 270481 138026 270533
rect 212662 270481 212714 270533
rect 280150 270481 280202 270533
rect 322390 270481 322442 270533
rect 348406 270481 348458 270533
rect 491350 270481 491402 270533
rect 134422 270407 134474 270459
rect 211894 270407 211946 270459
rect 253942 270407 253994 270459
rect 257302 270407 257354 270459
rect 262966 270407 263018 270459
rect 279766 270407 279818 270459
rect 280630 270407 280682 270459
rect 323542 270407 323594 270459
rect 350710 270407 350762 270459
rect 497302 270407 497354 270459
rect 121462 270333 121514 270385
rect 208342 270333 208394 270385
rect 209590 270333 209642 270385
rect 216886 270333 216938 270385
rect 262486 270333 262538 270385
rect 278614 270333 278666 270385
rect 284182 270333 284234 270385
rect 117910 270259 117962 270311
rect 207574 270259 207626 270311
rect 212566 270259 212618 270311
rect 225526 270259 225578 270311
rect 255286 270259 255338 270311
rect 260854 270259 260906 270311
rect 286294 270259 286346 270311
rect 114358 270185 114410 270237
rect 206422 270185 206474 270237
rect 209782 270185 209834 270237
rect 211414 270185 211466 270237
rect 212758 270185 212810 270237
rect 226678 270185 226730 270237
rect 261238 270185 261290 270237
rect 275062 270185 275114 270237
rect 284470 270185 284522 270237
rect 293974 270185 294026 270237
rect 109558 270111 109610 270163
rect 205270 270111 205322 270163
rect 209878 270111 209930 270163
rect 212374 270111 212426 270163
rect 212854 270111 212906 270163
rect 222838 270111 222890 270163
rect 265366 270111 265418 270163
rect 285718 270111 285770 270163
rect 287926 270111 287978 270163
rect 298198 270333 298250 270385
rect 319990 270333 320042 270385
rect 351286 270333 351338 270385
rect 498454 270333 498506 270385
rect 298294 270259 298346 270311
rect 330646 270259 330698 270311
rect 354070 270259 354122 270311
rect 505558 270259 505610 270311
rect 331798 270185 331850 270237
rect 353686 270185 353738 270237
rect 504406 270185 504458 270237
rect 102550 270037 102602 270089
rect 203350 270037 203402 270089
rect 212950 270037 213002 270089
rect 224758 270037 224810 270089
rect 264694 270037 264746 270089
rect 107254 269963 107306 270015
rect 204694 269963 204746 270015
rect 213046 269963 213098 270015
rect 221014 269963 221066 270015
rect 261814 269963 261866 270015
rect 276214 269963 276266 270015
rect 283318 269963 283370 270015
rect 100150 269889 100202 269941
rect 202870 269889 202922 269941
rect 205942 269889 205994 269941
rect 224086 269889 224138 269941
rect 256246 269889 256298 269941
rect 263254 269889 263306 269941
rect 264886 269889 264938 269941
rect 284566 269889 284618 269941
rect 95446 269815 95498 269867
rect 195190 269815 195242 269867
rect 205846 269815 205898 269867
rect 226006 269815 226058 269867
rect 260566 269815 260618 269867
rect 273910 269815 273962 269867
rect 93046 269741 93098 269793
rect 200950 269741 201002 269793
rect 205750 269741 205802 269793
rect 225238 269741 225290 269793
rect 259894 269741 259946 269793
rect 271510 269741 271562 269793
rect 90646 269667 90698 269719
rect 199702 269667 199754 269719
rect 201526 269667 201578 269719
rect 222358 269667 222410 269719
rect 258166 269667 258218 269719
rect 267958 269667 268010 269719
rect 268630 269667 268682 269719
rect 284470 269741 284522 269793
rect 271702 269667 271754 269719
rect 288022 270037 288074 270089
rect 286486 269963 286538 270015
rect 295222 269963 295274 270015
rect 334102 270111 334154 270163
rect 356758 270111 356810 270163
rect 511510 270111 511562 270163
rect 298198 270037 298250 270089
rect 342454 270037 342506 270089
rect 356950 270037 357002 270089
rect 512662 270037 512714 270089
rect 338134 269963 338186 270015
rect 359350 269963 359402 270015
rect 518518 269963 518570 270015
rect 290614 269889 290666 269941
rect 342742 269889 342794 269941
rect 359830 269889 359882 269941
rect 519766 269889 519818 269941
rect 291094 269815 291146 269867
rect 349558 269815 349610 269867
rect 362230 269815 362282 269867
rect 525622 269815 525674 269867
rect 293974 269741 294026 269793
rect 356662 269741 356714 269793
rect 362806 269741 362858 269793
rect 526870 269741 526922 269793
rect 293494 269667 293546 269719
rect 351382 269667 351434 269719
rect 365302 269667 365354 269719
rect 532726 269667 532778 269719
rect 83638 269593 83690 269645
rect 87190 269519 87242 269571
rect 185686 269519 185738 269571
rect 196342 269593 196394 269645
rect 220534 269593 220586 269645
rect 249046 269593 249098 269645
rect 250294 269593 250346 269645
rect 255766 269593 255818 269645
rect 262102 269593 262154 269645
rect 267766 269593 267818 269645
rect 291574 269593 291626 269645
rect 297046 269593 297098 269645
rect 363670 269593 363722 269645
rect 198070 269519 198122 269571
rect 206518 269519 206570 269571
rect 233398 269519 233450 269571
rect 258646 269519 258698 269571
rect 269110 269519 269162 269571
rect 271510 269519 271562 269571
rect 286486 269519 286538 269571
rect 288502 269519 288554 269571
rect 298198 269519 298250 269571
rect 299638 269519 299690 269571
rect 370774 269519 370826 269571
rect 371254 269519 371306 269571
rect 548086 269519 548138 269571
rect 81238 269445 81290 269497
rect 196822 269445 196874 269497
rect 204118 269445 204170 269497
rect 232150 269445 232202 269497
rect 260086 269445 260138 269497
rect 272662 269445 272714 269497
rect 272950 269445 273002 269497
rect 302422 269445 302474 269497
rect 302614 269445 302666 269497
rect 377878 269445 377930 269497
rect 379894 269445 379946 269497
rect 569398 269445 569450 269497
rect 82390 269371 82442 269423
rect 197398 269371 197450 269423
rect 202966 269371 203018 269423
rect 231958 269371 232010 269423
rect 266518 269371 266570 269423
rect 271702 269371 271754 269423
rect 274678 269371 274730 269423
rect 308182 269371 308234 269423
rect 308278 269371 308330 269423
rect 392086 269371 392138 269423
rect 394390 269371 394442 269423
rect 604822 269371 604874 269423
rect 74134 269297 74186 269349
rect 185590 269297 185642 269349
rect 185686 269297 185738 269349
rect 199030 269297 199082 269349
rect 200662 269297 200714 269349
rect 230998 269297 231050 269349
rect 257686 269297 257738 269349
rect 266806 269297 266858 269349
rect 67030 269223 67082 269275
rect 192598 269223 192650 269275
rect 197110 269223 197162 269275
rect 229558 269223 229610 269275
rect 145078 269149 145130 269201
rect 214486 269149 214538 269201
rect 262006 269149 262058 269201
rect 275830 269297 275882 269349
rect 277462 269223 277514 269275
rect 283702 269223 283754 269275
rect 298294 269223 298346 269275
rect 311158 269297 311210 269349
rect 399190 269297 399242 269349
rect 399958 269297 400010 269349
rect 619030 269297 619082 269349
rect 311734 269223 311786 269275
rect 314230 269223 314282 269275
rect 406294 269223 406346 269275
rect 406582 269223 406634 269275
rect 408598 269223 408650 269275
rect 269686 269149 269738 269201
rect 296374 269149 296426 269201
rect 303766 269149 303818 269201
rect 334294 269149 334346 269201
rect 345238 269149 345290 269201
rect 483094 269149 483146 269201
rect 148630 269075 148682 269127
rect 215734 269075 215786 269127
rect 253366 269075 253418 269127
rect 256150 269075 256202 269127
rect 266038 269075 266090 269127
rect 286870 269075 286922 269127
rect 302038 269075 302090 269127
rect 331222 269075 331274 269127
rect 342646 269075 342698 269127
rect 477142 269075 477194 269127
rect 149782 269001 149834 269053
rect 216214 269001 216266 269053
rect 281302 269001 281354 269053
rect 300118 269001 300170 269053
rect 384118 269001 384170 269053
rect 516310 269001 516362 269053
rect 152182 268927 152234 268979
rect 216694 268927 216746 268979
rect 259414 268927 259466 268979
rect 270358 268927 270410 268979
rect 155734 268853 155786 268905
rect 217366 268853 217418 268905
rect 263638 268853 263690 268905
rect 281014 268927 281066 268979
rect 282070 268927 282122 268979
rect 298102 268927 298154 268979
rect 300694 268927 300746 268979
rect 326134 268927 326186 268979
rect 339766 268927 339818 268979
rect 470134 268927 470186 268979
rect 156886 268779 156938 268831
rect 218134 268779 218186 268831
rect 257494 268779 257546 268831
rect 265654 268779 265706 268831
rect 278902 268779 278954 268831
rect 298390 268853 298442 268905
rect 336886 268853 336938 268905
rect 463030 268853 463082 268905
rect 289174 268779 289226 268831
rect 310582 268779 310634 268831
rect 334294 268779 334346 268831
rect 455926 268779 455978 268831
rect 162838 268705 162890 268757
rect 219286 268705 219338 268757
rect 268438 268705 268490 268757
rect 292822 268705 292874 268757
rect 295222 268705 295274 268757
rect 307030 268705 307082 268757
rect 331222 268705 331274 268757
rect 448822 268705 448874 268757
rect 163990 268631 164042 268683
rect 219958 268631 220010 268683
rect 254614 268631 254666 268683
rect 258550 268631 258602 268683
rect 277558 268631 277610 268683
rect 315286 268631 315338 268683
rect 328342 268631 328394 268683
rect 441718 268631 441770 268683
rect 42166 268557 42218 268609
rect 48214 268557 48266 268609
rect 171094 268557 171146 268609
rect 221782 268557 221834 268609
rect 266806 268557 266858 268609
rect 289270 268557 289322 268609
rect 325750 268557 325802 268609
rect 434614 268557 434666 268609
rect 169750 268483 169802 268535
rect 221206 268483 221258 268535
rect 253174 268483 253226 268535
rect 254998 268483 255050 268535
rect 257014 268483 257066 268535
rect 264406 268483 264458 268535
rect 267286 268483 267338 268535
rect 290422 268483 290474 268535
rect 322582 268483 322634 268535
rect 427510 268483 427562 268535
rect 185590 268409 185642 268461
rect 194998 268409 195050 268461
rect 176950 268261 177002 268313
rect 223414 268409 223466 268461
rect 319702 268409 319754 268461
rect 420502 268409 420554 268461
rect 195190 268335 195242 268387
rect 201142 268335 201194 268387
rect 219094 268335 219146 268387
rect 178198 268113 178250 268165
rect 223606 268261 223658 268313
rect 247894 268335 247946 268387
rect 249814 268335 249866 268387
rect 255094 268335 255146 268387
rect 259702 268335 259754 268387
rect 317110 268335 317162 268387
rect 408982 268335 409034 268387
rect 227830 268261 227882 268313
rect 312310 268261 312362 268313
rect 348502 268261 348554 268313
rect 195286 268187 195338 268239
rect 218614 268187 218666 268239
rect 222070 268187 222122 268239
rect 230038 268187 230090 268239
rect 309238 268187 309290 268239
rect 347062 268187 347114 268239
rect 408502 268187 408554 268239
rect 640342 268187 640394 268239
rect 190102 268039 190154 268091
rect 210742 268113 210794 268165
rect 221974 268113 222026 268165
rect 231478 268113 231530 268165
rect 305686 268113 305738 268165
rect 384982 268113 385034 268165
rect 218902 268039 218954 268091
rect 230518 268039 230570 268091
rect 252694 268039 252746 268091
rect 253750 268039 253802 268091
rect 264118 268039 264170 268091
rect 282166 268039 282218 268091
rect 342166 268039 342218 268091
rect 359446 268039 359498 268091
rect 365686 268039 365738 268091
rect 533878 268039 533930 268091
rect 218998 267965 219050 268017
rect 229078 267965 229130 268017
rect 336694 267965 336746 268017
rect 354262 267965 354314 268017
rect 209398 267891 209450 267943
rect 218902 267891 218954 267943
rect 222262 267891 222314 267943
rect 228406 267891 228458 267943
rect 333622 267891 333674 267943
rect 351382 267891 351434 267943
rect 199126 267817 199178 267869
rect 202294 267817 202346 267869
rect 207286 267817 207338 267869
rect 209494 267817 209546 267869
rect 222166 267817 222218 267869
rect 227638 267817 227690 267869
rect 282550 267817 282602 267869
rect 298006 267817 298058 267869
rect 339286 267817 339338 267869
rect 360406 267817 360458 267869
rect 401302 267817 401354 267869
rect 402838 267817 402890 267869
rect 409942 267817 409994 267869
rect 413686 267817 413738 267869
rect 351958 267743 352010 267795
rect 499606 267743 499658 267795
rect 354838 267669 354890 267721
rect 506710 267669 506762 267721
rect 357430 267595 357482 267647
rect 513814 267595 513866 267647
rect 360310 267521 360362 267573
rect 520918 267521 520970 267573
rect 363382 267447 363434 267499
rect 528022 267447 528074 267499
rect 365974 267373 366026 267425
rect 535126 267373 535178 267425
rect 368950 267299 369002 267351
rect 542230 267299 542282 267351
rect 372502 267225 372554 267277
rect 550486 267225 550538 267277
rect 384886 267151 384938 267203
rect 581206 267151 581258 267203
rect 386038 267077 386090 267129
rect 584758 267077 584810 267129
rect 387766 267003 387818 267055
rect 588310 267003 588362 267055
rect 301846 266929 301898 266981
rect 375286 266929 375338 266981
rect 394678 266929 394730 266981
rect 606070 266929 606122 266981
rect 305014 266855 305066 266907
rect 383830 266855 383882 266907
rect 393238 266855 393290 266907
rect 602518 266855 602570 266907
rect 306166 266781 306218 266833
rect 386134 266781 386186 266833
rect 397558 266781 397610 266833
rect 613078 266781 613130 266833
rect 308758 266707 308810 266759
rect 392950 266707 393002 266759
rect 398230 266707 398282 266759
rect 614326 266707 614378 266759
rect 308086 266633 308138 266685
rect 390934 266633 390986 266685
rect 400630 266633 400682 266685
rect 620182 266633 620234 266685
rect 310678 266559 310730 266611
rect 398038 266559 398090 266611
rect 403222 266559 403274 266611
rect 627286 266559 627338 266611
rect 313558 266485 313610 266537
rect 405046 266485 405098 266537
rect 406102 266485 406154 266537
rect 634390 266485 634442 266537
rect 187222 266411 187274 266463
rect 189718 266411 189770 266463
rect 313078 266411 313130 266463
rect 403894 266411 403946 266463
rect 409174 266411 409226 266463
rect 641494 266411 641546 266463
rect 44950 266337 45002 266389
rect 671638 266337 671690 266389
rect 348886 266263 348938 266315
rect 492598 266263 492650 266315
rect 346006 266189 346058 266241
rect 485494 266189 485546 266241
rect 343318 266115 343370 266167
rect 478390 266115 478442 266167
rect 340246 266041 340298 266093
rect 471286 266041 471338 266093
rect 337366 265967 337418 266019
rect 464182 265967 464234 266019
rect 334774 265893 334826 265945
rect 457078 265893 457130 265945
rect 331894 265819 331946 265871
rect 449974 265819 450026 265871
rect 327574 265745 327626 265797
rect 439318 265745 439370 265797
rect 324502 265671 324554 265723
rect 432310 265671 432362 265723
rect 321622 265597 321674 265649
rect 425206 265597 425258 265649
rect 408022 265523 408074 265575
rect 508246 265523 508298 265575
rect 319030 265449 319082 265501
rect 418102 265449 418154 265501
rect 656566 265375 656618 265427
rect 676054 265375 676106 265427
rect 656278 265227 656330 265279
rect 676246 265227 676298 265279
rect 673270 265153 673322 265205
rect 676054 265153 676106 265205
rect 656086 265079 656138 265131
rect 676150 265079 676202 265131
rect 23062 265005 23114 265057
rect 43510 265005 43562 265057
rect 671638 265005 671690 265057
rect 673366 265005 673418 265057
rect 676054 265005 676106 265057
rect 43222 264931 43274 264983
rect 44086 264931 44138 264983
rect 669814 264931 669866 264983
rect 43318 264857 43370 264909
rect 44182 264857 44234 264909
rect 669622 264857 669674 264909
rect 359446 264783 359498 264835
rect 475990 264783 476042 264835
rect 328054 264709 328106 264761
rect 440566 264709 440618 264761
rect 331126 264635 331178 264687
rect 447670 264635 447722 264687
rect 354262 264561 354314 264613
rect 461782 264561 461834 264613
rect 360406 264487 360458 264539
rect 468886 264487 468938 264539
rect 351382 264413 351434 264465
rect 454774 264413 454826 264465
rect 399382 264117 399434 264169
rect 410998 264117 411050 264169
rect 324982 264043 325034 264095
rect 433462 264043 433514 264095
rect 387958 263969 388010 264021
rect 589462 263969 589514 264021
rect 390838 263895 390890 263947
rect 596566 263895 596618 263947
rect 393910 263821 393962 263873
rect 603670 263821 603722 263873
rect 396790 263747 396842 263799
rect 610774 263747 610826 263799
rect 401110 263673 401162 263725
rect 23350 263599 23402 263651
rect 44182 263599 44234 263651
rect 403990 263599 404042 263651
rect 410998 263673 411050 263725
rect 617878 263673 617930 263725
rect 23254 263525 23306 263577
rect 44086 263525 44138 263577
rect 409654 263525 409706 263577
rect 621430 263599 621482 263651
rect 628438 263525 628490 263577
rect 642646 263451 642698 263503
rect 23158 262119 23210 262171
rect 43318 262119 43370 262171
rect 420406 262119 420458 262171
rect 606166 262119 606218 262171
rect 674710 259307 674762 259359
rect 675958 259307 676010 259359
rect 420406 259233 420458 259285
rect 606262 259233 606314 259285
rect 675190 259233 675242 259285
rect 676054 259233 676106 259285
rect 674614 256939 674666 256991
rect 676054 256939 676106 256991
rect 674806 256421 674858 256473
rect 676054 256421 676106 256473
rect 40246 256347 40298 256399
rect 59062 256347 59114 256399
rect 420406 256347 420458 256399
rect 606358 256347 606410 256399
rect 674902 256347 674954 256399
rect 676246 256347 676298 256399
rect 41782 255385 41834 255437
rect 53206 255385 53258 255437
rect 47830 255089 47882 255141
rect 186070 255089 186122 255141
rect 47446 255015 47498 255067
rect 185974 255015 186026 255067
rect 41782 254941 41834 254993
rect 43414 254941 43466 254993
rect 47926 254941 47978 254993
rect 186550 254941 186602 254993
rect 48022 254867 48074 254919
rect 186742 254867 186794 254919
rect 41782 254423 41834 254475
rect 43414 254423 43466 254475
rect 674998 253535 675050 253587
rect 676054 253535 676106 253587
rect 41590 253461 41642 253513
rect 56182 253461 56234 253513
rect 420406 253461 420458 253513
rect 603286 253461 603338 253513
rect 646678 253461 646730 253513
rect 679702 253461 679754 253513
rect 106486 252277 106538 252329
rect 156886 252277 156938 252329
rect 92086 252203 92138 252255
rect 145462 252203 145514 252255
rect 109366 252129 109418 252181
rect 171286 252129 171338 252181
rect 97846 252055 97898 252107
rect 182806 252055 182858 252107
rect 56086 251981 56138 252033
rect 186358 251981 186410 252033
rect 666646 250649 666698 250701
rect 675382 250649 675434 250701
rect 420406 250575 420458 250627
rect 603382 250575 603434 250627
rect 120886 249909 120938 249961
rect 145654 249909 145706 249961
rect 132406 249835 132458 249887
rect 159862 249835 159914 249887
rect 135286 249761 135338 249813
rect 168502 249761 168554 249813
rect 138166 249687 138218 249739
rect 171478 249687 171530 249739
rect 141046 249613 141098 249665
rect 180022 249613 180074 249665
rect 123766 249539 123818 249591
rect 165718 249539 165770 249591
rect 126646 249465 126698 249517
rect 177046 249465 177098 249517
rect 94966 249391 95018 249443
rect 154006 249391 154058 249443
rect 118006 249317 118058 249369
rect 182902 249317 182954 249369
rect 77686 249243 77738 249295
rect 145366 249243 145418 249295
rect 80566 249169 80618 249221
rect 162646 249169 162698 249221
rect 86326 249095 86378 249147
rect 174166 249095 174218 249147
rect 675190 247911 675242 247963
rect 675382 247911 675434 247963
rect 420310 247763 420362 247815
rect 603478 247763 603530 247815
rect 420406 247689 420458 247741
rect 629206 247689 629258 247741
rect 655894 247615 655946 247667
rect 666646 247615 666698 247667
rect 674710 247245 674762 247297
rect 675478 247245 675530 247297
rect 103606 246727 103658 246779
rect 165526 246727 165578 246779
rect 112246 246653 112298 246705
rect 185782 246653 185834 246705
rect 47638 246579 47690 246631
rect 186262 246579 186314 246631
rect 674614 246579 674666 246631
rect 675382 246579 675434 246631
rect 47542 246505 47594 246557
rect 186454 246505 186506 246557
rect 47734 246431 47786 246483
rect 186646 246431 186698 246483
rect 45814 246357 45866 246409
rect 187030 246357 187082 246409
rect 45430 246283 45482 246335
rect 186838 246283 186890 246335
rect 44566 246209 44618 246261
rect 186166 246209 186218 246261
rect 674902 246061 674954 246113
rect 675382 246061 675434 246113
rect 41590 244951 41642 245003
rect 145558 244951 145610 245003
rect 44758 244877 44810 244929
rect 186934 244877 186986 244929
rect 41782 244803 41834 244855
rect 145750 244803 145802 244855
rect 420406 244803 420458 244855
rect 629302 244803 629354 244855
rect 41494 244655 41546 244707
rect 42934 244655 42986 244707
rect 41398 244581 41450 244633
rect 42838 244581 42890 244633
rect 41302 244507 41354 244559
rect 43030 244507 43082 244559
rect 44854 242805 44906 242857
rect 185686 242805 185738 242857
rect 44662 242731 44714 242783
rect 185590 242731 185642 242783
rect 674806 242731 674858 242783
rect 675382 242731 675434 242783
rect 44566 242657 44618 242709
rect 185878 242657 185930 242709
rect 41590 242583 41642 242635
rect 142582 242583 142634 242635
rect 41686 241991 41738 242043
rect 42742 241991 42794 242043
rect 420310 241917 420362 241969
rect 600406 241917 600458 241969
rect 674998 241547 675050 241599
rect 675478 241547 675530 241599
rect 41878 240585 41930 240637
rect 41878 240363 41930 240415
rect 380854 239919 380906 239971
rect 412054 239919 412106 239971
rect 409558 239845 409610 239897
rect 412150 239845 412202 239897
rect 360022 239771 360074 239823
rect 434614 239771 434666 239823
rect 371446 239697 371498 239749
rect 446710 239697 446762 239749
rect 378838 239623 378890 239675
rect 458806 239623 458858 239675
rect 383062 239549 383114 239601
rect 470902 239549 470954 239601
rect 394774 239475 394826 239527
rect 532822 239475 532874 239527
rect 406198 239327 406250 239379
rect 411574 239401 411626 239453
rect 541462 239401 541514 239453
rect 550870 239327 550922 239379
rect 400438 239253 400490 239305
rect 411382 239253 411434 239305
rect 411478 239253 411530 239305
rect 412246 239253 412298 239305
rect 420310 239253 420362 239305
rect 599062 239253 599114 239305
rect 341206 239179 341258 239231
rect 488278 239179 488330 239231
rect 350422 239105 350474 239157
rect 508630 239105 508682 239157
rect 368566 239031 368618 239083
rect 544822 239031 544874 239083
rect 382774 238957 382826 239009
rect 414646 238957 414698 239009
rect 324406 238883 324458 238935
rect 455158 238883 455210 238935
rect 323926 238809 323978 238861
rect 455062 238809 455114 238861
rect 326710 238735 326762 238787
rect 462550 238735 462602 238787
rect 328918 238661 328970 238713
rect 464758 238661 464810 238713
rect 329878 238587 329930 238639
rect 468598 238587 468650 238639
rect 332662 238513 332714 238565
rect 474646 238513 474698 238565
rect 335734 238439 335786 238491
rect 478198 238439 478250 238491
rect 336694 238365 336746 238417
rect 378646 238365 378698 238417
rect 397078 238365 397130 238417
rect 397750 238365 397802 238417
rect 403414 238365 403466 238417
rect 478390 238365 478442 238417
rect 338998 238291 339050 238343
rect 486742 238291 486794 238343
rect 341782 238217 341834 238269
rect 492790 238217 492842 238269
rect 345334 238143 345386 238195
rect 500278 238143 500330 238195
rect 346678 238069 346730 238121
rect 503350 238069 503402 238121
rect 349942 237995 349994 238047
rect 509398 237995 509450 238047
rect 353494 237921 353546 237973
rect 378550 237921 378602 237973
rect 378646 237921 378698 237973
rect 403414 237921 403466 237973
rect 403510 237921 403562 237973
rect 403702 237921 403754 237973
rect 407446 237921 407498 237973
rect 512758 237921 512810 237973
rect 352726 237847 352778 237899
rect 513910 237847 513962 237899
rect 355702 237773 355754 237825
rect 521494 237773 521546 237825
rect 358582 237699 358634 237751
rect 526006 237699 526058 237751
rect 275350 237625 275402 237677
rect 359926 237625 359978 237677
rect 363094 237625 363146 237677
rect 535126 237625 535178 237677
rect 277078 237551 277130 237603
rect 363670 237551 363722 237603
rect 364438 237551 364490 237603
rect 535798 237551 535850 237603
rect 317590 237477 317642 237529
rect 444502 237477 444554 237529
rect 317110 237403 317162 237455
rect 441430 237403 441482 237455
rect 314806 237329 314858 237381
rect 438358 237329 438410 237381
rect 311542 237255 311594 237307
rect 432406 237255 432458 237307
rect 308566 237181 308618 237233
rect 426358 237181 426410 237233
rect 310774 237107 310826 237159
rect 411190 237107 411242 237159
rect 305782 237033 305834 237085
rect 420310 237107 420362 237159
rect 411382 237033 411434 237085
rect 413974 237033 414026 237085
rect 300214 236959 300266 237011
rect 406774 236959 406826 237011
rect 408790 236959 408842 237011
rect 414262 236959 414314 237011
rect 279862 236885 279914 236937
rect 368950 236885 369002 236937
rect 388438 236885 388490 236937
rect 397750 236885 397802 236937
rect 405910 236885 405962 236937
rect 414454 236885 414506 236937
rect 278422 236811 278474 236863
rect 366742 236811 366794 236863
rect 378550 236811 378602 236863
rect 407446 236811 407498 236863
rect 320854 236737 320906 236789
rect 411190 236811 411242 236863
rect 428662 236811 428714 236863
rect 450454 236737 450506 236789
rect 42166 236663 42218 236715
rect 42742 236663 42794 236715
rect 377782 236663 377834 236715
rect 388726 236663 388778 236715
rect 397462 236663 397514 236715
rect 413686 236663 413738 236715
rect 400342 236589 400394 236641
rect 42742 236515 42794 236567
rect 43030 236515 43082 236567
rect 397558 236515 397610 236567
rect 413398 236515 413450 236567
rect 511606 236515 511658 236567
rect 376534 236441 376586 236493
rect 397366 236441 397418 236493
rect 412054 236441 412106 236493
rect 430102 236441 430154 236493
rect 412726 236367 412778 236419
rect 442198 236367 442250 236419
rect 391606 236293 391658 236345
rect 492022 236293 492074 236345
rect 394582 236219 394634 236271
rect 505654 236219 505706 236271
rect 222358 236071 222410 236123
rect 243958 236071 244010 236123
rect 251062 236071 251114 236123
rect 273718 236071 273770 236123
rect 277558 236071 277610 236123
rect 313942 236071 313994 236123
rect 319894 236071 319946 236123
rect 371446 236071 371498 236123
rect 371830 236071 371882 236123
rect 406198 236071 406250 236123
rect 406294 236071 406346 236123
rect 411766 236071 411818 236123
rect 208438 235997 208490 236049
rect 223222 235997 223274 236049
rect 247990 235997 248042 236049
rect 273622 235997 273674 236049
rect 280630 235997 280682 236049
rect 322006 235997 322058 236049
rect 386710 235997 386762 236049
rect 411478 235997 411530 236049
rect 207478 235923 207530 235975
rect 223990 235923 224042 235975
rect 243286 235923 243338 235975
rect 271030 235923 271082 235975
rect 279286 235923 279338 235975
rect 319606 235923 319658 235975
rect 332566 235923 332618 235975
rect 472342 235923 472394 235975
rect 209686 235849 209738 235901
rect 226198 235849 226250 235901
rect 234262 235849 234314 235901
rect 264886 235849 264938 235901
rect 273046 235849 273098 235901
rect 305014 235849 305066 235901
rect 343510 235849 343562 235901
rect 495766 235849 495818 235901
rect 208918 235775 208970 235827
rect 226966 235775 227018 235827
rect 237526 235775 237578 235827
rect 268150 235775 268202 235827
rect 276118 235775 276170 235827
rect 308278 235775 308330 235827
rect 348886 235775 348938 235827
rect 394582 235775 394634 235827
rect 403606 235775 403658 235827
rect 588886 235775 588938 235827
rect 211222 235701 211274 235753
rect 229270 235701 229322 235753
rect 231190 235701 231242 235753
rect 259030 235701 259082 235753
rect 262870 235701 262922 235753
rect 305110 235701 305162 235753
rect 313846 235701 313898 235753
rect 360022 235701 360074 235753
rect 393430 235701 393482 235753
rect 587062 235701 587114 235753
rect 210646 235627 210698 235679
rect 230038 235627 230090 235679
rect 236470 235627 236522 235679
rect 282934 235627 282986 235679
rect 285142 235627 285194 235679
rect 323830 235627 323882 235679
rect 326134 235627 326186 235679
rect 378838 235627 378890 235679
rect 385846 235627 385898 235679
rect 580342 235627 580394 235679
rect 210070 235553 210122 235605
rect 227830 235553 227882 235605
rect 239350 235553 239402 235605
rect 285334 235553 285386 235605
rect 286678 235553 286730 235605
rect 326710 235553 326762 235605
rect 332182 235553 332234 235605
rect 383062 235553 383114 235605
rect 392182 235553 392234 235605
rect 586294 235553 586346 235605
rect 212950 235479 213002 235531
rect 232342 235479 232394 235531
rect 249718 235479 249770 235531
rect 302326 235479 302378 235531
rect 309334 235479 309386 235531
rect 362806 235479 362858 235531
rect 387670 235479 387722 235531
rect 583414 235479 583466 235531
rect 42166 235405 42218 235457
rect 42934 235405 42986 235457
rect 211990 235405 212042 235457
rect 233014 235405 233066 235457
rect 238006 235405 238058 235457
rect 285910 235405 285962 235457
rect 295222 235405 295274 235457
rect 348694 235405 348746 235457
rect 389878 235405 389930 235457
rect 587926 235405 587978 235457
rect 214198 235331 214250 235383
rect 235318 235331 235370 235383
rect 242134 235331 242186 235383
rect 293398 235331 293450 235383
rect 299830 235331 299882 235383
rect 356470 235331 356522 235383
rect 206998 235257 207050 235309
rect 221782 235257 221834 235309
rect 223894 235257 223946 235309
rect 244726 235257 244778 235309
rect 246646 235257 246698 235309
rect 299254 235257 299306 235309
rect 301750 235257 301802 235309
rect 358582 235257 358634 235309
rect 361366 235257 361418 235309
rect 385750 235331 385802 235383
rect 394870 235331 394922 235383
rect 597718 235331 597770 235383
rect 370198 235257 370250 235309
rect 385942 235257 385994 235309
rect 394966 235257 395018 235309
rect 598486 235257 598538 235309
rect 220630 235183 220682 235235
rect 240502 235183 240554 235235
rect 240598 235183 240650 235235
rect 290422 235183 290474 235235
rect 342550 235183 342602 235235
rect 391606 235183 391658 235235
rect 396310 235183 396362 235235
rect 600790 235183 600842 235235
rect 211606 235109 211658 235161
rect 230710 235109 230762 235161
rect 232918 235109 232970 235161
rect 262006 235109 262058 235161
rect 266134 235109 266186 235161
rect 324118 235109 324170 235161
rect 334966 235109 335018 235161
rect 391702 235109 391754 235161
rect 398998 235109 399050 235161
rect 605974 235109 606026 235161
rect 213430 235035 213482 235087
rect 211030 234961 211082 235013
rect 231574 234961 231626 235013
rect 235702 235035 235754 235087
rect 266422 235035 266474 235087
rect 268918 235035 268970 235087
rect 331414 235035 331466 235087
rect 333430 235035 333482 235087
rect 394678 235035 394730 235087
rect 398614 235035 398666 235087
rect 605302 235035 605354 235087
rect 235990 234961 236042 235013
rect 243862 234961 243914 235013
rect 296470 234961 296522 235013
rect 296566 234961 296618 235013
rect 360214 234961 360266 235013
rect 378454 234961 378506 235013
rect 399574 234961 399626 235013
rect 406678 234961 406730 235013
rect 621814 234961 621866 235013
rect 208822 234887 208874 234939
rect 224758 234887 224810 234939
rect 225526 234887 225578 234939
rect 260182 234887 260234 234939
rect 260278 234887 260330 234939
rect 325270 234887 325322 234939
rect 327670 234887 327722 234939
rect 392470 234887 392522 234939
rect 409174 234887 409226 234939
rect 626422 234887 626474 234939
rect 42166 234813 42218 234865
rect 42742 234813 42794 234865
rect 206518 234813 206570 234865
rect 222454 234813 222506 234865
rect 254230 234813 254282 234865
rect 306646 234813 306698 234865
rect 321622 234813 321674 234865
rect 370198 234813 370250 234865
rect 370294 234813 370346 234865
rect 386902 234813 386954 234865
rect 410806 234813 410858 234865
rect 630166 234813 630218 234865
rect 203254 234739 203306 234791
rect 205558 234665 205610 234717
rect 207286 234665 207338 234717
rect 209302 234739 209354 234791
rect 228502 234739 228554 234791
rect 229750 234739 229802 234791
rect 253558 234739 253610 234791
rect 257494 234739 257546 234791
rect 308182 234739 308234 234791
rect 315286 234739 315338 234791
rect 394870 234739 394922 234791
rect 410038 234739 410090 234791
rect 628630 234739 628682 234791
rect 215830 234665 215882 234717
rect 225142 234665 225194 234717
rect 247702 234665 247754 234717
rect 251158 234665 251210 234717
rect 304150 234665 304202 234717
rect 308470 234665 308522 234717
rect 411574 234665 411626 234717
rect 412150 234665 412202 234717
rect 632374 234665 632426 234717
rect 204790 234591 204842 234643
rect 211990 234591 212042 234643
rect 240214 234591 240266 234643
rect 264694 234591 264746 234643
rect 267478 234591 267530 234643
rect 285046 234591 285098 234643
rect 287062 234591 287114 234643
rect 318358 234591 318410 234643
rect 320278 234591 320330 234643
rect 448246 234591 448298 234643
rect 202870 234517 202922 234569
rect 214870 234517 214922 234569
rect 235606 234517 235658 234569
rect 250582 234517 250634 234569
rect 255286 234517 255338 234569
rect 278230 234517 278282 234569
rect 283894 234517 283946 234569
rect 320854 234517 320906 234569
rect 329302 234517 329354 234569
rect 449302 234517 449354 234569
rect 202006 234443 202058 234495
rect 213430 234443 213482 234495
rect 239830 234443 239882 234495
rect 260470 234443 260522 234495
rect 262486 234443 262538 234495
rect 290902 234443 290954 234495
rect 297142 234443 297194 234495
rect 319414 234443 319466 234495
rect 323542 234443 323594 234495
rect 434902 234443 434954 234495
rect 206134 234369 206186 234421
rect 221014 234369 221066 234421
rect 250486 234369 250538 234421
rect 267958 234369 268010 234421
rect 271606 234369 271658 234421
rect 302230 234369 302282 234421
rect 207862 234295 207914 234347
rect 200278 234221 200330 234273
rect 210358 234221 210410 234273
rect 200182 234147 200234 234199
rect 208822 234147 208874 234199
rect 237046 234295 237098 234347
rect 258454 234295 258506 234347
rect 261238 234295 261290 234347
rect 288022 234295 288074 234347
rect 292918 234295 292970 234347
rect 313846 234369 313898 234421
rect 314422 234369 314474 234421
rect 423382 234369 423434 234421
rect 312694 234295 312746 234347
rect 418294 234295 418346 234347
rect 211990 234221 212042 234273
rect 219382 234221 219434 234273
rect 256534 234221 256586 234273
rect 278134 234221 278186 234273
rect 290326 234221 290378 234273
rect 334294 234221 334346 234273
rect 339478 234221 339530 234273
rect 378646 234221 378698 234273
rect 378838 234221 378890 234273
rect 400054 234221 400106 234273
rect 403702 234221 403754 234273
rect 501046 234221 501098 234273
rect 225526 234147 225578 234199
rect 244342 234147 244394 234199
rect 263638 234147 263690 234199
rect 268534 234147 268586 234199
rect 293782 234147 293834 234199
rect 295702 234147 295754 234199
rect 342358 234147 342410 234199
rect 345910 234147 345962 234199
rect 400150 234147 400202 234199
rect 401782 234147 401834 234199
rect 484630 234147 484682 234199
rect 198742 234073 198794 234125
rect 207382 234073 207434 234125
rect 247414 234073 247466 234125
rect 266326 234073 266378 234125
rect 267094 234073 267146 234125
rect 290998 234073 291050 234125
rect 294454 234073 294506 234125
rect 331222 234073 331274 234125
rect 338038 234073 338090 234125
rect 378550 234073 378602 234125
rect 378646 234073 378698 234125
rect 394582 234073 394634 234125
rect 396694 234073 396746 234125
rect 475222 234073 475274 234125
rect 42070 233999 42122 234051
rect 42838 233999 42890 234051
rect 198358 233999 198410 234051
rect 205942 233999 205994 234051
rect 197494 233925 197546 233977
rect 204310 233925 204362 233977
rect 204406 233925 204458 233977
rect 217942 233999 217994 234051
rect 259798 233999 259850 234051
rect 282070 233999 282122 234051
rect 305206 233999 305258 234051
rect 351382 233999 351434 234051
rect 358006 233999 358058 234051
rect 378838 233999 378890 234051
rect 395926 233999 395978 234051
rect 398134 233999 398186 234051
rect 398230 233999 398282 234051
rect 405238 233999 405290 234051
rect 206902 233925 206954 233977
rect 220246 233925 220298 233977
rect 258358 233925 258410 233977
rect 277078 233925 277130 233977
rect 294838 233925 294890 233977
rect 339766 233925 339818 233977
rect 361270 233925 361322 233977
rect 432022 233925 432074 233977
rect 199126 233851 199178 233903
rect 205078 233851 205130 233903
rect 205174 233851 205226 233903
rect 196918 233777 196970 233829
rect 202870 233777 202922 233829
rect 204214 233777 204266 233829
rect 215542 233777 215594 233829
rect 196534 233703 196586 233755
rect 200566 233703 200618 233755
rect 201526 233703 201578 233755
rect 211894 233703 211946 233755
rect 215830 233851 215882 233903
rect 216502 233851 216554 233903
rect 253462 233851 253514 233903
rect 270838 233851 270890 233903
rect 296086 233851 296138 233903
rect 339094 233851 339146 233903
rect 352150 233851 352202 233903
rect 361078 233851 361130 233903
rect 378550 233851 378602 233903
rect 386806 233851 386858 233903
rect 386902 233851 386954 233903
rect 427894 233851 427946 233903
rect 306262 233777 306314 233829
rect 345526 233777 345578 233829
rect 354934 233777 354986 233829
rect 404662 233777 404714 233829
rect 217174 233703 217226 233755
rect 297238 233703 297290 233755
rect 328342 233703 328394 233755
rect 330742 233703 330794 233755
rect 371638 233703 371690 233755
rect 383638 233703 383690 233755
rect 407638 233703 407690 233755
rect 195670 233629 195722 233681
rect 201334 233629 201386 233681
rect 202486 233629 202538 233681
rect 212566 233629 212618 233681
rect 302902 233629 302954 233681
rect 334102 233629 334154 233681
rect 360310 233629 360362 233681
rect 360982 233629 361034 233681
rect 361078 233629 361130 233681
rect 400342 233629 400394 233681
rect 192886 233555 192938 233607
rect 195286 233555 195338 233607
rect 195574 233555 195626 233607
rect 199798 233555 199850 233607
rect 201046 233555 201098 233607
rect 209686 233555 209738 233607
rect 194230 233481 194282 233533
rect 198358 233481 198410 233533
rect 200662 233481 200714 233533
rect 208150 233481 208202 233533
rect 194614 233407 194666 233459
rect 196054 233407 196106 233459
rect 196150 233407 196202 233459
rect 199126 233407 199178 233459
rect 199702 233407 199754 233459
rect 206614 233407 206666 233459
rect 207286 233407 207338 233459
rect 218710 233555 218762 233607
rect 283990 233555 284042 233607
rect 311254 233555 311306 233607
rect 319510 233555 319562 233607
rect 328150 233555 328202 233607
rect 335350 233555 335402 233607
rect 463606 233555 463658 233607
rect 259894 233481 259946 233533
rect 267766 233481 267818 233533
rect 287446 233481 287498 233533
rect 311350 233481 311402 233533
rect 324790 233481 324842 233533
rect 325942 233481 325994 233533
rect 326230 233481 326282 233533
rect 460246 233481 460298 233533
rect 226678 233407 226730 233459
rect 236758 233407 236810 233459
rect 264406 233407 264458 233459
rect 272374 233407 272426 233459
rect 288406 233407 288458 233459
rect 311062 233407 311114 233459
rect 317206 233407 317258 233459
rect 412726 233407 412778 233459
rect 192406 233333 192458 233385
rect 193750 233333 193802 233385
rect 193846 233333 193898 233385
rect 196822 233333 196874 233385
rect 197974 233333 198026 233385
rect 203638 233333 203690 233385
rect 203926 233333 203978 233385
rect 214198 233333 214250 233385
rect 228406 233333 228458 233385
rect 238966 233333 239018 233385
rect 257974 233333 258026 233385
rect 269878 233333 269930 233385
rect 270550 233333 270602 233385
rect 274678 233333 274730 233385
rect 282550 233333 282602 233385
rect 299158 233333 299210 233385
rect 311158 233333 311210 233385
rect 412054 233333 412106 233385
rect 193462 233259 193514 233311
rect 194614 233259 194666 233311
rect 195190 233259 195242 233311
rect 197494 233259 197546 233311
rect 197878 233259 197930 233311
rect 202102 233259 202154 233311
rect 202390 233259 202442 233311
rect 211126 233259 211178 233311
rect 242902 233259 242954 233311
rect 259510 233259 259562 233311
rect 261622 233259 261674 233311
rect 269590 233259 269642 233311
rect 270262 233259 270314 233311
rect 273334 233259 273386 233311
rect 285334 233259 285386 233311
rect 287446 233259 287498 233311
rect 288886 233259 288938 233311
rect 346966 233259 347018 233311
rect 362518 233259 362570 233311
rect 394774 233259 394826 233311
rect 400246 233259 400298 233311
rect 479158 233259 479210 233311
rect 258742 233185 258794 233237
rect 326614 233185 326666 233237
rect 340822 233185 340874 233237
rect 491254 233185 491306 233237
rect 501046 233185 501098 233237
rect 614998 233185 615050 233237
rect 262102 233111 262154 233163
rect 334198 233111 334250 233163
rect 347062 233111 347114 233163
rect 260662 233037 260714 233089
rect 331318 233037 331370 233089
rect 350326 233037 350378 233089
rect 265750 232963 265802 233015
rect 338038 232963 338090 233015
rect 353110 232963 353162 233015
rect 500854 232963 500906 233015
rect 501046 233037 501098 233089
rect 507094 232963 507146 233015
rect 289942 232889 289994 232941
rect 382198 232889 382250 232941
rect 411766 232889 411818 232941
rect 572086 232889 572138 232941
rect 263926 232815 263978 232867
rect 337270 232815 337322 232867
rect 339190 232815 339242 232867
rect 356086 232815 356138 232867
rect 356278 232815 356330 232867
rect 519190 232815 519242 232867
rect 237622 232741 237674 232793
rect 284374 232741 284426 232793
rect 295318 232741 295370 232793
rect 397366 232741 397418 232793
rect 399574 232741 399626 232793
rect 566710 232741 566762 232793
rect 216598 232667 216650 232719
rect 242134 232667 242186 232719
rect 265174 232667 265226 232719
rect 340246 232667 340298 232719
rect 362134 232667 362186 232719
rect 531286 232667 531338 232719
rect 218038 232593 218090 232645
rect 245110 232593 245162 232645
rect 268438 232593 268490 232645
rect 346294 232593 346346 232645
rect 365398 232593 365450 232645
rect 537238 232593 537290 232645
rect 219766 232519 219818 232571
rect 248086 232519 248138 232571
rect 266614 232519 266666 232571
rect 221110 232445 221162 232497
rect 251158 232445 251210 232497
rect 271222 232445 271274 232497
rect 339286 232445 339338 232497
rect 339478 232519 339530 232571
rect 361366 232519 361418 232571
rect 368182 232519 368234 232571
rect 543382 232519 543434 232571
rect 343222 232445 343274 232497
rect 344182 232445 344234 232497
rect 355318 232445 355370 232497
rect 365014 232445 365066 232497
rect 539542 232445 539594 232497
rect 222550 232371 222602 232423
rect 254230 232371 254282 232423
rect 269686 232371 269738 232423
rect 349366 232371 349418 232423
rect 366262 232371 366314 232423
rect 542614 232371 542666 232423
rect 222934 232297 222986 232349
rect 255670 232297 255722 232349
rect 274870 232297 274922 232349
rect 339190 232297 339242 232349
rect 339286 232297 339338 232349
rect 352342 232297 352394 232349
rect 371158 232297 371210 232349
rect 549430 232297 549482 232349
rect 224278 232223 224330 232275
rect 257206 232223 257258 232275
rect 272950 232223 273002 232275
rect 344182 232223 344234 232275
rect 344278 232223 344330 232275
rect 358486 232223 358538 232275
rect 369526 232223 369578 232275
rect 548566 232223 548618 232275
rect 147862 232149 147914 232201
rect 154102 232149 154154 232201
rect 226294 232149 226346 232201
rect 261718 232149 261770 232201
rect 274198 232149 274250 232201
rect 227062 232075 227114 232127
rect 263254 232075 263306 232127
rect 275734 232075 275786 232127
rect 339478 232075 339530 232127
rect 356470 232149 356522 232201
rect 365206 232149 365258 232201
rect 368086 232149 368138 232201
rect 545590 232149 545642 232201
rect 358198 232075 358250 232127
rect 358582 232075 358634 232127
rect 362230 232075 362282 232127
rect 233878 232001 233930 232053
rect 274486 232001 274538 232053
rect 277462 232001 277514 232053
rect 364438 232001 364490 232053
rect 233206 231927 233258 231979
rect 275350 231927 275402 231979
rect 280246 231927 280298 231979
rect 370390 232075 370442 232127
rect 372694 232075 372746 232127
rect 552406 232075 552458 232127
rect 234838 231853 234890 231905
rect 278326 231853 278378 231905
rect 278998 231853 279050 231905
rect 367414 231853 367466 231905
rect 236086 231779 236138 231831
rect 281302 231779 281354 231831
rect 281974 231779 282026 231831
rect 373462 232001 373514 232053
rect 372310 231927 372362 231979
rect 554710 232001 554762 232053
rect 375766 231927 375818 231979
rect 558454 231927 558506 231979
rect 374518 231853 374570 231905
rect 557014 231853 557066 231905
rect 374038 231779 374090 231831
rect 557686 231779 557738 231831
rect 259126 231705 259178 231757
rect 328054 231705 328106 231757
rect 358486 231705 358538 231757
rect 495094 231705 495146 231757
rect 500854 231705 500906 231757
rect 513142 231705 513194 231757
rect 257590 231631 257642 231683
rect 325174 231631 325226 231683
rect 337558 231631 337610 231683
rect 485206 231631 485258 231683
rect 256150 231557 256202 231609
rect 322102 231557 322154 231609
rect 328150 231557 328202 231609
rect 448918 231557 448970 231609
rect 248374 231483 248426 231535
rect 305494 231483 305546 231535
rect 312214 231483 312266 231535
rect 433846 231483 433898 231535
rect 281206 231409 281258 231461
rect 289654 231409 289706 231461
rect 292534 231409 292586 231461
rect 379990 231409 380042 231461
rect 402550 231409 402602 231461
rect 520726 231409 520778 231461
rect 290806 231335 290858 231387
rect 374614 231335 374666 231387
rect 400150 231335 400202 231387
rect 499606 231335 499658 231387
rect 293110 231261 293162 231313
rect 372790 231261 372842 231313
rect 394582 231261 394634 231313
rect 485974 231261 486026 231313
rect 255766 231187 255818 231239
rect 320662 231187 320714 231239
rect 334102 231187 334154 231239
rect 415702 231187 415754 231239
rect 293494 231113 293546 231165
rect 364054 231113 364106 231165
rect 394678 231113 394730 231165
rect 473878 231113 473930 231165
rect 252982 231039 253034 231091
rect 314518 231039 314570 231091
rect 345526 231039 345578 231091
rect 419254 231039 419306 231091
rect 245206 230965 245258 231017
rect 299446 230965 299498 231017
rect 308182 230965 308234 231017
rect 323638 230965 323690 231017
rect 328342 230965 328394 231017
rect 401398 230965 401450 231017
rect 411574 230965 411626 231017
rect 424054 230965 424106 231017
rect 325270 230891 325322 230943
rect 329590 230891 329642 230943
rect 331222 230891 331274 230943
rect 395350 230891 395402 230943
rect 326710 230817 326762 230869
rect 352726 230817 352778 230869
rect 358774 230817 358826 230869
rect 377110 230817 377162 230869
rect 385942 230817 385994 230869
rect 449686 230817 449738 230869
rect 319606 230743 319658 230795
rect 358582 230743 358634 230795
rect 358870 230743 358922 230795
rect 365110 230743 365162 230795
rect 365206 230743 365258 230795
rect 409654 230743 409706 230795
rect 320854 230669 320906 230721
rect 290614 230595 290666 230647
rect 297334 230595 297386 230647
rect 302326 230595 302378 230647
rect 308566 230595 308618 230647
rect 313942 230595 313994 230647
rect 358390 230595 358442 230647
rect 306646 230521 306698 230573
rect 317590 230521 317642 230573
rect 323830 230521 323882 230573
rect 359062 230669 359114 230721
rect 380278 230669 380330 230721
rect 358582 230595 358634 230647
rect 362134 230595 362186 230647
rect 362230 230595 362282 230647
rect 410518 230595 410570 230647
rect 149398 230447 149450 230499
rect 156982 230447 157034 230499
rect 299254 230447 299306 230499
rect 302518 230447 302570 230499
rect 304150 230447 304202 230499
rect 311638 230447 311690 230499
rect 322006 230447 322058 230499
rect 358294 230447 358346 230499
rect 374230 230521 374282 230573
rect 358678 230447 358730 230499
rect 358774 230447 358826 230499
rect 368182 230447 368234 230499
rect 423382 230447 423434 230499
rect 436150 230447 436202 230499
rect 241078 230373 241130 230425
rect 291958 230373 292010 230425
rect 314902 230373 314954 230425
rect 439990 230373 440042 230425
rect 245782 230299 245834 230351
rect 300982 230299 301034 230351
rect 321238 230299 321290 230351
rect 248950 230225 249002 230277
rect 304822 230225 304874 230277
rect 305014 230225 305066 230277
rect 326806 230225 326858 230277
rect 329206 230299 329258 230351
rect 445942 230299 445994 230351
rect 449302 230299 449354 230351
rect 466390 230299 466442 230351
rect 451990 230225 452042 230277
rect 228886 230151 228938 230203
rect 267862 230151 267914 230203
rect 269878 230151 269930 230203
rect 322966 230151 323018 230203
rect 325750 230151 325802 230203
rect 461014 230151 461066 230203
rect 463606 230151 463658 230203
rect 478294 230151 478346 230203
rect 248758 230077 248810 230129
rect 307030 230077 307082 230129
rect 324022 230077 324074 230129
rect 458038 230077 458090 230129
rect 466486 230077 466538 230129
rect 484438 230077 484490 230129
rect 227446 230003 227498 230055
rect 264790 230003 264842 230055
rect 290902 230003 290954 230055
rect 331894 230003 331946 230055
rect 475222 230003 475274 230055
rect 601462 230003 601514 230055
rect 251926 229929 251978 229981
rect 310774 229929 310826 229981
rect 317974 229929 318026 229981
rect 329206 229929 329258 229981
rect 331606 229929 331658 229981
rect 473110 229929 473162 229981
rect 479158 229929 479210 229981
rect 609046 229929 609098 229981
rect 250294 229855 250346 229907
rect 310006 229855 310058 229907
rect 336310 229855 336362 229907
rect 482134 229855 482186 229907
rect 484630 229855 484682 229907
rect 612118 229855 612170 229907
rect 146902 229781 146954 229833
rect 151222 229781 151274 229833
rect 251542 229781 251594 229833
rect 313078 229781 313130 229833
rect 328534 229781 328586 229833
rect 331126 229781 331178 229833
rect 348502 229781 348554 229833
rect 504022 229781 504074 229833
rect 506806 229781 506858 229833
rect 622678 229781 622730 229833
rect 244246 229707 244298 229759
rect 298006 229707 298058 229759
rect 298582 229707 298634 229759
rect 406774 229707 406826 229759
rect 411478 229707 411530 229759
rect 565942 229707 565994 229759
rect 215254 229633 215306 229685
rect 239062 229633 239114 229685
rect 253078 229633 253130 229685
rect 316150 229633 316202 229685
rect 351766 229633 351818 229685
rect 510166 229633 510218 229685
rect 220150 229559 220202 229611
rect 249718 229559 249770 229611
rect 255190 229559 255242 229611
rect 316822 229559 316874 229611
rect 354838 229559 354890 229611
rect 516118 229559 516170 229611
rect 221590 229485 221642 229537
rect 252598 229485 252650 229537
rect 254806 229485 254858 229537
rect 319126 229485 319178 229537
rect 357622 229485 357674 229537
rect 522166 229485 522218 229537
rect 264310 229411 264362 229463
rect 334966 229411 335018 229463
rect 366646 229411 366698 229463
rect 230614 229337 230666 229389
rect 270742 229337 270794 229389
rect 273334 229337 273386 229389
rect 347062 229337 347114 229389
rect 230326 229263 230378 229315
rect 269302 229263 269354 229315
rect 283510 229263 283562 229315
rect 367030 229337 367082 229389
rect 369910 229411 369962 229463
rect 371446 229411 371498 229463
rect 377206 229411 377258 229463
rect 538870 229411 538922 229463
rect 540310 229337 540362 229389
rect 233494 229189 233546 229241
rect 276790 229189 276842 229241
rect 282166 229189 282218 229241
rect 371254 229263 371306 229315
rect 371446 229263 371498 229315
rect 546358 229263 546410 229315
rect 231958 229115 232010 229167
rect 273814 229115 273866 229167
rect 284758 229115 284810 229167
rect 371542 229189 371594 229241
rect 374326 229189 374378 229241
rect 555382 229189 555434 229241
rect 235222 229041 235274 229093
rect 279862 229041 279914 229093
rect 286294 229041 286346 229093
rect 374518 229115 374570 229167
rect 377014 229115 377066 229167
rect 561430 229115 561482 229167
rect 380470 229041 380522 229093
rect 567478 229041 567530 229093
rect 238390 228967 238442 229019
rect 283606 228967 283658 229019
rect 287926 228967 287978 229019
rect 374422 228967 374474 229019
rect 379894 228967 379946 229019
rect 569782 228967 569834 229019
rect 246166 228893 246218 228945
rect 298678 228893 298730 228945
rect 308950 228893 309002 228945
rect 427798 228893 427850 228945
rect 427894 228893 427946 228945
rect 547894 228893 547946 228945
rect 242518 228819 242570 228871
rect 294934 228819 294986 228871
rect 310678 228819 310730 228871
rect 430870 228819 430922 228871
rect 432022 228819 432074 228871
rect 529750 228819 529802 228871
rect 241654 228745 241706 228797
rect 289750 228745 289802 228797
rect 304438 228745 304490 228797
rect 418774 228745 418826 228797
rect 434902 228745 434954 228797
rect 454294 228745 454346 228797
rect 239734 228671 239786 228723
rect 288886 228671 288938 228723
rect 306166 228671 306218 228723
rect 421846 228671 421898 228723
rect 231862 228597 231914 228649
rect 272278 228597 272330 228649
rect 291190 228597 291242 228649
rect 382966 228597 383018 228649
rect 404662 228597 404714 228649
rect 517654 228597 517706 228649
rect 190198 228523 190250 228575
rect 192310 228523 192362 228575
rect 228790 228523 228842 228575
rect 266230 228523 266282 228575
rect 266326 228523 266378 228575
rect 301750 228523 301802 228575
rect 303478 228523 303530 228575
rect 413494 228523 413546 228575
rect 455062 228523 455114 228575
rect 456502 228523 456554 228575
rect 478198 228523 478250 228575
rect 480694 228523 480746 228575
rect 512758 228523 512810 228575
rect 514678 228523 514730 228575
rect 535798 228523 535850 228575
rect 538006 228523 538058 228575
rect 544342 228523 544394 228575
rect 547126 228523 547178 228575
rect 567382 228523 567434 228575
rect 569014 228523 569066 228575
rect 224374 228449 224426 228501
rect 258742 228449 258794 228501
rect 260470 228449 260522 228501
rect 286678 228449 286730 228501
rect 289366 228449 289418 228501
rect 380086 228449 380138 228501
rect 407446 228449 407498 228501
rect 502582 228449 502634 228501
rect 250582 228375 250634 228427
rect 276502 228375 276554 228427
rect 288022 228375 288074 228427
rect 328918 228375 328970 228427
rect 331126 228375 331178 228427
rect 467062 228375 467114 228427
rect 535798 228375 535850 228427
rect 537910 228375 537962 228427
rect 259510 228301 259562 228353
rect 292630 228301 292682 228353
rect 293878 228301 293930 228353
rect 380758 228301 380810 228353
rect 391702 228301 391754 228353
rect 476950 228301 477002 228353
rect 270838 228227 270890 228279
rect 313846 228227 313898 228279
rect 313942 228227 313994 228279
rect 392374 228227 392426 228279
rect 392470 228227 392522 228279
rect 461878 228227 461930 228279
rect 267958 228153 268010 228205
rect 307702 228153 307754 228205
rect 311062 228153 311114 228205
rect 383254 228153 383306 228205
rect 394870 228153 394922 228205
rect 437686 228153 437738 228205
rect 293782 228079 293834 228131
rect 343990 228079 344042 228131
rect 345334 228079 345386 228131
rect 412726 228079 412778 228131
rect 258454 228005 258506 228057
rect 280630 228005 280682 228057
rect 298102 228005 298154 228057
rect 362806 228005 362858 228057
rect 362902 228005 362954 228057
rect 425590 228005 425642 228057
rect 290998 227931 291050 227983
rect 341014 227931 341066 227983
rect 342358 227931 342410 227983
rect 398326 227931 398378 227983
rect 247030 227857 247082 227909
rect 303958 227857 304010 227909
rect 308278 227857 308330 227909
rect 359158 227857 359210 227909
rect 263638 227783 263690 227835
rect 295702 227783 295754 227835
rect 302230 227783 302282 227835
rect 350038 227783 350090 227835
rect 319414 227709 319466 227761
rect 282070 227635 282122 227687
rect 325846 227635 325898 227687
rect 149398 227561 149450 227613
rect 174262 227561 174314 227613
rect 278134 227561 278186 227613
rect 319894 227561 319946 227613
rect 326806 227709 326858 227761
rect 353110 227709 353162 227761
rect 387766 227635 387818 227687
rect 396406 227635 396458 227687
rect 403702 227561 403754 227613
rect 418294 227561 418346 227613
rect 433174 227561 433226 227613
rect 187126 227487 187178 227539
rect 190774 227487 190826 227539
rect 216118 227487 216170 227539
rect 239830 227487 239882 227539
rect 249334 227487 249386 227539
rect 306262 227487 306314 227539
rect 311254 227487 311306 227539
rect 375766 227487 375818 227539
rect 389494 227487 389546 227539
rect 587158 227487 587210 227539
rect 588886 227487 588938 227539
rect 615862 227487 615914 227539
rect 238774 227413 238826 227465
rect 252022 227413 252074 227465
rect 253846 227413 253898 227465
rect 315382 227413 315434 227465
rect 318358 227413 318410 227465
rect 381814 227413 381866 227465
rect 390070 227413 390122 227465
rect 588598 227413 588650 227465
rect 588982 227413 589034 227465
rect 618838 227413 618890 227465
rect 217078 227339 217130 227391
rect 243574 227339 243626 227391
rect 311350 227339 311402 227391
rect 384022 227339 384074 227391
rect 392278 227339 392330 227391
rect 593110 227339 593162 227391
rect 606262 227339 606314 227391
rect 639190 227339 639242 227391
rect 236758 227265 236810 227317
rect 261046 227265 261098 227317
rect 274678 227265 274730 227317
rect 348598 227265 348650 227317
rect 390838 227265 390890 227317
rect 590134 227265 590186 227317
rect 599062 227265 599114 227317
rect 633142 227265 633194 227317
rect 217846 227191 217898 227243
rect 242902 227191 242954 227243
rect 253558 227191 253610 227243
rect 266998 227191 267050 227243
rect 271990 227191 272042 227243
rect 351574 227191 351626 227243
rect 388534 227191 388586 227243
rect 585622 227191 585674 227243
rect 587350 227191 587402 227243
rect 616630 227191 616682 227243
rect 215734 227117 215786 227169
rect 238390 227117 238442 227169
rect 238966 227117 239018 227169
rect 264022 227117 264074 227169
rect 264694 227117 264746 227169
rect 288118 227117 288170 227169
rect 289654 227117 289706 227169
rect 369622 227117 369674 227169
rect 385654 227117 385706 227169
rect 398806 227117 398858 227169
rect 398902 227117 398954 227169
rect 584854 227117 584906 227169
rect 587446 227117 587498 227169
rect 619606 227117 619658 227169
rect 219478 227043 219530 227095
rect 245878 227043 245930 227095
rect 276694 227043 276746 227095
rect 360598 227043 360650 227095
rect 390454 227043 390506 227095
rect 589366 227043 589418 227095
rect 606358 227043 606410 227095
rect 638518 227043 638570 227095
rect 149398 226969 149450 227021
rect 159766 226969 159818 227021
rect 213814 226969 213866 227021
rect 237526 226969 237578 227021
rect 240502 226969 240554 227021
rect 248854 226969 248906 227021
rect 275254 226969 275306 227021
rect 357622 226969 357674 227021
rect 392662 226969 392714 227021
rect 593974 226969 594026 227021
rect 603478 226969 603530 227021
rect 636214 226969 636266 227021
rect 221686 226895 221738 226947
rect 250390 226895 250442 226947
rect 273430 226895 273482 226947
rect 354550 226895 354602 226947
rect 359830 226895 359882 226947
rect 393142 226895 393194 226947
rect 395542 226895 395594 226947
rect 599158 226895 599210 226947
rect 600406 226895 600458 226947
rect 634678 226895 634730 226947
rect 223318 226821 223370 226873
rect 253462 226821 253514 226873
rect 324118 226821 324170 226873
rect 339478 226821 339530 226873
rect 364054 226821 364106 226873
rect 396118 226821 396170 226873
rect 399382 226821 399434 226873
rect 419350 226821 419402 226873
rect 419446 226821 419498 226873
rect 603670 226821 603722 226873
rect 606166 226821 606218 226873
rect 639958 226821 640010 226873
rect 224950 226747 225002 226799
rect 256438 226747 256490 226799
rect 257110 226747 257162 226799
rect 273238 226747 273290 226799
rect 279766 226747 279818 226799
rect 298198 226747 298250 226799
rect 298390 226747 298442 226799
rect 366742 226747 366794 226799
rect 374614 226747 374666 226799
rect 391510 226747 391562 226799
rect 397174 226747 397226 226799
rect 227926 226673 227978 226725
rect 262486 226673 262538 226725
rect 284662 226673 284714 226725
rect 298102 226673 298154 226725
rect 299158 226673 299210 226725
rect 372694 226673 372746 226725
rect 372790 226673 372842 226725
rect 393814 226673 393866 226725
rect 400822 226673 400874 226725
rect 602998 226747 603050 226799
rect 603382 226747 603434 226799
rect 636886 226747 636938 226799
rect 226582 226599 226634 226651
rect 259414 226599 259466 226651
rect 268150 226599 268202 226651
rect 282070 226599 282122 226651
rect 285718 226599 285770 226651
rect 378742 226599 378794 226651
rect 379990 226599 380042 226651
rect 394582 226599 394634 226651
rect 397654 226599 397706 226651
rect 418678 226599 418730 226651
rect 419638 226673 419690 226725
rect 606742 226673 606794 226725
rect 609814 226599 609866 226651
rect 629302 226599 629354 226651
rect 634006 226599 634058 226651
rect 229558 226525 229610 226577
rect 265558 226525 265610 226577
rect 271030 226525 271082 226577
rect 294262 226525 294314 226577
rect 297334 226525 297386 226577
rect 390070 226525 390122 226577
rect 401206 226525 401258 226577
rect 610486 226525 610538 226577
rect 231094 226451 231146 226503
rect 268534 226451 268586 226503
rect 288502 226451 288554 226503
rect 232534 226377 232586 226429
rect 271606 226377 271658 226429
rect 298102 226377 298154 226429
rect 378070 226377 378122 226429
rect 380566 226451 380618 226503
rect 387766 226451 387818 226503
rect 388150 226451 388202 226503
rect 398902 226451 398954 226503
rect 402166 226451 402218 226503
rect 612790 226451 612842 226503
rect 384790 226377 384842 226429
rect 385846 226377 385898 226429
rect 388822 226377 388874 226429
rect 388918 226377 388970 226429
rect 402838 226377 402890 226429
rect 404950 226377 405002 226429
rect 618070 226377 618122 226429
rect 212374 226303 212426 226355
rect 234550 226303 234602 226355
rect 243958 226303 244010 226355
rect 251926 226303 251978 226355
rect 252022 226303 252074 226355
rect 285142 226303 285194 226355
rect 291574 226303 291626 226355
rect 390838 226303 390890 226355
rect 398710 226303 398762 226355
rect 220342 226229 220394 226281
rect 247414 226229 247466 226281
rect 215638 226155 215690 226207
rect 240598 226155 240650 226207
rect 245014 226155 245066 226207
rect 297238 226229 297290 226281
rect 297622 226229 297674 226281
rect 388918 226229 388970 226281
rect 389014 226229 389066 226281
rect 398998 226229 399050 226281
rect 404374 226303 404426 226355
rect 617302 226303 617354 226355
rect 404470 226229 404522 226281
rect 407734 226229 407786 226281
rect 624118 226229 624170 226281
rect 151126 226081 151178 226133
rect 187126 226081 187178 226133
rect 214582 226007 214634 226059
rect 236854 226007 236906 226059
rect 241846 226007 241898 226059
rect 291190 226155 291242 226207
rect 300694 226155 300746 226207
rect 408982 226155 409034 226207
rect 418678 226155 418730 226207
rect 419446 226155 419498 226207
rect 213046 225933 213098 225985
rect 233782 225933 233834 225985
rect 246550 225933 246602 225985
rect 300214 226081 300266 226133
rect 301270 226081 301322 226133
rect 411286 226081 411338 226133
rect 411670 226081 411722 226133
rect 631702 226081 631754 226133
rect 264886 226007 264938 226059
rect 276118 226007 276170 226059
rect 334294 226007 334346 226059
rect 380566 226007 380618 226059
rect 267766 225933 267818 225985
rect 217462 225859 217514 225911
rect 241270 225859 241322 225911
rect 262006 225859 262058 225911
rect 273046 225859 273098 225911
rect 273238 225933 273290 225985
rect 321334 225933 321386 225985
rect 386998 226007 387050 226059
rect 388822 226007 388874 226059
rect 398710 226007 398762 226059
rect 398806 226007 398858 226059
rect 327382 225859 327434 225911
rect 331414 225859 331466 225911
rect 345526 225859 345578 225911
rect 346966 225859 347018 225911
rect 380758 225933 380810 225985
rect 386422 225933 386474 225985
rect 386614 225933 386666 225985
rect 398998 226007 399050 226059
rect 586390 226007 586442 226059
rect 587830 226007 587882 226059
rect 594646 226007 594698 226059
rect 603286 226007 603338 226059
rect 637750 226007 637802 226059
rect 374422 225859 374474 225911
rect 385558 225859 385610 225911
rect 387286 225859 387338 225911
rect 398614 225859 398666 225911
rect 218806 225785 218858 225837
rect 244342 225785 244394 225837
rect 269590 225785 269642 225837
rect 330454 225785 330506 225837
rect 374518 225785 374570 225837
rect 382582 225785 382634 225837
rect 382966 225785 383018 225837
rect 389302 225785 389354 225837
rect 579574 225933 579626 225985
rect 587062 225933 587114 225985
rect 595414 225933 595466 225985
rect 398902 225859 398954 225911
rect 582646 225859 582698 225911
rect 629206 225859 629258 225911
rect 635446 225859 635498 225911
rect 581110 225785 581162 225837
rect 218326 225711 218378 225763
rect 246646 225711 246698 225763
rect 247702 225711 247754 225763
rect 257974 225711 258026 225763
rect 266422 225711 266474 225763
rect 279094 225711 279146 225763
rect 285046 225711 285098 225763
rect 342550 225711 342602 225763
rect 371542 225711 371594 225763
rect 379510 225711 379562 225763
rect 380086 225711 380138 225763
rect 388630 225711 388682 225763
rect 396406 225711 396458 225763
rect 584086 225711 584138 225763
rect 278230 225637 278282 225689
rect 318358 225637 318410 225689
rect 321718 225637 321770 225689
rect 451222 225637 451274 225689
rect 244726 225563 244778 225615
rect 254902 225563 254954 225615
rect 259030 225563 259082 225615
rect 269974 225563 270026 225615
rect 273718 225563 273770 225615
rect 309334 225563 309386 225615
rect 315766 225563 315818 225615
rect 439126 225563 439178 225615
rect 273622 225489 273674 225541
rect 303190 225489 303242 225541
rect 309910 225489 309962 225541
rect 427030 225489 427082 225541
rect 306742 225415 306794 225467
rect 420982 225415 421034 225467
rect 303862 225341 303914 225393
rect 415030 225341 415082 225393
rect 302134 225267 302186 225319
rect 411958 225267 412010 225319
rect 277078 225193 277130 225245
rect 324406 225193 324458 225245
rect 351382 225193 351434 225245
rect 418006 225193 418058 225245
rect 305110 225119 305162 225171
rect 333526 225119 333578 225171
rect 339094 225119 339146 225171
rect 399958 225119 400010 225171
rect 410422 225119 410474 225171
rect 629398 225119 629450 225171
rect 252694 225045 252746 225097
rect 312310 225045 312362 225097
rect 339766 225045 339818 225097
rect 396790 225045 396842 225097
rect 272374 224971 272426 225023
rect 336406 224971 336458 225023
rect 354358 224971 354410 225023
rect 408214 225045 408266 225097
rect 348694 224897 348746 224949
rect 394390 224897 394442 224949
rect 362806 224823 362858 224875
rect 405142 224971 405194 225023
rect 147094 224749 147146 224801
rect 151318 224749 151370 224801
rect 360310 224749 360362 224801
rect 149494 224675 149546 224727
rect 162742 224675 162794 224727
rect 277942 224675 277994 224727
rect 363766 224675 363818 224727
rect 367030 224749 367082 224801
rect 376438 224749 376490 224801
rect 402166 224823 402218 224875
rect 382198 224675 382250 224727
rect 386326 224675 386378 224727
rect 386422 224675 386474 224727
rect 397654 224749 397706 224801
rect 586294 224749 586346 224801
rect 592342 224749 592394 224801
rect 397462 224675 397514 224727
rect 400630 224675 400682 224727
rect 316342 224601 316394 224653
rect 441430 224601 441482 224653
rect 323158 224527 323210 224579
rect 452758 224527 452810 224579
rect 319318 224453 319370 224505
rect 447478 224453 447530 224505
rect 322294 224379 322346 224431
rect 453430 224379 453482 224431
rect 325366 224305 325418 224357
rect 459574 224305 459626 224357
rect 328246 224231 328298 224283
rect 465622 224231 465674 224283
rect 331510 224157 331562 224209
rect 471574 224157 471626 224209
rect 334486 224083 334538 224135
rect 477622 224083 477674 224135
rect 337174 224009 337226 224061
rect 483766 224009 483818 224061
rect 340438 223935 340490 223987
rect 489718 223935 489770 223987
rect 343606 223861 343658 223913
rect 497302 223861 497354 223913
rect 261910 223787 261962 223839
rect 332662 223787 332714 223839
rect 346582 223787 346634 223839
rect 501814 223787 501866 223839
rect 263542 223713 263594 223765
rect 335734 223713 335786 223765
rect 348118 223713 348170 223765
rect 506326 223713 506378 223765
rect 266518 223639 266570 223691
rect 341782 223639 341834 223691
rect 349558 223639 349610 223691
rect 507862 223639 507914 223691
rect 264598 223565 264650 223617
rect 338710 223565 338762 223617
rect 351190 223565 351242 223617
rect 512374 223565 512426 223617
rect 268054 223491 268106 223543
rect 344854 223491 344906 223543
rect 348022 223491 348074 223543
rect 504790 223491 504842 223543
rect 270934 223417 270986 223469
rect 350806 223417 350858 223469
rect 351094 223417 351146 223469
rect 510838 223417 510890 223469
rect 269398 223343 269450 223395
rect 347734 223343 347786 223395
rect 352534 223343 352586 223395
rect 514006 223343 514058 223395
rect 355606 223269 355658 223321
rect 519862 223269 519914 223321
rect 354070 223195 354122 223247
rect 516982 223195 517034 223247
rect 318550 223121 318602 223173
rect 443734 223121 443786 223173
rect 313366 223047 313418 223099
rect 435382 223047 435434 223099
rect 310294 222973 310346 223025
rect 429334 222973 429386 223025
rect 307990 222899 308042 222951
rect 422518 222899 422570 222951
rect 312598 222825 312650 222877
rect 431542 222825 431594 222877
rect 307222 222751 307274 222803
rect 423286 222751 423338 222803
rect 304246 222677 304298 222729
rect 417238 222677 417290 222729
rect 302806 222603 302858 222655
rect 414262 222603 414314 222655
rect 304918 222529 304970 222581
rect 416470 222529 416522 222581
rect 286198 222455 286250 222507
rect 381046 222455 381098 222507
rect 396982 222455 397034 222507
rect 496534 222455 496586 222507
rect 272566 222381 272618 222433
rect 353878 222381 353930 222433
rect 371638 222381 371690 222433
rect 467830 222381 467882 222433
rect 283126 222307 283178 222359
rect 374998 222307 375050 222359
rect 386806 222307 386858 222359
rect 482902 222307 482954 222359
rect 281590 222233 281642 222285
rect 371926 222233 371978 222285
rect 394390 222233 394442 222285
rect 399094 222233 399146 222285
rect 274102 222159 274154 222211
rect 356854 222159 356906 222211
rect 149398 221863 149450 221915
rect 168406 221863 168458 221915
rect 149494 221789 149546 221841
rect 171382 221789 171434 221841
rect 656182 221789 656234 221841
rect 676246 221789 676298 221841
rect 42070 221715 42122 221767
rect 50326 221715 50378 221767
rect 145750 221715 145802 221767
rect 184342 221715 184394 221767
rect 276406 221715 276458 221767
rect 277558 221715 277610 221767
rect 478486 221715 478538 221767
rect 479974 221715 480026 221767
rect 513814 221715 513866 221767
rect 515398 221715 515450 221767
rect 147286 220753 147338 220805
rect 151414 220753 151466 220805
rect 673270 220605 673322 220657
rect 676054 220605 676106 220657
rect 673366 219495 673418 219547
rect 676054 219495 676106 219547
rect 655990 219199 656042 219251
rect 676246 219199 676298 219251
rect 655798 219051 655850 219103
rect 676150 219051 676202 219103
rect 149494 218977 149546 219029
rect 165622 218977 165674 219029
rect 149398 218903 149450 218955
rect 179926 218903 179978 218955
rect 143062 218829 143114 218881
rect 184342 218829 184394 218881
rect 149494 216091 149546 216143
rect 174358 216091 174410 216143
rect 149398 216017 149450 216069
rect 177142 216017 177194 216069
rect 149398 214685 149450 214737
rect 159958 214685 160010 214737
rect 147286 214019 147338 214071
rect 151798 214019 151850 214071
rect 41782 213279 41834 213331
rect 45718 213279 45770 213331
rect 675094 213205 675146 213257
rect 675958 213205 676010 213257
rect 675286 213131 675338 213183
rect 676054 213131 676106 213183
rect 41590 212909 41642 212961
rect 45622 212909 45674 212961
rect 146902 212835 146954 212887
rect 152086 212835 152138 212887
rect 41782 212169 41834 212221
rect 45526 212169 45578 212221
rect 674710 212095 674762 212147
rect 676054 212095 676106 212147
rect 41782 211725 41834 211777
rect 43414 211725 43466 211777
rect 41590 211429 41642 211481
rect 44854 211429 44906 211481
rect 147094 211281 147146 211333
rect 151702 211281 151754 211333
rect 41782 210689 41834 210741
rect 50614 210689 50666 210741
rect 674806 210393 674858 210445
rect 675958 210393 676010 210445
rect 147478 210319 147530 210371
rect 151606 210319 151658 210371
rect 674902 210319 674954 210371
rect 676246 210319 676298 210371
rect 674998 210245 675050 210297
rect 676054 210245 676106 210297
rect 41782 210171 41834 210223
rect 43318 210171 43370 210223
rect 41590 209949 41642 210001
rect 50422 209949 50474 210001
rect 41590 209357 41642 209409
rect 43510 209357 43562 209409
rect 147190 207877 147242 207929
rect 151510 207877 151562 207929
rect 146902 207359 146954 207411
rect 151990 207359 152042 207411
rect 646774 207359 646826 207411
rect 679798 207359 679850 207411
rect 675766 206101 675818 206153
rect 675094 205657 675146 205709
rect 675478 205657 675530 205709
rect 675766 205583 675818 205635
rect 147094 204547 147146 204599
rect 151894 204547 151946 204599
rect 149398 204473 149450 204525
rect 182998 204473 183050 204525
rect 675190 201883 675242 201935
rect 675478 201883 675530 201935
rect 149398 201735 149450 201787
rect 174454 201735 174506 201787
rect 41878 201661 41930 201713
rect 44758 201661 44810 201713
rect 149494 201661 149546 201713
rect 177238 201661 177290 201713
rect 149302 201587 149354 201639
rect 180118 201587 180170 201639
rect 143062 201513 143114 201565
rect 184342 201513 184394 201565
rect 655606 201513 655658 201565
rect 675094 201513 675146 201565
rect 41494 201439 41546 201491
rect 42934 201439 42986 201491
rect 41878 201365 41930 201417
rect 44566 201365 44618 201417
rect 41494 200921 41546 200973
rect 44662 200921 44714 200973
rect 674998 200847 675050 200899
rect 675382 200847 675434 200899
rect 41590 198923 41642 198975
rect 42742 198923 42794 198975
rect 41686 198849 41738 198901
rect 42838 198849 42890 198901
rect 41782 198775 41834 198827
rect 43030 198775 43082 198827
rect 147478 198775 147530 198827
rect 154198 198775 154250 198827
rect 149398 198701 149450 198753
rect 162838 198701 162890 198753
rect 181366 198627 181418 198679
rect 184438 198627 184490 198679
rect 178294 198553 178346 198605
rect 184342 198553 184394 198605
rect 674902 197739 674954 197791
rect 675382 197739 675434 197791
rect 41974 197369 42026 197421
rect 41974 197147 42026 197199
rect 674710 196999 674762 197051
rect 675478 196999 675530 197051
rect 674806 196555 674858 196607
rect 675382 196555 675434 196607
rect 149398 195963 149450 196015
rect 168598 195963 168650 196015
rect 149494 195889 149546 195941
rect 171574 195889 171626 195941
rect 149398 195815 149450 195867
rect 183094 195815 183146 195867
rect 166966 195741 167018 195793
rect 184534 195741 184586 195793
rect 169846 195667 169898 195719
rect 184438 195667 184490 195719
rect 172726 195593 172778 195645
rect 184342 195593 184394 195645
rect 42070 193447 42122 193499
rect 42838 193447 42890 193499
rect 149398 193151 149450 193203
rect 160054 193151 160106 193203
rect 149494 193003 149546 193055
rect 165814 193003 165866 193055
rect 152374 192929 152426 192981
rect 184630 192929 184682 192981
rect 155446 192855 155498 192907
rect 184534 192855 184586 192907
rect 158134 192781 158186 192833
rect 184342 192781 184394 192833
rect 163894 192707 163946 192759
rect 184438 192707 184490 192759
rect 42166 192189 42218 192241
rect 42742 192189 42794 192241
rect 42070 191449 42122 191501
rect 43030 191449 43082 191501
rect 42166 191005 42218 191057
rect 42934 191005 42986 191057
rect 147382 190191 147434 190243
rect 154294 190191 154346 190243
rect 149398 190117 149450 190169
rect 157078 190117 157130 190169
rect 143926 190043 143978 190095
rect 184534 190043 184586 190095
rect 149686 189969 149738 190021
rect 184342 189969 184394 190021
rect 171478 189895 171530 189947
rect 184438 189895 184490 189947
rect 180022 189821 180074 189873
rect 184342 189821 184394 189873
rect 159862 187157 159914 187209
rect 184438 187157 184490 187209
rect 165718 187083 165770 187135
rect 184534 187083 184586 187135
rect 168502 187009 168554 187061
rect 184342 187009 184394 187061
rect 177046 186935 177098 186987
rect 184630 186935 184682 186987
rect 149398 185751 149450 185803
rect 185974 185751 186026 185803
rect 145654 184271 145706 184323
rect 184342 184271 184394 184323
rect 171286 184197 171338 184249
rect 184438 184197 184490 184249
rect 182902 184123 182954 184175
rect 186742 184123 186794 184175
rect 645142 183087 645194 183139
rect 649366 183087 649418 183139
rect 149302 182939 149354 182991
rect 186262 182939 186314 182991
rect 149494 182865 149546 182917
rect 186070 182865 186122 182917
rect 42166 182199 42218 182251
rect 48118 182199 48170 182251
rect 149398 181459 149450 181511
rect 171478 181459 171530 181511
rect 182806 181385 182858 181437
rect 184630 181385 184682 181437
rect 156886 181311 156938 181363
rect 184342 181311 184394 181363
rect 165526 181237 165578 181289
rect 184438 181237 184490 181289
rect 154006 181163 154058 181215
rect 184534 181163 184586 181215
rect 149590 180053 149642 180105
rect 185494 180053 185546 180105
rect 149206 179979 149258 180031
rect 186454 179979 186506 180031
rect 645142 179387 645194 179439
rect 649462 179387 649514 179439
rect 149398 178721 149450 178773
rect 162934 178721 162986 178773
rect 149494 178647 149546 178699
rect 165718 178647 165770 178699
rect 149302 178573 149354 178625
rect 168502 178573 168554 178625
rect 145462 178499 145514 178551
rect 184438 178499 184490 178551
rect 162646 178425 162698 178477
rect 184534 178425 184586 178477
rect 174166 178351 174218 178403
rect 184342 178351 184394 178403
rect 149398 177241 149450 177293
rect 156886 177241 156938 177293
rect 655702 176131 655754 176183
rect 676246 176131 676298 176183
rect 147766 175983 147818 176035
rect 154006 175983 154058 176035
rect 655510 175983 655562 176035
rect 676342 175983 676394 176035
rect 655414 175835 655466 175887
rect 676150 175835 676202 175887
rect 145366 175613 145418 175665
rect 184342 175613 184394 175665
rect 145558 175539 145610 175591
rect 184438 175539 184490 175591
rect 645142 174873 645194 174925
rect 649558 174873 649610 174925
rect 149206 174207 149258 174259
rect 186166 174207 186218 174259
rect 149398 172801 149450 172853
rect 182806 172801 182858 172853
rect 148342 172727 148394 172779
rect 184534 172727 184586 172779
rect 149014 172653 149066 172705
rect 184630 172653 184682 172705
rect 148726 172579 148778 172631
rect 184342 172579 184394 172631
rect 148534 172505 148586 172557
rect 184438 172505 184490 172557
rect 645142 171025 645194 171077
rect 649654 171025 649706 171077
rect 675286 169989 675338 170041
rect 676246 169989 676298 170041
rect 675094 169915 675146 169967
rect 676054 169915 676106 169967
rect 148438 169841 148490 169893
rect 184534 169841 184586 169893
rect 148246 169767 148298 169819
rect 184342 169767 184394 169819
rect 149302 169693 149354 169745
rect 184630 169693 184682 169745
rect 148918 169619 148970 169671
rect 184438 169619 184490 169671
rect 645142 168213 645194 168265
rect 649846 168213 649898 168265
rect 674902 167103 674954 167155
rect 676246 167103 676298 167155
rect 674998 167029 675050 167081
rect 676054 167029 676106 167081
rect 148822 166955 148874 167007
rect 184342 166955 184394 167007
rect 148630 166881 148682 166933
rect 184438 166881 184490 166933
rect 154102 166807 154154 166859
rect 184534 166807 184586 166859
rect 674134 166215 674186 166267
rect 676054 166215 676106 166267
rect 646870 164365 646922 164417
rect 676054 164365 676106 164417
rect 647062 164291 647114 164343
rect 676246 164291 676298 164343
rect 646966 164217 647018 164269
rect 676150 164217 676202 164269
rect 151222 164069 151274 164121
rect 184534 164069 184586 164121
rect 156982 163995 157034 164047
rect 184342 163995 184394 164047
rect 159766 163921 159818 163973
rect 184438 163921 184490 163973
rect 174262 163847 174314 163899
rect 184342 163847 184394 163899
rect 645142 163329 645194 163381
rect 649942 163329 649994 163381
rect 151318 161183 151370 161235
rect 184438 161183 184490 161235
rect 162742 161109 162794 161161
rect 184534 161109 184586 161161
rect 168406 161035 168458 161087
rect 184630 161035 184682 161087
rect 171382 160961 171434 161013
rect 184342 160961 184394 161013
rect 675094 160591 675146 160643
rect 675382 160591 675434 160643
rect 645142 159703 645194 159755
rect 650038 159703 650090 159755
rect 147478 158889 147530 158941
rect 152182 158889 152234 158941
rect 151414 158371 151466 158423
rect 184342 158371 184394 158423
rect 165622 158297 165674 158349
rect 184438 158297 184490 158349
rect 179926 158223 179978 158275
rect 184534 158223 184586 158275
rect 177142 158149 177194 158201
rect 184630 158149 184682 158201
rect 674998 157039 675050 157091
rect 675478 157039 675530 157091
rect 674902 156299 674954 156351
rect 675382 156299 675434 156351
rect 146902 156151 146954 156203
rect 151222 156151 151274 156203
rect 645142 156003 645194 156055
rect 650134 156003 650186 156055
rect 149302 155707 149354 155759
rect 180022 155707 180074 155759
rect 149398 155633 149450 155685
rect 177046 155633 177098 155685
rect 151798 155485 151850 155537
rect 184534 155485 184586 155537
rect 658006 155485 658058 155537
rect 675094 155485 675146 155537
rect 152086 155411 152138 155463
rect 184630 155411 184682 155463
rect 159958 155337 160010 155389
rect 184438 155337 184490 155389
rect 174358 155263 174410 155315
rect 184342 155263 184394 155315
rect 149398 152747 149450 152799
rect 174166 152747 174218 152799
rect 149302 152673 149354 152725
rect 182902 152673 182954 152725
rect 151990 152599 152042 152651
rect 184534 152599 184586 152651
rect 151606 152525 151658 152577
rect 184438 152525 184490 152577
rect 645142 152525 645194 152577
rect 650230 152525 650282 152577
rect 151702 152451 151754 152503
rect 184342 152451 184394 152503
rect 674134 151415 674186 151467
rect 675382 151415 675434 151467
rect 149302 149935 149354 149987
rect 171382 149935 171434 149987
rect 149398 149861 149450 149913
rect 174262 149861 174314 149913
rect 149206 149787 149258 149839
rect 180214 149787 180266 149839
rect 182998 149713 183050 149765
rect 184726 149713 184778 149765
rect 151894 149639 151946 149691
rect 184438 149639 184490 149691
rect 180118 149565 180170 149617
rect 184534 149565 184586 149617
rect 151510 149491 151562 149543
rect 184342 149491 184394 149543
rect 645142 148159 645194 148211
rect 650326 148159 650378 148211
rect 149398 146975 149450 147027
rect 168406 146975 168458 147027
rect 149302 146901 149354 146953
rect 177142 146901 177194 146953
rect 154198 146827 154250 146879
rect 184534 146827 184586 146879
rect 162838 146753 162890 146805
rect 184438 146753 184490 146805
rect 174454 146679 174506 146731
rect 184342 146679 184394 146731
rect 177238 146605 177290 146657
rect 184630 146605 184682 146657
rect 147670 145717 147722 145769
rect 165526 145717 165578 145769
rect 147478 144015 147530 144067
rect 162742 144015 162794 144067
rect 183094 143941 183146 143993
rect 184630 143941 184682 143993
rect 168598 143867 168650 143919
rect 184438 143867 184490 143919
rect 171574 143793 171626 143845
rect 184342 143793 184394 143845
rect 165814 143719 165866 143771
rect 184534 143719 184586 143771
rect 147478 143349 147530 143401
rect 159862 143349 159914 143401
rect 147670 142387 147722 142439
rect 156982 142387 157034 142439
rect 149686 141203 149738 141255
rect 154102 141203 154154 141255
rect 154294 141055 154346 141107
rect 184534 141055 184586 141107
rect 157078 140981 157130 141033
rect 184438 140981 184490 141033
rect 160054 140907 160106 140959
rect 184342 140907 184394 140959
rect 147478 140315 147530 140367
rect 151126 140315 151178 140367
rect 147478 138243 147530 138295
rect 159766 138243 159818 138295
rect 148054 137059 148106 137111
rect 148438 137059 148490 137111
rect 148246 136985 148298 137037
rect 148726 136985 148778 137037
rect 148438 136911 148490 136963
rect 148630 136911 148682 136963
rect 148918 136911 148970 136963
rect 148726 136689 148778 136741
rect 149686 135431 149738 135483
rect 171286 135431 171338 135483
rect 149590 135357 149642 135409
rect 179926 135357 179978 135409
rect 168502 135283 168554 135335
rect 184438 135283 184490 135335
rect 171478 135209 171530 135261
rect 184342 135209 184394 135261
rect 177142 132545 177194 132597
rect 184726 132545 184778 132597
rect 149686 132471 149738 132523
rect 182998 132471 183050 132523
rect 154006 132397 154058 132449
rect 184630 132397 184682 132449
rect 156886 132323 156938 132375
rect 184534 132323 184586 132375
rect 162934 132249 162986 132301
rect 184438 132249 184490 132301
rect 165718 132175 165770 132227
rect 184342 132175 184394 132227
rect 180214 132027 180266 132079
rect 185590 132027 185642 132079
rect 655318 130103 655370 130155
rect 676150 130103 676202 130155
rect 655222 129955 655274 130007
rect 676246 129955 676298 130007
rect 655126 129807 655178 129859
rect 676342 129807 676394 129859
rect 147478 129659 147530 129711
rect 165622 129659 165674 129711
rect 149686 129585 149738 129637
rect 168502 129585 168554 129637
rect 645718 129585 645770 129637
rect 676246 129585 676298 129637
rect 182806 129511 182858 129563
rect 186742 129511 186794 129563
rect 149494 129437 149546 129489
rect 184438 129437 184490 129489
rect 149398 129363 149450 129415
rect 184534 129363 184586 129415
rect 149110 129289 149162 129341
rect 184342 129289 184394 129341
rect 147478 127809 147530 127861
rect 162646 127809 162698 127861
rect 646486 126921 646538 126973
rect 676246 126921 676298 126973
rect 646582 126773 646634 126825
rect 676150 126773 676202 126825
rect 674326 126699 674378 126751
rect 676054 126699 676106 126751
rect 148342 126625 148394 126677
rect 184534 126625 184586 126677
rect 148534 126551 148586 126603
rect 184438 126551 184490 126603
rect 148918 126477 148970 126529
rect 184342 126477 184394 126529
rect 149398 124183 149450 124235
rect 156886 124183 156938 124235
rect 674614 124183 674666 124235
rect 676054 124183 676106 124235
rect 674806 123961 674858 124013
rect 676054 123961 676106 124013
rect 675286 123887 675338 123939
rect 676246 123887 676298 123939
rect 148150 123813 148202 123865
rect 184630 123813 184682 123865
rect 148726 123739 148778 123791
rect 184534 123739 184586 123791
rect 148054 123665 148106 123717
rect 184438 123665 184490 123717
rect 148246 123591 148298 123643
rect 184342 123591 184394 123643
rect 174262 122407 174314 122459
rect 186166 122407 186218 122459
rect 675094 122111 675146 122163
rect 676054 122111 676106 122163
rect 674710 121149 674762 121201
rect 675958 121149 676010 121201
rect 674902 121075 674954 121127
rect 676246 121075 676298 121127
rect 674998 121001 675050 121053
rect 676054 121001 676106 121053
rect 148630 120927 148682 120979
rect 184534 120927 184586 120979
rect 148438 120853 148490 120905
rect 184342 120853 184394 120905
rect 171382 120779 171434 120831
rect 184438 120779 184490 120831
rect 147862 120483 147914 120535
rect 154486 120483 154538 120535
rect 647830 118337 647882 118389
rect 676246 118337 676298 118389
rect 149398 118189 149450 118241
rect 168598 118189 168650 118241
rect 647926 118189 647978 118241
rect 676150 118189 676202 118241
rect 149494 118115 149546 118167
rect 174262 118115 174314 118167
rect 645238 118115 645290 118167
rect 676054 118115 676106 118167
rect 159862 118041 159914 118093
rect 184630 118041 184682 118093
rect 162742 117967 162794 118019
rect 184534 117967 184586 118019
rect 165526 117893 165578 117945
rect 184438 117893 184490 117945
rect 168406 117819 168458 117871
rect 184342 117819 184394 117871
rect 675574 115969 675626 116021
rect 149398 115303 149450 115355
rect 162838 115303 162890 115355
rect 675574 115303 675626 115355
rect 149494 115229 149546 115281
rect 165718 115229 165770 115281
rect 647926 115229 647978 115281
rect 665302 115229 665354 115281
rect 670390 115229 670442 115281
rect 675478 115229 675530 115281
rect 152182 115155 152234 115207
rect 184534 115155 184586 115207
rect 154102 115081 154154 115133
rect 184438 115081 184490 115133
rect 156982 115007 157034 115059
rect 184342 115007 184394 115059
rect 180022 114119 180074 114171
rect 184630 114119 184682 114171
rect 674326 114119 674378 114171
rect 675382 114119 675434 114171
rect 149398 114045 149450 114097
rect 159862 114045 159914 114097
rect 663766 112935 663818 112987
rect 665206 112935 665258 112987
rect 674614 112491 674666 112543
rect 675382 112491 675434 112543
rect 149398 112343 149450 112395
rect 177142 112343 177194 112395
rect 151222 112269 151274 112321
rect 184342 112269 184394 112321
rect 665206 112269 665258 112321
rect 670390 112269 670442 112321
rect 182902 112195 182954 112247
rect 184534 112195 184586 112247
rect 177046 112121 177098 112173
rect 184438 112121 184490 112173
rect 674806 111825 674858 111877
rect 675382 111825 675434 111877
rect 675190 111159 675242 111211
rect 675382 111159 675434 111211
rect 674998 110641 675050 110693
rect 675382 110641 675434 110693
rect 148630 109531 148682 109583
rect 154006 109531 154058 109583
rect 149398 109457 149450 109509
rect 156982 109457 157034 109509
rect 159766 109383 159818 109435
rect 184438 109383 184490 109435
rect 174166 109309 174218 109361
rect 184342 109309 184394 109361
rect 147190 108273 147242 108325
rect 151126 108273 151178 108325
rect 674902 107533 674954 107585
rect 675382 107533 675434 107585
rect 182998 106497 183050 106549
rect 184534 106497 184586 106549
rect 171286 106423 171338 106475
rect 184342 106423 184394 106475
rect 179926 106349 179978 106401
rect 185302 106349 185354 106401
rect 674806 106349 674858 106401
rect 675382 106349 675434 106401
rect 149494 106275 149546 106327
rect 184438 106275 184490 106327
rect 154486 105091 154538 105143
rect 184726 105091 184778 105143
rect 647926 103907 647978 103959
rect 661174 103907 661226 103959
rect 645910 103685 645962 103737
rect 657526 103685 657578 103737
rect 149014 103611 149066 103663
rect 184438 103611 184490 103663
rect 149110 103537 149162 103589
rect 184630 103537 184682 103589
rect 165622 103463 165674 103515
rect 184534 103463 184586 103515
rect 168502 103389 168554 103441
rect 184342 103389 184394 103441
rect 645142 102057 645194 102109
rect 652438 102057 652490 102109
rect 149398 100799 149450 100851
rect 171286 100799 171338 100851
rect 149590 100725 149642 100777
rect 184630 100725 184682 100777
rect 149302 100651 149354 100703
rect 184438 100651 184490 100703
rect 156886 100577 156938 100629
rect 184534 100577 184586 100629
rect 162646 100503 162698 100555
rect 184342 100503 184394 100555
rect 149398 97987 149450 98039
rect 184246 97987 184298 98039
rect 149494 97913 149546 97965
rect 186166 97913 186218 97965
rect 647926 97913 647978 97965
rect 662518 97913 662570 97965
rect 148342 97839 148394 97891
rect 184342 97839 184394 97891
rect 148534 97765 148586 97817
rect 184438 97765 184490 97817
rect 642262 96433 642314 96485
rect 665206 96433 665258 96485
rect 645430 95915 645482 95967
rect 653686 95915 653738 95967
rect 149494 95101 149546 95153
rect 168214 95101 168266 95153
rect 149398 95027 149450 95079
rect 179926 95027 179978 95079
rect 162838 94953 162890 95005
rect 184630 94953 184682 95005
rect 165718 94879 165770 94931
rect 184534 94879 184586 94931
rect 168598 94805 168650 94857
rect 184438 94805 184490 94857
rect 174262 94731 174314 94783
rect 184342 94731 184394 94783
rect 646774 92659 646826 92711
rect 663094 92659 663146 92711
rect 646486 92363 646538 92415
rect 660694 92363 660746 92415
rect 645526 92289 645578 92341
rect 661750 92289 661802 92341
rect 149398 92215 149450 92267
rect 162454 92215 162506 92267
rect 646870 92215 646922 92267
rect 659830 92215 659882 92267
rect 149494 92141 149546 92193
rect 165238 92141 165290 92193
rect 646966 92141 647018 92193
rect 658870 92141 658922 92193
rect 148246 92067 148298 92119
rect 184438 92067 184490 92119
rect 156982 91993 157034 92045
rect 184534 91993 184586 92045
rect 159862 91919 159914 91971
rect 184342 91919 184394 91971
rect 177142 91845 177194 91897
rect 184630 91845 184682 91897
rect 149398 90069 149450 90121
rect 159766 90069 159818 90121
rect 148438 89181 148490 89233
rect 184534 89181 184586 89233
rect 148822 89107 148874 89159
rect 184630 89107 184682 89159
rect 151126 89033 151178 89085
rect 184438 89033 184490 89085
rect 154006 88959 154058 89011
rect 184342 88959 184394 89011
rect 645910 87479 645962 87531
rect 650902 87479 650954 87531
rect 647926 87257 647978 87309
rect 658006 87257 658058 87309
rect 647062 87035 647114 87087
rect 663286 87035 663338 87087
rect 149494 86739 149546 86791
rect 156502 86739 156554 86791
rect 148822 86443 148874 86495
rect 154102 86443 154154 86495
rect 148630 86369 148682 86421
rect 184342 86369 184394 86421
rect 148726 86295 148778 86347
rect 184438 86295 184490 86347
rect 148918 86221 148970 86273
rect 184534 86221 184586 86273
rect 645910 84149 645962 84201
rect 657046 84149 657098 84201
rect 147094 83557 147146 83609
rect 151126 83557 151178 83609
rect 646774 83557 646826 83609
rect 651766 83557 651818 83609
rect 168214 83483 168266 83535
rect 184438 83483 184490 83535
rect 640726 83483 640778 83535
rect 642262 83483 642314 83535
rect 171286 83409 171338 83461
rect 184342 83409 184394 83461
rect 647926 81855 647978 81907
rect 663286 81855 663338 81907
rect 647830 81781 647882 81833
rect 663382 81781 663434 81833
rect 657046 81633 657098 81685
rect 658582 81633 658634 81685
rect 647734 81559 647786 81611
rect 662422 81559 662474 81611
rect 647926 80745 647978 80797
rect 662518 80745 662570 80797
rect 659446 80671 659498 80723
rect 659542 80671 659594 80723
rect 149590 80597 149642 80649
rect 184438 80597 184490 80649
rect 162454 80523 162506 80575
rect 184534 80523 184586 80575
rect 165238 80449 165290 80501
rect 184342 80449 184394 80501
rect 179926 80375 179978 80427
rect 184630 80375 184682 80427
rect 149302 77711 149354 77763
rect 184438 77711 184490 77763
rect 647158 77711 647210 77763
rect 658294 77711 658346 77763
rect 149398 77637 149450 77689
rect 184534 77637 184586 77689
rect 646582 77637 646634 77689
rect 659446 77637 659498 77689
rect 156502 77563 156554 77615
rect 184630 77563 184682 77615
rect 646678 77563 646730 77615
rect 661750 77563 661802 77615
rect 159766 77489 159818 77541
rect 184342 77489 184394 77541
rect 647926 77489 647978 77541
rect 656950 77489 657002 77541
rect 646006 76083 646058 76135
rect 657526 76083 657578 76135
rect 647062 74899 647114 74951
rect 660118 74899 660170 74951
rect 148822 74825 148874 74877
rect 184534 74825 184586 74877
rect 149110 74751 149162 74803
rect 184630 74751 184682 74803
rect 151126 74677 151178 74729
rect 184438 74677 184490 74729
rect 154102 74603 154154 74655
rect 184342 74603 184394 74655
rect 647926 72161 647978 72213
rect 660694 72161 660746 72213
rect 148438 71939 148490 71991
rect 184438 71939 184490 71991
rect 149686 71865 149738 71917
rect 184534 71865 184586 71917
rect 149590 71791 149642 71843
rect 184342 71791 184394 71843
rect 647926 69571 647978 69623
rect 661462 69571 661514 69623
rect 149590 69053 149642 69105
rect 184534 69053 184586 69105
rect 148918 68979 148970 69031
rect 184342 68979 184394 69031
rect 149206 68905 149258 68957
rect 184438 68905 184490 68957
rect 149302 68831 149354 68883
rect 184342 68831 184394 68883
rect 149110 66167 149162 66219
rect 184534 66167 184586 66219
rect 646006 66167 646058 66219
rect 652342 66167 652394 66219
rect 149398 66093 149450 66145
rect 184630 66093 184682 66145
rect 149494 66019 149546 66071
rect 184438 66019 184490 66071
rect 149014 65945 149066 65997
rect 184342 65945 184394 65997
rect 647926 63577 647978 63629
rect 663190 63577 663242 63629
rect 149206 63281 149258 63333
rect 184438 63281 184490 63333
rect 149494 63207 149546 63259
rect 184534 63207 184586 63259
rect 149398 63133 149450 63185
rect 184630 63133 184682 63185
rect 149590 63059 149642 63111
rect 184342 63059 184394 63111
rect 647926 60987 647978 61039
rect 663478 60987 663530 61039
rect 149302 60395 149354 60447
rect 184438 60395 184490 60447
rect 149494 60321 149546 60373
rect 184534 60321 184586 60373
rect 149398 60247 149450 60299
rect 184342 60247 184394 60299
rect 646006 59063 646058 59115
rect 652246 59063 652298 59115
rect 149398 58989 149450 59041
rect 184342 58989 184394 59041
rect 149398 57509 149450 57561
rect 184342 57509 184394 57561
rect 149398 56177 149450 56229
rect 184438 56177 184490 56229
rect 149494 56103 149546 56155
rect 184342 56103 184394 56155
rect 149686 54623 149738 54675
rect 184342 54623 184394 54675
rect 149398 53217 149450 53269
rect 184342 53217 184394 53269
rect 175606 53143 175658 53195
rect 668278 53143 668330 53195
rect 633622 48999 633674 49051
rect 640726 48999 640778 49051
rect 480982 48111 481034 48163
rect 527926 48111 527978 48163
rect 460342 48037 460394 48089
rect 510358 48037 510410 48089
rect 417526 47963 417578 48015
rect 492982 47963 493034 48015
rect 311062 47889 311114 47941
rect 371926 47889 371978 47941
rect 405526 47889 405578 47941
rect 441334 47889 441386 47941
rect 472246 47889 472298 47941
rect 562486 47889 562538 47941
rect 302902 47815 302954 47867
rect 506806 47815 506858 47867
rect 320182 47741 320234 47793
rect 529270 47741 529322 47793
rect 233686 47667 233738 47719
rect 475510 47667 475562 47719
rect 268534 47593 268586 47645
rect 520630 47593 520682 47645
rect 250966 47519 251018 47571
rect 521206 47519 521258 47571
rect 418870 47445 418922 47497
rect 424054 47445 424106 47497
rect 145366 47075 145418 47127
rect 199126 47075 199178 47127
rect 331222 46557 331274 46609
rect 337462 46557 337514 46609
rect 464854 46409 464906 46461
rect 475702 46409 475754 46461
rect 539734 46187 539786 46239
rect 545206 46187 545258 46239
rect 207382 46113 207434 46165
rect 216406 46113 216458 46165
rect 402166 46113 402218 46165
rect 406774 46113 406826 46165
rect 506806 44855 506858 44907
rect 512182 44855 512234 44907
rect 175606 44140 175658 44192
rect 285814 43227 285866 43279
rect 518710 43227 518762 43279
rect 629014 43227 629066 43279
rect 633622 43227 633674 43279
rect 403510 43153 403562 43205
rect 418870 43153 418922 43205
rect 444886 43153 444938 43205
rect 458614 43153 458666 43205
rect 302902 42117 302954 42169
rect 311158 42117 311210 42169
rect 357718 42117 357770 42169
rect 307222 42043 307274 42095
rect 311062 42043 311114 42095
rect 335446 42043 335498 42095
rect 354838 42043 354890 42095
rect 362038 42043 362090 42095
rect 365974 42043 366026 42095
rect 402166 42043 402218 42095
rect 471670 42043 471722 42095
rect 480982 42043 481034 42095
rect 186262 41969 186314 42021
rect 187030 41969 187082 42021
rect 194326 41969 194378 42021
rect 629014 41969 629066 42021
rect 514006 41747 514058 41799
rect 514870 41747 514922 41799
rect 186262 41451 186314 41503
rect 207382 41451 207434 41503
rect 365878 37381 365930 37433
rect 403510 37455 403562 37507
rect 475510 37381 475562 37433
rect 514006 37381 514058 37433
rect 365974 37307 366026 37359
rect 389206 37307 389258 37359
rect 420790 34495 420842 34547
rect 444886 34495 444938 34547
rect 328342 31609 328394 31661
rect 335446 31609 335498 31661
<< metal2 >>
rect 81140 1002358 81196 1002367
rect 80578 1002316 81140 1002344
rect 80578 982979 80606 1002316
rect 184052 1002358 184108 1002367
rect 81140 1002293 81196 1002302
rect 181462 1002319 181514 1002325
rect 184052 1002293 184054 1002302
rect 181462 1002261 181514 1002267
rect 184106 1002293 184108 1002302
rect 482612 1002358 482668 1002367
rect 482612 1002293 482614 1002302
rect 184054 1002261 184106 1002267
rect 482666 1002293 482668 1002302
rect 483862 1002319 483914 1002325
rect 482614 1002261 482666 1002267
rect 483862 1002261 483914 1002267
rect 181474 1002196 181502 1002261
rect 181378 1002168 181502 1002196
rect 132404 997178 132460 997187
rect 132404 997113 132460 997122
rect 132418 982979 132446 997113
rect 181378 992261 181406 1002168
rect 394580 997770 394636 997779
rect 181366 992255 181418 992261
rect 181366 992197 181418 992203
rect 184246 992255 184298 992261
rect 184246 992197 184298 992203
rect 184258 982979 184286 992197
rect 233218 982979 233246 997742
rect 241172 997178 241228 997187
rect 241172 997113 241228 997122
rect 240886 983005 240938 983011
rect 80564 982970 80620 982979
rect 80564 982905 80620 982914
rect 132404 982970 132460 982979
rect 132404 982905 132460 982914
rect 184244 982970 184300 982979
rect 184244 982905 184300 982914
rect 233204 982970 233260 982979
rect 233204 982905 233260 982914
rect 240884 982970 240886 982979
rect 241186 982979 241214 997113
rect 241954 983011 241982 997742
rect 241942 983005 241994 983011
rect 240938 982970 240940 982979
rect 240884 982905 240940 982914
rect 241172 982970 241228 982979
rect 285058 982979 285086 997742
rect 290804 997178 290860 997187
rect 290804 997113 290860 997122
rect 290818 983275 290846 997113
rect 290804 983266 290860 983275
rect 290804 983201 290860 983210
rect 292162 983127 292190 997742
rect 394580 997705 394636 997714
rect 394594 991521 394622 997705
rect 394582 991515 394634 991521
rect 394582 991457 394634 991463
rect 397462 991515 397514 991521
rect 397462 991457 397514 991463
rect 397474 983275 397502 991457
rect 397460 983266 397516 983275
rect 397460 983201 397516 983210
rect 292148 983118 292204 983127
rect 292148 983053 292204 983062
rect 483874 982979 483902 1002261
rect 535700 997770 535756 997779
rect 535700 997705 535756 997714
rect 636500 997770 636556 997779
rect 636500 997705 636556 997714
rect 535714 992187 535742 997705
rect 535702 992181 535754 992187
rect 535702 992123 535754 992129
rect 538582 992181 538634 992187
rect 538582 992123 538634 992129
rect 538594 982979 538622 992123
rect 636514 983127 636542 997705
rect 636500 983118 636556 983127
rect 636500 983053 636556 983062
rect 656662 983005 656714 983011
rect 241942 982947 241994 982953
rect 285044 982970 285100 982979
rect 241172 982905 241228 982914
rect 285044 982905 285100 982914
rect 391604 982970 391660 982979
rect 391604 982905 391606 982914
rect 391658 982905 391660 982914
rect 394580 982970 394636 982979
rect 394580 982905 394636 982914
rect 483860 982970 483916 982979
rect 483860 982905 483916 982914
rect 538580 982970 538636 982979
rect 656662 982947 656714 982953
rect 538580 982905 538636 982914
rect 649462 982931 649514 982937
rect 391606 982873 391658 982879
rect 394594 982863 394622 982905
rect 649462 982873 649514 982879
rect 394582 982857 394634 982863
rect 394582 982799 394634 982805
rect 649474 982049 649502 982873
rect 649462 982043 649514 982049
rect 649462 981985 649514 981991
rect 652246 982043 652298 982049
rect 652246 981985 652298 981991
rect 652258 979237 652286 981985
rect 656674 979311 656702 982947
rect 656662 979305 656714 979311
rect 656662 979247 656714 979253
rect 679702 979305 679754 979311
rect 679702 979247 679754 979253
rect 652246 979231 652298 979237
rect 652246 979173 652298 979179
rect 677590 979231 677642 979237
rect 677590 979173 677642 979179
rect 677494 967687 677546 967693
rect 677494 967629 677546 967635
rect 40148 959290 40204 959299
rect 40148 959225 40204 959234
rect 40162 959109 40190 959225
rect 60020 959142 60076 959151
rect 40150 959103 40202 959109
rect 60020 959077 60022 959086
rect 40150 959045 40202 959051
rect 60074 959077 60076 959086
rect 653780 959142 653836 959151
rect 653780 959077 653836 959086
rect 60022 959045 60074 959051
rect 653794 950377 653822 959077
rect 677506 957500 677534 967629
rect 677602 967402 677630 979173
rect 679714 967693 679742 979247
rect 679702 967687 679754 967693
rect 679702 967629 679754 967635
rect 677506 957472 677616 957500
rect 676820 950410 676876 950419
rect 653782 950371 653834 950377
rect 676820 950345 676822 950354
rect 653782 950313 653834 950319
rect 676874 950345 676876 950354
rect 676822 950313 676874 950319
rect 676148 894170 676204 894179
rect 676148 894105 676204 894114
rect 676052 893430 676108 893439
rect 676052 893365 676108 893374
rect 655414 893021 655466 893027
rect 655414 892963 655466 892969
rect 655222 892947 655274 892953
rect 655222 892889 655274 892895
rect 655126 892873 655178 892879
rect 655126 892815 655178 892821
rect 649462 881477 649514 881483
rect 649462 881419 649514 881425
rect 649474 861134 649502 881419
rect 654166 872671 654218 872677
rect 654166 872613 654218 872619
rect 653782 864013 653834 864019
rect 654178 863987 654206 872613
rect 655138 866503 655166 892815
rect 655234 868871 655262 892889
rect 655318 881403 655370 881409
rect 655318 881345 655370 881351
rect 655220 868862 655276 868871
rect 655220 868797 655276 868806
rect 655124 866494 655180 866503
rect 655124 866429 655180 866438
rect 655330 865319 655358 881345
rect 655426 867687 655454 892963
rect 676066 892879 676094 893365
rect 676162 893027 676190 894105
rect 676244 893578 676300 893587
rect 676244 893513 676300 893522
rect 676150 893021 676202 893027
rect 676150 892963 676202 892969
rect 676258 892953 676286 893513
rect 676246 892947 676298 892953
rect 676246 892889 676298 892895
rect 676054 892873 676106 892879
rect 676054 892815 676106 892821
rect 676052 892468 676108 892477
rect 673366 892429 673418 892435
rect 676052 892403 676054 892412
rect 673366 892371 673418 892377
rect 676106 892403 676108 892412
rect 676054 892371 676106 892377
rect 670966 891467 671018 891473
rect 670966 891409 671018 891415
rect 670870 890431 670922 890437
rect 670870 890373 670922 890379
rect 655412 867678 655468 867687
rect 655412 867613 655468 867622
rect 655316 865310 655372 865319
rect 655316 865245 655372 865254
rect 653782 863955 653834 863961
rect 654164 863978 654220 863987
rect 653794 862951 653822 863955
rect 654164 863913 654220 863922
rect 653780 862942 653836 862951
rect 653780 862877 653836 862886
rect 649378 861106 649502 861134
rect 41782 817985 41834 817991
rect 41780 817950 41782 817959
rect 47446 817985 47498 817991
rect 41834 817950 41836 817959
rect 47446 817927 47498 817933
rect 41780 817885 41836 817894
rect 41780 817358 41836 817367
rect 41780 817293 41782 817302
rect 41834 817293 41836 817302
rect 44854 817319 44906 817325
rect 41782 817261 41834 817267
rect 44854 817261 44906 817267
rect 41588 816618 41644 816627
rect 41588 816553 41590 816562
rect 41642 816553 41644 816562
rect 41590 816521 41642 816527
rect 41780 815878 41836 815887
rect 41780 815813 41782 815822
rect 41834 815813 41836 815822
rect 43222 815839 43274 815845
rect 41782 815781 41834 815787
rect 43222 815781 43274 815787
rect 41780 814916 41836 814925
rect 41780 814851 41782 814860
rect 41834 814851 41836 814860
rect 41782 814819 41834 814825
rect 41588 813658 41644 813667
rect 41588 813593 41590 813602
rect 41642 813593 41644 813602
rect 41590 813561 41642 813567
rect 41588 813214 41644 813223
rect 41588 813149 41644 813158
rect 40244 812474 40300 812483
rect 41602 812441 41630 813149
rect 42548 812918 42604 812927
rect 42548 812853 42604 812862
rect 40244 812409 40300 812418
rect 41590 812435 41642 812441
rect 28820 805666 28876 805675
rect 28820 805601 28876 805610
rect 28834 805231 28862 805601
rect 28820 805222 28876 805231
rect 28820 805157 28876 805166
rect 40258 802123 40286 812409
rect 41590 812377 41642 812383
rect 41588 811734 41644 811743
rect 41588 811669 41644 811678
rect 41602 809925 41630 811669
rect 41972 811364 42028 811373
rect 41972 811299 42028 811308
rect 41876 810846 41932 810855
rect 41876 810781 41932 810790
rect 41590 809919 41642 809925
rect 41590 809861 41642 809867
rect 41780 809884 41836 809893
rect 41780 809819 41782 809828
rect 41834 809819 41836 809828
rect 41782 809787 41834 809793
rect 41780 808922 41836 808931
rect 41780 808857 41836 808866
rect 41794 808667 41822 808857
rect 41782 808661 41834 808667
rect 41782 808603 41834 808609
rect 41684 808182 41740 808191
rect 41684 808117 41740 808126
rect 41588 806702 41644 806711
rect 41588 806637 41590 806646
rect 41642 806637 41644 806646
rect 41590 806605 41642 806611
rect 41588 806110 41644 806119
rect 41588 806045 41644 806054
rect 41602 805231 41630 806045
rect 41588 805222 41644 805231
rect 41588 805157 41590 805166
rect 41642 805157 41644 805166
rect 41590 805125 41642 805131
rect 40244 802114 40300 802123
rect 40244 802049 40300 802058
rect 41698 800495 41726 808117
rect 41780 807442 41836 807451
rect 41780 807377 41782 807386
rect 41834 807377 41836 807386
rect 41782 807345 41834 807351
rect 41684 800486 41740 800495
rect 41684 800421 41740 800430
rect 41890 800231 41918 810781
rect 41986 800347 42014 811299
rect 42068 809366 42124 809375
rect 42068 809301 42124 809310
rect 42082 800495 42110 809301
rect 42164 807886 42220 807895
rect 42164 807821 42220 807830
rect 42068 800486 42124 800495
rect 42068 800421 42124 800430
rect 41972 800338 42028 800347
rect 41972 800273 42028 800282
rect 42178 800231 42206 807821
rect 41878 800225 41930 800231
rect 41878 800167 41930 800173
rect 42166 800225 42218 800231
rect 42166 800167 42218 800173
rect 41878 800003 41930 800009
rect 41878 799945 41930 799951
rect 41890 799422 41918 799945
rect 42562 798159 42590 812853
rect 42934 812435 42986 812441
rect 42934 812377 42986 812383
rect 42838 809919 42890 809925
rect 42838 809861 42890 809867
rect 42742 809845 42794 809851
rect 42742 809787 42794 809793
rect 42646 807403 42698 807409
rect 42646 807345 42698 807351
rect 42166 798153 42218 798159
rect 42166 798095 42218 798101
rect 42550 798153 42602 798159
rect 42550 798095 42602 798101
rect 42178 797605 42206 798095
rect 42658 797937 42686 807345
rect 42754 800939 42782 809787
rect 42740 800930 42796 800939
rect 42740 800865 42796 800874
rect 42850 800823 42878 809861
rect 42838 800817 42890 800823
rect 42838 800759 42890 800765
rect 42742 800743 42794 800749
rect 42742 800685 42794 800691
rect 42646 797931 42698 797937
rect 42646 797873 42698 797879
rect 42754 797345 42782 800685
rect 42838 800669 42890 800675
rect 42838 800611 42890 800617
rect 42070 797339 42122 797345
rect 42070 797281 42122 797287
rect 42742 797339 42794 797345
rect 42742 797281 42794 797287
rect 42082 796980 42110 797281
rect 42742 796895 42794 796901
rect 42742 796837 42794 796843
rect 42166 796303 42218 796309
rect 42166 796245 42218 796251
rect 42178 795765 42206 796245
rect 42070 795637 42122 795643
rect 42070 795579 42122 795585
rect 42082 795130 42110 795579
rect 42166 794823 42218 794829
rect 42166 794765 42218 794771
rect 42178 794569 42206 794765
rect 41780 794270 41836 794279
rect 41780 794205 41836 794214
rect 41794 793946 41822 794205
rect 42754 793645 42782 796837
rect 42850 795643 42878 800611
rect 42838 795637 42890 795643
rect 42838 795579 42890 795585
rect 42166 793639 42218 793645
rect 42166 793581 42218 793587
rect 42742 793639 42794 793645
rect 42742 793581 42794 793587
rect 42178 793280 42206 793581
rect 42740 793530 42796 793539
rect 42740 793465 42796 793474
rect 41972 792938 42028 792947
rect 41972 792873 42028 792882
rect 41986 792729 42014 792873
rect 42166 790679 42218 790685
rect 42166 790621 42218 790627
rect 42178 790246 42206 790621
rect 42164 790126 42220 790135
rect 42164 790061 42220 790070
rect 42178 789580 42206 790061
rect 42754 789501 42782 793465
rect 42946 792165 42974 812377
rect 43126 808661 43178 808667
rect 43126 808603 43178 808609
rect 43030 806663 43082 806669
rect 43030 806605 43082 806611
rect 43042 794829 43070 806605
rect 43138 796309 43166 808603
rect 43234 796309 43262 815781
rect 44662 814877 44714 814883
rect 44662 814819 44714 814825
rect 44566 805183 44618 805189
rect 44566 805125 44618 805131
rect 43510 800817 43562 800823
rect 43510 800759 43562 800765
rect 43318 800225 43370 800231
rect 43318 800167 43370 800173
rect 43126 796303 43178 796309
rect 43126 796245 43178 796251
rect 43222 796303 43274 796309
rect 43222 796245 43274 796251
rect 43330 796180 43358 800167
rect 43138 796152 43358 796180
rect 43030 794823 43082 794829
rect 43030 794765 43082 794771
rect 43030 794675 43082 794681
rect 43030 794617 43082 794623
rect 42934 792159 42986 792165
rect 42934 792101 42986 792107
rect 42166 789495 42218 789501
rect 42166 789437 42218 789443
rect 42742 789495 42794 789501
rect 42742 789437 42794 789443
rect 42178 788957 42206 789437
rect 42836 789386 42892 789395
rect 42836 789321 42892 789330
rect 42740 789238 42796 789247
rect 42740 789173 42796 789182
rect 42166 788755 42218 788761
rect 42166 788697 42218 788703
rect 42178 788396 42206 788697
rect 42166 786905 42218 786911
rect 42166 786847 42218 786853
rect 42178 786546 42206 786847
rect 42754 786467 42782 789173
rect 42166 786461 42218 786467
rect 42166 786403 42218 786409
rect 42742 786461 42794 786467
rect 42742 786403 42794 786409
rect 42178 785921 42206 786403
rect 42850 785653 42878 789321
rect 42934 789199 42986 789205
rect 42934 789141 42986 789147
rect 42070 785647 42122 785653
rect 42070 785589 42122 785595
rect 42838 785647 42890 785653
rect 42838 785589 42890 785595
rect 42082 785288 42110 785589
rect 42946 785061 42974 789141
rect 43042 788761 43070 794617
rect 43138 790685 43166 796152
rect 43222 796081 43274 796087
rect 43222 796023 43274 796029
rect 43234 790852 43262 796023
rect 43522 794681 43550 800759
rect 43510 794675 43562 794681
rect 43510 794617 43562 794623
rect 43510 792159 43562 792165
rect 43510 792101 43562 792107
rect 43234 790824 43454 790852
rect 43126 790679 43178 790685
rect 43126 790621 43178 790627
rect 43126 790531 43178 790537
rect 43126 790473 43178 790479
rect 43030 788755 43082 788761
rect 43030 788697 43082 788703
rect 43138 786911 43166 790473
rect 43126 786905 43178 786911
rect 43126 786847 43178 786853
rect 42166 785055 42218 785061
rect 42166 784997 42218 785003
rect 42934 785055 42986 785061
rect 42934 784997 42986 785003
rect 42178 784725 42206 784997
rect 41780 774734 41836 774743
rect 41780 774669 41782 774678
rect 41834 774669 41836 774678
rect 41782 774637 41834 774643
rect 41588 773994 41644 774003
rect 41588 773929 41590 773938
rect 41642 773929 41644 773938
rect 41590 773897 41642 773903
rect 41588 773402 41644 773411
rect 41588 773337 41590 773346
rect 41642 773337 41644 773346
rect 41590 773305 41642 773311
rect 43426 773295 43454 790824
rect 43522 790537 43550 792101
rect 43510 790531 43562 790537
rect 43510 790473 43562 790479
rect 41782 773289 41834 773295
rect 41780 773254 41782 773263
rect 43414 773289 43466 773295
rect 41834 773254 41836 773263
rect 43414 773231 43466 773237
rect 41780 773189 41836 773198
rect 41588 772958 41644 772967
rect 41588 772893 41644 772902
rect 41602 771889 41630 772893
rect 41780 772662 41836 772671
rect 41780 772597 41782 772606
rect 41834 772597 41836 772606
rect 43318 772623 43370 772629
rect 41782 772565 41834 772571
rect 43318 772565 43370 772571
rect 42742 771957 42794 771963
rect 42740 771922 42742 771931
rect 42794 771922 42796 771931
rect 41590 771883 41642 771889
rect 42740 771857 42796 771866
rect 41590 771825 41642 771831
rect 41602 770895 41630 771825
rect 41588 770886 41644 770895
rect 41588 770821 41644 770830
rect 41396 769998 41452 770007
rect 41396 769933 41452 769942
rect 40244 768962 40300 768971
rect 40244 768897 40300 768906
rect 28820 762450 28876 762459
rect 28820 762385 28876 762394
rect 28834 762015 28862 762385
rect 28820 762006 28876 762015
rect 28820 761941 28876 761950
rect 40258 759943 40286 768897
rect 40244 759934 40300 759943
rect 40244 759869 40300 759878
rect 41410 757385 41438 769933
rect 41972 769702 42028 769711
rect 41972 769637 42028 769646
rect 41684 768518 41740 768527
rect 41684 768453 41740 768462
rect 41492 766446 41548 766455
rect 41492 766381 41548 766390
rect 41398 757379 41450 757385
rect 41398 757321 41450 757327
rect 41506 757311 41534 766381
rect 41588 763486 41644 763495
rect 41588 763421 41590 763430
rect 41642 763421 41644 763430
rect 41590 763389 41642 763395
rect 41698 757427 41726 768453
rect 41780 768222 41836 768231
rect 41780 768157 41782 768166
rect 41834 768157 41836 768166
rect 41782 768125 41834 768131
rect 41876 767630 41932 767639
rect 41876 767565 41932 767574
rect 41780 765188 41836 765197
rect 41780 765123 41782 765132
rect 41834 765123 41836 765132
rect 41782 765091 41834 765097
rect 41780 764226 41836 764235
rect 41780 764161 41782 764170
rect 41834 764161 41836 764170
rect 41782 764129 41834 764135
rect 41780 762154 41836 762163
rect 41780 762089 41782 762098
rect 41834 762089 41836 762098
rect 41782 762057 41834 762063
rect 41684 757418 41740 757427
rect 41684 757353 41740 757362
rect 41494 757305 41546 757311
rect 41494 757247 41546 757253
rect 41890 757015 41918 767565
rect 41986 757131 42014 769637
rect 42838 768183 42890 768189
rect 42838 768125 42890 768131
rect 42068 766150 42124 766159
rect 42068 766085 42124 766094
rect 42082 757279 42110 766085
rect 42164 765706 42220 765715
rect 42164 765641 42220 765650
rect 42178 757404 42206 765641
rect 42850 757871 42878 768125
rect 42934 765149 42986 765155
rect 42934 765091 42986 765097
rect 42836 757862 42892 757871
rect 42836 757797 42892 757806
rect 42946 757681 42974 765091
rect 43030 764187 43082 764193
rect 43030 764129 43082 764135
rect 42934 757675 42986 757681
rect 42934 757617 42986 757623
rect 42934 757527 42986 757533
rect 42934 757469 42986 757475
rect 42178 757376 42398 757404
rect 42068 757270 42124 757279
rect 42068 757205 42124 757214
rect 41972 757122 42028 757131
rect 41972 757057 42028 757066
rect 41878 757009 41930 757015
rect 41878 756951 41930 756957
rect 41878 756787 41930 756793
rect 41878 756729 41930 756735
rect 41890 756245 41918 756729
rect 41972 754902 42028 754911
rect 41972 754837 42028 754846
rect 41986 754430 42014 754837
rect 42166 754271 42218 754277
rect 42166 754213 42218 754219
rect 42178 753764 42206 754213
rect 42370 753093 42398 757376
rect 42946 754277 42974 757469
rect 42934 754271 42986 754277
rect 42934 754213 42986 754219
rect 42070 753087 42122 753093
rect 42070 753029 42122 753035
rect 42358 753087 42410 753093
rect 42358 753029 42410 753035
rect 42082 752580 42110 753029
rect 43042 752945 43070 764129
rect 43126 763447 43178 763453
rect 43126 763389 43178 763395
rect 42358 752939 42410 752945
rect 42358 752881 42410 752887
rect 43030 752939 43082 752945
rect 43030 752881 43082 752887
rect 42082 751835 42110 751914
rect 42070 751829 42122 751835
rect 42070 751771 42122 751777
rect 42070 751533 42122 751539
rect 42070 751475 42122 751481
rect 42082 751396 42110 751475
rect 42070 751163 42122 751169
rect 42070 751105 42122 751111
rect 42082 750730 42110 751105
rect 42370 750651 42398 752881
rect 43138 752816 43166 763389
rect 43222 757675 43274 757681
rect 43222 757617 43274 757623
rect 42946 752788 43166 752816
rect 42946 751539 42974 752788
rect 43234 752668 43262 757617
rect 43138 752640 43262 752668
rect 42934 751533 42986 751539
rect 42934 751475 42986 751481
rect 42932 751350 42988 751359
rect 42932 751285 42988 751294
rect 42166 750645 42218 750651
rect 42166 750587 42218 750593
rect 42358 750645 42410 750651
rect 42358 750587 42410 750593
rect 42178 750064 42206 750587
rect 42946 749837 42974 751285
rect 43138 751169 43166 752640
rect 43222 751829 43274 751835
rect 43222 751771 43274 751777
rect 43126 751163 43178 751169
rect 43126 751105 43178 751111
rect 43126 751015 43178 751021
rect 43126 750957 43178 750963
rect 42070 749831 42122 749837
rect 42070 749773 42122 749779
rect 42934 749831 42986 749837
rect 42934 749773 42986 749779
rect 42082 749546 42110 749773
rect 42934 749683 42986 749689
rect 42934 749625 42986 749631
rect 42452 747798 42508 747807
rect 42452 747733 42508 747742
rect 41780 747502 41836 747511
rect 41780 747437 41836 747446
rect 41794 747030 41822 747437
rect 42164 746910 42220 746919
rect 42164 746845 42220 746854
rect 42178 746401 42206 746845
rect 42356 746614 42412 746623
rect 42356 746549 42412 746558
rect 42070 746131 42122 746137
rect 42070 746073 42122 746079
rect 42082 745772 42110 746073
rect 42166 745539 42218 745545
rect 42166 745481 42218 745487
rect 42178 745180 42206 745481
rect 42370 745416 42398 746549
rect 42466 745545 42494 747733
rect 42946 747340 42974 749625
rect 42946 747312 43070 747340
rect 42932 747206 42988 747215
rect 42932 747141 42988 747150
rect 42454 745539 42506 745545
rect 42454 745481 42506 745487
rect 42370 745388 42494 745416
rect 42166 743615 42218 743621
rect 42166 743557 42218 743563
rect 42178 743365 42206 743557
rect 42070 743245 42122 743251
rect 42070 743187 42122 743193
rect 42082 742738 42110 743187
rect 42466 742659 42494 745388
rect 42946 743251 42974 747141
rect 43042 743621 43070 747312
rect 43138 746137 43166 750957
rect 43126 746131 43178 746137
rect 43126 746073 43178 746079
rect 43126 745983 43178 745989
rect 43126 745925 43178 745931
rect 43030 743615 43082 743621
rect 43030 743557 43082 743563
rect 42934 743245 42986 743251
rect 42934 743187 42986 743193
rect 42166 742653 42218 742659
rect 42166 742595 42218 742601
rect 42454 742653 42506 742659
rect 42454 742595 42506 742601
rect 42178 742072 42206 742595
rect 43138 741993 43166 745925
rect 43234 745323 43262 751771
rect 43222 745317 43274 745323
rect 43222 745259 43274 745265
rect 42166 741987 42218 741993
rect 42166 741929 42218 741935
rect 43126 741987 43178 741993
rect 43126 741929 43178 741935
rect 42178 741525 42206 741929
rect 41780 731518 41836 731527
rect 41780 731453 41782 731462
rect 41834 731453 41836 731462
rect 41782 731421 41834 731427
rect 41588 730778 41644 730787
rect 41588 730713 41590 730722
rect 41642 730713 41644 730722
rect 41590 730681 41642 730687
rect 41780 730408 41836 730417
rect 41780 730343 41782 730352
rect 41834 730343 41836 730352
rect 41782 730311 41834 730317
rect 43330 730227 43358 772565
rect 43606 757379 43658 757385
rect 43606 757321 43658 757327
rect 43510 757305 43562 757311
rect 43510 757247 43562 757253
rect 43522 751021 43550 757247
rect 43510 751015 43562 751021
rect 43510 750957 43562 750963
rect 43618 749689 43646 757321
rect 43606 749683 43658 749689
rect 43606 749625 43658 749631
rect 41590 730221 41642 730227
rect 41588 730186 41590 730195
rect 43318 730221 43370 730227
rect 41642 730186 41644 730195
rect 43318 730163 43370 730169
rect 41588 730121 41644 730130
rect 41396 729298 41452 729307
rect 41396 729233 41452 729242
rect 41588 729298 41644 729307
rect 41588 729233 41590 729242
rect 40438 728741 40490 728747
rect 40436 728706 40438 728715
rect 40490 728706 40492 728715
rect 41410 728673 41438 729233
rect 41642 729233 41644 729242
rect 43894 729259 43946 729265
rect 41590 729201 41642 729207
rect 43894 729201 43946 729207
rect 41780 728854 41836 728863
rect 41780 728789 41782 728798
rect 41834 728789 41836 728798
rect 43798 728815 43850 728821
rect 41782 728757 41834 728763
rect 43798 728757 43850 728763
rect 40436 728641 40492 728650
rect 41398 728667 41450 728673
rect 41398 728609 41450 728615
rect 41780 727966 41836 727975
rect 41780 727901 41782 727910
rect 41834 727901 41836 727910
rect 43702 727927 43754 727933
rect 41782 727869 41834 727875
rect 43702 727869 43754 727875
rect 41492 726782 41548 726791
rect 41492 726717 41548 726726
rect 34388 725746 34444 725755
rect 34388 725681 34444 725690
rect 28820 719234 28876 719243
rect 28820 719169 28876 719178
rect 28834 718799 28862 719169
rect 28820 718790 28876 718799
rect 28820 718725 28876 718734
rect 34402 716727 34430 725681
rect 34484 723822 34540 723831
rect 34484 723757 34540 723766
rect 34388 716718 34444 716727
rect 34388 716653 34444 716662
rect 34498 716135 34526 723757
rect 34484 716126 34540 716135
rect 34484 716061 34540 716070
rect 41506 714211 41534 726717
rect 42068 726486 42124 726495
rect 42068 726421 42124 726430
rect 41972 725524 42028 725533
rect 41972 725459 42028 725468
rect 41780 724414 41836 724423
rect 41780 724349 41836 724358
rect 41684 722342 41740 722351
rect 41684 722277 41740 722286
rect 41588 721750 41644 721759
rect 41588 721685 41644 721694
rect 41602 720459 41630 721685
rect 41590 720453 41642 720459
rect 41590 720395 41642 720401
rect 41588 720270 41644 720279
rect 41588 720205 41590 720214
rect 41642 720205 41644 720214
rect 41590 720173 41642 720179
rect 41588 718790 41644 718799
rect 41588 718725 41590 718734
rect 41642 718725 41644 718734
rect 41590 718693 41642 718699
rect 41492 714202 41548 714211
rect 41492 714137 41548 714146
rect 41698 714095 41726 722277
rect 41686 714089 41738 714095
rect 41686 714031 41738 714037
rect 41794 713873 41822 724349
rect 41878 722969 41930 722975
rect 41876 722934 41878 722943
rect 41930 722934 41932 722943
rect 41876 722869 41932 722878
rect 41986 714063 42014 725459
rect 41972 714054 42028 714063
rect 41972 713989 42028 713998
rect 42082 713915 42110 726421
rect 42164 725006 42220 725015
rect 42164 724941 42220 724950
rect 42178 713947 42206 724941
rect 42452 723526 42508 723535
rect 42452 723461 42508 723470
rect 42166 713941 42218 713947
rect 42068 713906 42124 713915
rect 41782 713867 41834 713873
rect 42166 713883 42218 713889
rect 42068 713841 42124 713850
rect 41782 713809 41834 713815
rect 41782 713571 41834 713577
rect 41782 713513 41834 713519
rect 41794 713064 41822 713513
rect 42466 712287 42494 723461
rect 42934 722969 42986 722975
rect 42934 722911 42986 722917
rect 42452 712278 42508 712287
rect 42452 712213 42508 712222
rect 42454 712017 42506 712023
rect 42454 711959 42506 711965
rect 42068 711686 42124 711695
rect 42068 711621 42124 711630
rect 42082 711214 42110 711621
rect 42466 710913 42494 711959
rect 42946 711547 42974 722911
rect 43030 720453 43082 720459
rect 43030 720395 43082 720401
rect 43042 711695 43070 720395
rect 43126 720231 43178 720237
rect 43126 720173 43178 720179
rect 43028 711686 43084 711695
rect 43028 711621 43084 711630
rect 43030 711573 43082 711579
rect 42932 711538 42988 711547
rect 43030 711515 43082 711521
rect 42932 711473 42988 711482
rect 42932 711242 42988 711251
rect 43042 711209 43070 711515
rect 42932 711177 42988 711186
rect 43030 711203 43082 711209
rect 42166 710907 42218 710913
rect 42166 710849 42218 710855
rect 42454 710907 42506 710913
rect 42454 710849 42506 710855
rect 42178 710548 42206 710849
rect 42166 709945 42218 709951
rect 42166 709887 42218 709893
rect 42178 709364 42206 709887
rect 42452 708874 42508 708883
rect 42452 708809 42508 708818
rect 42082 708545 42110 708698
rect 42070 708539 42122 708545
rect 42070 708481 42122 708487
rect 42070 708391 42122 708397
rect 42070 708333 42122 708339
rect 42082 708180 42110 708333
rect 42166 708095 42218 708101
rect 42166 708037 42218 708043
rect 42178 707514 42206 708037
rect 41780 707394 41836 707403
rect 41780 707329 41836 707338
rect 41794 706881 41822 707329
rect 42166 706615 42218 706621
rect 42166 706557 42218 706563
rect 42178 706330 42206 706557
rect 42466 704993 42494 708809
rect 42946 708101 42974 711177
rect 43030 711145 43082 711151
rect 43028 711094 43084 711103
rect 43028 711029 43084 711038
rect 42934 708095 42986 708101
rect 42934 708037 42986 708043
rect 42932 707986 42988 707995
rect 42932 707921 42988 707930
rect 42946 706473 42974 707921
rect 42934 706467 42986 706473
rect 42934 706409 42986 706415
rect 42932 705174 42988 705183
rect 42932 705109 42988 705118
rect 42454 704987 42506 704993
rect 42454 704929 42506 704935
rect 42356 704878 42412 704887
rect 42356 704813 42412 704822
rect 42166 704321 42218 704327
rect 42166 704263 42218 704269
rect 42178 703845 42206 704263
rect 42070 703729 42122 703735
rect 42070 703671 42122 703677
rect 42082 703222 42110 703671
rect 42370 702699 42398 704813
rect 42166 702693 42218 702699
rect 42166 702635 42218 702641
rect 42358 702693 42410 702699
rect 42358 702635 42410 702641
rect 42178 702556 42206 702635
rect 42166 702323 42218 702329
rect 42166 702265 42218 702271
rect 42178 702005 42206 702265
rect 42070 700547 42122 700553
rect 42070 700489 42122 700495
rect 42082 700188 42110 700489
rect 41780 699994 41836 700003
rect 41780 699929 41836 699938
rect 41794 699522 41822 699929
rect 42946 699443 42974 705109
rect 43042 703735 43070 711029
rect 43138 708397 43166 720173
rect 43222 714311 43274 714317
rect 43222 714253 43274 714259
rect 43234 712023 43262 714253
rect 43510 714089 43562 714095
rect 43510 714031 43562 714037
rect 43414 713941 43466 713947
rect 43414 713883 43466 713889
rect 43222 712017 43274 712023
rect 43222 711959 43274 711965
rect 43222 711869 43274 711875
rect 43222 711811 43274 711817
rect 43126 708391 43178 708397
rect 43126 708333 43178 708339
rect 43126 708243 43178 708249
rect 43126 708185 43178 708191
rect 43138 706621 43166 708185
rect 43126 706615 43178 706621
rect 43126 706557 43178 706563
rect 43126 706467 43178 706473
rect 43126 706409 43178 706415
rect 43030 703729 43082 703735
rect 43030 703671 43082 703677
rect 43028 703546 43084 703555
rect 43028 703481 43084 703490
rect 43042 700553 43070 703481
rect 43138 702329 43166 706409
rect 43126 702323 43178 702329
rect 43126 702265 43178 702271
rect 43030 700547 43082 700553
rect 43030 700489 43082 700495
rect 42166 699437 42218 699443
rect 42166 699379 42218 699385
rect 42934 699437 42986 699443
rect 42934 699379 42986 699385
rect 42178 698856 42206 699379
rect 42070 698771 42122 698777
rect 42070 698713 42122 698719
rect 42082 698338 42110 698713
rect 41780 688302 41836 688311
rect 41780 688237 41782 688246
rect 41834 688237 41836 688246
rect 41782 688205 41834 688211
rect 41588 687562 41644 687571
rect 41588 687497 41590 687506
rect 41642 687497 41644 687506
rect 41590 687465 41642 687471
rect 41780 687266 41836 687275
rect 41780 687201 41782 687210
rect 41834 687201 41836 687210
rect 41782 687169 41834 687175
rect 41590 687005 41642 687011
rect 41588 686970 41590 686979
rect 41642 686970 41644 686979
rect 41588 686905 41644 686914
rect 41588 686082 41644 686091
rect 41588 686017 41590 686026
rect 41642 686017 41644 686026
rect 41590 685985 41642 685991
rect 43234 685383 43262 711811
rect 43426 711579 43454 713883
rect 43414 711573 43466 711579
rect 43414 711515 43466 711521
rect 43414 711425 43466 711431
rect 43316 711390 43372 711399
rect 43414 711367 43466 711373
rect 43316 711325 43372 711334
rect 41782 685377 41834 685383
rect 41780 685342 41782 685351
rect 43222 685377 43274 685383
rect 41834 685342 41836 685351
rect 43222 685319 43274 685325
rect 41780 685277 41836 685286
rect 43330 684199 43358 711325
rect 43426 687011 43454 711367
rect 43522 709951 43550 714031
rect 43714 711399 43742 727869
rect 43810 711875 43838 728757
rect 43798 711869 43850 711875
rect 43798 711811 43850 711817
rect 43906 711431 43934 729201
rect 43894 711425 43946 711431
rect 43700 711390 43756 711399
rect 43894 711367 43946 711373
rect 43700 711325 43756 711334
rect 43606 711129 43658 711135
rect 43606 711071 43658 711077
rect 43510 709945 43562 709951
rect 43510 709887 43562 709893
rect 43510 708539 43562 708545
rect 43510 708481 43562 708487
rect 43522 702699 43550 708481
rect 43618 708249 43646 711071
rect 43606 708243 43658 708249
rect 43606 708185 43658 708191
rect 43510 702693 43562 702699
rect 43510 702635 43562 702641
rect 43414 687005 43466 687011
rect 43414 686947 43466 686953
rect 43510 686043 43562 686049
rect 43510 685985 43562 685991
rect 41782 684193 41834 684199
rect 41780 684158 41782 684167
rect 43318 684193 43370 684199
rect 41834 684158 41836 684167
rect 43318 684135 43370 684141
rect 41780 684093 41836 684102
rect 41972 683862 42028 683871
rect 41972 683797 42028 683806
rect 41780 683270 41836 683279
rect 41780 683205 41836 683214
rect 41794 683089 41822 683205
rect 41782 683083 41834 683089
rect 41782 683025 41834 683031
rect 34388 682530 34444 682539
rect 34388 682465 34444 682474
rect 28820 676018 28876 676027
rect 28820 675953 28876 675962
rect 28834 675583 28862 675953
rect 28820 675574 28876 675583
rect 28820 675509 28876 675518
rect 34402 672475 34430 682465
rect 37364 682086 37420 682095
rect 37364 682021 37420 682030
rect 34484 679570 34540 679579
rect 34484 679505 34540 679514
rect 34498 672507 34526 679505
rect 34486 672501 34538 672507
rect 34388 672466 34444 672475
rect 34486 672443 34538 672449
rect 34388 672401 34444 672410
rect 37378 671323 37406 682021
rect 41876 681790 41932 681799
rect 41876 681725 41932 681734
rect 41780 681198 41836 681207
rect 41780 681133 41836 681142
rect 39764 680606 39820 680615
rect 39764 680541 39820 680550
rect 37366 671317 37418 671323
rect 37366 671259 37418 671265
rect 39778 671143 39806 680541
rect 39860 680014 39916 680023
rect 39860 679949 39916 679958
rect 39874 671249 39902 679949
rect 41588 679126 41644 679135
rect 41588 679061 41644 679070
rect 41602 677317 41630 679061
rect 41684 677646 41740 677655
rect 41684 677581 41740 677590
rect 41590 677311 41642 677317
rect 41590 677253 41642 677259
rect 41588 677054 41644 677063
rect 41588 676989 41590 676998
rect 41642 676989 41644 676998
rect 41590 676957 41642 676963
rect 41588 675574 41644 675583
rect 41588 675509 41590 675518
rect 41642 675509 41644 675518
rect 41590 675477 41642 675483
rect 40342 672501 40394 672507
rect 40342 672443 40394 672449
rect 39862 671243 39914 671249
rect 39862 671185 39914 671191
rect 40354 671175 40382 672443
rect 40342 671169 40394 671175
rect 39764 671134 39820 671143
rect 40342 671111 40394 671117
rect 39764 671069 39820 671078
rect 41698 670879 41726 677581
rect 41686 670873 41738 670879
rect 41686 670815 41738 670821
rect 41794 670657 41822 681133
rect 41890 670657 41918 681725
rect 41986 670699 42014 683797
rect 42934 683083 42986 683089
rect 42934 683025 42986 683031
rect 42068 678830 42124 678839
rect 42068 678765 42124 678774
rect 42082 670731 42110 678765
rect 42260 678238 42316 678247
rect 42260 678173 42316 678182
rect 42274 670805 42302 678173
rect 42742 671095 42794 671101
rect 42742 671037 42794 671043
rect 42262 670799 42314 670805
rect 42262 670741 42314 670747
rect 42070 670725 42122 670731
rect 41972 670690 42028 670699
rect 41782 670651 41834 670657
rect 41782 670593 41834 670599
rect 41878 670651 41930 670657
rect 42070 670667 42122 670673
rect 41972 670625 42028 670634
rect 41878 670593 41930 670599
rect 41782 670355 41834 670361
rect 41782 670297 41834 670303
rect 41794 669848 41822 670297
rect 42166 668579 42218 668585
rect 42166 668521 42218 668527
rect 42178 667998 42206 668521
rect 42754 667919 42782 671037
rect 42838 670873 42890 670879
rect 42838 670815 42890 670821
rect 42166 667913 42218 667919
rect 42166 667855 42218 667861
rect 42742 667913 42794 667919
rect 42742 667855 42794 667861
rect 42178 667361 42206 667855
rect 42742 667765 42794 667771
rect 42742 667707 42794 667713
rect 42166 666729 42218 666735
rect 42166 666671 42218 666677
rect 42178 666148 42206 666671
rect 42178 665329 42206 665521
rect 42166 665323 42218 665329
rect 42166 665265 42218 665271
rect 42754 665181 42782 667707
rect 42166 665175 42218 665181
rect 42166 665117 42218 665123
rect 42742 665175 42794 665181
rect 42742 665117 42794 665123
rect 42178 664964 42206 665117
rect 42740 665066 42796 665075
rect 42740 665001 42796 665010
rect 42166 664879 42218 664885
rect 42166 664821 42218 664827
rect 42178 664298 42206 664821
rect 42070 664213 42122 664219
rect 42070 664155 42122 664161
rect 42082 663706 42110 664155
rect 42166 663399 42218 663405
rect 42166 663341 42218 663347
rect 42178 663114 42206 663341
rect 42070 660957 42122 660963
rect 42070 660899 42122 660905
rect 42082 660672 42110 660899
rect 42070 660439 42122 660445
rect 42070 660381 42122 660387
rect 42082 660006 42110 660381
rect 42166 659699 42218 659705
rect 42166 659641 42218 659647
rect 42178 659340 42206 659641
rect 42166 659255 42218 659261
rect 42166 659197 42218 659203
rect 42178 659132 42206 659197
rect 42082 659104 42206 659132
rect 42082 658822 42110 659104
rect 42754 657411 42782 665001
rect 42850 664219 42878 670815
rect 42946 668585 42974 683025
rect 43126 677311 43178 677317
rect 43126 677253 43178 677259
rect 43030 677015 43082 677021
rect 43030 676957 43082 676963
rect 43042 670879 43070 676957
rect 43030 670873 43082 670879
rect 43030 670815 43082 670821
rect 43138 670824 43166 677253
rect 43318 671169 43370 671175
rect 43318 671111 43370 671117
rect 43330 671054 43358 671111
rect 43330 671026 43454 671054
rect 43522 671027 43550 685985
rect 43702 671317 43754 671323
rect 43702 671259 43754 671265
rect 43606 671243 43658 671249
rect 43606 671185 43658 671191
rect 43318 670873 43370 670879
rect 43138 670796 43262 670824
rect 43318 670815 43370 670821
rect 43426 670824 43454 671026
rect 43510 671021 43562 671027
rect 43510 670963 43562 670969
rect 43618 670972 43646 671185
rect 43714 671054 43742 671259
rect 43714 671026 43838 671054
rect 43618 670944 43742 670972
rect 43126 670725 43178 670731
rect 43126 670667 43178 670673
rect 43030 670651 43082 670657
rect 43030 670593 43082 670599
rect 42934 668579 42986 668585
rect 42934 668521 42986 668527
rect 42934 668431 42986 668437
rect 42934 668373 42986 668379
rect 42946 666735 42974 668373
rect 42934 666729 42986 666735
rect 42934 666671 42986 666677
rect 42934 666581 42986 666587
rect 42934 666523 42986 666529
rect 42838 664213 42890 664219
rect 42838 664155 42890 664161
rect 42836 662402 42892 662411
rect 42836 662337 42892 662346
rect 42070 657405 42122 657411
rect 42070 657347 42122 657353
rect 42742 657405 42794 657411
rect 42742 657347 42794 657353
rect 42082 656972 42110 657347
rect 42850 656745 42878 662337
rect 42946 660963 42974 666523
rect 43042 663405 43070 670593
rect 43138 664885 43166 670667
rect 43234 668437 43262 670796
rect 43222 668431 43274 668437
rect 43222 668373 43274 668379
rect 43330 667771 43358 670815
rect 43426 670796 43646 670824
rect 43414 670725 43466 670731
rect 43414 670667 43466 670673
rect 43510 670725 43562 670731
rect 43510 670667 43562 670673
rect 43318 667765 43370 667771
rect 43318 667707 43370 667713
rect 43426 666587 43454 670667
rect 43414 666581 43466 666587
rect 43414 666523 43466 666529
rect 43222 665323 43274 665329
rect 43222 665265 43274 665271
rect 43126 664879 43178 664885
rect 43126 664821 43178 664827
rect 43126 664731 43178 664737
rect 43126 664673 43178 664679
rect 43030 663399 43082 663405
rect 43030 663341 43082 663347
rect 43030 663251 43082 663257
rect 43030 663193 43082 663199
rect 42934 660957 42986 660963
rect 42934 660899 42986 660905
rect 42932 660774 42988 660783
rect 42932 660709 42988 660718
rect 42166 656739 42218 656745
rect 42166 656681 42218 656687
rect 42838 656739 42890 656745
rect 42838 656681 42890 656687
rect 42178 656306 42206 656681
rect 42946 656227 42974 660709
rect 43042 659705 43070 663193
rect 43138 660445 43166 664673
rect 43126 660439 43178 660445
rect 43126 660381 43178 660387
rect 43030 659699 43082 659705
rect 43030 659641 43082 659647
rect 43234 659483 43262 665265
rect 43222 659477 43274 659483
rect 43222 659419 43274 659425
rect 43028 658850 43084 658859
rect 43028 658785 43084 658794
rect 42166 656221 42218 656227
rect 42166 656163 42218 656169
rect 42934 656221 42986 656227
rect 42934 656163 42986 656169
rect 42178 655677 42206 656163
rect 43042 655561 43070 658785
rect 42166 655555 42218 655561
rect 42166 655497 42218 655503
rect 43030 655555 43082 655561
rect 43030 655497 43082 655503
rect 42178 655122 42206 655497
rect 41588 644938 41644 644947
rect 41588 644873 41590 644882
rect 41642 644873 41644 644882
rect 41590 644841 41642 644847
rect 41492 644790 41548 644799
rect 41492 644725 41548 644734
rect 41506 642537 41534 644725
rect 41588 644346 41644 644355
rect 41588 644281 41590 644290
rect 41642 644281 41644 644290
rect 41590 644249 41642 644255
rect 41780 644050 41836 644059
rect 41780 643985 41782 643994
rect 41834 643985 41836 643994
rect 41782 643953 41834 643959
rect 43522 643795 43550 670667
rect 43618 664737 43646 670796
rect 43606 664731 43658 664737
rect 43606 664673 43658 664679
rect 43714 663257 43742 670944
rect 43702 663251 43754 663257
rect 43702 663193 43754 663199
rect 43810 659261 43838 671026
rect 43798 659255 43850 659261
rect 43798 659197 43850 659203
rect 41590 643789 41642 643795
rect 41588 643754 41590 643763
rect 43510 643789 43562 643795
rect 41642 643754 41644 643763
rect 43510 643731 43562 643737
rect 41588 643689 41644 643698
rect 41588 642866 41644 642875
rect 41588 642801 41590 642810
rect 41642 642801 41644 642810
rect 43606 642827 43658 642833
rect 41590 642769 41642 642775
rect 43606 642769 43658 642775
rect 41494 642531 41546 642537
rect 41494 642473 41546 642479
rect 41506 641247 41534 642473
rect 41588 641386 41644 641395
rect 41588 641321 41590 641330
rect 41642 641321 41644 641330
rect 43510 641347 43562 641353
rect 41590 641289 41642 641295
rect 43510 641289 43562 641295
rect 41492 641238 41548 641247
rect 41492 641173 41548 641182
rect 37364 640350 37420 640359
rect 37364 640285 37420 640294
rect 34484 639314 34540 639323
rect 34484 639249 34540 639258
rect 34388 636798 34444 636807
rect 34388 636733 34444 636742
rect 28820 632802 28876 632811
rect 28820 632737 28876 632746
rect 28834 632367 28862 632737
rect 28820 632358 28876 632367
rect 28820 632293 28876 632302
rect 34402 629291 34430 636733
rect 34390 629285 34442 629291
rect 34498 629259 34526 639249
rect 34390 629227 34442 629233
rect 34484 629250 34540 629259
rect 34484 629185 34540 629194
rect 37378 627959 37406 640285
rect 41972 640054 42028 640063
rect 41972 639989 42028 639998
rect 40148 638870 40204 638879
rect 40148 638805 40204 638814
rect 40162 630697 40190 638805
rect 41684 638722 41740 638731
rect 41684 638657 41740 638666
rect 40244 637390 40300 637399
rect 40244 637325 40300 637334
rect 40150 630691 40202 630697
rect 40150 630633 40202 630639
rect 40258 628371 40286 637325
rect 41588 635318 41644 635327
rect 41588 635253 41644 635262
rect 41602 634545 41630 635253
rect 41590 634539 41642 634545
rect 41590 634481 41642 634487
rect 41588 634430 41644 634439
rect 41588 634365 41644 634374
rect 41602 634175 41630 634365
rect 41590 634169 41642 634175
rect 41590 634111 41642 634117
rect 41698 633824 41726 638657
rect 41876 637982 41932 637991
rect 41876 637917 41932 637926
rect 41780 636132 41836 636141
rect 41780 636067 41836 636076
rect 41794 634249 41822 636067
rect 41782 634243 41834 634249
rect 41782 634185 41834 634191
rect 41780 634134 41836 634143
rect 41780 634069 41836 634078
rect 41794 633953 41822 634069
rect 41782 633947 41834 633953
rect 41782 633889 41834 633895
rect 41698 633796 41822 633824
rect 41588 632358 41644 632367
rect 41588 632293 41590 632302
rect 41642 632293 41644 632302
rect 41590 632261 41642 632267
rect 40438 629285 40490 629291
rect 40438 629227 40490 629233
rect 40244 628362 40300 628371
rect 40244 628297 40300 628306
rect 37366 627953 37418 627959
rect 37366 627895 37418 627901
rect 40450 627885 40478 629227
rect 40438 627879 40490 627885
rect 40438 627821 40490 627827
rect 41794 627483 41822 633796
rect 41780 627474 41836 627483
rect 41890 627441 41918 637917
rect 41986 632103 42014 639989
rect 42164 636502 42220 636511
rect 42164 636437 42220 636446
rect 41974 632097 42026 632103
rect 41974 632039 42026 632045
rect 42070 630691 42122 630697
rect 42070 630633 42122 630639
rect 42082 627631 42110 630633
rect 42068 627622 42124 627631
rect 42068 627557 42124 627566
rect 42178 627483 42206 636437
rect 42260 635022 42316 635031
rect 42260 634957 42316 634966
rect 42164 627474 42220 627483
rect 41780 627409 41836 627418
rect 41878 627435 41930 627441
rect 42274 627441 42302 634957
rect 43126 634539 43178 634545
rect 43126 634481 43178 634487
rect 42934 634243 42986 634249
rect 42934 634185 42986 634191
rect 42838 633947 42890 633953
rect 42838 633889 42890 633895
rect 42742 632097 42794 632103
rect 42742 632039 42794 632045
rect 42164 627409 42220 627418
rect 42262 627435 42314 627441
rect 41878 627377 41930 627383
rect 42262 627377 42314 627383
rect 41878 627213 41930 627219
rect 41878 627155 41930 627161
rect 41890 626632 41918 627155
rect 42754 625369 42782 632039
rect 42166 625363 42218 625369
rect 42166 625305 42218 625311
rect 42742 625363 42794 625369
rect 42742 625305 42794 625311
rect 42178 624782 42206 625305
rect 42740 625254 42796 625263
rect 42740 625189 42796 625198
rect 42178 624037 42206 624161
rect 42166 624031 42218 624037
rect 42166 623973 42218 623979
rect 42166 623513 42218 623519
rect 42166 623455 42218 623461
rect 42178 622965 42206 623455
rect 42082 622113 42110 622340
rect 42166 622255 42218 622261
rect 42166 622197 42218 622203
rect 42070 622107 42122 622113
rect 42070 622049 42122 622055
rect 42178 621748 42206 622197
rect 42166 621663 42218 621669
rect 42166 621605 42218 621611
rect 42178 621125 42206 621605
rect 42070 620997 42122 621003
rect 42070 620939 42122 620945
rect 42082 620490 42110 620939
rect 42754 620189 42782 625189
rect 42850 622261 42878 633889
rect 42946 623519 42974 634185
rect 43030 634169 43082 634175
rect 43030 634111 43082 634117
rect 42934 623513 42986 623519
rect 42934 623455 42986 623461
rect 42934 623365 42986 623371
rect 42934 623307 42986 623313
rect 42838 622255 42890 622261
rect 42838 622197 42890 622203
rect 42836 622146 42892 622155
rect 42836 622081 42892 622090
rect 42850 620504 42878 622081
rect 42946 620652 42974 623307
rect 43042 621003 43070 634111
rect 43138 621669 43166 634481
rect 43222 627879 43274 627885
rect 43222 627821 43274 627827
rect 43126 621663 43178 621669
rect 43126 621605 43178 621611
rect 43234 621540 43262 627821
rect 43318 627435 43370 627441
rect 43318 627377 43370 627383
rect 43330 623371 43358 627377
rect 43318 623365 43370 623371
rect 43318 623307 43370 623313
rect 43138 621512 43262 621540
rect 43030 620997 43082 621003
rect 43030 620939 43082 620945
rect 42946 620624 43070 620652
rect 42850 620476 42974 620504
rect 42166 620183 42218 620189
rect 42166 620125 42218 620131
rect 42742 620183 42794 620189
rect 42742 620125 42794 620131
rect 42178 619929 42206 620125
rect 42836 619186 42892 619195
rect 42836 619121 42892 619130
rect 42070 617889 42122 617895
rect 42070 617831 42122 617837
rect 42082 617456 42110 617831
rect 42166 617223 42218 617229
rect 42166 617165 42218 617171
rect 42178 616790 42206 617165
rect 42166 616705 42218 616711
rect 42166 616647 42218 616653
rect 42178 616157 42206 616647
rect 42740 616522 42796 616531
rect 42740 616457 42796 616466
rect 42356 616374 42412 616383
rect 42356 616309 42412 616318
rect 42166 615891 42218 615897
rect 42166 615833 42218 615839
rect 42178 615606 42206 615833
rect 42166 614189 42218 614195
rect 42166 614131 42218 614137
rect 42178 613756 42206 614131
rect 42166 613671 42218 613677
rect 42166 613613 42218 613619
rect 42178 613121 42206 613613
rect 42370 612863 42398 616309
rect 42754 613677 42782 616457
rect 42850 615897 42878 619121
rect 42946 617229 42974 620476
rect 43042 617895 43070 620624
rect 43030 617889 43082 617895
rect 43030 617831 43082 617837
rect 43030 617741 43082 617747
rect 43030 617683 43082 617689
rect 42934 617223 42986 617229
rect 42934 617165 42986 617171
rect 42934 616409 42986 616415
rect 42934 616351 42986 616357
rect 42838 615891 42890 615897
rect 42838 615833 42890 615839
rect 42742 613671 42794 613677
rect 42742 613613 42794 613619
rect 42070 612857 42122 612863
rect 42070 612799 42122 612805
rect 42358 612857 42410 612863
rect 42358 612799 42410 612805
rect 42082 612498 42110 612799
rect 42946 612197 42974 616351
rect 43042 614195 43070 617683
rect 43138 616711 43166 621512
rect 43222 620405 43274 620411
rect 43222 620347 43274 620353
rect 43126 616705 43178 616711
rect 43126 616647 43178 616653
rect 43030 614189 43082 614195
rect 43030 614131 43082 614137
rect 42166 612191 42218 612197
rect 42166 612133 42218 612139
rect 42934 612191 42986 612197
rect 42934 612133 42986 612139
rect 42178 611906 42206 612133
rect 40340 601722 40396 601731
rect 40340 601657 40396 601666
rect 41588 601722 41644 601731
rect 41588 601657 41590 601666
rect 40354 599511 40382 601657
rect 41642 601657 41644 601666
rect 41590 601625 41642 601631
rect 41780 601426 41836 601435
rect 41780 601361 41782 601370
rect 41834 601361 41836 601370
rect 41782 601329 41834 601335
rect 41780 600834 41836 600843
rect 41780 600769 41782 600778
rect 41834 600769 41836 600778
rect 41782 600737 41834 600743
rect 43234 600431 43262 620347
rect 43522 619214 43550 641289
rect 43618 620411 43646 642769
rect 43702 627953 43754 627959
rect 43702 627895 43754 627901
rect 43606 620405 43658 620411
rect 43606 620347 43658 620353
rect 43714 619214 43742 627895
rect 43330 619186 43550 619214
rect 43618 619186 43742 619214
rect 41782 600425 41834 600431
rect 41780 600390 41782 600399
rect 43222 600425 43274 600431
rect 41834 600390 41836 600399
rect 43222 600367 43274 600373
rect 41780 600325 41836 600334
rect 41780 599872 41836 599881
rect 41780 599807 41782 599816
rect 41834 599807 41836 599816
rect 43222 599833 43274 599839
rect 41782 599775 41834 599781
rect 43222 599775 43274 599781
rect 40340 599502 40396 599511
rect 40340 599437 40396 599446
rect 40354 598771 40382 599437
rect 41780 599354 41836 599363
rect 41780 599289 41782 599298
rect 41834 599289 41836 599298
rect 41782 599257 41834 599263
rect 40340 598762 40396 598771
rect 40340 598697 40396 598706
rect 41780 598392 41836 598401
rect 41780 598327 41782 598336
rect 41834 598327 41836 598336
rect 41782 598295 41834 598301
rect 41782 597909 41834 597915
rect 41780 597874 41782 597883
rect 41834 597874 41836 597883
rect 41780 597809 41836 597818
rect 37364 597134 37420 597143
rect 37364 597069 37420 597078
rect 34292 596098 34348 596107
rect 34292 596033 34348 596042
rect 28820 589586 28876 589595
rect 28820 589521 28876 589530
rect 28834 589151 28862 589521
rect 28820 589142 28876 589151
rect 28820 589077 28876 589086
rect 34306 585303 34334 596033
rect 34388 594174 34444 594183
rect 34388 594109 34444 594118
rect 34402 585747 34430 594109
rect 34484 593138 34540 593147
rect 34484 593073 34540 593082
rect 34388 585738 34444 585747
rect 34388 585673 34444 585682
rect 34292 585294 34348 585303
rect 34292 585229 34348 585238
rect 34498 584817 34526 593073
rect 37378 585039 37406 597069
rect 41588 596690 41644 596699
rect 41588 596625 41590 596634
rect 41642 596625 41644 596634
rect 43126 596651 43178 596657
rect 41590 596593 41642 596599
rect 43126 596593 43178 596599
rect 40148 595654 40204 595663
rect 40148 595589 40204 595598
rect 37366 585033 37418 585039
rect 37366 584975 37418 584981
rect 40162 584891 40190 595589
rect 41972 595358 42028 595367
rect 41972 595293 42028 595302
rect 41780 594840 41836 594849
rect 41780 594775 41836 594784
rect 40244 593730 40300 593739
rect 40244 593665 40300 593674
rect 40150 584885 40202 584891
rect 40150 584827 40202 584833
rect 34486 584811 34538 584817
rect 34486 584753 34538 584759
rect 40258 584743 40286 593665
rect 41588 591066 41644 591075
rect 41588 591001 41590 591010
rect 41642 591001 41644 591010
rect 41590 590969 41642 590975
rect 41588 589142 41644 589151
rect 41588 589077 41644 589086
rect 41602 587555 41630 589077
rect 41590 587549 41642 587555
rect 41590 587491 41642 587497
rect 40246 584737 40298 584743
rect 40246 584679 40298 584685
rect 41794 584225 41822 594775
rect 41876 592990 41932 592999
rect 41876 592925 41932 592934
rect 41890 590441 41918 592925
rect 41878 590435 41930 590441
rect 41878 590377 41930 590383
rect 41878 584885 41930 584891
rect 41878 584827 41930 584833
rect 41890 584267 41918 584827
rect 41876 584258 41932 584267
rect 41782 584219 41834 584225
rect 41986 584225 42014 595293
rect 42068 592398 42124 592407
rect 42068 592333 42124 592342
rect 42082 584891 42110 592333
rect 42260 591806 42316 591815
rect 42260 591741 42316 591750
rect 42164 591362 42220 591371
rect 42164 591297 42220 591306
rect 42070 584885 42122 584891
rect 42070 584827 42122 584833
rect 42178 584299 42206 591297
rect 42274 584859 42302 591741
rect 43030 591027 43082 591033
rect 43030 590969 43082 590975
rect 42934 590435 42986 590441
rect 42934 590377 42986 590383
rect 42550 584885 42602 584891
rect 42260 584850 42316 584859
rect 42602 584833 42686 584836
rect 42550 584827 42686 584833
rect 42562 584808 42686 584827
rect 42260 584785 42316 584794
rect 42262 584737 42314 584743
rect 42262 584679 42314 584685
rect 42550 584737 42602 584743
rect 42550 584679 42602 584685
rect 42166 584293 42218 584299
rect 42274 584267 42302 584679
rect 42166 584235 42218 584241
rect 42260 584258 42316 584267
rect 41876 584193 41932 584202
rect 41974 584219 42026 584225
rect 41782 584161 41834 584167
rect 42260 584193 42316 584202
rect 41974 584161 42026 584167
rect 41782 583997 41834 584003
rect 41782 583939 41834 583945
rect 41794 583445 41822 583939
rect 42166 582147 42218 582153
rect 42166 582089 42218 582095
rect 42178 581605 42206 582089
rect 42562 581487 42590 584679
rect 42070 581481 42122 581487
rect 42070 581423 42122 581429
rect 42550 581481 42602 581487
rect 42550 581423 42602 581429
rect 42082 580974 42110 581423
rect 42658 581284 42686 584808
rect 42946 584392 42974 590377
rect 43042 584521 43070 590969
rect 43030 584515 43082 584521
rect 43030 584457 43082 584463
rect 43138 584447 43166 596593
rect 43126 584441 43178 584447
rect 42946 584364 43070 584392
rect 43126 584383 43178 584389
rect 42934 584219 42986 584225
rect 42934 584161 42986 584167
rect 42562 581256 42686 581284
rect 42070 580297 42122 580303
rect 42070 580239 42122 580245
rect 42082 579790 42110 580239
rect 42166 579335 42218 579341
rect 42166 579277 42218 579283
rect 42178 579124 42206 579277
rect 42166 578891 42218 578897
rect 42166 578833 42218 578839
rect 42178 578569 42206 578833
rect 42562 578453 42590 581256
rect 42070 578447 42122 578453
rect 42070 578389 42122 578395
rect 42550 578447 42602 578453
rect 42550 578389 42602 578395
rect 42082 577940 42110 578389
rect 42548 578338 42604 578347
rect 42548 578273 42604 578282
rect 42166 577707 42218 577713
rect 42166 577649 42218 577655
rect 42178 577274 42206 577649
rect 42070 577189 42122 577195
rect 42070 577131 42122 577137
rect 42082 576756 42110 577131
rect 42356 575378 42412 575387
rect 42356 575313 42412 575322
rect 42166 574673 42218 574679
rect 42166 574615 42218 574621
rect 42178 574240 42206 574615
rect 42166 574155 42218 574161
rect 42166 574097 42218 574103
rect 42178 573574 42206 574097
rect 42070 573489 42122 573495
rect 42070 573431 42122 573437
rect 42082 572982 42110 573431
rect 41876 572714 41932 572723
rect 41876 572649 41932 572658
rect 41890 572390 41918 572649
rect 42370 572163 42398 575313
rect 42562 573495 42590 578273
rect 42946 577195 42974 584161
rect 43042 580303 43070 584364
rect 43126 584293 43178 584299
rect 43126 584235 43178 584241
rect 43030 580297 43082 580303
rect 43030 580239 43082 580245
rect 43030 580149 43082 580155
rect 43030 580091 43082 580097
rect 43042 578897 43070 580091
rect 43030 578891 43082 578897
rect 43030 578833 43082 578839
rect 43028 578782 43084 578791
rect 43028 578717 43084 578726
rect 42934 577189 42986 577195
rect 42934 577131 42986 577137
rect 42934 577041 42986 577047
rect 42934 576983 42986 576989
rect 42946 574476 42974 576983
rect 43042 574679 43070 578717
rect 43138 577713 43166 584235
rect 43126 577707 43178 577713
rect 43126 577649 43178 577655
rect 43126 577559 43178 577565
rect 43126 577501 43178 577507
rect 43030 574673 43082 574679
rect 43030 574615 43082 574621
rect 42946 574448 43070 574476
rect 42550 573489 42602 573495
rect 42550 573431 42602 573437
rect 42934 573193 42986 573199
rect 42934 573135 42986 573141
rect 42358 572157 42410 572163
rect 42358 572099 42410 572105
rect 42838 572157 42890 572163
rect 42838 572099 42890 572105
rect 42166 571047 42218 571053
rect 42166 570989 42218 570995
rect 42178 570540 42206 570989
rect 42850 570905 42878 572099
rect 42838 570899 42890 570905
rect 42838 570841 42890 570847
rect 42166 570455 42218 570461
rect 42166 570397 42218 570403
rect 42178 570254 42206 570397
rect 42082 570226 42206 570254
rect 42082 569948 42110 570226
rect 42070 569789 42122 569795
rect 42070 569731 42122 569737
rect 42082 569282 42110 569731
rect 42946 569203 42974 573135
rect 43042 571053 43070 574448
rect 43138 574161 43166 577501
rect 43126 574155 43178 574161
rect 43126 574097 43178 574103
rect 43124 574046 43180 574055
rect 43124 573981 43180 573990
rect 43030 571047 43082 571053
rect 43030 570989 43082 570995
rect 43030 570899 43082 570905
rect 43030 570841 43082 570847
rect 43042 569795 43070 570841
rect 43138 570461 43166 573981
rect 43126 570455 43178 570461
rect 43126 570397 43178 570403
rect 43030 569789 43082 569795
rect 43030 569731 43082 569737
rect 42166 569197 42218 569203
rect 42166 569139 42218 569145
rect 42934 569197 42986 569203
rect 42934 569139 42986 569145
rect 42178 568725 42206 569139
rect 43030 541595 43082 541601
rect 43030 541537 43082 541543
rect 42934 541521 42986 541527
rect 42934 541463 42986 541469
rect 41794 539867 41822 540245
rect 41780 539858 41836 539867
rect 41780 539793 41836 539802
rect 41794 538091 41822 538424
rect 42166 538191 42218 538197
rect 42166 538133 42218 538139
rect 41780 538082 41836 538091
rect 41780 538017 41836 538026
rect 42178 537758 42206 538133
rect 41794 536315 41822 536574
rect 42946 536495 42974 541463
rect 43042 538197 43070 541537
rect 43030 538191 43082 538197
rect 43030 538133 43082 538139
rect 42166 536489 42218 536495
rect 42166 536431 42218 536437
rect 42934 536489 42986 536495
rect 42934 536431 42986 536437
rect 41780 536306 41836 536315
rect 41780 536241 41836 536250
rect 42178 535908 42206 536431
rect 41794 535131 41822 535390
rect 41780 535122 41836 535131
rect 41780 535057 41836 535066
rect 41794 534243 41822 534724
rect 41780 534234 41836 534243
rect 41780 534169 41836 534178
rect 41794 533947 41822 534058
rect 41780 533938 41836 533947
rect 41780 533873 41836 533882
rect 41794 533207 41822 533540
rect 41780 533198 41836 533207
rect 41780 533133 41836 533142
rect 41794 530839 41822 531024
rect 41780 530830 41836 530839
rect 41780 530765 41836 530774
rect 41890 530099 41918 530401
rect 41876 530090 41932 530099
rect 41876 530025 41932 530034
rect 42934 529977 42986 529983
rect 42934 529919 42986 529925
rect 42082 529359 42110 529766
rect 42068 529350 42124 529359
rect 42068 529285 42124 529294
rect 42178 528767 42206 529205
rect 42164 528758 42220 528767
rect 42164 528693 42220 528702
rect 42178 527139 42206 527365
rect 42164 527130 42220 527139
rect 42164 527065 42220 527074
rect 42178 526431 42206 526732
rect 42166 526425 42218 526431
rect 42166 526367 42218 526373
rect 42550 526425 42602 526431
rect 42550 526367 42602 526373
rect 42082 525691 42110 526066
rect 42070 525685 42122 525691
rect 42070 525627 42122 525633
rect 42358 525685 42410 525691
rect 42358 525627 42410 525633
rect 42178 525469 42206 525548
rect 42166 525463 42218 525469
rect 42166 525405 42218 525411
rect 41782 476105 41834 476111
rect 41780 476070 41782 476079
rect 41834 476070 41836 476079
rect 41780 476005 41836 476014
rect 41782 475587 41834 475593
rect 41780 475552 41782 475561
rect 41834 475552 41836 475561
rect 41780 475487 41836 475496
rect 42370 475297 42398 525627
rect 37366 475291 37418 475297
rect 37366 475233 37418 475239
rect 42358 475291 42410 475297
rect 42358 475233 42410 475239
rect 37378 470751 37406 475233
rect 41780 475034 41836 475043
rect 41780 474969 41836 474978
rect 40436 473850 40492 473859
rect 40436 473785 40492 473794
rect 39668 473258 39724 473267
rect 39668 473193 39724 473202
rect 37364 470742 37420 470751
rect 37364 470677 37420 470686
rect 34484 464378 34540 464387
rect 34484 464313 34540 464322
rect 23060 463786 23116 463795
rect 23060 463721 23116 463730
rect 23074 463351 23102 463721
rect 34498 463605 34526 464313
rect 34486 463599 34538 463605
rect 34486 463541 34538 463547
rect 23060 463342 23116 463351
rect 23060 463277 23116 463286
rect 23062 437847 23114 437853
rect 23062 437789 23114 437795
rect 23074 422757 23102 437789
rect 39682 437724 39710 473193
rect 39764 472370 39820 472379
rect 39764 472305 39820 472314
rect 39778 437853 39806 472305
rect 39766 437847 39818 437853
rect 39766 437789 39818 437795
rect 39862 437847 39914 437853
rect 39862 437789 39914 437795
rect 39874 437724 39902 437789
rect 39682 437696 39902 437724
rect 39682 424279 39710 437696
rect 40450 425315 40478 473785
rect 41590 472479 41642 472485
rect 41590 472421 41642 472427
rect 41602 472231 41630 472421
rect 41794 472411 41822 474969
rect 41878 474625 41930 474631
rect 41876 474590 41878 474599
rect 41930 474590 41932 474599
rect 41876 474525 41932 474534
rect 41782 472405 41834 472411
rect 41782 472347 41834 472353
rect 41588 472222 41644 472231
rect 41588 472157 41644 472166
rect 42562 469377 42590 526367
rect 42946 525469 42974 529919
rect 42934 525463 42986 525469
rect 42934 525405 42986 525411
rect 43234 474631 43262 599775
rect 43330 597915 43358 619186
rect 43618 617747 43646 619186
rect 43606 617741 43658 617747
rect 43606 617683 43658 617689
rect 43414 599315 43466 599321
rect 43414 599257 43466 599263
rect 43318 597909 43370 597915
rect 43318 597851 43370 597857
rect 43330 596213 43358 597851
rect 43318 596207 43370 596213
rect 43318 596149 43370 596155
rect 43318 584441 43370 584447
rect 43318 584383 43370 584389
rect 43330 582153 43358 584383
rect 43318 582147 43370 582153
rect 43318 582089 43370 582095
rect 43222 474625 43274 474631
rect 43222 474567 43274 474573
rect 43426 473119 43454 599257
rect 43894 598353 43946 598359
rect 43894 598295 43946 598301
rect 43798 585033 43850 585039
rect 43798 584975 43850 584981
rect 43606 584811 43658 584817
rect 43606 584753 43658 584759
rect 43510 584515 43562 584521
rect 43510 584457 43562 584463
rect 43522 580155 43550 584457
rect 43510 580149 43562 580155
rect 43510 580091 43562 580097
rect 43618 577565 43646 584753
rect 43606 577559 43658 577565
rect 43606 577501 43658 577507
rect 43810 577047 43838 584975
rect 43798 577041 43850 577047
rect 43798 576983 43850 576989
rect 43906 570254 43934 598295
rect 43522 570226 43934 570254
rect 43412 473110 43468 473119
rect 43412 473045 43468 473054
rect 43522 472485 43550 570226
rect 43510 472479 43562 472485
rect 43510 472421 43562 472427
rect 41590 469371 41642 469377
rect 41590 469313 41642 469319
rect 42550 469371 42602 469377
rect 42550 469313 42602 469319
rect 41602 468827 41630 469313
rect 41588 468818 41644 468827
rect 41588 468753 41644 468762
rect 41780 463638 41836 463647
rect 41780 463573 41782 463582
rect 41834 463573 41836 463582
rect 41782 463541 41834 463547
rect 41588 426934 41644 426943
rect 41588 426869 41590 426878
rect 41642 426869 41644 426878
rect 41590 426837 41642 426843
rect 41780 426564 41836 426573
rect 41780 426499 41782 426508
rect 41834 426499 41836 426508
rect 41782 426467 41834 426473
rect 41780 426046 41836 426055
rect 41780 425981 41782 425990
rect 41834 425981 41836 425990
rect 41782 425949 41834 425955
rect 40436 425306 40492 425315
rect 40436 425241 40492 425250
rect 41588 424862 41644 424871
rect 41588 424797 41590 424806
rect 41642 424797 41644 424806
rect 43318 424823 43370 424829
rect 41590 424765 41642 424771
rect 43318 424765 43370 424771
rect 34484 424270 34540 424279
rect 34484 424205 34540 424214
rect 39668 424270 39724 424279
rect 39668 424205 39724 424214
rect 23062 422751 23114 422757
rect 23062 422693 23114 422699
rect 34498 421763 34526 424205
rect 41780 423530 41836 423539
rect 41780 423465 41782 423474
rect 41834 423465 41836 423474
rect 43222 423491 43274 423497
rect 41782 423433 41834 423439
rect 43222 423433 43274 423439
rect 41588 422790 41644 422799
rect 41588 422725 41590 422734
rect 41642 422725 41644 422734
rect 41590 422693 41642 422699
rect 34484 421754 34540 421763
rect 34484 421689 34540 421698
rect 39764 420866 39820 420875
rect 39764 420801 39820 420810
rect 39668 419238 39724 419247
rect 39668 419173 39724 419182
rect 39682 416435 39710 419173
rect 39668 416426 39724 416435
rect 39668 416361 39724 416370
rect 39778 414955 39806 420801
rect 41602 420537 41630 422693
rect 41590 420531 41642 420537
rect 41590 420473 41642 420479
rect 39956 420274 40012 420283
rect 39956 420209 40012 420218
rect 39860 419830 39916 419839
rect 39860 419765 39916 419774
rect 39874 417577 39902 419765
rect 39862 417571 39914 417577
rect 39862 417513 39914 417519
rect 39970 416879 39998 420209
rect 40244 418794 40300 418803
rect 40244 418729 40300 418738
rect 40052 418350 40108 418359
rect 40052 418285 40108 418294
rect 39956 416870 40012 416879
rect 39956 416805 40012 416814
rect 40066 416287 40094 418285
rect 40148 417906 40204 417915
rect 40148 417841 40204 417850
rect 40162 417503 40190 417841
rect 40150 417497 40202 417503
rect 40150 417439 40202 417445
rect 40258 417323 40286 418729
rect 41782 417571 41834 417577
rect 41782 417513 41834 417519
rect 40244 417314 40300 417323
rect 40244 417249 40300 417258
rect 41588 416426 41644 416435
rect 41588 416361 41644 416370
rect 40052 416278 40108 416287
rect 40052 416213 40108 416222
rect 41602 415209 41630 416361
rect 41590 415203 41642 415209
rect 41590 415145 41642 415151
rect 39764 414946 39820 414955
rect 39764 414881 39820 414890
rect 23060 414798 23116 414807
rect 23060 414733 23116 414742
rect 23074 414363 23102 414733
rect 23060 414354 23116 414363
rect 23060 414289 23116 414298
rect 41588 414354 41644 414363
rect 41588 414289 41590 414298
rect 41642 414289 41644 414298
rect 41590 414257 41642 414263
rect 41794 413433 41822 417513
rect 42934 417497 42986 417503
rect 42934 417439 42986 417445
rect 41876 416130 41932 416139
rect 41876 416065 41932 416074
rect 41890 414765 41918 416065
rect 41878 414759 41930 414765
rect 41878 414701 41930 414707
rect 41782 413427 41834 413433
rect 41782 413369 41834 413375
rect 41782 413205 41834 413211
rect 41782 413147 41834 413153
rect 41794 412624 41822 413147
rect 41876 411246 41932 411255
rect 41876 411181 41932 411190
rect 41890 410805 41918 411181
rect 42178 409733 42206 410182
rect 42166 409727 42218 409733
rect 42166 409669 42218 409675
rect 42838 409727 42890 409733
rect 42838 409669 42890 409675
rect 42166 409505 42218 409511
rect 42166 409447 42218 409453
rect 42178 408965 42206 409447
rect 42850 408974 42878 409669
rect 42946 409511 42974 417439
rect 43126 415203 43178 415209
rect 43126 415145 43178 415151
rect 43030 414759 43082 414765
rect 43030 414701 43082 414707
rect 42934 409505 42986 409511
rect 42934 409447 42986 409453
rect 42850 408946 42974 408974
rect 42082 408031 42110 408332
rect 42166 408247 42218 408253
rect 42166 408189 42218 408195
rect 42070 408025 42122 408031
rect 42070 407967 42122 407973
rect 42178 407769 42206 408189
rect 42838 408025 42890 408031
rect 42838 407967 42890 407973
rect 41780 407694 41836 407703
rect 41780 407629 41836 407638
rect 41794 407148 41822 407629
rect 42166 406915 42218 406921
rect 42166 406857 42218 406863
rect 42178 406482 42206 406857
rect 42068 406066 42124 406075
rect 42068 406001 42124 406010
rect 42082 405929 42110 406001
rect 41780 403846 41836 403855
rect 41780 403781 41836 403790
rect 41794 403448 41822 403781
rect 42164 403106 42220 403115
rect 42164 403041 42220 403050
rect 42178 402782 42206 403041
rect 41876 402662 41932 402671
rect 42850 402629 42878 407967
rect 42946 406107 42974 408946
rect 43042 408253 43070 414701
rect 43030 408247 43082 408253
rect 43030 408189 43082 408195
rect 43138 406921 43166 415145
rect 43126 406915 43178 406921
rect 43126 406857 43178 406863
rect 42934 406101 42986 406107
rect 42934 406043 42986 406049
rect 41876 402597 41932 402606
rect 42838 402623 42890 402629
rect 41890 402157 41918 402597
rect 42838 402565 42890 402571
rect 41780 401922 41836 401931
rect 41780 401857 41836 401866
rect 41794 401598 41822 401857
rect 41780 400146 41836 400155
rect 41780 400081 41836 400090
rect 41794 399748 41822 400081
rect 41780 399406 41836 399415
rect 41780 399341 41836 399350
rect 41794 399121 41822 399341
rect 41780 398814 41836 398823
rect 41780 398749 41836 398758
rect 41794 398490 41822 398749
rect 42082 394563 42110 397898
rect 42070 394557 42122 394563
rect 42070 394499 42122 394505
rect 41780 388750 41836 388759
rect 41780 388685 41836 388694
rect 41794 386391 41822 388685
rect 41780 386382 41836 386391
rect 41780 386317 41836 386326
rect 41590 385973 41642 385979
rect 41588 385938 41590 385947
rect 41642 385938 41644 385947
rect 41588 385873 41644 385882
rect 41588 385346 41644 385355
rect 41588 385281 41590 385290
rect 41642 385281 41644 385290
rect 41590 385249 41642 385255
rect 41590 384789 41642 384795
rect 41588 384754 41590 384763
rect 41642 384754 41644 384763
rect 41588 384689 41644 384698
rect 41588 383866 41644 383875
rect 41588 383801 41590 383810
rect 41642 383801 41644 383810
rect 41590 383769 41642 383775
rect 34484 383274 34540 383283
rect 34484 383209 34540 383218
rect 34498 378843 34526 383209
rect 41794 383135 41822 386317
rect 41876 385050 41932 385059
rect 41876 384985 41878 384994
rect 41930 384985 41932 384994
rect 41878 384953 41930 384959
rect 41780 383126 41836 383135
rect 41780 383061 41836 383070
rect 41588 382386 41644 382395
rect 41588 382321 41590 382330
rect 41642 382321 41644 382330
rect 41590 382289 41642 382295
rect 43234 382057 43262 423433
rect 43330 384795 43358 424765
rect 43318 384789 43370 384795
rect 43318 384731 43370 384737
rect 43414 383827 43466 383833
rect 43414 383769 43466 383775
rect 41782 382051 41834 382057
rect 41780 382016 41782 382025
rect 43222 382051 43274 382057
rect 41834 382016 41836 382025
rect 43222 381993 43274 381999
rect 41780 381951 41836 381960
rect 39188 381350 39244 381359
rect 39188 381285 39244 381294
rect 34484 378834 34540 378843
rect 34484 378769 34540 378778
rect 28820 373802 28876 373811
rect 28820 373737 28876 373746
rect 28834 373367 28862 373737
rect 28820 373358 28876 373367
rect 28820 373293 28876 373302
rect 39202 372331 39230 381285
rect 39284 380906 39340 380915
rect 39284 380841 39340 380850
rect 39298 373811 39326 380841
rect 39476 379278 39532 379287
rect 39476 379213 39532 379222
rect 39490 374361 39518 379213
rect 40052 378390 40108 378399
rect 40052 378325 40108 378334
rect 39764 377798 39820 377807
rect 39764 377733 39820 377742
rect 39478 374355 39530 374361
rect 39478 374297 39530 374303
rect 39284 373802 39340 373811
rect 39284 373737 39340 373746
rect 39778 373219 39806 377733
rect 39956 377354 40012 377363
rect 39956 377289 40012 377298
rect 39970 373367 39998 377289
rect 40066 373959 40094 378325
rect 42452 376910 42508 376919
rect 42452 376845 42508 376854
rect 41492 376318 41548 376327
rect 41492 376253 41548 376262
rect 41506 374287 41534 376253
rect 41684 375282 41740 375291
rect 41684 375217 41740 375226
rect 41588 374838 41644 374847
rect 41588 374773 41644 374782
rect 41494 374281 41546 374287
rect 41494 374223 41546 374229
rect 40052 373950 40108 373959
rect 40052 373885 40108 373894
rect 39956 373358 40012 373367
rect 39956 373293 40012 373302
rect 39764 373210 39820 373219
rect 39764 373145 39820 373154
rect 39188 372322 39244 372331
rect 39188 372257 39244 372266
rect 41602 371993 41630 374773
rect 41590 371987 41642 371993
rect 41590 371929 41642 371935
rect 41698 371845 41726 375217
rect 41780 374542 41836 374551
rect 41780 374477 41836 374486
rect 41794 373589 41822 374477
rect 41878 374355 41930 374361
rect 41878 374297 41930 374303
rect 41780 373580 41836 373589
rect 41780 373515 41782 373524
rect 41834 373515 41836 373524
rect 41782 373483 41834 373489
rect 41686 371839 41738 371845
rect 41686 371781 41738 371787
rect 41890 370217 41918 374297
rect 41878 370211 41930 370217
rect 41878 370153 41930 370159
rect 41878 369989 41930 369995
rect 41878 369931 41930 369937
rect 41890 369445 41918 369931
rect 41780 368178 41836 368187
rect 41780 368113 41836 368122
rect 41794 367632 41822 368113
rect 42178 366591 42206 366966
rect 42466 366739 42494 376845
rect 43030 374281 43082 374287
rect 43030 374223 43082 374229
rect 42838 371987 42890 371993
rect 42838 371929 42890 371935
rect 42454 366733 42506 366739
rect 42454 366675 42506 366681
rect 42166 366585 42218 366591
rect 42166 366527 42218 366533
rect 42454 366585 42506 366591
rect 42454 366527 42506 366533
rect 42070 366289 42122 366295
rect 42070 366231 42122 366237
rect 42082 365782 42110 366231
rect 42082 364741 42110 365116
rect 42166 365031 42218 365037
rect 42166 364973 42218 364979
rect 42070 364735 42122 364741
rect 42070 364677 42122 364683
rect 42178 364569 42206 364973
rect 42070 364291 42122 364297
rect 42070 364233 42122 364239
rect 42082 363932 42110 364233
rect 42166 363847 42218 363853
rect 42166 363789 42218 363795
rect 42178 363266 42206 363789
rect 41780 362850 41836 362859
rect 41780 362785 41836 362794
rect 41794 362748 41822 362785
rect 42466 362003 42494 366527
rect 42850 365037 42878 371929
rect 42934 371839 42986 371845
rect 42934 371781 42986 371787
rect 42838 365031 42890 365037
rect 42838 364973 42890 364979
rect 42838 364735 42890 364741
rect 42838 364677 42890 364683
rect 42454 361997 42506 362003
rect 42454 361939 42506 361945
rect 41780 360630 41836 360639
rect 41780 360565 41836 360574
rect 41794 360232 41822 360565
rect 42850 360005 42878 364677
rect 42946 363853 42974 371781
rect 43042 364297 43070 374223
rect 43030 364291 43082 364297
rect 43030 364233 43082 364239
rect 42934 363847 42986 363853
rect 42934 363789 42986 363795
rect 42838 359999 42890 360005
rect 42838 359941 42890 359947
rect 41972 359890 42028 359899
rect 41972 359825 42028 359834
rect 41986 359601 42014 359825
rect 42068 359298 42124 359307
rect 42068 359233 42124 359242
rect 42082 358974 42110 359233
rect 41780 358854 41836 358863
rect 41780 358789 41836 358798
rect 41794 358382 41822 358789
rect 41876 356930 41932 356939
rect 41876 356865 41932 356874
rect 41890 356565 41918 356865
rect 41780 356190 41836 356199
rect 41780 356125 41836 356134
rect 41794 355940 41822 356125
rect 42164 355598 42220 355607
rect 42164 355533 42220 355542
rect 42178 355274 42206 355533
rect 42178 351347 42206 354725
rect 42166 351341 42218 351347
rect 42166 351283 42218 351289
rect 41684 343166 41740 343175
rect 41684 343101 41740 343110
rect 41588 340650 41644 340659
rect 41588 340585 41590 340594
rect 41642 340585 41644 340594
rect 41590 340553 41642 340559
rect 41698 340067 41726 343101
rect 41780 342870 41836 342879
rect 41780 342805 41782 342814
rect 41834 342805 41836 342814
rect 41782 342773 41834 342779
rect 41780 342352 41836 342361
rect 41780 342287 41782 342296
rect 41834 342287 41836 342296
rect 41782 342255 41834 342261
rect 41780 341834 41836 341843
rect 41780 341769 41782 341778
rect 41834 341769 41836 341778
rect 41782 341737 41834 341743
rect 43426 341431 43454 383769
rect 43510 382347 43562 382353
rect 43510 382289 43562 382295
rect 41782 341425 41834 341431
rect 41780 341390 41782 341399
rect 43414 341425 43466 341431
rect 41834 341390 41836 341399
rect 43414 341367 43466 341373
rect 41780 341325 41836 341334
rect 43222 340611 43274 340617
rect 43222 340553 43274 340559
rect 41780 340354 41836 340363
rect 41780 340289 41782 340298
rect 41834 340289 41836 340298
rect 41782 340257 41834 340263
rect 41684 340058 41740 340067
rect 41684 339993 41740 340002
rect 41782 339501 41834 339507
rect 41782 339443 41834 339449
rect 41588 339170 41644 339179
rect 41588 339105 41590 339114
rect 41642 339105 41644 339114
rect 41590 339073 41642 339079
rect 41794 338883 41822 339443
rect 41780 338874 41836 338883
rect 41780 338809 41836 338818
rect 28724 338134 28780 338143
rect 28724 338069 28780 338078
rect 28738 329115 28766 338069
rect 39764 337690 39820 337699
rect 39764 337625 39820 337634
rect 39284 337098 39340 337107
rect 39284 337033 39340 337042
rect 39298 330743 39326 337033
rect 39778 331187 39806 337625
rect 41780 335766 41836 335775
rect 41780 335701 41836 335710
rect 41492 333694 41548 333703
rect 41492 333629 41548 333638
rect 41396 333102 41452 333111
rect 41396 333037 41452 333046
rect 41410 331219 41438 333037
rect 41398 331213 41450 331219
rect 39764 331178 39820 331187
rect 41398 331155 41450 331161
rect 41506 331145 41534 333629
rect 41588 331622 41644 331631
rect 41588 331557 41644 331566
rect 39764 331113 39820 331122
rect 41494 331139 41546 331145
rect 41494 331081 41546 331087
rect 39284 330734 39340 330743
rect 39284 330669 39340 330678
rect 28820 330586 28876 330595
rect 28820 330521 28876 330530
rect 28834 330151 28862 330521
rect 28820 330142 28876 330151
rect 28820 330077 28876 330086
rect 28724 329106 28780 329115
rect 28724 329041 28780 329050
rect 41602 328851 41630 331557
rect 41590 328845 41642 328851
rect 41590 328787 41642 328793
rect 41794 327075 41822 335701
rect 41876 331326 41932 331335
rect 41876 331261 41932 331270
rect 41890 330447 41918 331261
rect 42742 331213 42794 331219
rect 42742 331155 42794 331161
rect 41876 330438 41932 330447
rect 41876 330373 41878 330382
rect 41930 330373 41932 330382
rect 41878 330341 41930 330347
rect 42754 328334 42782 331155
rect 43030 331139 43082 331145
rect 43030 331081 43082 331087
rect 42934 328845 42986 328851
rect 42934 328787 42986 328793
rect 42754 328306 42878 328334
rect 41782 327069 41834 327075
rect 41782 327011 41834 327017
rect 41782 326773 41834 326779
rect 41782 326715 41834 326721
rect 41794 326266 41822 326715
rect 42850 325688 42878 328306
rect 42946 325817 42974 328787
rect 42934 325811 42986 325817
rect 42934 325753 42986 325759
rect 42850 325660 42974 325688
rect 41780 324962 41836 324971
rect 41780 324897 41836 324906
rect 41794 324416 41822 324897
rect 42082 323375 42110 323750
rect 42070 323369 42122 323375
rect 42070 323311 42122 323317
rect 42454 323369 42506 323375
rect 42454 323311 42506 323317
rect 42166 323147 42218 323153
rect 42166 323089 42218 323095
rect 42178 322566 42206 323089
rect 42082 321692 42110 321900
rect 41974 321667 42026 321673
rect 42082 321664 42206 321692
rect 41974 321609 42026 321615
rect 41986 321382 42014 321609
rect 42178 321525 42206 321664
rect 42166 321519 42218 321525
rect 42166 321461 42218 321467
rect 42166 321297 42218 321303
rect 42166 321239 42218 321245
rect 42178 320716 42206 321239
rect 41780 320522 41836 320531
rect 41780 320457 41836 320466
rect 41794 320081 41822 320457
rect 41780 319782 41836 319791
rect 41780 319717 41836 319726
rect 41794 319532 41822 319717
rect 42466 319675 42494 323311
rect 42946 321692 42974 325660
rect 43042 323153 43070 331081
rect 43126 325811 43178 325817
rect 43126 325753 43178 325759
rect 43030 323147 43082 323153
rect 43030 323089 43082 323095
rect 42946 321664 43070 321692
rect 43138 321673 43166 325753
rect 43042 321303 43070 321664
rect 43126 321667 43178 321673
rect 43126 321609 43178 321615
rect 43126 321519 43178 321525
rect 43126 321461 43178 321467
rect 43030 321297 43082 321303
rect 43030 321239 43082 321245
rect 42454 319669 42506 319675
rect 42454 319611 42506 319617
rect 41876 317414 41932 317423
rect 41876 317349 41932 317358
rect 41890 317045 41918 317349
rect 43138 316789 43166 321461
rect 43126 316783 43178 316789
rect 43126 316725 43178 316731
rect 41780 316674 41836 316683
rect 41780 316609 41836 316618
rect 41794 316424 41822 316609
rect 41780 316230 41836 316239
rect 41780 316165 41836 316174
rect 41794 315758 41822 316165
rect 41780 315490 41836 315499
rect 41780 315425 41836 315434
rect 41794 315205 41822 315425
rect 42068 313714 42124 313723
rect 42068 313649 42124 313658
rect 42082 313390 42110 313649
rect 41780 313122 41836 313131
rect 41780 313057 41836 313066
rect 41794 312724 41822 313057
rect 42164 312530 42220 312539
rect 42164 312465 42220 312474
rect 42178 312058 42206 312465
rect 42178 308131 42206 311540
rect 42166 308125 42218 308131
rect 42166 308067 42218 308073
rect 39766 299689 39818 299695
rect 39766 299631 39818 299637
rect 41780 299654 41836 299663
rect 39668 298766 39724 298775
rect 39668 298701 39724 298710
rect 28724 294918 28780 294927
rect 28724 294853 28780 294862
rect 28738 285159 28766 294853
rect 39682 293775 39710 298701
rect 39778 296555 39806 299631
rect 41780 299589 41782 299598
rect 41834 299589 41836 299598
rect 41782 299557 41834 299563
rect 41780 299210 41836 299219
rect 41780 299145 41782 299154
rect 41834 299145 41836 299154
rect 41782 299113 41834 299119
rect 43234 298215 43262 340553
rect 43318 340315 43370 340321
rect 43318 340257 43370 340263
rect 43330 300953 43358 340257
rect 43522 339507 43550 382289
rect 43510 339501 43562 339507
rect 43510 339443 43562 339449
rect 43414 339131 43466 339137
rect 43414 339073 43466 339079
rect 43426 328334 43454 339073
rect 43426 328306 43550 328334
rect 43318 300947 43370 300953
rect 43318 300889 43370 300895
rect 43330 299695 43358 300889
rect 43318 299689 43370 299695
rect 43318 299631 43370 299637
rect 41782 298209 41834 298215
rect 41780 298174 41782 298183
rect 43222 298209 43274 298215
rect 41834 298174 41836 298183
rect 43222 298151 43274 298157
rect 43522 298141 43550 328306
rect 41780 298109 41836 298118
rect 43510 298135 43562 298141
rect 43510 298077 43562 298083
rect 41780 297656 41836 297665
rect 41780 297591 41782 297600
rect 41834 297591 41836 297600
rect 43414 297617 43466 297623
rect 41782 297559 41834 297565
rect 43414 297559 43466 297565
rect 41780 297138 41836 297147
rect 41780 297073 41782 297082
rect 41834 297073 41836 297082
rect 43318 297099 43370 297105
rect 41782 297041 41834 297047
rect 43318 297041 43370 297047
rect 39958 296729 40010 296735
rect 39958 296671 40010 296677
rect 39764 296546 39820 296555
rect 39764 296481 39820 296490
rect 39970 295963 39998 296671
rect 39956 295954 40012 295963
rect 39956 295889 40012 295898
rect 41588 295954 41644 295963
rect 41588 295889 41590 295898
rect 41642 295889 41644 295898
rect 43222 295915 43274 295921
rect 41590 295857 41642 295863
rect 43222 295857 43274 295863
rect 39670 293769 39722 293775
rect 39670 293711 39722 293717
rect 41780 292624 41836 292633
rect 41780 292559 41836 292568
rect 41492 290478 41548 290487
rect 41492 290413 41548 290422
rect 28820 287370 28876 287379
rect 28820 287305 28876 287314
rect 28834 286935 28862 287305
rect 28820 286926 28876 286935
rect 28820 286861 28876 286870
rect 41506 285339 41534 290413
rect 41684 288850 41740 288859
rect 41684 288785 41740 288794
rect 41588 288406 41644 288415
rect 41588 288341 41644 288350
rect 41494 285333 41546 285339
rect 41494 285275 41546 285281
rect 41602 285191 41630 288341
rect 41698 285265 41726 288785
rect 41686 285259 41738 285265
rect 41686 285201 41738 285207
rect 41590 285185 41642 285191
rect 28724 285150 28780 285159
rect 41590 285127 41642 285133
rect 28724 285085 28780 285094
rect 41794 283859 41822 292559
rect 42452 290182 42508 290191
rect 42452 290117 42508 290126
rect 42466 288014 42494 290117
rect 42466 287986 42590 288014
rect 41876 287222 41932 287231
rect 41876 287157 41878 287166
rect 41930 287157 41932 287166
rect 41878 287125 41930 287131
rect 41782 283853 41834 283859
rect 41782 283795 41834 283801
rect 41782 283557 41834 283563
rect 41782 283499 41834 283505
rect 41794 283050 41822 283499
rect 42562 282254 42590 287986
rect 43126 285333 43178 285339
rect 43126 285275 43178 285281
rect 43030 285259 43082 285265
rect 43030 285201 43082 285207
rect 42934 285185 42986 285191
rect 42934 285127 42986 285133
rect 42466 282226 42590 282254
rect 41876 281746 41932 281755
rect 41876 281681 41932 281690
rect 41890 281200 41918 281681
rect 42466 281607 42494 282226
rect 42452 281598 42508 281607
rect 42452 281533 42508 281542
rect 42082 280159 42110 280534
rect 42070 280153 42122 280159
rect 42070 280095 42122 280101
rect 42838 280153 42890 280159
rect 42838 280095 42890 280101
rect 42166 279931 42218 279937
rect 42166 279873 42218 279879
rect 42178 279350 42206 279873
rect 42082 278531 42110 278721
rect 42166 278599 42218 278605
rect 42166 278541 42218 278547
rect 42070 278525 42122 278531
rect 42070 278467 42122 278473
rect 42178 278166 42206 278541
rect 42164 278046 42220 278055
rect 42164 277981 42220 277990
rect 42178 277500 42206 277981
rect 42070 277415 42122 277421
rect 42070 277357 42122 277363
rect 42082 276908 42110 277357
rect 41780 276566 41836 276575
rect 41780 276501 41836 276510
rect 41794 276316 41822 276501
rect 42850 276459 42878 280095
rect 42946 278605 42974 285127
rect 42934 278599 42986 278605
rect 42934 278541 42986 278547
rect 43042 277421 43070 285201
rect 43138 279937 43166 285275
rect 43126 279931 43178 279937
rect 43126 279873 43178 279879
rect 43126 278525 43178 278531
rect 43126 278467 43178 278473
rect 43030 277415 43082 277421
rect 43030 277357 43082 277363
rect 42838 276453 42890 276459
rect 42838 276395 42890 276401
rect 41780 274198 41836 274207
rect 41780 274133 41836 274142
rect 41794 273845 41822 274133
rect 41780 273606 41836 273615
rect 43138 273573 43166 278467
rect 41780 273541 41836 273550
rect 43126 273567 43178 273573
rect 41794 273208 41822 273541
rect 43126 273509 43178 273515
rect 41780 272866 41836 272875
rect 41780 272801 41836 272810
rect 41794 272542 41822 272801
rect 41780 272422 41836 272431
rect 41780 272357 41836 272366
rect 41794 272024 41822 272357
rect 42068 270646 42124 270655
rect 42068 270581 42124 270590
rect 42082 270174 42110 270581
rect 41780 270054 41836 270063
rect 41780 269989 41836 269998
rect 41794 269508 41822 269989
rect 41876 269314 41932 269323
rect 41876 269249 41932 269258
rect 41890 268877 41918 269249
rect 42166 268609 42218 268615
rect 42166 268551 42218 268557
rect 42178 268324 42206 268551
rect 23062 265057 23114 265063
rect 23062 264999 23114 265005
rect 23074 253339 23102 264999
rect 43234 264989 43262 295857
rect 43222 264983 43274 264989
rect 43222 264925 43274 264931
rect 43330 264915 43358 297041
rect 43318 264909 43370 264915
rect 43318 264851 43370 264857
rect 23350 263651 23402 263657
rect 23350 263593 23402 263599
rect 23254 263577 23306 263583
rect 23254 263519 23306 263525
rect 23158 262171 23210 262177
rect 23158 262113 23210 262119
rect 23170 254227 23198 262113
rect 23156 254218 23212 254227
rect 23156 254153 23212 254162
rect 23060 253330 23116 253339
rect 23060 253265 23116 253274
rect 23266 252747 23294 263519
rect 23362 253339 23390 263593
rect 43316 263542 43372 263551
rect 43316 263477 43372 263486
rect 43330 262177 43358 263477
rect 43318 262171 43370 262177
rect 43318 262113 43370 262119
rect 40246 256399 40298 256405
rect 40246 256341 40298 256347
rect 40258 256299 40286 256341
rect 40244 256290 40300 256299
rect 40244 256225 40300 256234
rect 41588 255698 41644 255707
rect 41588 255633 41644 255642
rect 41602 253519 41630 255633
rect 41782 255437 41834 255443
rect 41780 255402 41782 255411
rect 41834 255402 41836 255411
rect 41780 255337 41836 255346
rect 41782 254993 41834 254999
rect 41780 254958 41782 254967
rect 41834 254958 41836 254967
rect 41780 254893 41836 254902
rect 41780 254514 41836 254523
rect 41780 254449 41782 254458
rect 41834 254449 41836 254458
rect 41782 254417 41834 254423
rect 41590 253513 41642 253519
rect 41590 253455 41642 253461
rect 23348 253330 23404 253339
rect 23348 253265 23404 253274
rect 23252 252738 23308 252747
rect 23252 252673 23308 252682
rect 41876 249482 41932 249491
rect 41876 249417 41932 249426
rect 41684 247262 41740 247271
rect 41684 247197 41740 247206
rect 41300 246818 41356 246827
rect 41300 246753 41356 246762
rect 41314 244565 41342 246753
rect 41396 245634 41452 245643
rect 41396 245569 41452 245578
rect 41410 244639 41438 245569
rect 41492 245190 41548 245199
rect 41492 245125 41548 245134
rect 41506 244713 41534 245125
rect 41590 245003 41642 245009
rect 41590 244945 41642 244951
rect 41602 244755 41630 244945
rect 41588 244746 41644 244755
rect 41494 244707 41546 244713
rect 41588 244681 41644 244690
rect 41494 244649 41546 244655
rect 41398 244633 41450 244639
rect 41398 244575 41450 244581
rect 41302 244559 41354 244565
rect 41302 244501 41354 244507
rect 41588 243710 41644 243719
rect 41588 243645 41644 243654
rect 41602 242641 41630 243645
rect 41590 242635 41642 242641
rect 41590 242577 41642 242583
rect 41698 242049 41726 247197
rect 41780 244894 41836 244903
rect 41780 244829 41782 244838
rect 41834 244829 41836 244838
rect 41782 244797 41834 244803
rect 41686 242043 41738 242049
rect 41686 241985 41738 241991
rect 41890 240643 41918 249417
rect 42934 244707 42986 244713
rect 42934 244649 42986 244655
rect 42838 244633 42890 244639
rect 42838 244575 42890 244581
rect 42742 242043 42794 242049
rect 42742 241985 42794 241991
rect 41878 240637 41930 240643
rect 41878 240579 41930 240585
rect 41878 240415 41930 240421
rect 41878 240357 41930 240363
rect 41890 239834 41918 240357
rect 41794 237947 41822 237984
rect 41780 237938 41836 237947
rect 41780 237873 41836 237882
rect 42754 236721 42782 241985
rect 42166 236715 42218 236721
rect 42166 236657 42218 236663
rect 42742 236715 42794 236721
rect 42742 236657 42794 236663
rect 42178 236165 42206 236657
rect 42742 236567 42794 236573
rect 42742 236509 42794 236515
rect 42166 235457 42218 235463
rect 42166 235399 42218 235405
rect 42178 234950 42206 235399
rect 42754 234871 42782 236509
rect 42166 234865 42218 234871
rect 42166 234807 42218 234813
rect 42742 234865 42794 234871
rect 42742 234807 42794 234813
rect 42178 234325 42206 234807
rect 42850 234057 42878 244575
rect 42946 235463 42974 244649
rect 43030 244559 43082 244565
rect 43030 244501 43082 244507
rect 43042 236573 43070 244501
rect 43030 236567 43082 236573
rect 43030 236509 43082 236515
rect 42934 235457 42986 235463
rect 42934 235399 42986 235405
rect 42070 234051 42122 234057
rect 42070 233993 42122 233999
rect 42838 234051 42890 234057
rect 42838 233993 42890 233999
rect 42082 233692 42110 233993
rect 41780 233350 41836 233359
rect 41780 233285 41836 233294
rect 41794 233129 41822 233285
rect 41780 231130 41836 231139
rect 41780 231065 41836 231074
rect 41794 230658 41822 231065
rect 41780 230390 41836 230399
rect 41780 230325 41836 230334
rect 41794 229992 41822 230325
rect 41780 229798 41836 229807
rect 41780 229733 41836 229742
rect 41794 229357 41822 229733
rect 41780 229058 41836 229067
rect 41780 228993 41836 229002
rect 41794 228808 41822 228993
rect 41780 227430 41836 227439
rect 41780 227365 41836 227374
rect 41794 226958 41822 227365
rect 41780 226690 41836 226699
rect 41780 226625 41836 226634
rect 41794 226321 41822 226625
rect 42068 226246 42124 226255
rect 42068 226181 42124 226190
rect 42082 225700 42110 226181
rect 42082 221773 42110 225108
rect 42070 221767 42122 221773
rect 42070 221709 42122 221715
rect 41782 213331 41834 213337
rect 41780 213296 41782 213305
rect 41834 213296 41836 213305
rect 41780 213231 41836 213240
rect 41590 212961 41642 212967
rect 41588 212926 41590 212935
rect 41642 212926 41644 212935
rect 41588 212861 41644 212870
rect 41782 212221 41834 212227
rect 41780 212186 41782 212195
rect 41834 212186 41836 212195
rect 41780 212121 41836 212130
rect 41782 211777 41834 211783
rect 41780 211742 41782 211751
rect 41834 211742 41836 211751
rect 41780 211677 41836 211686
rect 41590 211481 41642 211487
rect 41588 211446 41590 211455
rect 41642 211446 41644 211455
rect 41588 211381 41644 211390
rect 41782 210741 41834 210747
rect 41780 210706 41782 210715
rect 41834 210706 41836 210715
rect 41780 210641 41836 210650
rect 41780 210262 41836 210271
rect 43330 210229 43358 262113
rect 43426 254999 43454 297559
rect 43522 296735 43550 298077
rect 43510 296729 43562 296735
rect 43510 296671 43562 296677
rect 43508 266946 43564 266955
rect 43508 266881 43564 266890
rect 43522 265063 43550 266881
rect 43510 265057 43562 265063
rect 43510 264999 43562 265005
rect 43414 254993 43466 254999
rect 43414 254935 43466 254941
rect 43414 254475 43466 254481
rect 43414 254417 43466 254423
rect 43426 211783 43454 254417
rect 43414 211777 43466 211783
rect 43414 211719 43466 211725
rect 41780 210197 41782 210206
rect 41834 210197 41836 210206
rect 43318 210223 43370 210229
rect 41782 210165 41834 210171
rect 43318 210165 43370 210171
rect 41590 210001 41642 210007
rect 41588 209966 41590 209975
rect 41642 209966 41644 209975
rect 41588 209901 41644 209910
rect 43522 209415 43550 264999
rect 44086 264983 44138 264989
rect 44086 264925 44138 264931
rect 44098 263583 44126 264925
rect 44182 264909 44234 264915
rect 44182 264851 44234 264857
rect 44194 263657 44222 264851
rect 44182 263651 44234 263657
rect 44182 263593 44234 263599
rect 44086 263577 44138 263583
rect 44086 263519 44138 263525
rect 44578 246267 44606 805125
rect 44674 267103 44702 814819
rect 44758 813619 44810 813625
rect 44758 813561 44810 813567
rect 44770 275391 44798 813561
rect 44866 785579 44894 817261
rect 44950 816579 45002 816585
rect 44950 816521 45002 816527
rect 44962 789131 44990 816521
rect 44950 789125 45002 789131
rect 44950 789067 45002 789073
rect 44854 785573 44906 785579
rect 44854 785515 44906 785521
rect 47458 785431 47486 817927
rect 57718 800743 57770 800749
rect 57718 800685 57770 800691
rect 57622 800669 57674 800675
rect 57622 800611 57674 800617
rect 57634 789691 57662 800611
rect 57730 790875 57758 800685
rect 57716 790866 57772 790875
rect 57716 790801 57772 790810
rect 57620 789682 57676 789691
rect 57620 789617 57676 789626
rect 58198 789199 58250 789205
rect 58198 789141 58250 789147
rect 58210 788507 58238 789141
rect 58390 789125 58442 789131
rect 58390 789067 58442 789073
rect 58196 788498 58252 788507
rect 58196 788433 58252 788442
rect 58402 787323 58430 789067
rect 58388 787314 58444 787323
rect 58388 787249 58444 787258
rect 59158 785573 59210 785579
rect 59158 785515 59210 785521
rect 59636 785538 59692 785547
rect 47446 785425 47498 785431
rect 47446 785367 47498 785373
rect 59170 784955 59198 785515
rect 59636 785473 59692 785482
rect 59650 785431 59678 785473
rect 59638 785425 59690 785431
rect 59638 785367 59690 785373
rect 59156 784946 59212 784955
rect 59156 784881 59212 784890
rect 47542 774695 47594 774701
rect 47542 774637 47594 774643
rect 44854 773955 44906 773961
rect 44854 773897 44906 773903
rect 44866 742955 44894 773897
rect 44950 773363 45002 773369
rect 44950 773305 45002 773311
rect 44962 745175 44990 773305
rect 47446 762115 47498 762121
rect 47446 762057 47498 762063
rect 44950 745169 45002 745175
rect 44950 745111 45002 745117
rect 44854 742949 44906 742955
rect 44854 742891 44906 742897
rect 44854 730739 44906 730745
rect 44854 730681 44906 730687
rect 44866 699739 44894 730681
rect 44950 730369 45002 730375
rect 44950 730311 45002 730317
rect 44962 702625 44990 730311
rect 44950 702619 45002 702625
rect 44950 702561 45002 702567
rect 45236 702066 45292 702075
rect 45236 702001 45292 702010
rect 44854 699733 44906 699739
rect 44854 699675 44906 699681
rect 45250 698777 45278 702001
rect 45238 698771 45290 698777
rect 45238 698713 45290 698719
rect 45046 687227 45098 687233
rect 45046 687169 45098 687175
rect 44950 685377 45002 685383
rect 44950 685319 45002 685325
rect 44854 684193 44906 684199
rect 44854 684135 44906 684141
rect 44756 275382 44812 275391
rect 44756 275317 44812 275326
rect 44660 267094 44716 267103
rect 44660 267029 44716 267038
rect 44866 263107 44894 684135
rect 44962 266395 44990 685319
rect 45058 659409 45086 687169
rect 45046 659403 45098 659409
rect 45046 659345 45098 659351
rect 45046 596207 45098 596213
rect 45046 596149 45098 596155
rect 45058 274207 45086 596149
rect 45236 473110 45292 473119
rect 45236 473045 45292 473054
rect 45142 472479 45194 472485
rect 45142 472421 45194 472427
rect 45154 278351 45182 472421
rect 45140 278342 45196 278351
rect 45140 278277 45196 278286
rect 45250 276279 45278 473045
rect 45334 382051 45386 382057
rect 45334 381993 45386 381999
rect 45236 276270 45292 276279
rect 45236 276205 45292 276214
rect 45044 274198 45100 274207
rect 45044 274133 45100 274142
rect 45346 273615 45374 381993
rect 45430 330399 45482 330405
rect 45430 330341 45482 330347
rect 45332 273606 45388 273615
rect 45332 273541 45388 273550
rect 44950 266389 45002 266395
rect 44950 266331 45002 266337
rect 44852 263098 44908 263107
rect 44852 263033 44908 263042
rect 45442 246341 45470 330341
rect 45814 287183 45866 287189
rect 45814 287125 45866 287131
rect 45526 282373 45578 282379
rect 45526 282315 45578 282321
rect 45430 246335 45482 246341
rect 45430 246277 45482 246283
rect 44566 246261 44618 246267
rect 44566 246203 44618 246209
rect 44758 244929 44810 244935
rect 44758 244871 44810 244877
rect 44662 242783 44714 242789
rect 44662 242725 44714 242731
rect 44566 242709 44618 242715
rect 44566 242651 44618 242657
rect 41590 209409 41642 209415
rect 41588 209374 41590 209383
rect 43510 209409 43562 209415
rect 41642 209374 41644 209383
rect 43510 209351 43562 209357
rect 41588 209309 41644 209318
rect 25556 208486 25612 208495
rect 25556 208421 25612 208430
rect 25570 200059 25598 208421
rect 25748 208042 25804 208051
rect 25748 207977 25804 207986
rect 25652 206414 25708 206423
rect 25652 206349 25708 206358
rect 25556 200050 25612 200059
rect 25556 199985 25612 199994
rect 25666 199615 25694 206349
rect 25762 200503 25790 207977
rect 25844 207894 25900 207903
rect 25844 207829 25900 207838
rect 25858 200947 25886 207829
rect 41972 206266 42028 206275
rect 41972 206201 42028 206210
rect 41684 204046 41740 204055
rect 41684 203981 41740 203990
rect 41492 202566 41548 202575
rect 41492 202501 41548 202510
rect 41506 201497 41534 202501
rect 41588 202122 41644 202131
rect 41588 202057 41644 202066
rect 41494 201491 41546 201497
rect 41494 201433 41546 201439
rect 41494 200973 41546 200979
rect 25844 200938 25900 200947
rect 25844 200873 25900 200882
rect 41492 200938 41494 200947
rect 41546 200938 41548 200947
rect 41492 200873 41548 200882
rect 25748 200494 25804 200503
rect 25748 200429 25804 200438
rect 25652 199606 25708 199615
rect 25652 199541 25708 199550
rect 41602 198981 41630 202057
rect 41590 198975 41642 198981
rect 41590 198917 41642 198923
rect 41698 198907 41726 203981
rect 41780 203750 41836 203759
rect 41780 203685 41836 203694
rect 41686 198901 41738 198907
rect 41686 198843 41738 198849
rect 41794 198833 41822 203685
rect 41878 201713 41930 201719
rect 41876 201678 41878 201687
rect 41930 201678 41932 201687
rect 41876 201613 41932 201622
rect 41878 201417 41930 201423
rect 41876 201382 41878 201391
rect 41930 201382 41932 201391
rect 41876 201317 41932 201326
rect 41782 198827 41834 198833
rect 41782 198769 41834 198775
rect 41986 197427 42014 206201
rect 42934 201491 42986 201497
rect 42934 201433 42986 201439
rect 42742 198975 42794 198981
rect 42742 198917 42794 198923
rect 41974 197421 42026 197427
rect 41974 197363 42026 197369
rect 41974 197199 42026 197205
rect 41974 197141 42026 197147
rect 41986 196618 42014 197141
rect 41780 195314 41836 195323
rect 41780 195249 41836 195258
rect 41794 194805 41822 195249
rect 42070 193499 42122 193505
rect 42070 193441 42122 193447
rect 42082 192992 42110 193441
rect 42754 192247 42782 198917
rect 42838 198901 42890 198907
rect 42838 198843 42890 198849
rect 42850 193505 42878 198843
rect 42838 193499 42890 193505
rect 42838 193441 42890 193447
rect 42166 192241 42218 192247
rect 42166 192183 42218 192189
rect 42742 192241 42794 192247
rect 42742 192183 42794 192189
rect 42178 191769 42206 192183
rect 42070 191501 42122 191507
rect 42070 191443 42122 191449
rect 42082 191142 42110 191443
rect 42946 191063 42974 201433
rect 44578 201423 44606 242651
rect 44566 201417 44618 201423
rect 44566 201359 44618 201365
rect 44674 200979 44702 242725
rect 44770 201719 44798 244871
rect 44854 242857 44906 242863
rect 44854 242799 44906 242805
rect 44866 211487 44894 242799
rect 45538 212227 45566 282315
rect 45718 279487 45770 279493
rect 45718 279429 45770 279435
rect 45622 279413 45674 279419
rect 45622 279355 45674 279361
rect 45634 212967 45662 279355
rect 45730 213337 45758 279429
rect 45826 246415 45854 287125
rect 47458 255073 47486 762057
rect 47554 743029 47582 774637
rect 62038 771957 62090 771963
rect 62038 771899 62090 771905
rect 61846 771883 61898 771889
rect 61846 771825 61898 771831
rect 58678 757527 58730 757533
rect 58678 757469 58730 757475
rect 58690 747659 58718 757469
rect 58676 747650 58732 747659
rect 58676 747585 58732 747594
rect 54740 746022 54796 746031
rect 54646 745983 54698 745989
rect 54740 745957 54742 745966
rect 54646 745925 54698 745931
rect 54794 745957 54796 745966
rect 57622 745983 57674 745989
rect 54742 745925 54794 745931
rect 57622 745925 57674 745931
rect 54658 745883 54686 745925
rect 54644 745874 54700 745883
rect 54644 745809 54700 745818
rect 57634 745291 57662 745925
rect 59636 745430 59692 745439
rect 59636 745365 59692 745374
rect 59650 745323 59678 745365
rect 59638 745317 59690 745323
rect 57620 745282 57676 745291
rect 59638 745259 59690 745265
rect 57620 745217 57676 745226
rect 58198 745169 58250 745175
rect 58198 745111 58250 745117
rect 58210 744107 58238 745111
rect 58196 744098 58252 744107
rect 58196 744033 58252 744042
rect 47542 743023 47594 743029
rect 47542 742965 47594 742971
rect 59638 743023 59690 743029
rect 59638 742965 59690 742971
rect 59650 742923 59678 742965
rect 59734 742949 59786 742955
rect 59636 742914 59692 742923
rect 59734 742891 59786 742897
rect 59636 742849 59692 742858
rect 59746 741739 59774 742891
rect 59732 741730 59788 741739
rect 59732 741665 59788 741674
rect 47638 731479 47690 731485
rect 47638 731421 47690 731427
rect 47542 718751 47594 718757
rect 47542 718693 47594 718699
rect 47446 255067 47498 255073
rect 47446 255009 47498 255015
rect 47554 246563 47582 718693
rect 47650 699813 47678 731421
rect 59638 714311 59690 714317
rect 59638 714253 59690 714259
rect 59650 704443 59678 714253
rect 59636 704434 59692 704443
rect 59636 704369 59692 704378
rect 58774 702693 58826 702699
rect 58772 702658 58774 702667
rect 58826 702658 58828 702667
rect 58678 702619 58730 702625
rect 58772 702593 58828 702602
rect 58678 702561 58730 702567
rect 58690 700891 58718 702561
rect 58676 700882 58732 700891
rect 58676 700817 58732 700826
rect 47638 699807 47690 699813
rect 47638 699749 47690 699755
rect 59254 699807 59306 699813
rect 59254 699749 59306 699755
rect 58870 699733 58922 699739
rect 59266 699707 59294 699749
rect 58870 699675 58922 699681
rect 59252 699698 59308 699707
rect 58882 698523 58910 699675
rect 59252 699633 59308 699642
rect 58868 698514 58924 698523
rect 58868 698449 58924 698458
rect 50326 688263 50378 688269
rect 50326 688205 50378 688211
rect 47734 687523 47786 687529
rect 47734 687465 47786 687471
rect 47638 675535 47690 675541
rect 47638 675477 47690 675483
rect 47650 246637 47678 675477
rect 47746 656597 47774 687465
rect 50338 656671 50366 688205
rect 59638 671095 59690 671101
rect 59638 671037 59690 671043
rect 59650 661227 59678 671037
rect 59636 661218 59692 661227
rect 59636 661153 59692 661162
rect 58774 659477 58826 659483
rect 58772 659442 58774 659451
rect 58826 659442 58828 659451
rect 58678 659403 58730 659409
rect 58772 659377 58828 659386
rect 58678 659345 58730 659351
rect 58690 657675 58718 659345
rect 58676 657666 58732 657675
rect 58676 657601 58732 657610
rect 50326 656665 50378 656671
rect 50326 656607 50378 656613
rect 58198 656665 58250 656671
rect 58198 656607 58250 656613
rect 47734 656591 47786 656597
rect 47734 656533 47786 656539
rect 58210 656491 58238 656607
rect 58390 656591 58442 656597
rect 58390 656533 58442 656539
rect 58196 656482 58252 656491
rect 58196 656417 58252 656426
rect 58402 655307 58430 656533
rect 58388 655298 58444 655307
rect 58388 655233 58444 655242
rect 50326 644899 50378 644905
rect 50326 644841 50378 644847
rect 47830 644307 47882 644313
rect 47830 644249 47882 644255
rect 47734 632319 47786 632325
rect 47734 632261 47786 632267
rect 47638 246631 47690 246637
rect 47638 246573 47690 246579
rect 47542 246557 47594 246563
rect 47542 246499 47594 246505
rect 47746 246489 47774 632261
rect 47842 613381 47870 644249
rect 47926 644011 47978 644017
rect 47926 643953 47978 643959
rect 47938 616341 47966 643953
rect 48022 622107 48074 622113
rect 48022 622049 48074 622055
rect 47926 616335 47978 616341
rect 47926 616277 47978 616283
rect 48034 616267 48062 622049
rect 48022 616261 48074 616267
rect 48022 616203 48074 616209
rect 50338 613455 50366 644841
rect 58966 624031 59018 624037
rect 58966 623973 59018 623979
rect 58978 618011 59006 623973
rect 58964 618002 59020 618011
rect 58964 617937 59020 617946
rect 58198 616409 58250 616415
rect 58198 616351 58250 616357
rect 58210 615643 58238 616351
rect 58966 616335 59018 616341
rect 58966 616277 59018 616283
rect 58196 615634 58252 615643
rect 58196 615569 58252 615578
rect 58978 614459 59006 616277
rect 59638 616261 59690 616267
rect 59636 616226 59638 616235
rect 59690 616226 59692 616235
rect 59636 616161 59692 616170
rect 58964 614450 59020 614459
rect 58964 614385 59020 614394
rect 50326 613449 50378 613455
rect 50326 613391 50378 613397
rect 59638 613449 59690 613455
rect 59638 613391 59690 613397
rect 47830 613375 47882 613381
rect 47830 613317 47882 613323
rect 59542 613375 59594 613381
rect 59542 613317 59594 613323
rect 59554 612091 59582 613317
rect 59650 613275 59678 613391
rect 59636 613266 59692 613275
rect 59636 613201 59692 613210
rect 59540 612082 59596 612091
rect 59540 612017 59596 612026
rect 50326 601683 50378 601689
rect 50326 601625 50378 601631
rect 47830 601387 47882 601393
rect 47830 601329 47882 601335
rect 47842 570165 47870 601329
rect 47926 600795 47978 600801
rect 47926 600737 47978 600743
rect 47938 573125 47966 600737
rect 48022 579335 48074 579341
rect 48022 579277 48074 579283
rect 47926 573119 47978 573125
rect 47926 573061 47978 573067
rect 48034 573051 48062 579277
rect 48022 573045 48074 573051
rect 48022 572987 48074 572993
rect 50338 570239 50366 601625
rect 56086 587549 56138 587555
rect 56086 587491 56138 587497
rect 50326 570233 50378 570239
rect 50326 570175 50378 570181
rect 47830 570159 47882 570165
rect 47830 570101 47882 570107
rect 50326 524353 50378 524359
rect 50326 524295 50378 524301
rect 47830 524279 47882 524285
rect 47830 524221 47882 524227
rect 47842 475593 47870 524221
rect 50338 476111 50366 524295
rect 50326 476105 50378 476111
rect 50326 476047 50378 476053
rect 47830 475587 47882 475593
rect 47830 475529 47882 475535
rect 47830 463599 47882 463605
rect 47830 463541 47882 463547
rect 47842 255147 47870 463541
rect 53206 426895 53258 426901
rect 53206 426837 53258 426843
rect 50326 426525 50378 426531
rect 50326 426467 50378 426473
rect 48022 426007 48074 426013
rect 48022 425949 48074 425955
rect 47926 414315 47978 414321
rect 47926 414257 47978 414263
rect 47830 255141 47882 255147
rect 47830 255083 47882 255089
rect 47938 254999 47966 414257
rect 48034 400187 48062 425949
rect 50338 400261 50366 426467
rect 53218 400335 53246 426837
rect 53206 400329 53258 400335
rect 53206 400271 53258 400277
rect 50326 400255 50378 400261
rect 50326 400197 50378 400203
rect 48022 400181 48074 400187
rect 48022 400123 48074 400129
rect 53206 385973 53258 385979
rect 53206 385915 53258 385921
rect 50326 385307 50378 385313
rect 50326 385249 50378 385255
rect 48118 385011 48170 385017
rect 48118 384953 48170 384959
rect 48022 373541 48074 373547
rect 48022 373483 48074 373489
rect 47926 254993 47978 254999
rect 47926 254935 47978 254941
rect 48034 254925 48062 373483
rect 48130 357045 48158 384953
rect 48118 357039 48170 357045
rect 48118 356981 48170 356987
rect 50338 356971 50366 385249
rect 53218 357119 53246 385915
rect 53206 357113 53258 357119
rect 53206 357055 53258 357061
rect 50326 356965 50378 356971
rect 50326 356907 50378 356913
rect 53206 342831 53258 342837
rect 53206 342773 53258 342779
rect 50326 342313 50378 342319
rect 50326 342255 50378 342261
rect 48118 341795 48170 341801
rect 48118 341737 48170 341743
rect 48130 313829 48158 341737
rect 48118 313823 48170 313829
rect 48118 313765 48170 313771
rect 50338 313755 50366 342255
rect 53218 313903 53246 342773
rect 53206 313897 53258 313903
rect 53206 313839 53258 313845
rect 50326 313749 50378 313755
rect 50326 313691 50378 313697
rect 51766 299171 51818 299177
rect 51766 299113 51818 299119
rect 48214 290957 48266 290963
rect 48214 290899 48266 290905
rect 48118 282595 48170 282601
rect 48118 282537 48170 282543
rect 48022 254919 48074 254925
rect 48022 254861 48074 254867
rect 47734 246483 47786 246489
rect 47734 246425 47786 246431
rect 45814 246409 45866 246415
rect 45814 246351 45866 246357
rect 45718 213331 45770 213337
rect 45718 213273 45770 213279
rect 45622 212961 45674 212967
rect 45622 212903 45674 212909
rect 45526 212221 45578 212227
rect 45526 212163 45578 212169
rect 44854 211481 44906 211487
rect 44854 211423 44906 211429
rect 44758 201713 44810 201719
rect 44758 201655 44810 201661
rect 44662 200973 44714 200979
rect 44662 200915 44714 200921
rect 43030 198827 43082 198833
rect 43030 198769 43082 198775
rect 43042 191507 43070 198769
rect 43030 191501 43082 191507
rect 43030 191443 43082 191449
rect 42166 191057 42218 191063
rect 42166 190999 42218 191005
rect 42934 191057 42986 191063
rect 42934 190999 42986 191005
rect 42178 190476 42206 190999
rect 41780 190134 41836 190143
rect 41780 190069 41836 190078
rect 41794 189929 41822 190069
rect 41876 187914 41932 187923
rect 41876 187849 41932 187858
rect 41890 187442 41918 187849
rect 42164 187174 42220 187183
rect 42164 187109 42220 187118
rect 42178 186776 42206 187109
rect 41780 186434 41836 186443
rect 41780 186369 41836 186378
rect 41794 186184 41822 186369
rect 41780 185842 41836 185851
rect 41780 185777 41836 185786
rect 41794 185592 41822 185777
rect 41780 184214 41836 184223
rect 41780 184149 41836 184158
rect 41794 183742 41822 184149
rect 41780 183474 41836 183483
rect 41780 183409 41836 183418
rect 41794 183121 41822 183409
rect 42068 183030 42124 183039
rect 42068 182965 42124 182974
rect 42082 182484 42110 182965
rect 48130 182257 48158 282537
rect 48226 268615 48254 290899
rect 51778 289557 51806 299113
rect 53302 293917 53354 293923
rect 53302 293859 53354 293865
rect 51766 289551 51818 289557
rect 51766 289493 51818 289499
rect 50326 288071 50378 288077
rect 50326 288013 50378 288019
rect 48214 268609 48266 268615
rect 48214 268551 48266 268557
rect 50338 221773 50366 288013
rect 53206 285185 53258 285191
rect 53206 285127 53258 285133
rect 50420 275234 50476 275243
rect 50420 275169 50476 275178
rect 50326 221767 50378 221773
rect 50326 221709 50378 221715
rect 50434 210007 50462 275169
rect 50612 275086 50668 275095
rect 50612 275021 50668 275030
rect 50626 210747 50654 275021
rect 53218 255443 53246 285127
rect 53314 276459 53342 293859
rect 53302 276453 53354 276459
rect 53302 276395 53354 276401
rect 53206 255437 53258 255443
rect 53206 255379 53258 255385
rect 56098 252039 56126 587491
rect 58966 584737 59018 584743
rect 58966 584679 59018 584685
rect 58978 574795 59006 584679
rect 58964 574786 59020 574795
rect 58964 574721 59020 574730
rect 58198 573193 58250 573199
rect 58198 573135 58250 573141
rect 58210 572427 58238 573135
rect 58966 573119 59018 573125
rect 58966 573061 59018 573067
rect 58196 572418 58252 572427
rect 58196 572353 58252 572362
rect 58978 571243 59006 573061
rect 59638 573045 59690 573051
rect 59636 573010 59638 573019
rect 59690 573010 59692 573019
rect 59636 572945 59692 572954
rect 58964 571234 59020 571243
rect 58964 571169 59020 571178
rect 59350 570233 59402 570239
rect 59350 570175 59402 570181
rect 59362 570059 59390 570175
rect 59542 570159 59594 570165
rect 59542 570101 59594 570107
rect 59348 570050 59404 570059
rect 59348 569985 59404 569994
rect 59554 568875 59582 570101
rect 59540 568866 59596 568875
rect 59540 568801 59596 568810
rect 57718 541595 57770 541601
rect 57718 541537 57770 541543
rect 57622 541521 57674 541527
rect 57622 541463 57674 541469
rect 57634 530543 57662 541463
rect 57730 531727 57758 541537
rect 57716 531718 57772 531727
rect 57716 531653 57772 531662
rect 57620 530534 57676 530543
rect 57620 530469 57676 530478
rect 58198 529977 58250 529983
rect 58198 529919 58250 529925
rect 58210 529359 58238 529919
rect 58196 529350 58252 529359
rect 58196 529285 58252 529294
rect 58964 527130 59020 527139
rect 58964 527065 59020 527074
rect 58580 525946 58636 525955
rect 58580 525881 58636 525890
rect 58594 524359 58622 525881
rect 58582 524353 58634 524359
rect 58582 524295 58634 524301
rect 58978 472411 59006 527065
rect 59348 524762 59404 524771
rect 59348 524697 59404 524706
rect 59362 524285 59390 524697
rect 59350 524279 59402 524285
rect 59350 524221 59402 524227
rect 58966 472405 59018 472411
rect 58966 472347 59018 472353
rect 58486 406101 58538 406107
rect 58486 406043 58538 406049
rect 58498 404151 58526 406043
rect 58484 404142 58540 404151
rect 58484 404077 58540 404086
rect 59350 402623 59402 402629
rect 59350 402565 59402 402571
rect 59362 402375 59390 402565
rect 59348 402366 59404 402375
rect 59348 402301 59404 402310
rect 57716 400590 57772 400599
rect 57716 400525 57772 400534
rect 57730 394563 57758 400525
rect 59734 400329 59786 400335
rect 59734 400271 59786 400277
rect 59542 400255 59594 400261
rect 59542 400197 59594 400203
rect 59554 398231 59582 400197
rect 59638 400181 59690 400187
rect 59638 400123 59690 400129
rect 59650 400007 59678 400123
rect 59636 399998 59692 400007
rect 59636 399933 59692 399942
rect 59746 399415 59774 400271
rect 59732 399406 59788 399415
rect 59732 399341 59788 399350
rect 59540 398222 59596 398231
rect 59540 398157 59596 398166
rect 57718 394557 57770 394563
rect 57718 394499 57770 394505
rect 59254 361997 59306 362003
rect 59254 361939 59306 361945
rect 59266 360935 59294 361939
rect 59252 360926 59308 360935
rect 59252 360861 59308 360870
rect 59158 359999 59210 360005
rect 59158 359941 59210 359947
rect 59170 359751 59198 359941
rect 59156 359742 59212 359751
rect 59156 359677 59212 359686
rect 57620 357522 57676 357531
rect 57620 357457 57676 357466
rect 57634 351347 57662 357457
rect 58198 357113 58250 357119
rect 58198 357055 58250 357061
rect 58210 356199 58238 357055
rect 59638 357039 59690 357045
rect 59638 356981 59690 356987
rect 58582 356965 58634 356971
rect 58582 356907 58634 356913
rect 58196 356190 58252 356199
rect 58196 356125 58252 356134
rect 58594 355015 58622 356907
rect 59650 356791 59678 356981
rect 59636 356782 59692 356791
rect 59636 356717 59692 356726
rect 58580 355006 58636 355015
rect 58580 354941 58636 354950
rect 57622 351341 57674 351347
rect 57622 351283 57674 351289
rect 58486 319669 58538 319675
rect 58486 319611 58538 319617
rect 58498 317719 58526 319611
rect 58484 317710 58540 317719
rect 58484 317645 58540 317654
rect 59158 316783 59210 316789
rect 59158 316725 59210 316731
rect 59170 316535 59198 316725
rect 59156 316526 59212 316535
rect 59156 316461 59212 316470
rect 59348 314158 59404 314167
rect 59348 314093 59404 314102
rect 58198 313897 58250 313903
rect 58198 313839 58250 313845
rect 58210 312983 58238 313839
rect 58196 312974 58252 312983
rect 58196 312909 58252 312918
rect 59362 308131 59390 314093
rect 59638 313823 59690 313829
rect 59638 313765 59690 313771
rect 59650 313575 59678 313765
rect 59734 313749 59786 313755
rect 59734 313691 59786 313697
rect 59636 313566 59692 313575
rect 59636 313501 59692 313510
rect 59746 311799 59774 313691
rect 59732 311790 59788 311799
rect 59732 311725 59788 311734
rect 59350 308125 59402 308131
rect 59350 308067 59402 308073
rect 60214 299615 60266 299621
rect 60214 299557 60266 299563
rect 59636 295214 59692 295223
rect 59636 295149 59692 295158
rect 59650 293923 59678 295149
rect 59638 293917 59690 293923
rect 59638 293859 59690 293865
rect 56278 293843 56330 293849
rect 56278 293785 56330 293791
rect 56182 282299 56234 282305
rect 56182 282241 56234 282247
rect 56194 253519 56222 282241
rect 56290 273573 56318 293785
rect 58774 293769 58826 293775
rect 58774 293711 58826 293717
rect 58388 292846 58444 292855
rect 58388 292781 58444 292790
rect 58402 290963 58430 292781
rect 58786 292707 58814 293711
rect 58772 292698 58828 292707
rect 58772 292633 58828 292642
rect 60226 291523 60254 299557
rect 60308 294030 60364 294039
rect 60308 293965 60364 293974
rect 60322 293849 60350 293965
rect 60310 293843 60362 293849
rect 60310 293785 60362 293791
rect 60212 291514 60268 291523
rect 60212 291449 60268 291458
rect 58390 290957 58442 290963
rect 58390 290899 58442 290905
rect 58004 289590 58060 289599
rect 58004 289525 58006 289534
rect 58058 289525 58060 289534
rect 58006 289493 58058 289499
rect 59636 288110 59692 288119
rect 59636 288045 59638 288054
rect 59690 288045 59692 288054
rect 59638 288013 59690 288019
rect 58964 286926 59020 286935
rect 58964 286861 59020 286870
rect 58978 285191 59006 286861
rect 59060 285742 59116 285751
rect 59060 285677 59116 285686
rect 58966 285185 59018 285191
rect 58966 285127 59018 285133
rect 57620 284558 57676 284567
rect 57620 284493 57676 284502
rect 57634 282305 57662 284493
rect 58964 282486 59020 282495
rect 58964 282421 59020 282430
rect 58978 282379 59006 282421
rect 58966 282373 59018 282379
rect 58966 282315 59018 282321
rect 57622 282299 57674 282305
rect 57622 282241 57674 282247
rect 56278 273567 56330 273573
rect 56278 273509 56330 273515
rect 59074 256405 59102 285677
rect 59636 283374 59692 283383
rect 59636 283309 59692 283318
rect 59650 282601 59678 283309
rect 59638 282595 59690 282601
rect 59638 282537 59690 282543
rect 59540 281006 59596 281015
rect 59540 280941 59596 280950
rect 59348 279822 59404 279831
rect 59348 279757 59404 279766
rect 59362 279419 59390 279757
rect 59554 279493 59582 280941
rect 59542 279487 59594 279493
rect 59542 279429 59594 279435
rect 59350 279413 59402 279419
rect 59350 279355 59402 279361
rect 61858 266363 61886 771825
rect 61942 642531 61994 642537
rect 61942 642473 61994 642479
rect 61954 278203 61982 642473
rect 61940 278194 61996 278203
rect 61940 278129 61996 278138
rect 62050 266659 62078 771899
rect 62230 728741 62282 728747
rect 62230 728683 62282 728689
rect 62132 537046 62188 537055
rect 62132 536981 62188 536990
rect 62146 276131 62174 536981
rect 62132 276122 62188 276131
rect 62132 276057 62188 276066
rect 62036 266650 62092 266659
rect 62036 266585 62092 266594
rect 62242 266511 62270 728683
rect 62422 728667 62474 728673
rect 62422 728609 62474 728615
rect 62326 437847 62378 437853
rect 62326 437789 62378 437795
rect 62338 277907 62366 437789
rect 62324 277898 62380 277907
rect 62324 277833 62380 277842
rect 62434 266807 62462 728609
rect 62518 420531 62570 420537
rect 62518 420473 62570 420479
rect 62530 270655 62558 420473
rect 64724 386382 64780 386391
rect 64724 386317 64780 386326
rect 62612 343166 62668 343175
rect 62612 343101 62668 343110
rect 62626 278055 62654 343101
rect 62806 300947 62858 300953
rect 62806 300889 62858 300895
rect 62612 278046 62668 278055
rect 62612 277981 62668 277990
rect 62818 277759 62846 300889
rect 62998 298135 63050 298141
rect 62998 298077 63050 298083
rect 62804 277750 62860 277759
rect 62804 277685 62860 277694
rect 63010 277611 63038 298077
rect 62996 277602 63052 277611
rect 62996 277537 63052 277546
rect 64738 277463 64766 386317
rect 408322 278309 408624 278328
rect 314902 278303 314954 278309
rect 314902 278245 314954 278251
rect 408310 278303 408624 278309
rect 408362 278300 408624 278303
rect 408310 278245 408362 278251
rect 64724 277454 64780 277463
rect 64724 277389 64780 277398
rect 62516 270646 62572 270655
rect 62516 270581 62572 270590
rect 65890 269323 65918 278018
rect 65876 269314 65932 269323
rect 67042 269281 67070 278018
rect 68290 273277 68318 278018
rect 68278 273271 68330 273277
rect 68278 273213 68330 273219
rect 69442 269619 69470 278018
rect 70594 272135 70622 278018
rect 70580 272126 70636 272135
rect 70580 272061 70636 272070
rect 69428 269610 69484 269619
rect 69428 269545 69484 269554
rect 71746 269471 71774 278018
rect 72994 272283 73022 278018
rect 72980 272274 73036 272283
rect 72980 272209 73036 272218
rect 71732 269462 71788 269471
rect 71732 269397 71788 269406
rect 74146 269355 74174 278018
rect 75298 271649 75326 278018
rect 76546 272315 76574 278018
rect 77698 276494 77726 278018
rect 77602 276466 77726 276494
rect 76534 272309 76586 272315
rect 76534 272251 76586 272257
rect 75286 271643 75338 271649
rect 75286 271585 75338 271591
rect 77602 269767 77630 276466
rect 78850 272431 78878 278018
rect 80112 278004 80606 278032
rect 78836 272422 78892 272431
rect 78836 272357 78892 272366
rect 77686 271643 77738 271649
rect 77686 271585 77738 271591
rect 77588 269758 77644 269767
rect 77588 269693 77644 269702
rect 74134 269349 74186 269355
rect 74134 269291 74186 269297
rect 65876 269249 65932 269258
rect 67030 269275 67082 269281
rect 67030 269217 67082 269223
rect 62420 266798 62476 266807
rect 62420 266733 62476 266742
rect 62228 266502 62284 266511
rect 62228 266437 62284 266446
rect 61844 266354 61900 266363
rect 61844 266289 61900 266298
rect 59062 256399 59114 256405
rect 59062 256341 59114 256347
rect 56182 253513 56234 253519
rect 56182 253455 56234 253461
rect 56086 252033 56138 252039
rect 56086 251975 56138 251981
rect 77698 249301 77726 271585
rect 77686 249295 77738 249301
rect 77686 249237 77738 249243
rect 80578 249227 80606 278004
rect 81250 269503 81278 278018
rect 81238 269497 81290 269503
rect 81238 269439 81290 269445
rect 82402 269429 82430 278018
rect 83650 269651 83678 278018
rect 84802 272241 84830 278018
rect 84790 272235 84842 272241
rect 84790 272177 84842 272183
rect 85954 271131 85982 278018
rect 86326 272235 86378 272241
rect 86326 272177 86378 272183
rect 85942 271125 85994 271131
rect 85942 271067 85994 271073
rect 83638 269645 83690 269651
rect 83638 269587 83690 269593
rect 82390 269423 82442 269429
rect 82390 269365 82442 269371
rect 80566 249221 80618 249227
rect 80566 249163 80618 249169
rect 86338 249153 86366 272177
rect 87202 269577 87230 278018
rect 88354 272579 88382 278018
rect 88340 272570 88396 272579
rect 88340 272505 88396 272514
rect 89506 271575 89534 278018
rect 89494 271569 89546 271575
rect 89494 271511 89546 271517
rect 90658 269725 90686 278018
rect 91906 272727 91934 278018
rect 91892 272718 91948 272727
rect 91892 272653 91948 272662
rect 92086 271569 92138 271575
rect 92086 271511 92138 271517
rect 90646 269719 90698 269725
rect 90646 269661 90698 269667
rect 87190 269571 87242 269577
rect 87190 269513 87242 269519
rect 92098 252261 92126 271511
rect 93058 269799 93086 278018
rect 94210 270761 94238 278018
rect 94198 270755 94250 270761
rect 94198 270697 94250 270703
rect 94966 270755 95018 270761
rect 94966 270697 95018 270703
rect 93046 269793 93098 269799
rect 93046 269735 93098 269741
rect 92086 252255 92138 252261
rect 92086 252197 92138 252203
rect 94978 249449 95006 270697
rect 95458 269873 95486 278018
rect 96610 272611 96638 278018
rect 97776 278004 97886 278032
rect 96598 272605 96650 272611
rect 96598 272547 96650 272553
rect 95446 269867 95498 269873
rect 95446 269809 95498 269815
rect 97858 252113 97886 278004
rect 99010 272389 99038 278018
rect 98998 272383 99050 272389
rect 98998 272325 99050 272331
rect 100162 269947 100190 278018
rect 101314 270761 101342 278018
rect 101302 270755 101354 270761
rect 101302 270697 101354 270703
rect 102562 270095 102590 278018
rect 103714 272537 103742 278018
rect 103702 272531 103754 272537
rect 103702 272473 103754 272479
rect 104866 272241 104894 278018
rect 106114 272463 106142 278018
rect 106678 272605 106730 272611
rect 106678 272547 106730 272553
rect 106102 272457 106154 272463
rect 106102 272399 106154 272405
rect 106690 272315 106718 272547
rect 106678 272309 106730 272315
rect 106678 272251 106730 272257
rect 104854 272235 104906 272241
rect 104854 272177 104906 272183
rect 106486 272235 106538 272241
rect 106486 272177 106538 272183
rect 103606 270755 103658 270761
rect 103606 270697 103658 270703
rect 102550 270089 102602 270095
rect 102550 270031 102602 270037
rect 100150 269941 100202 269947
rect 100150 269883 100202 269889
rect 97846 252107 97898 252113
rect 97846 252049 97898 252055
rect 94966 249443 95018 249449
rect 94966 249385 95018 249391
rect 86326 249147 86378 249153
rect 86326 249089 86378 249095
rect 103618 246785 103646 270697
rect 106498 252335 106526 272177
rect 107266 270021 107294 278018
rect 108418 273425 108446 278018
rect 108406 273419 108458 273425
rect 108406 273361 108458 273367
rect 109366 273419 109418 273425
rect 109366 273361 109418 273367
rect 107254 270015 107306 270021
rect 107254 269957 107306 269963
rect 106486 252329 106538 252335
rect 106486 252271 106538 252277
rect 109378 252187 109406 273361
rect 109570 270169 109598 278018
rect 110818 272611 110846 278018
rect 111984 278004 112286 278032
rect 110806 272605 110858 272611
rect 110806 272547 110858 272553
rect 109558 270163 109610 270169
rect 109558 270105 109610 270111
rect 109366 252181 109418 252187
rect 109366 252123 109418 252129
rect 103606 246779 103658 246785
rect 103606 246721 103658 246727
rect 112258 246711 112286 278004
rect 113122 272685 113150 278018
rect 113110 272679 113162 272685
rect 113110 272621 113162 272627
rect 114370 270243 114398 278018
rect 115522 270761 115550 278018
rect 116674 272759 116702 278018
rect 116662 272753 116714 272759
rect 116662 272695 116714 272701
rect 115510 270755 115562 270761
rect 115510 270697 115562 270703
rect 117922 270317 117950 278018
rect 119074 272093 119102 278018
rect 120226 272833 120254 278018
rect 120214 272827 120266 272833
rect 120214 272769 120266 272775
rect 119062 272087 119114 272093
rect 119062 272029 119114 272035
rect 120886 272087 120938 272093
rect 120886 272029 120938 272035
rect 118006 270755 118058 270761
rect 118006 270697 118058 270703
rect 117910 270311 117962 270317
rect 117910 270253 117962 270259
rect 114358 270237 114410 270243
rect 114358 270179 114410 270185
rect 118018 249375 118046 270697
rect 120898 249967 120926 272029
rect 121474 270391 121502 278018
rect 122626 273425 122654 278018
rect 123778 276494 123806 278018
rect 123682 276466 123806 276494
rect 122614 273419 122666 273425
rect 122614 273361 122666 273367
rect 123682 272907 123710 276466
rect 123766 273419 123818 273425
rect 123766 273361 123818 273367
rect 123670 272901 123722 272907
rect 123670 272843 123722 272849
rect 121462 270385 121514 270391
rect 121462 270327 121514 270333
rect 120886 249961 120938 249967
rect 120886 249903 120938 249909
rect 123778 249597 123806 273361
rect 125026 272981 125054 278018
rect 126192 278004 126686 278032
rect 125014 272975 125066 272981
rect 125014 272917 125066 272923
rect 123766 249591 123818 249597
rect 123766 249533 123818 249539
rect 126658 249523 126686 278004
rect 127330 273129 127358 278018
rect 127318 273123 127370 273129
rect 127318 273065 127370 273071
rect 128482 273055 128510 278018
rect 128470 273049 128522 273055
rect 128470 272991 128522 272997
rect 129730 271649 129758 278018
rect 130882 273499 130910 278018
rect 130870 273493 130922 273499
rect 130870 273435 130922 273441
rect 132034 273203 132062 278018
rect 132022 273197 132074 273203
rect 132022 273139 132074 273145
rect 129718 271643 129770 271649
rect 129718 271585 129770 271591
rect 132406 271643 132458 271649
rect 132406 271585 132458 271591
rect 132418 249893 132446 271585
rect 133282 270761 133310 278018
rect 133270 270755 133322 270761
rect 133270 270697 133322 270703
rect 134434 270465 134462 278018
rect 135586 273351 135614 278018
rect 135574 273345 135626 273351
rect 135574 273287 135626 273293
rect 136834 270761 136862 278018
rect 135286 270755 135338 270761
rect 135286 270697 135338 270703
rect 136822 270755 136874 270761
rect 136822 270697 136874 270703
rect 134422 270459 134474 270465
rect 134422 270401 134474 270407
rect 132406 249887 132458 249893
rect 132406 249829 132458 249835
rect 135298 249819 135326 270697
rect 137986 270539 138014 278018
rect 138166 270755 138218 270761
rect 138166 270697 138218 270703
rect 137974 270533 138026 270539
rect 137974 270475 138026 270481
rect 135286 249813 135338 249819
rect 135286 249755 135338 249761
rect 138178 249745 138206 270697
rect 139138 269915 139166 278018
rect 140400 278004 141086 278032
rect 139124 269906 139180 269915
rect 139124 269841 139180 269850
rect 138166 249739 138218 249745
rect 138166 249681 138218 249687
rect 141058 249671 141086 278004
rect 141538 270613 141566 278018
rect 142690 273425 142718 278018
rect 142678 273419 142730 273425
rect 142678 273361 142730 273367
rect 142486 273271 142538 273277
rect 142486 273213 142538 273219
rect 141526 270607 141578 270613
rect 141526 270549 141578 270555
rect 141046 249665 141098 249671
rect 141046 249607 141098 249613
rect 126646 249517 126698 249523
rect 126646 249459 126698 249465
rect 118006 249369 118058 249375
rect 118006 249311 118058 249317
rect 112246 246705 112298 246711
rect 112246 246647 112298 246653
rect 142498 216014 142526 273213
rect 142582 242635 142634 242641
rect 142582 242577 142634 242583
rect 142594 236174 142622 242577
rect 142594 236146 143102 236174
rect 143074 218887 143102 236146
rect 143062 218881 143114 218887
rect 143062 218823 143114 218829
rect 142498 215986 143102 216014
rect 50614 210741 50666 210747
rect 50614 210683 50666 210689
rect 50422 210001 50474 210007
rect 50422 209943 50474 209949
rect 143074 201571 143102 215986
rect 143062 201565 143114 201571
rect 143062 201507 143114 201513
rect 143938 190101 143966 278018
rect 145090 269207 145118 278018
rect 146242 270687 146270 278018
rect 147394 271797 147422 278018
rect 147382 271791 147434 271797
rect 147382 271733 147434 271739
rect 146230 270681 146282 270687
rect 146230 270623 146282 270629
rect 145078 269201 145130 269207
rect 145078 269143 145130 269149
rect 148642 269133 148670 278018
rect 149686 271791 149738 271797
rect 149686 271733 149738 271739
rect 148630 269127 148682 269133
rect 148630 269069 148682 269075
rect 145462 252255 145514 252261
rect 145462 252197 145514 252203
rect 145366 249295 145418 249301
rect 145366 249237 145418 249243
rect 143926 190095 143978 190101
rect 143926 190037 143978 190043
rect 42166 182251 42218 182257
rect 42166 182193 42218 182199
rect 48118 182251 48170 182257
rect 48118 182193 48170 182199
rect 42178 181925 42206 182193
rect 145378 175671 145406 249237
rect 145474 178557 145502 252197
rect 145654 249961 145706 249967
rect 145654 249903 145706 249909
rect 145558 245003 145610 245009
rect 145558 244945 145610 244951
rect 145462 178551 145514 178557
rect 145462 178493 145514 178499
rect 145366 175665 145418 175671
rect 145366 175607 145418 175613
rect 145570 175597 145598 244945
rect 145666 184329 145694 249903
rect 145750 244855 145802 244861
rect 145750 244797 145802 244803
rect 145762 221773 145790 244797
rect 148340 244598 148396 244607
rect 148340 244533 148396 244542
rect 148244 239714 148300 239723
rect 148244 239649 148300 239658
rect 147860 232314 147916 232323
rect 147860 232249 147916 232258
rect 147874 232207 147902 232249
rect 147862 232201 147914 232207
rect 147862 232143 147914 232149
rect 146900 229946 146956 229955
rect 146900 229881 146956 229890
rect 146914 229839 146942 229881
rect 146902 229833 146954 229839
rect 146902 229775 146954 229781
rect 147092 226394 147148 226403
rect 147092 226329 147148 226338
rect 147106 224807 147134 226329
rect 147094 224801 147146 224807
rect 147094 224743 147146 224749
rect 145750 221767 145802 221773
rect 145750 221709 145802 221715
rect 147284 221510 147340 221519
rect 147284 221445 147340 221454
rect 147298 220811 147326 221445
rect 147286 220805 147338 220811
rect 147286 220747 147338 220753
rect 147284 214110 147340 214119
rect 147284 214045 147286 214054
rect 147338 214045 147340 214054
rect 147286 214013 147338 214019
rect 146900 212926 146956 212935
rect 146900 212861 146902 212870
rect 146954 212861 146956 212870
rect 146902 212829 146954 212835
rect 147092 211742 147148 211751
rect 147092 211677 147148 211686
rect 147106 211339 147134 211677
rect 147094 211333 147146 211339
rect 147094 211275 147146 211281
rect 147476 210410 147532 210419
rect 147476 210345 147478 210354
rect 147530 210345 147532 210354
rect 147478 210313 147530 210319
rect 146900 209226 146956 209235
rect 146900 209161 146956 209170
rect 146914 207417 146942 209161
rect 147188 208042 147244 208051
rect 147188 207977 147244 207986
rect 147202 207935 147230 207977
rect 147190 207929 147242 207935
rect 147190 207871 147242 207877
rect 146902 207411 146954 207417
rect 146902 207353 146954 207359
rect 147092 206414 147148 206423
rect 147092 206349 147148 206358
rect 147106 204605 147134 206349
rect 147094 204599 147146 204605
rect 147094 204541 147146 204547
rect 147476 199606 147532 199615
rect 147476 199541 147532 199550
rect 147490 198833 147518 199541
rect 147478 198827 147530 198833
rect 147478 198769 147530 198775
rect 147380 191022 147436 191031
rect 147380 190957 147436 190966
rect 147394 190249 147422 190957
rect 147382 190243 147434 190249
rect 147382 190185 147434 190191
rect 145654 184323 145706 184329
rect 145654 184265 145706 184271
rect 147764 176518 147820 176527
rect 147764 176453 147820 176462
rect 147778 176041 147806 176453
rect 147766 176035 147818 176041
rect 147766 175977 147818 175983
rect 145558 175591 145610 175597
rect 145558 175533 145610 175539
rect 148258 169825 148286 239649
rect 148354 172785 148382 244533
rect 148724 243414 148780 243423
rect 148724 243349 148780 243358
rect 148532 242082 148588 242091
rect 148532 242017 148588 242026
rect 148436 238530 148492 238539
rect 148436 238465 148492 238474
rect 148342 172779 148394 172785
rect 148342 172721 148394 172727
rect 148450 169899 148478 238465
rect 148546 172563 148574 242017
rect 148628 233646 148684 233655
rect 148628 233581 148684 233590
rect 148534 172557 148586 172563
rect 148534 172499 148586 172505
rect 148438 169893 148490 169899
rect 148438 169835 148490 169841
rect 148246 169819 148298 169825
rect 148246 169761 148298 169767
rect 148532 169118 148588 169127
rect 148532 169053 148588 169062
rect 148340 168082 148396 168091
rect 148340 168017 148396 168026
rect 148244 164382 148300 164391
rect 148244 164317 148300 164326
rect 147476 159498 147532 159507
rect 147476 159433 147532 159442
rect 147490 158947 147518 159433
rect 147478 158941 147530 158947
rect 147478 158883 147530 158889
rect 146900 156982 146956 156991
rect 146900 156917 146956 156926
rect 146914 156209 146942 156917
rect 146902 156203 146954 156209
rect 146902 156145 146954 156151
rect 148258 155534 148286 164317
rect 148162 155506 148286 155534
rect 147668 146178 147724 146187
rect 147668 146113 147724 146122
rect 147682 145775 147710 146113
rect 147670 145769 147722 145775
rect 147670 145711 147722 145717
rect 147476 144550 147532 144559
rect 147476 144485 147532 144494
rect 147490 144073 147518 144485
rect 147478 144067 147530 144073
rect 147478 144009 147530 144015
rect 147476 143662 147532 143671
rect 147476 143597 147532 143606
rect 147490 143407 147518 143597
rect 147478 143401 147530 143407
rect 147478 143343 147530 143349
rect 147668 142478 147724 142487
rect 147668 142413 147670 142422
rect 147722 142413 147724 142422
rect 147670 142381 147722 142387
rect 147478 140367 147530 140373
rect 147478 140309 147530 140315
rect 147490 139971 147518 140309
rect 147476 139962 147532 139971
rect 147476 139897 147532 139906
rect 147476 138778 147532 138787
rect 147476 138713 147532 138722
rect 147490 138301 147518 138713
rect 147478 138295 147530 138301
rect 147478 138237 147530 138243
rect 148054 137111 148106 137117
rect 148054 137053 148106 137059
rect 147476 130342 147532 130351
rect 147476 130277 147532 130286
rect 147490 129717 147518 130277
rect 147478 129711 147530 129717
rect 147478 129653 147530 129659
rect 147476 127974 147532 127983
rect 147476 127909 147532 127918
rect 147490 127867 147518 127909
rect 147478 127861 147530 127867
rect 147478 127803 147530 127809
rect 148066 123723 148094 137053
rect 148162 123871 148190 155506
rect 148246 137037 148298 137043
rect 148246 136979 148298 136985
rect 148150 123865 148202 123871
rect 148150 123807 148202 123813
rect 148054 123717 148106 123723
rect 148054 123659 148106 123665
rect 148258 123649 148286 136979
rect 148354 126683 148382 168017
rect 148436 166306 148492 166315
rect 148436 166241 148492 166250
rect 148450 137117 148478 166241
rect 148438 137111 148490 137117
rect 148438 137053 148490 137059
rect 148438 136963 148490 136969
rect 148438 136905 148490 136911
rect 148342 126677 148394 126683
rect 148342 126619 148394 126625
rect 148246 123643 148298 123649
rect 148246 123585 148298 123591
rect 148340 122498 148396 122507
rect 148340 122433 148396 122442
rect 147860 120574 147916 120583
rect 147860 120509 147862 120518
rect 147914 120509 147916 120518
rect 147862 120477 147914 120483
rect 148244 111990 148300 111999
rect 148244 111925 148300 111934
rect 147188 108438 147244 108447
rect 147188 108373 147244 108382
rect 147202 108331 147230 108373
rect 147190 108325 147242 108331
rect 147190 108267 147242 108273
rect 148258 92125 148286 111925
rect 148354 97897 148382 122433
rect 148450 120911 148478 136905
rect 148546 126609 148574 169053
rect 148642 166939 148670 233581
rect 148738 172637 148766 243349
rect 149012 240898 149068 240907
rect 149012 240833 149068 240842
rect 148916 236754 148972 236763
rect 148916 236689 148972 236698
rect 148820 234830 148876 234839
rect 148820 234765 148876 234774
rect 148726 172631 148778 172637
rect 148726 172573 148778 172579
rect 148834 167013 148862 234765
rect 148930 169677 148958 236689
rect 149026 172711 149054 240833
rect 149108 236014 149164 236023
rect 149108 235949 149164 235958
rect 149122 174136 149150 235949
rect 149396 231130 149452 231139
rect 149396 231065 149452 231074
rect 149410 230505 149438 231065
rect 149398 230499 149450 230505
rect 149398 230441 149450 230447
rect 149396 228170 149452 228179
rect 149396 228105 149452 228114
rect 149410 227619 149438 228105
rect 149398 227613 149450 227619
rect 149398 227555 149450 227561
rect 149396 227430 149452 227439
rect 149396 227365 149452 227374
rect 149410 227027 149438 227365
rect 149398 227021 149450 227027
rect 149398 226963 149450 226969
rect 149492 225210 149548 225219
rect 149492 225145 149548 225154
rect 149506 224733 149534 225145
rect 149494 224727 149546 224733
rect 149494 224669 149546 224675
rect 149492 223878 149548 223887
rect 149492 223813 149548 223822
rect 149396 222694 149452 222703
rect 149396 222629 149452 222638
rect 149410 221921 149438 222629
rect 149398 221915 149450 221921
rect 149398 221857 149450 221863
rect 149506 221847 149534 223813
rect 149494 221841 149546 221847
rect 149494 221783 149546 221789
rect 149492 219734 149548 219743
rect 149492 219669 149548 219678
rect 149506 219035 149534 219669
rect 149494 219029 149546 219035
rect 149396 218994 149452 219003
rect 149494 218971 149546 218977
rect 149396 218929 149398 218938
rect 149450 218929 149452 218938
rect 149398 218897 149450 218903
rect 149396 217810 149452 217819
rect 149396 217745 149452 217754
rect 149410 216075 149438 217745
rect 149492 216626 149548 216635
rect 149492 216561 149548 216570
rect 149506 216149 149534 216561
rect 149494 216143 149546 216149
rect 149494 216085 149546 216091
rect 149398 216069 149450 216075
rect 149398 216011 149450 216017
rect 149396 214998 149452 215007
rect 149396 214933 149452 214942
rect 149410 214743 149438 214933
rect 149398 214737 149450 214743
rect 149398 214679 149450 214685
rect 149396 205674 149452 205683
rect 149396 205609 149452 205618
rect 149410 204531 149438 205609
rect 149398 204525 149450 204531
rect 149300 204490 149356 204499
rect 149398 204467 149450 204473
rect 149300 204425 149356 204434
rect 149314 201645 149342 204425
rect 149492 203306 149548 203315
rect 149492 203241 149548 203250
rect 149396 201974 149452 201983
rect 149396 201909 149452 201918
rect 149410 201793 149438 201909
rect 149398 201787 149450 201793
rect 149398 201729 149450 201735
rect 149506 201719 149534 203241
rect 149494 201713 149546 201719
rect 149494 201655 149546 201661
rect 149302 201639 149354 201645
rect 149302 201581 149354 201587
rect 149396 200790 149452 200799
rect 149396 200725 149452 200734
rect 149410 198759 149438 200725
rect 149398 198753 149450 198759
rect 149398 198695 149450 198701
rect 149492 198422 149548 198431
rect 149492 198357 149548 198366
rect 149396 197090 149452 197099
rect 149396 197025 149452 197034
rect 149410 196021 149438 197025
rect 149398 196015 149450 196021
rect 149398 195957 149450 195963
rect 149506 195947 149534 198357
rect 149494 195941 149546 195947
rect 149396 195906 149452 195915
rect 149494 195883 149546 195889
rect 149396 195841 149398 195850
rect 149450 195841 149452 195850
rect 149398 195809 149450 195815
rect 149492 194722 149548 194731
rect 149492 194657 149548 194666
rect 149396 193390 149452 193399
rect 149396 193325 149452 193334
rect 149410 193209 149438 193325
rect 149398 193203 149450 193209
rect 149398 193145 149450 193151
rect 149506 193061 149534 194657
rect 149494 193055 149546 193061
rect 149494 192997 149546 193003
rect 149396 192206 149452 192215
rect 149396 192141 149452 192150
rect 149410 190175 149438 192141
rect 149398 190169 149450 190175
rect 149398 190111 149450 190117
rect 149698 190027 149726 271733
rect 149794 269059 149822 278018
rect 150946 271575 150974 278018
rect 150934 271569 150986 271575
rect 150934 271511 150986 271517
rect 149782 269053 149834 269059
rect 149782 268995 149834 269001
rect 152194 268985 152222 278018
rect 153346 273277 153374 278018
rect 153334 273271 153386 273277
rect 153334 273213 153386 273219
rect 152374 271569 152426 271575
rect 152374 271511 152426 271517
rect 152182 268979 152234 268985
rect 152182 268921 152234 268927
rect 151222 229833 151274 229839
rect 151222 229775 151274 229781
rect 151126 226133 151178 226139
rect 151126 226075 151178 226081
rect 149686 190021 149738 190027
rect 149686 189963 149738 189969
rect 149396 189838 149452 189847
rect 149396 189773 149452 189782
rect 149300 187470 149356 187479
rect 149300 187405 149356 187414
rect 149204 186286 149260 186295
rect 149204 186221 149260 186230
rect 149218 180037 149246 186221
rect 149314 182997 149342 187405
rect 149410 185809 149438 189773
rect 149492 188062 149548 188071
rect 149492 187997 149548 188006
rect 149398 185803 149450 185809
rect 149398 185745 149450 185751
rect 149396 183770 149452 183779
rect 149396 183705 149452 183714
rect 149302 182991 149354 182997
rect 149302 182933 149354 182939
rect 149410 181517 149438 183705
rect 149506 182923 149534 187997
rect 149588 184510 149644 184519
rect 149588 184445 149644 184454
rect 149494 182917 149546 182923
rect 149494 182859 149546 182865
rect 149492 182586 149548 182595
rect 149492 182521 149548 182530
rect 149398 181511 149450 181517
rect 149398 181453 149450 181459
rect 149300 181402 149356 181411
rect 149300 181337 149356 181346
rect 149206 180031 149258 180037
rect 149206 179973 149258 179979
rect 149314 178631 149342 181337
rect 149506 179908 149534 182521
rect 149602 180111 149630 184445
rect 149590 180105 149642 180111
rect 149590 180047 149642 180053
rect 149506 179880 149630 179908
rect 149492 179626 149548 179635
rect 149492 179561 149548 179570
rect 149396 178886 149452 178895
rect 149396 178821 149452 178830
rect 149410 178779 149438 178821
rect 149398 178773 149450 178779
rect 149398 178715 149450 178721
rect 149506 178705 149534 179561
rect 149494 178699 149546 178705
rect 149494 178641 149546 178647
rect 149302 178625 149354 178631
rect 149302 178567 149354 178573
rect 149396 177702 149452 177711
rect 149396 177637 149452 177646
rect 149410 177299 149438 177637
rect 149398 177293 149450 177299
rect 149398 177235 149450 177241
rect 149602 175694 149630 179880
rect 149218 175666 149630 175694
rect 149218 174265 149246 175666
rect 149396 175186 149452 175195
rect 149396 175121 149452 175130
rect 149206 174259 149258 174265
rect 149206 174201 149258 174207
rect 149122 174108 149342 174136
rect 149108 174002 149164 174011
rect 149108 173937 149164 173946
rect 149014 172705 149066 172711
rect 149014 172647 149066 172653
rect 149012 170302 149068 170311
rect 149012 170237 149068 170246
rect 148918 169671 148970 169677
rect 148918 169613 148970 169619
rect 148822 167007 148874 167013
rect 148822 166949 148874 166955
rect 148630 166933 148682 166939
rect 148630 166875 148682 166881
rect 148724 165566 148780 165575
rect 148724 165501 148780 165510
rect 148628 161866 148684 161875
rect 148628 161801 148684 161810
rect 148642 136969 148670 161801
rect 148738 137043 148766 165501
rect 148916 163198 148972 163207
rect 148916 163133 148972 163142
rect 148820 160682 148876 160691
rect 148820 160617 148876 160626
rect 148726 137037 148778 137043
rect 148726 136979 148778 136985
rect 148630 136963 148682 136969
rect 148630 136905 148682 136911
rect 148834 136840 148862 160617
rect 148930 136969 148958 163133
rect 148918 136963 148970 136969
rect 148918 136905 148970 136911
rect 149026 136840 149054 170237
rect 149122 155636 149150 173937
rect 149314 169751 149342 174108
rect 149410 172859 149438 175121
rect 149398 172853 149450 172859
rect 149398 172795 149450 172801
rect 149588 172818 149644 172827
rect 149588 172753 149644 172762
rect 149492 171042 149548 171051
rect 149492 170977 149548 170986
rect 149302 169745 149354 169751
rect 149302 169687 149354 169693
rect 149300 157722 149356 157731
rect 149300 157657 149356 157666
rect 149314 155765 149342 157657
rect 149396 155798 149452 155807
rect 149302 155759 149354 155765
rect 149396 155733 149452 155742
rect 149302 155701 149354 155707
rect 149410 155691 149438 155733
rect 149398 155685 149450 155691
rect 149122 155608 149342 155636
rect 149398 155627 149450 155633
rect 149314 155534 149342 155608
rect 148642 136812 148862 136840
rect 148930 136812 149054 136840
rect 149122 155506 149342 155534
rect 148534 126603 148586 126609
rect 148534 126545 148586 126551
rect 148532 121758 148588 121767
rect 148532 121693 148588 121702
rect 148438 120905 148490 120911
rect 148438 120847 148490 120853
rect 148436 107254 148492 107263
rect 148436 107189 148492 107198
rect 148342 97891 148394 97897
rect 148342 97833 148394 97839
rect 148246 92119 148298 92125
rect 148246 92061 148298 92067
rect 148450 89239 148478 107189
rect 148546 97823 148574 121693
rect 148642 120985 148670 136812
rect 148726 136741 148778 136747
rect 148726 136683 148778 136689
rect 148738 123797 148766 136683
rect 148820 133894 148876 133903
rect 148820 133829 148876 133838
rect 148726 123791 148778 123797
rect 148726 123733 148778 123739
rect 148630 120979 148682 120985
rect 148630 120921 148682 120927
rect 148834 115255 148862 133829
rect 148930 126535 148958 136812
rect 149012 132710 149068 132719
rect 149012 132645 149068 132654
rect 148918 126529 148970 126535
rect 148918 126471 148970 126477
rect 148820 115246 148876 115255
rect 148820 115181 148876 115190
rect 148628 109622 148684 109631
rect 148628 109557 148630 109566
rect 148682 109557 148684 109566
rect 148630 109525 148682 109531
rect 148820 106070 148876 106079
rect 148820 106005 148876 106014
rect 148628 104738 148684 104747
rect 148628 104673 148684 104682
rect 148534 97817 148586 97823
rect 148534 97759 148586 97765
rect 148438 89233 148490 89239
rect 148438 89175 148490 89181
rect 148642 86427 148670 104673
rect 148724 103554 148780 103563
rect 148724 103489 148780 103498
rect 148630 86421 148682 86427
rect 148630 86363 148682 86369
rect 148738 86353 148766 103489
rect 148834 89165 148862 106005
rect 149026 103669 149054 132645
rect 149122 129347 149150 155506
rect 149300 154614 149356 154623
rect 149300 154549 149356 154558
rect 149314 152731 149342 154549
rect 149396 153134 149452 153143
rect 149396 153069 149452 153078
rect 149410 152805 149438 153069
rect 149398 152799 149450 152805
rect 149398 152741 149450 152747
rect 149302 152725 149354 152731
rect 149302 152667 149354 152673
rect 149204 152098 149260 152107
rect 149204 152033 149260 152042
rect 149218 149845 149246 152033
rect 149396 150914 149452 150923
rect 149396 150849 149452 150858
rect 149302 149987 149354 149993
rect 149302 149929 149354 149935
rect 149314 149887 149342 149929
rect 149410 149919 149438 150849
rect 149398 149913 149450 149919
rect 149300 149878 149356 149887
rect 149206 149839 149258 149845
rect 149398 149855 149450 149861
rect 149300 149813 149356 149822
rect 149206 149781 149258 149787
rect 149300 148546 149356 148555
rect 149300 148481 149356 148490
rect 149314 146959 149342 148481
rect 149396 147362 149452 147371
rect 149396 147297 149452 147306
rect 149410 147033 149438 147297
rect 149398 147027 149450 147033
rect 149398 146969 149450 146975
rect 149302 146953 149354 146959
rect 149302 146895 149354 146901
rect 149506 146894 149534 170977
rect 149410 146866 149534 146894
rect 149410 129421 149438 146866
rect 149602 137728 149630 172753
rect 149684 141294 149740 141303
rect 149684 141229 149686 141238
rect 149738 141229 149740 141238
rect 149686 141197 149738 141203
rect 151138 140373 151166 226075
rect 151234 164127 151262 229775
rect 151318 224801 151370 224807
rect 151318 224743 151370 224749
rect 151222 164121 151274 164127
rect 151222 164063 151274 164069
rect 151330 161241 151358 224743
rect 151414 220805 151466 220811
rect 151414 220747 151466 220753
rect 151318 161235 151370 161241
rect 151318 161177 151370 161183
rect 151426 158429 151454 220747
rect 151798 214071 151850 214077
rect 151798 214013 151850 214019
rect 151702 211333 151754 211339
rect 151702 211275 151754 211281
rect 151606 210371 151658 210377
rect 151606 210313 151658 210319
rect 151510 207929 151562 207935
rect 151510 207871 151562 207877
rect 151414 158423 151466 158429
rect 151414 158365 151466 158371
rect 151222 156203 151274 156209
rect 151222 156145 151274 156151
rect 151126 140367 151178 140373
rect 151126 140309 151178 140315
rect 149506 137700 149630 137728
rect 149506 129495 149534 137700
rect 149588 137594 149644 137603
rect 149588 137529 149644 137538
rect 149602 135415 149630 137529
rect 149684 135966 149740 135975
rect 149684 135901 149740 135910
rect 149698 135489 149726 135901
rect 149686 135483 149738 135489
rect 149686 135425 149738 135431
rect 149590 135409 149642 135415
rect 149590 135351 149642 135357
rect 149684 135078 149740 135087
rect 149684 135013 149740 135022
rect 149698 132529 149726 135013
rect 149686 132523 149738 132529
rect 149686 132465 149738 132471
rect 149684 130934 149740 130943
rect 149684 130869 149740 130878
rect 149698 129643 149726 130869
rect 149686 129637 149738 129643
rect 149686 129579 149738 129585
rect 149494 129489 149546 129495
rect 149494 129431 149546 129437
rect 149398 129415 149450 129421
rect 149398 129357 149450 129363
rect 149110 129341 149162 129347
rect 149110 129283 149162 129289
rect 149108 129158 149164 129167
rect 149108 129093 149164 129102
rect 149014 103663 149066 103669
rect 149014 103605 149066 103611
rect 149122 103595 149150 129093
rect 149300 126642 149356 126651
rect 149300 126577 149356 126586
rect 149110 103589 149162 103595
rect 149110 103531 149162 103537
rect 148916 102370 148972 102379
rect 148916 102305 148972 102314
rect 148822 89159 148874 89165
rect 148822 89101 148874 89107
rect 148820 86534 148876 86543
rect 148820 86469 148822 86478
rect 148874 86469 148876 86478
rect 148822 86437 148874 86443
rect 148726 86347 148778 86353
rect 148726 86289 148778 86295
rect 148930 86279 148958 102305
rect 149314 100709 149342 126577
rect 149588 125458 149644 125467
rect 149588 125393 149644 125402
rect 149396 124274 149452 124283
rect 149396 124209 149398 124218
rect 149450 124209 149452 124218
rect 149398 124177 149450 124183
rect 149492 119390 149548 119399
rect 149492 119325 149548 119334
rect 149398 118241 149450 118247
rect 149396 118206 149398 118215
rect 149450 118206 149452 118215
rect 149506 118173 149534 119325
rect 149396 118141 149452 118150
rect 149494 118167 149546 118173
rect 149494 118109 149546 118115
rect 149492 116874 149548 116883
rect 149492 116809 149548 116818
rect 149396 115690 149452 115699
rect 149396 115625 149452 115634
rect 149410 115361 149438 115625
rect 149398 115355 149450 115361
rect 149398 115297 149450 115303
rect 149506 115287 149534 116809
rect 149494 115281 149546 115287
rect 149396 115246 149452 115255
rect 149494 115223 149546 115229
rect 149396 115181 149452 115190
rect 149410 114640 149438 115181
rect 149410 114612 149534 114640
rect 149396 114506 149452 114515
rect 149396 114441 149452 114450
rect 149410 114103 149438 114441
rect 149398 114097 149450 114103
rect 149398 114039 149450 114045
rect 149396 113174 149452 113183
rect 149396 113109 149452 113118
rect 149410 112401 149438 113109
rect 149398 112395 149450 112401
rect 149398 112337 149450 112343
rect 149396 110954 149452 110963
rect 149396 110889 149452 110898
rect 149410 109515 149438 110889
rect 149398 109509 149450 109515
rect 149398 109451 149450 109457
rect 149506 106333 149534 114612
rect 149494 106327 149546 106333
rect 149494 106269 149546 106275
rect 149396 100890 149452 100899
rect 149396 100825 149398 100834
rect 149450 100825 149452 100834
rect 149398 100793 149450 100799
rect 149602 100783 149630 125393
rect 151234 112327 151262 156145
rect 151522 149549 151550 207871
rect 151618 152583 151646 210313
rect 151606 152577 151658 152583
rect 151606 152519 151658 152525
rect 151714 152509 151742 211275
rect 151810 155543 151838 214013
rect 152086 212887 152138 212893
rect 152086 212829 152138 212835
rect 151990 207411 152042 207417
rect 151990 207353 152042 207359
rect 151894 204599 151946 204605
rect 151894 204541 151946 204547
rect 151798 155537 151850 155543
rect 151798 155479 151850 155485
rect 151702 152503 151754 152509
rect 151702 152445 151754 152451
rect 151906 149697 151934 204541
rect 152002 152657 152030 207353
rect 152098 155469 152126 212829
rect 152386 192987 152414 271511
rect 154498 270761 154526 278018
rect 154486 270755 154538 270761
rect 154486 270697 154538 270703
rect 155446 270755 155498 270761
rect 155446 270697 155498 270703
rect 154006 249443 154058 249449
rect 154006 249385 154058 249391
rect 152374 192981 152426 192987
rect 152374 192923 152426 192929
rect 154018 181221 154046 249385
rect 154102 232201 154154 232207
rect 154102 232143 154154 232149
rect 154006 181215 154058 181221
rect 154006 181157 154058 181163
rect 154006 176035 154058 176041
rect 154006 175977 154058 175983
rect 152182 158941 152234 158947
rect 152182 158883 152234 158889
rect 152086 155463 152138 155469
rect 152086 155405 152138 155411
rect 151990 152651 152042 152657
rect 151990 152593 152042 152599
rect 151894 149691 151946 149697
rect 151894 149633 151946 149639
rect 151510 149543 151562 149549
rect 151510 149485 151562 149491
rect 152194 115213 152222 158883
rect 154018 132455 154046 175977
rect 154114 166865 154142 232143
rect 154198 198827 154250 198833
rect 154198 198769 154250 198775
rect 154102 166859 154154 166865
rect 154102 166801 154154 166807
rect 154210 146885 154238 198769
rect 155458 192913 155486 270697
rect 155746 268911 155774 278018
rect 155734 268905 155786 268911
rect 155734 268847 155786 268853
rect 156898 268837 156926 278018
rect 158050 276494 158078 278018
rect 158050 276466 158174 276494
rect 156886 268831 156938 268837
rect 156886 268773 156938 268779
rect 156886 252329 156938 252335
rect 156886 252271 156938 252277
rect 155446 192907 155498 192913
rect 155446 192849 155498 192855
rect 154294 190243 154346 190249
rect 154294 190185 154346 190191
rect 154198 146879 154250 146885
rect 154198 146821 154250 146827
rect 154102 141255 154154 141261
rect 154102 141197 154154 141203
rect 154006 132449 154058 132455
rect 154006 132391 154058 132397
rect 152182 115207 152234 115213
rect 152182 115149 152234 115155
rect 154114 115139 154142 141197
rect 154306 141113 154334 190185
rect 156898 181369 156926 252271
rect 156982 230499 157034 230505
rect 156982 230441 157034 230447
rect 156886 181363 156938 181369
rect 156886 181305 156938 181311
rect 156886 177293 156938 177299
rect 156886 177235 156938 177241
rect 154294 141107 154346 141113
rect 154294 141049 154346 141055
rect 156898 132381 156926 177235
rect 156994 164053 157022 230441
rect 158146 192839 158174 276466
rect 159298 271945 159326 278018
rect 160450 273573 160478 278018
rect 160438 273567 160490 273573
rect 160438 273509 160490 273515
rect 159286 271939 159338 271945
rect 159286 271881 159338 271887
rect 161602 271279 161630 278018
rect 161590 271273 161642 271279
rect 161590 271215 161642 271221
rect 162850 268763 162878 278018
rect 163894 271273 163946 271279
rect 163894 271215 163946 271221
rect 162838 268757 162890 268763
rect 162838 268699 162890 268705
rect 159862 249887 159914 249893
rect 159862 249829 159914 249835
rect 159766 227021 159818 227027
rect 159766 226963 159818 226969
rect 158134 192833 158186 192839
rect 158134 192775 158186 192781
rect 157078 190169 157130 190175
rect 157078 190111 157130 190117
rect 156982 164047 157034 164053
rect 156982 163989 157034 163995
rect 156982 142439 157034 142445
rect 156982 142381 157034 142387
rect 156886 132375 156938 132381
rect 156886 132317 156938 132323
rect 156886 124235 156938 124241
rect 156886 124177 156938 124183
rect 154486 120535 154538 120541
rect 154486 120477 154538 120483
rect 154102 115133 154154 115139
rect 154102 115075 154154 115081
rect 151222 112321 151274 112327
rect 151222 112263 151274 112269
rect 154006 109583 154058 109589
rect 154006 109525 154058 109531
rect 151126 108325 151178 108331
rect 151126 108267 151178 108273
rect 149590 100777 149642 100783
rect 149590 100719 149642 100725
rect 149302 100703 149354 100709
rect 149302 100645 149354 100651
rect 149492 99854 149548 99863
rect 149492 99789 149548 99798
rect 149396 98670 149452 98679
rect 149396 98605 149452 98614
rect 149410 98045 149438 98605
rect 149398 98039 149450 98045
rect 149398 97981 149450 97987
rect 149506 97971 149534 99789
rect 149494 97965 149546 97971
rect 149494 97907 149546 97913
rect 149492 97486 149548 97495
rect 149492 97421 149548 97430
rect 149396 95710 149452 95719
rect 149396 95645 149452 95654
rect 149410 95085 149438 95645
rect 149506 95159 149534 97421
rect 149494 95153 149546 95159
rect 149494 95095 149546 95101
rect 149398 95079 149450 95085
rect 149398 95021 149450 95027
rect 149588 94970 149644 94979
rect 149588 94905 149644 94914
rect 149492 93786 149548 93795
rect 149492 93721 149548 93730
rect 149396 92602 149452 92611
rect 149396 92537 149452 92546
rect 149410 92273 149438 92537
rect 149398 92267 149450 92273
rect 149398 92209 149450 92215
rect 149506 92199 149534 93721
rect 149494 92193 149546 92199
rect 149494 92135 149546 92141
rect 149300 91418 149356 91427
rect 149300 91353 149356 91362
rect 148918 86273 148970 86279
rect 148918 86215 148970 86221
rect 148820 85350 148876 85359
rect 148820 85285 148876 85294
rect 147092 84166 147148 84175
rect 147092 84101 147148 84110
rect 147106 83615 147134 84101
rect 147094 83609 147146 83615
rect 147094 83551 147146 83557
rect 148436 81650 148492 81659
rect 148436 81585 148492 81594
rect 148450 71997 148478 81585
rect 148834 74883 148862 85285
rect 149108 82390 149164 82399
rect 149108 82325 149164 82334
rect 148916 77950 148972 77959
rect 148916 77885 148972 77894
rect 148822 74877 148874 74883
rect 148822 74819 148874 74825
rect 148438 71991 148490 71997
rect 148438 71933 148490 71939
rect 148930 69037 148958 77885
rect 149122 74809 149150 82325
rect 149314 77769 149342 91353
rect 149396 90234 149452 90243
rect 149396 90169 149452 90178
rect 149410 90127 149438 90169
rect 149398 90121 149450 90127
rect 149398 90063 149450 90069
rect 149396 89050 149452 89059
rect 149396 88985 149452 88994
rect 149302 77763 149354 77769
rect 149302 77705 149354 77711
rect 149410 77695 149438 88985
rect 149492 87274 149548 87283
rect 149492 87209 149548 87218
rect 149506 86797 149534 87209
rect 149494 86791 149546 86797
rect 149494 86733 149546 86739
rect 149602 80655 149630 94905
rect 151138 89091 151166 108267
rect 151126 89085 151178 89091
rect 151126 89027 151178 89033
rect 154018 89017 154046 109525
rect 154498 105149 154526 120477
rect 154486 105143 154538 105149
rect 154486 105085 154538 105091
rect 156898 100635 156926 124177
rect 156994 115065 157022 142381
rect 157090 141039 157118 190111
rect 159778 163979 159806 226963
rect 159874 187215 159902 249829
rect 162646 249221 162698 249227
rect 162646 249163 162698 249169
rect 159958 214737 160010 214743
rect 159958 214679 160010 214685
rect 159862 187209 159914 187215
rect 159862 187151 159914 187157
rect 159766 163973 159818 163979
rect 159766 163915 159818 163921
rect 159970 155395 159998 214679
rect 160054 193203 160106 193209
rect 160054 193145 160106 193151
rect 159958 155389 160010 155395
rect 159958 155331 160010 155337
rect 159862 143401 159914 143407
rect 159862 143343 159914 143349
rect 157078 141033 157130 141039
rect 157078 140975 157130 140981
rect 159766 138295 159818 138301
rect 159766 138237 159818 138243
rect 156982 115059 157034 115065
rect 156982 115001 157034 115007
rect 156982 109509 157034 109515
rect 156982 109451 157034 109457
rect 156886 100629 156938 100635
rect 156886 100571 156938 100577
rect 156994 92051 157022 109451
rect 159778 109441 159806 138237
rect 159874 118099 159902 143343
rect 160066 140965 160094 193145
rect 162658 178483 162686 249163
rect 162742 224727 162794 224733
rect 162742 224669 162794 224675
rect 162646 178477 162698 178483
rect 162646 178419 162698 178425
rect 162754 161167 162782 224669
rect 162838 198753 162890 198759
rect 162838 198695 162890 198701
rect 162742 161161 162794 161167
rect 162742 161103 162794 161109
rect 162850 146811 162878 198695
rect 163906 192765 163934 271215
rect 164002 268689 164030 278018
rect 165154 272093 165182 278018
rect 165142 272087 165194 272093
rect 165142 272029 165194 272035
rect 166306 271723 166334 278018
rect 167554 272093 167582 278018
rect 166966 272087 167018 272093
rect 166966 272029 167018 272035
rect 167542 272087 167594 272093
rect 167542 272029 167594 272035
rect 166294 271717 166346 271723
rect 166294 271659 166346 271665
rect 163990 268683 164042 268689
rect 163990 268625 164042 268631
rect 165718 249591 165770 249597
rect 165718 249533 165770 249539
rect 165526 246779 165578 246785
rect 165526 246721 165578 246727
rect 163894 192759 163946 192765
rect 163894 192701 163946 192707
rect 165538 181295 165566 246721
rect 165622 219029 165674 219035
rect 165622 218971 165674 218977
rect 165526 181289 165578 181295
rect 165526 181231 165578 181237
rect 162934 178773 162986 178779
rect 162934 178715 162986 178721
rect 162838 146805 162890 146811
rect 162838 146747 162890 146753
rect 162742 144067 162794 144073
rect 162742 144009 162794 144015
rect 160054 140959 160106 140965
rect 160054 140901 160106 140907
rect 162646 127861 162698 127867
rect 162646 127803 162698 127809
rect 159862 118093 159914 118099
rect 159862 118035 159914 118041
rect 159862 114097 159914 114103
rect 159862 114039 159914 114045
rect 159766 109435 159818 109441
rect 159766 109377 159818 109383
rect 156982 92045 157034 92051
rect 156982 91987 157034 91993
rect 159874 91977 159902 114039
rect 162658 100561 162686 127803
rect 162754 118025 162782 144009
rect 162946 132307 162974 178715
rect 165634 158355 165662 218971
rect 165730 187141 165758 249533
rect 166978 195799 167006 272029
rect 168706 270761 168734 278018
rect 169762 278004 169872 278032
rect 168694 270755 168746 270761
rect 168694 270697 168746 270703
rect 169762 268541 169790 278004
rect 169846 270755 169898 270761
rect 169846 270697 169898 270703
rect 169750 268535 169802 268541
rect 169750 268477 169802 268483
rect 168502 249813 168554 249819
rect 168502 249755 168554 249761
rect 168406 221915 168458 221921
rect 168406 221857 168458 221863
rect 166966 195793 167018 195799
rect 166966 195735 167018 195741
rect 165814 193055 165866 193061
rect 165814 192997 165866 193003
rect 165718 187135 165770 187141
rect 165718 187077 165770 187083
rect 165718 178699 165770 178705
rect 165718 178641 165770 178647
rect 165622 158349 165674 158355
rect 165622 158291 165674 158297
rect 165526 145769 165578 145775
rect 165526 145711 165578 145717
rect 162934 132301 162986 132307
rect 162934 132243 162986 132249
rect 162742 118019 162794 118025
rect 162742 117961 162794 117967
rect 165538 117951 165566 145711
rect 165730 132233 165758 178641
rect 165826 143777 165854 192997
rect 168418 161093 168446 221857
rect 168514 187067 168542 249755
rect 168598 196015 168650 196021
rect 168598 195957 168650 195963
rect 168502 187061 168554 187067
rect 168502 187003 168554 187009
rect 168502 178625 168554 178631
rect 168502 178567 168554 178573
rect 168406 161087 168458 161093
rect 168406 161029 168458 161035
rect 168406 147027 168458 147033
rect 168406 146969 168458 146975
rect 165814 143771 165866 143777
rect 165814 143713 165866 143719
rect 165718 132227 165770 132233
rect 165718 132169 165770 132175
rect 165622 129711 165674 129717
rect 165622 129653 165674 129659
rect 165526 117945 165578 117951
rect 165526 117887 165578 117893
rect 162838 115355 162890 115361
rect 162838 115297 162890 115303
rect 162646 100555 162698 100561
rect 162646 100497 162698 100503
rect 162850 95011 162878 115297
rect 165634 103521 165662 129653
rect 168418 117877 168446 146969
rect 168514 135341 168542 178567
rect 168610 143925 168638 195957
rect 169858 195725 169886 270697
rect 171106 268615 171134 278018
rect 172272 278004 172766 278032
rect 171094 268609 171146 268615
rect 171094 268551 171146 268557
rect 171286 252181 171338 252187
rect 171286 252123 171338 252129
rect 169846 195719 169898 195725
rect 169846 195661 169898 195667
rect 171298 184255 171326 252123
rect 171478 249739 171530 249745
rect 171478 249681 171530 249687
rect 171382 221841 171434 221847
rect 171382 221783 171434 221789
rect 171286 184249 171338 184255
rect 171286 184191 171338 184197
rect 171394 161019 171422 221783
rect 171490 189953 171518 249681
rect 171574 195941 171626 195947
rect 171574 195883 171626 195889
rect 171478 189947 171530 189953
rect 171478 189889 171530 189895
rect 171478 181511 171530 181517
rect 171478 181453 171530 181459
rect 171382 161013 171434 161019
rect 171382 160955 171434 160961
rect 171382 149987 171434 149993
rect 171382 149929 171434 149935
rect 168598 143919 168650 143925
rect 168598 143861 168650 143867
rect 171286 135483 171338 135489
rect 171286 135425 171338 135431
rect 168502 135335 168554 135341
rect 168502 135277 168554 135283
rect 168502 129637 168554 129643
rect 168502 129579 168554 129585
rect 168406 117871 168458 117877
rect 168406 117813 168458 117819
rect 165718 115281 165770 115287
rect 165718 115223 165770 115229
rect 165622 103515 165674 103521
rect 165622 103457 165674 103463
rect 162838 95005 162890 95011
rect 162838 94947 162890 94953
rect 165730 94937 165758 115223
rect 168514 103447 168542 129579
rect 168598 118241 168650 118247
rect 168598 118183 168650 118189
rect 168502 103441 168554 103447
rect 168502 103383 168554 103389
rect 168214 95153 168266 95159
rect 168214 95095 168266 95101
rect 165718 94931 165770 94937
rect 165718 94873 165770 94879
rect 162454 92267 162506 92273
rect 162454 92209 162506 92215
rect 159862 91971 159914 91977
rect 159862 91913 159914 91919
rect 159766 90121 159818 90127
rect 159766 90063 159818 90069
rect 154006 89011 154058 89017
rect 154006 88953 154058 88959
rect 156502 86791 156554 86797
rect 156502 86733 156554 86739
rect 154102 86495 154154 86501
rect 154102 86437 154154 86443
rect 151126 83609 151178 83615
rect 151126 83551 151178 83557
rect 149590 80649 149642 80655
rect 149590 80591 149642 80597
rect 149588 80466 149644 80475
rect 149588 80401 149644 80410
rect 149398 77689 149450 77695
rect 149398 77631 149450 77637
rect 149396 76766 149452 76775
rect 149396 76701 149452 76710
rect 149204 75582 149260 75591
rect 149204 75517 149260 75526
rect 149110 74803 149162 74809
rect 149110 74745 149162 74751
rect 149012 73066 149068 73075
rect 149012 73001 149068 73010
rect 148918 69031 148970 69037
rect 148918 68973 148970 68979
rect 149026 66003 149054 73001
rect 149108 72030 149164 72039
rect 149108 71965 149164 71974
rect 149122 66225 149150 71965
rect 149218 68963 149246 75517
rect 149410 74894 149438 76701
rect 149410 74866 149534 74894
rect 149300 73806 149356 73815
rect 149300 73741 149356 73750
rect 149206 68957 149258 68963
rect 149206 68899 149258 68905
rect 149314 68889 149342 73741
rect 149506 70980 149534 74866
rect 149602 71849 149630 80401
rect 149684 79282 149740 79291
rect 149684 79217 149740 79226
rect 149698 71923 149726 79217
rect 151138 74735 151166 83551
rect 151126 74729 151178 74735
rect 151126 74671 151178 74677
rect 154114 74661 154142 86437
rect 156514 77621 156542 86733
rect 156502 77615 156554 77621
rect 156502 77557 156554 77563
rect 159778 77547 159806 90063
rect 162466 80581 162494 92209
rect 165238 92193 165290 92199
rect 165238 92135 165290 92141
rect 162454 80575 162506 80581
rect 162454 80517 162506 80523
rect 165250 80507 165278 92135
rect 168226 83541 168254 95095
rect 168610 94863 168638 118183
rect 171298 106481 171326 135425
rect 171394 120837 171422 149929
rect 171490 135267 171518 181453
rect 171586 143851 171614 195883
rect 172738 195651 172766 278004
rect 173410 271501 173438 278018
rect 174658 272019 174686 278018
rect 174646 272013 174698 272019
rect 174646 271955 174698 271961
rect 173398 271495 173450 271501
rect 173398 271437 173450 271443
rect 175810 271205 175838 278018
rect 175798 271199 175850 271205
rect 175798 271141 175850 271147
rect 176962 268319 176990 278018
rect 176950 268313 177002 268319
rect 176950 268255 177002 268261
rect 178210 268171 178238 278018
rect 178294 271199 178346 271205
rect 178294 271141 178346 271147
rect 178198 268165 178250 268171
rect 178198 268107 178250 268113
rect 177046 249517 177098 249523
rect 177046 249459 177098 249465
rect 174166 249147 174218 249153
rect 174166 249089 174218 249095
rect 172726 195645 172778 195651
rect 172726 195587 172778 195593
rect 174178 178409 174206 249089
rect 174262 227613 174314 227619
rect 174262 227555 174314 227561
rect 174166 178403 174218 178409
rect 174166 178345 174218 178351
rect 174274 163905 174302 227555
rect 174358 216143 174410 216149
rect 174358 216085 174410 216091
rect 174262 163899 174314 163905
rect 174262 163841 174314 163847
rect 174370 155321 174398 216085
rect 174454 201787 174506 201793
rect 174454 201729 174506 201735
rect 174358 155315 174410 155321
rect 174358 155257 174410 155263
rect 174166 152799 174218 152805
rect 174166 152741 174218 152747
rect 171574 143845 171626 143851
rect 171574 143787 171626 143793
rect 171478 135261 171530 135267
rect 171478 135203 171530 135209
rect 171382 120831 171434 120837
rect 171382 120773 171434 120779
rect 174178 109367 174206 152741
rect 174262 149913 174314 149919
rect 174262 149855 174314 149861
rect 174274 122465 174302 149855
rect 174466 146737 174494 201729
rect 177058 186993 177086 249459
rect 177142 216069 177194 216075
rect 177142 216011 177194 216017
rect 177046 186987 177098 186993
rect 177046 186929 177098 186935
rect 177154 158207 177182 216011
rect 177238 201713 177290 201719
rect 177238 201655 177290 201661
rect 177142 158201 177194 158207
rect 177142 158143 177194 158149
rect 177046 155685 177098 155691
rect 177046 155627 177098 155633
rect 174454 146731 174506 146737
rect 174454 146673 174506 146679
rect 174262 122459 174314 122465
rect 174262 122401 174314 122407
rect 174262 118167 174314 118173
rect 174262 118109 174314 118115
rect 174166 109361 174218 109367
rect 174166 109303 174218 109309
rect 171286 106475 171338 106481
rect 171286 106417 171338 106423
rect 171286 100851 171338 100857
rect 171286 100793 171338 100799
rect 168598 94857 168650 94863
rect 168598 94799 168650 94805
rect 168214 83535 168266 83541
rect 168214 83477 168266 83483
rect 171298 83467 171326 100793
rect 174274 94789 174302 118109
rect 177058 112179 177086 155627
rect 177142 146953 177194 146959
rect 177142 146895 177194 146901
rect 177154 132603 177182 146895
rect 177250 146663 177278 201655
rect 178306 198611 178334 271141
rect 179362 270761 179390 278018
rect 180514 271427 180542 278018
rect 181762 271649 181790 278018
rect 181750 271643 181802 271649
rect 181750 271585 181802 271591
rect 180502 271421 180554 271427
rect 180502 271363 180554 271369
rect 182914 270761 182942 278018
rect 184066 271279 184094 278018
rect 185218 271575 185246 278018
rect 185206 271569 185258 271575
rect 185206 271511 185258 271517
rect 184054 271273 184106 271279
rect 184054 271215 184106 271221
rect 186466 270761 186494 278018
rect 187618 271205 187646 278018
rect 188770 271353 188798 278018
rect 189730 278004 190032 278032
rect 188758 271347 188810 271353
rect 188758 271289 188810 271295
rect 187606 271199 187658 271205
rect 187606 271141 187658 271147
rect 179350 270755 179402 270761
rect 179350 270697 179402 270703
rect 181366 270755 181418 270761
rect 181366 270697 181418 270703
rect 182902 270755 182954 270761
rect 182902 270697 182954 270703
rect 184246 270755 184298 270761
rect 184246 270697 184298 270703
rect 185494 270755 185546 270761
rect 185494 270697 185546 270703
rect 186454 270755 186506 270761
rect 186454 270697 186506 270703
rect 180022 249665 180074 249671
rect 180022 249607 180074 249613
rect 179926 218955 179978 218961
rect 179926 218897 179978 218903
rect 178294 198605 178346 198611
rect 178294 198547 178346 198553
rect 179938 158281 179966 218897
rect 180034 189879 180062 249607
rect 180118 201639 180170 201645
rect 180118 201581 180170 201587
rect 180022 189873 180074 189879
rect 180022 189815 180074 189821
rect 179926 158275 179978 158281
rect 179926 158217 179978 158223
rect 180022 155759 180074 155765
rect 180022 155701 180074 155707
rect 177238 146657 177290 146663
rect 177238 146599 177290 146605
rect 179926 135409 179978 135415
rect 179926 135351 179978 135357
rect 177142 132597 177194 132603
rect 177142 132539 177194 132545
rect 177142 112395 177194 112401
rect 177142 112337 177194 112343
rect 177046 112173 177098 112179
rect 177046 112115 177098 112121
rect 174262 94783 174314 94789
rect 174262 94725 174314 94731
rect 177154 91903 177182 112337
rect 179938 106407 179966 135351
rect 180034 114177 180062 155701
rect 180130 149623 180158 201581
rect 181378 198685 181406 270697
rect 182806 252107 182858 252113
rect 182806 252049 182858 252055
rect 181366 198679 181418 198685
rect 181366 198621 181418 198627
rect 182818 181443 182846 252049
rect 182902 249369 182954 249375
rect 182902 249311 182954 249317
rect 182914 184181 182942 249311
rect 182998 204525 183050 204531
rect 182998 204467 183050 204473
rect 182902 184175 182954 184181
rect 182902 184117 182954 184123
rect 182806 181437 182858 181443
rect 182806 181379 182858 181385
rect 182806 172853 182858 172859
rect 182806 172795 182858 172801
rect 180214 149839 180266 149845
rect 180214 149781 180266 149787
rect 180118 149617 180170 149623
rect 180118 149559 180170 149565
rect 180226 132085 180254 149781
rect 180214 132079 180266 132085
rect 180214 132021 180266 132027
rect 182818 129569 182846 172795
rect 182902 152725 182954 152731
rect 182902 152667 182954 152673
rect 182806 129563 182858 129569
rect 182806 129505 182858 129511
rect 180022 114171 180074 114177
rect 180022 114113 180074 114119
rect 182914 112253 182942 152667
rect 183010 149771 183038 204467
rect 184258 197691 184286 270697
rect 184342 221767 184394 221773
rect 184342 221709 184394 221715
rect 184354 219595 184382 221709
rect 184340 219586 184396 219595
rect 184340 219521 184396 219530
rect 184342 218881 184394 218887
rect 184340 218846 184342 218855
rect 184394 218846 184396 218855
rect 184340 218781 184396 218790
rect 184342 201565 184394 201571
rect 184342 201507 184394 201513
rect 184354 199763 184382 201507
rect 184340 199754 184396 199763
rect 184340 199689 184396 199698
rect 184438 198679 184490 198685
rect 184438 198621 184490 198627
rect 184342 198605 184394 198611
rect 184342 198547 184394 198553
rect 184244 197682 184300 197691
rect 184244 197617 184300 197626
rect 184354 196063 184382 198547
rect 184450 196803 184478 198621
rect 185506 198283 185534 270697
rect 185686 269571 185738 269577
rect 185686 269513 185738 269519
rect 185698 269355 185726 269513
rect 185590 269349 185642 269355
rect 185590 269291 185642 269297
rect 185686 269349 185738 269355
rect 185686 269291 185738 269297
rect 185602 268467 185630 269291
rect 185590 268461 185642 268467
rect 185590 268403 185642 268409
rect 189730 266469 189758 278004
rect 190102 273493 190154 273499
rect 190102 273435 190154 273441
rect 190114 268097 190142 273435
rect 191170 271871 191198 278018
rect 191158 271865 191210 271871
rect 191158 271807 191210 271813
rect 192322 271797 192350 278018
rect 193570 273499 193598 278018
rect 193558 273493 193610 273499
rect 193558 273435 193610 273441
rect 194420 272274 194476 272283
rect 194420 272209 194476 272218
rect 193748 272126 193804 272135
rect 193748 272061 193804 272070
rect 192310 271791 192362 271797
rect 192310 271733 192362 271739
rect 193076 269610 193132 269619
rect 193076 269545 193132 269554
rect 192404 269314 192460 269323
rect 192404 269249 192460 269258
rect 192598 269275 192650 269281
rect 190102 268091 190154 268097
rect 190102 268033 190154 268039
rect 187222 266463 187274 266469
rect 187222 266405 187274 266411
rect 189718 266463 189770 266469
rect 189718 266405 189770 266411
rect 186070 255141 186122 255147
rect 186070 255083 186122 255089
rect 185974 255067 186026 255073
rect 185974 255009 186026 255015
rect 185782 246705 185834 246711
rect 185782 246647 185834 246653
rect 185686 242857 185738 242863
rect 185686 242799 185738 242805
rect 185590 242783 185642 242789
rect 185590 242725 185642 242731
rect 185602 220335 185630 242725
rect 185588 220326 185644 220335
rect 185588 220261 185644 220270
rect 185492 198274 185548 198283
rect 185492 198209 185548 198218
rect 184436 196794 184492 196803
rect 184436 196729 184492 196738
rect 184340 196054 184396 196063
rect 184340 195989 184396 195998
rect 183094 195867 183146 195873
rect 183094 195809 183146 195815
rect 182998 149765 183050 149771
rect 182998 149707 183050 149713
rect 183106 143999 183134 195809
rect 184534 195793 184586 195799
rect 184534 195735 184586 195741
rect 184438 195719 184490 195725
rect 184438 195661 184490 195667
rect 184342 195645 184394 195651
rect 184342 195587 184394 195593
rect 184354 195323 184382 195587
rect 184340 195314 184396 195323
rect 184340 195249 184396 195258
rect 184450 194435 184478 195661
rect 184436 194426 184492 194435
rect 184436 194361 184492 194370
rect 184546 193843 184574 195735
rect 184532 193834 184588 193843
rect 184532 193769 184588 193778
rect 184630 192981 184682 192987
rect 184436 192946 184492 192955
rect 184630 192923 184682 192929
rect 184436 192881 184492 192890
rect 184534 192907 184586 192913
rect 184342 192833 184394 192839
rect 184342 192775 184394 192781
rect 184354 192363 184382 192775
rect 184450 192765 184478 192881
rect 184534 192849 184586 192855
rect 184438 192759 184490 192765
rect 184438 192701 184490 192707
rect 184340 192354 184396 192363
rect 184340 192289 184396 192298
rect 184546 191475 184574 192849
rect 184532 191466 184588 191475
rect 184532 191401 184588 191410
rect 184642 190735 184670 192923
rect 184628 190726 184684 190735
rect 184628 190661 184684 190670
rect 184534 190095 184586 190101
rect 184534 190037 184586 190043
rect 184342 190021 184394 190027
rect 184340 189986 184342 189995
rect 184394 189986 184396 189995
rect 184340 189921 184396 189930
rect 184438 189947 184490 189953
rect 184438 189889 184490 189895
rect 184342 189873 184394 189879
rect 184342 189815 184394 189821
rect 184354 188515 184382 189815
rect 184340 188506 184396 188515
rect 184340 188441 184396 188450
rect 184450 187627 184478 189889
rect 184546 189255 184574 190037
rect 184532 189246 184588 189255
rect 184532 189181 184588 189190
rect 184436 187618 184492 187627
rect 184436 187553 184492 187562
rect 184438 187209 184490 187215
rect 184438 187151 184490 187157
rect 184342 187061 184394 187067
rect 184342 187003 184394 187009
rect 184354 186887 184382 187003
rect 184340 186878 184396 186887
rect 184340 186813 184396 186822
rect 184450 186147 184478 187151
rect 184534 187135 184586 187141
rect 184534 187077 184586 187083
rect 184436 186138 184492 186147
rect 184436 186073 184492 186082
rect 184546 184667 184574 187077
rect 184630 186987 184682 186993
rect 184630 186929 184682 186935
rect 184642 185407 184670 186929
rect 184628 185398 184684 185407
rect 184628 185333 184684 185342
rect 184532 184658 184588 184667
rect 184532 184593 184588 184602
rect 184342 184323 184394 184329
rect 184342 184265 184394 184271
rect 184354 183927 184382 184265
rect 184438 184249 184490 184255
rect 184438 184191 184490 184197
rect 184340 183918 184396 183927
rect 184340 183853 184396 183862
rect 184450 181559 184478 184191
rect 184436 181550 184492 181559
rect 184436 181485 184492 181494
rect 184630 181437 184682 181443
rect 184630 181379 184682 181385
rect 184342 181363 184394 181369
rect 184342 181305 184394 181311
rect 184354 180819 184382 181305
rect 184438 181289 184490 181295
rect 184438 181231 184490 181237
rect 184340 180810 184396 180819
rect 184340 180745 184396 180754
rect 184450 180079 184478 181231
rect 184534 181215 184586 181221
rect 184534 181157 184586 181163
rect 184436 180070 184492 180079
rect 184436 180005 184492 180014
rect 184546 178599 184574 181157
rect 184642 179339 184670 181379
rect 185494 180105 185546 180111
rect 185494 180047 185546 180053
rect 184628 179330 184684 179339
rect 184628 179265 184684 179274
rect 184532 178590 184588 178599
rect 184438 178551 184490 178557
rect 184532 178525 184588 178534
rect 184438 178493 184490 178499
rect 184342 178403 184394 178409
rect 184342 178345 184394 178351
rect 184354 177119 184382 178345
rect 184450 177711 184478 178493
rect 184534 178477 184586 178483
rect 184534 178419 184586 178425
rect 184436 177702 184492 177711
rect 184436 177637 184492 177646
rect 184340 177110 184396 177119
rect 184340 177045 184396 177054
rect 184546 176231 184574 178419
rect 184532 176222 184588 176231
rect 184532 176157 184588 176166
rect 184342 175665 184394 175671
rect 184340 175630 184342 175639
rect 184394 175630 184396 175639
rect 184340 175565 184396 175574
rect 184438 175591 184490 175597
rect 184438 175533 184490 175539
rect 184450 174011 184478 175533
rect 184436 174002 184492 174011
rect 184436 173937 184492 173946
rect 184534 172779 184586 172785
rect 184534 172721 184586 172727
rect 184342 172631 184394 172637
rect 184342 172573 184394 172579
rect 184354 171791 184382 172573
rect 184438 172557 184490 172563
rect 184546 172531 184574 172721
rect 184630 172705 184682 172711
rect 184630 172647 184682 172653
rect 184438 172499 184490 172505
rect 184532 172522 184588 172531
rect 184340 171782 184396 171791
rect 184340 171717 184396 171726
rect 184450 170903 184478 172499
rect 184532 172457 184588 172466
rect 184436 170894 184492 170903
rect 184436 170829 184492 170838
rect 184642 170311 184670 172647
rect 184628 170302 184684 170311
rect 184628 170237 184684 170246
rect 184534 169893 184586 169899
rect 184534 169835 184586 169841
rect 184342 169819 184394 169825
rect 184342 169761 184394 169767
rect 184354 169423 184382 169761
rect 184438 169671 184490 169677
rect 184438 169613 184490 169619
rect 184340 169414 184396 169423
rect 184340 169349 184396 169358
rect 184450 167943 184478 169613
rect 184546 168683 184574 169835
rect 184630 169745 184682 169751
rect 184630 169687 184682 169693
rect 184532 168674 184588 168683
rect 184532 168609 184588 168618
rect 184436 167934 184492 167943
rect 184436 167869 184492 167878
rect 184642 167203 184670 169687
rect 184628 167194 184684 167203
rect 184628 167129 184684 167138
rect 184342 167007 184394 167013
rect 184342 166949 184394 166955
rect 184354 166463 184382 166949
rect 184438 166933 184490 166939
rect 184438 166875 184490 166881
rect 184340 166454 184396 166463
rect 184340 166389 184396 166398
rect 184450 165723 184478 166875
rect 184534 166859 184586 166865
rect 184534 166801 184586 166807
rect 184436 165714 184492 165723
rect 184436 165649 184492 165658
rect 184546 164835 184574 166801
rect 184532 164826 184588 164835
rect 184532 164761 184588 164770
rect 184534 164121 184586 164127
rect 184340 164086 184396 164095
rect 184534 164063 184586 164069
rect 184340 164021 184342 164030
rect 184394 164021 184396 164030
rect 184342 163989 184394 163995
rect 184438 163973 184490 163979
rect 184438 163915 184490 163921
rect 184342 163899 184394 163905
rect 184342 163841 184394 163847
rect 184354 162615 184382 163841
rect 184340 162606 184396 162615
rect 184340 162541 184396 162550
rect 184450 161875 184478 163915
rect 184546 163355 184574 164063
rect 184532 163346 184588 163355
rect 184532 163281 184588 163290
rect 184436 161866 184492 161875
rect 184436 161801 184492 161810
rect 184438 161235 184490 161241
rect 184438 161177 184490 161183
rect 184342 161013 184394 161019
rect 184450 160987 184478 161177
rect 184534 161161 184586 161167
rect 184534 161103 184586 161109
rect 184342 160955 184394 160961
rect 184436 160978 184492 160987
rect 184354 159507 184382 160955
rect 184436 160913 184492 160922
rect 184546 160395 184574 161103
rect 184630 161087 184682 161093
rect 184630 161029 184682 161035
rect 184532 160386 184588 160395
rect 184532 160321 184588 160330
rect 184340 159498 184396 159507
rect 184340 159433 184396 159442
rect 184642 158915 184670 161029
rect 184628 158906 184684 158915
rect 184628 158841 184684 158850
rect 184342 158423 184394 158429
rect 184342 158365 184394 158371
rect 184354 158027 184382 158365
rect 184438 158349 184490 158355
rect 184438 158291 184490 158297
rect 184340 158018 184396 158027
rect 184340 157953 184396 157962
rect 184450 157435 184478 158291
rect 184534 158275 184586 158281
rect 184534 158217 184586 158223
rect 184436 157426 184492 157435
rect 184436 157361 184492 157370
rect 184546 156547 184574 158217
rect 184630 158201 184682 158207
rect 184630 158143 184682 158149
rect 184532 156538 184588 156547
rect 184532 156473 184588 156482
rect 184642 155659 184670 158143
rect 184628 155650 184684 155659
rect 184628 155585 184684 155594
rect 184534 155537 184586 155543
rect 185506 155534 185534 180047
rect 185698 174751 185726 242799
rect 185794 182447 185822 246647
rect 185878 242709 185930 242715
rect 185878 242651 185930 242657
rect 185890 195854 185918 242651
rect 185986 204351 186014 255009
rect 186082 212047 186110 255083
rect 186550 254993 186602 254999
rect 186550 254935 186602 254941
rect 186358 252033 186410 252039
rect 186358 251975 186410 251981
rect 186262 246631 186314 246637
rect 186262 246573 186314 246579
rect 186166 246261 186218 246267
rect 186166 246203 186218 246209
rect 186068 212038 186124 212047
rect 186068 211973 186124 211982
rect 185972 204342 186028 204351
rect 185972 204277 186028 204286
rect 186178 202871 186206 246203
rect 186274 207311 186302 246573
rect 186370 210567 186398 251975
rect 186454 246557 186506 246563
rect 186454 246499 186506 246505
rect 186356 210558 186412 210567
rect 186356 210493 186412 210502
rect 186260 207302 186316 207311
rect 186260 207237 186316 207246
rect 186466 205979 186494 246499
rect 186562 213527 186590 254935
rect 186742 254919 186794 254925
rect 186742 254861 186794 254867
rect 186646 246483 186698 246489
rect 186646 246425 186698 246431
rect 186548 213518 186604 213527
rect 186548 213453 186604 213462
rect 186658 209087 186686 246425
rect 186754 215007 186782 254861
rect 187030 246409 187082 246415
rect 187030 246351 187082 246357
rect 186838 246335 186890 246341
rect 186838 246277 186890 246283
rect 186850 216487 186878 246277
rect 186934 244929 186986 244935
rect 186934 244871 186986 244877
rect 186946 221075 186974 244871
rect 186932 221066 186988 221075
rect 186932 221001 186988 221010
rect 187042 218115 187070 246351
rect 187124 243414 187180 243423
rect 187124 243349 187180 243358
rect 187138 227545 187166 243349
rect 187126 227539 187178 227545
rect 187126 227481 187178 227487
rect 187138 226139 187166 227481
rect 187126 226133 187178 226139
rect 187126 226075 187178 226081
rect 187028 218106 187084 218115
rect 187028 218041 187084 218050
rect 186836 216478 186892 216487
rect 186836 216413 186892 216422
rect 186740 214998 186796 215007
rect 186740 214933 186796 214942
rect 186644 209078 186700 209087
rect 186644 209013 186700 209022
rect 186452 205970 186508 205979
rect 186452 205905 186508 205914
rect 186164 202862 186220 202871
rect 186164 202797 186220 202806
rect 187234 199171 187262 266405
rect 192418 263810 192446 269249
rect 192598 269217 192650 269223
rect 192610 263824 192638 269217
rect 193090 263824 193118 269545
rect 192610 263796 192864 263824
rect 193090 263796 193344 263824
rect 193762 263810 193790 272061
rect 194228 269462 194284 269471
rect 194228 269397 194284 269406
rect 194242 263810 194270 269397
rect 194434 263824 194462 272209
rect 194722 272167 194750 278018
rect 195670 272235 195722 272241
rect 195670 272177 195722 272183
rect 194710 272161 194762 272167
rect 194710 272103 194762 272109
rect 195286 271939 195338 271945
rect 195286 271881 195338 271887
rect 195190 269867 195242 269873
rect 195190 269809 195242 269815
rect 194998 268461 195050 268467
rect 194998 268403 195050 268409
rect 195010 263824 195038 268403
rect 195202 268393 195230 269809
rect 195190 268387 195242 268393
rect 195190 268329 195242 268335
rect 195298 268245 195326 271881
rect 195286 268239 195338 268245
rect 195286 268181 195338 268187
rect 194434 263796 194736 263824
rect 195010 263796 195264 263824
rect 195682 263810 195710 272177
rect 195874 271945 195902 278018
rect 196628 272422 196684 272431
rect 196628 272357 196684 272366
rect 195862 271939 195914 271945
rect 195862 271881 195914 271887
rect 196342 271717 196394 271723
rect 196342 271659 196394 271665
rect 196148 269758 196204 269767
rect 196148 269693 196204 269702
rect 196162 263810 196190 269693
rect 196354 269651 196382 271659
rect 196342 269645 196394 269651
rect 196342 269587 196394 269593
rect 196642 263810 196670 272357
rect 196822 269497 196874 269503
rect 196822 269439 196874 269445
rect 196834 263824 196862 269439
rect 197122 269281 197150 278018
rect 198274 272241 198302 278018
rect 199220 272570 199276 272579
rect 199220 272505 199276 272514
rect 199126 272383 199178 272389
rect 199126 272325 199178 272331
rect 198262 272235 198314 272241
rect 198262 272177 198314 272183
rect 198550 271125 198602 271131
rect 198550 271067 198602 271073
rect 198070 269571 198122 269577
rect 198070 269513 198122 269519
rect 197398 269423 197450 269429
rect 197398 269365 197450 269371
rect 197110 269275 197162 269281
rect 197110 269217 197162 269223
rect 197410 263824 197438 269365
rect 196834 263796 197088 263824
rect 197410 263796 197664 263824
rect 198082 263810 198110 269513
rect 198562 263810 198590 271067
rect 199030 269349 199082 269355
rect 199030 269291 199082 269297
rect 199042 263810 199070 269291
rect 199138 267875 199166 272325
rect 199126 267869 199178 267875
rect 199126 267811 199178 267817
rect 199234 263824 199262 272505
rect 199426 271723 199454 278018
rect 200468 272718 200524 272727
rect 200468 272653 200524 272662
rect 199414 271717 199466 271723
rect 199414 271659 199466 271665
rect 199702 269719 199754 269725
rect 199702 269661 199754 269667
rect 199714 263824 199742 269661
rect 199234 263796 199488 263824
rect 199714 263796 199968 263824
rect 200482 263810 200510 272653
rect 200674 269355 200702 278018
rect 201622 272309 201674 272315
rect 201622 272251 201674 272257
rect 201526 271495 201578 271501
rect 201526 271437 201578 271443
rect 200950 269793 201002 269799
rect 200950 269735 201002 269741
rect 200662 269349 200714 269355
rect 200662 269291 200714 269297
rect 200962 263810 200990 269735
rect 201538 269725 201566 271437
rect 201526 269719 201578 269725
rect 201526 269661 201578 269667
rect 201142 268387 201194 268393
rect 201142 268329 201194 268335
rect 201154 263824 201182 268329
rect 201634 263824 201662 272251
rect 201826 271501 201854 278018
rect 201814 271495 201866 271501
rect 201814 271437 201866 271443
rect 202870 269941 202922 269947
rect 202870 269883 202922 269889
rect 202294 267869 202346 267875
rect 202294 267811 202346 267817
rect 201154 263796 201408 263824
rect 201634 263796 201888 263824
rect 202306 263810 202334 267811
rect 202882 263810 202910 269883
rect 202978 269429 203006 278018
rect 203542 272531 203594 272537
rect 203542 272473 203594 272479
rect 203350 270089 203402 270095
rect 203350 270031 203402 270037
rect 202966 269423 203018 269429
rect 202966 269365 203018 269371
rect 203362 263810 203390 270031
rect 203554 263824 203582 272473
rect 204022 272457 204074 272463
rect 204022 272399 204074 272405
rect 204034 263824 204062 272399
rect 204130 269503 204158 278018
rect 205378 272463 205406 278018
rect 206038 272679 206090 272685
rect 206038 272621 206090 272627
rect 205462 272605 205514 272611
rect 205462 272547 205514 272553
rect 205366 272457 205418 272463
rect 205366 272399 205418 272405
rect 205270 270163 205322 270169
rect 205270 270105 205322 270111
rect 204694 270015 204746 270021
rect 204694 269957 204746 269963
rect 204118 269497 204170 269503
rect 204118 269439 204170 269445
rect 203554 263796 203808 263824
rect 204034 263796 204288 263824
rect 204706 263810 204734 269957
rect 205282 263810 205310 270105
rect 205474 263824 205502 272547
rect 205942 271421 205994 271427
rect 205942 271363 205994 271369
rect 205750 271273 205802 271279
rect 205750 271215 205802 271221
rect 205762 269799 205790 271215
rect 205846 271199 205898 271205
rect 205846 271141 205898 271147
rect 205858 269873 205886 271141
rect 205954 269947 205982 271363
rect 205942 269941 205994 269947
rect 205942 269883 205994 269889
rect 205846 269867 205898 269873
rect 205846 269809 205898 269815
rect 205750 269793 205802 269799
rect 205750 269735 205802 269741
rect 206050 263824 206078 272621
rect 206422 270237 206474 270243
rect 206422 270179 206474 270185
rect 206434 263824 206462 270179
rect 206530 269577 206558 278018
rect 207286 272975 207338 272981
rect 207286 272917 207338 272923
rect 207094 272753 207146 272759
rect 207094 272695 207146 272701
rect 206518 269571 206570 269577
rect 206518 269513 206570 269519
rect 205474 263796 205776 263824
rect 206050 263796 206208 263824
rect 206434 263796 206688 263824
rect 207106 263810 207134 272695
rect 207298 267875 207326 272917
rect 207682 272389 207710 278018
rect 207862 272827 207914 272833
rect 207862 272769 207914 272775
rect 207670 272383 207722 272389
rect 207670 272325 207722 272331
rect 207574 270311 207626 270317
rect 207574 270253 207626 270259
rect 207286 267869 207338 267875
rect 207286 267811 207338 267817
rect 207586 263810 207614 270253
rect 207874 263824 207902 272769
rect 208930 272315 208958 278018
rect 209398 273567 209450 273573
rect 209398 273509 209450 273515
rect 209014 272901 209066 272907
rect 209014 272843 209066 272849
rect 208918 272309 208970 272315
rect 208918 272251 208970 272257
rect 208342 270385 208394 270391
rect 208342 270327 208394 270333
rect 208354 263824 208382 270327
rect 207874 263796 208128 263824
rect 208354 263796 208608 263824
rect 209026 263810 209054 272843
rect 209410 267949 209438 273509
rect 209686 273419 209738 273425
rect 209686 273361 209738 273367
rect 209590 273271 209642 273277
rect 209590 273213 209642 273219
rect 209602 270391 209630 273213
rect 209698 270507 209726 273361
rect 209878 273345 209930 273351
rect 209878 273287 209930 273293
rect 209782 273197 209834 273203
rect 209782 273139 209834 273145
rect 209684 270498 209740 270507
rect 209684 270433 209740 270442
rect 209590 270385 209642 270391
rect 209590 270327 209642 270333
rect 209794 270243 209822 273139
rect 209782 270237 209834 270243
rect 209782 270179 209834 270185
rect 209890 270169 209918 273287
rect 209974 273123 210026 273129
rect 209974 273065 210026 273071
rect 209878 270163 209930 270169
rect 209878 270105 209930 270111
rect 209398 267943 209450 267949
rect 209398 267885 209450 267891
rect 209494 267869 209546 267875
rect 209494 267811 209546 267817
rect 209506 263810 209534 267811
rect 209986 263810 210014 273065
rect 210082 272537 210110 278018
rect 210166 273049 210218 273055
rect 210166 272991 210218 272997
rect 210070 272531 210122 272537
rect 210070 272473 210122 272479
rect 210178 267854 210206 272991
rect 211234 272833 211262 278018
rect 211222 272827 211274 272833
rect 211222 272769 211274 272775
rect 212482 271427 212510 278018
rect 213634 272685 213662 278018
rect 213622 272679 213674 272685
rect 213622 272621 213674 272627
rect 214786 272611 214814 278018
rect 216034 272981 216062 278018
rect 217186 273129 217214 278018
rect 217174 273123 217226 273129
rect 217174 273065 217226 273071
rect 218338 273055 218366 278018
rect 219094 273493 219146 273499
rect 219094 273435 219146 273441
rect 218326 273049 218378 273055
rect 218326 272991 218378 272997
rect 216022 272975 216074 272981
rect 216022 272917 216074 272923
rect 214774 272605 214826 272611
rect 214774 272547 214826 272553
rect 213046 272087 213098 272093
rect 213046 272029 213098 272035
rect 212854 272013 212906 272019
rect 212854 271955 212906 271961
rect 212566 271569 212618 271575
rect 212566 271511 212618 271517
rect 212470 271421 212522 271427
rect 212470 271363 212522 271369
rect 211894 270459 211946 270465
rect 211894 270401 211946 270407
rect 211414 270237 211466 270243
rect 211414 270179 211466 270185
rect 210742 268165 210794 268171
rect 210742 268107 210794 268113
rect 210178 267826 210302 267854
rect 210274 263824 210302 267826
rect 210754 263824 210782 268107
rect 210274 263796 210528 263824
rect 210754 263796 211008 263824
rect 211426 263810 211454 270179
rect 211906 263810 211934 270401
rect 212578 270317 212606 271511
rect 212758 271347 212810 271353
rect 212758 271289 212810 271295
rect 212662 270533 212714 270539
rect 212662 270475 212714 270481
rect 212566 270311 212618 270317
rect 212566 270253 212618 270259
rect 212374 270163 212426 270169
rect 212374 270105 212426 270111
rect 212386 263810 212414 270105
rect 212674 263824 212702 270475
rect 212770 270243 212798 271289
rect 212758 270237 212810 270243
rect 212758 270179 212810 270185
rect 212866 270169 212894 271955
rect 212950 271643 213002 271649
rect 212950 271585 213002 271591
rect 212854 270163 212906 270169
rect 212854 270105 212906 270111
rect 212962 270095 212990 271585
rect 212950 270089 213002 270095
rect 212950 270031 213002 270037
rect 213058 270021 213086 272029
rect 218998 271939 219050 271945
rect 218998 271881 219050 271887
rect 218902 271717 218954 271723
rect 218902 271659 218954 271665
rect 214966 270681 215018 270687
rect 214966 270623 215018 270629
rect 213814 270607 213866 270613
rect 213814 270549 213866 270555
rect 213046 270015 213098 270021
rect 213046 269957 213098 269963
rect 213332 269906 213388 269915
rect 213332 269841 213388 269850
rect 212674 263796 212928 263824
rect 213346 263810 213374 269841
rect 213826 263810 213854 270549
rect 214292 270498 214348 270507
rect 214292 270433 214348 270442
rect 214306 263810 214334 270433
rect 214486 269201 214538 269207
rect 214486 269143 214538 269149
rect 214498 263824 214526 269143
rect 214978 263824 215006 270623
rect 216886 270385 216938 270391
rect 216886 270327 216938 270333
rect 215734 269127 215786 269133
rect 215734 269069 215786 269075
rect 214498 263796 214752 263824
rect 214978 263796 215232 263824
rect 215746 263810 215774 269069
rect 216214 269053 216266 269059
rect 216214 268995 216266 269001
rect 216226 263810 216254 268995
rect 216694 268979 216746 268985
rect 216694 268921 216746 268927
rect 216706 263810 216734 268921
rect 216898 263824 216926 270327
rect 217366 268905 217418 268911
rect 217366 268847 217418 268853
rect 217378 263824 217406 268847
rect 218134 268831 218186 268837
rect 218134 268773 218186 268779
rect 216898 263796 217152 263824
rect 217378 263796 217632 263824
rect 218146 263810 218174 268773
rect 218614 268239 218666 268245
rect 218614 268181 218666 268187
rect 218626 263810 218654 268181
rect 218914 268097 218942 271659
rect 218902 268091 218954 268097
rect 218902 268033 218954 268039
rect 219010 268023 219038 271881
rect 219106 268393 219134 273435
rect 219586 273351 219614 278018
rect 219574 273345 219626 273351
rect 219574 273287 219626 273293
rect 220738 272907 220766 278018
rect 220726 272901 220778 272907
rect 220726 272843 220778 272849
rect 221890 271057 221918 278018
rect 222070 272235 222122 272241
rect 222070 272177 222122 272183
rect 221974 271495 222026 271501
rect 221974 271437 222026 271443
rect 221878 271051 221930 271057
rect 221878 270993 221930 270999
rect 221014 270015 221066 270021
rect 221014 269957 221066 269963
rect 220534 269645 220586 269651
rect 220534 269587 220586 269593
rect 219286 268757 219338 268763
rect 219286 268699 219338 268705
rect 219094 268387 219146 268393
rect 219094 268329 219146 268335
rect 218998 268017 219050 268023
rect 218998 267959 219050 267965
rect 218902 267943 218954 267949
rect 218902 267885 218954 267891
rect 218914 263824 218942 267885
rect 219298 263824 219326 268699
rect 219958 268683 220010 268689
rect 219958 268625 220010 268631
rect 218914 263796 219072 263824
rect 219298 263796 219552 263824
rect 219970 263810 219998 268625
rect 220546 263810 220574 269587
rect 221026 263810 221054 269957
rect 221782 268609 221834 268615
rect 221782 268551 221834 268557
rect 221206 268535 221258 268541
rect 221206 268477 221258 268483
rect 221218 263824 221246 268477
rect 221794 263824 221822 268551
rect 221986 268171 222014 271437
rect 222082 268245 222110 272177
rect 222262 272161 222314 272167
rect 222262 272103 222314 272109
rect 222166 271791 222218 271797
rect 222166 271733 222218 271739
rect 222070 268239 222122 268245
rect 222070 268181 222122 268187
rect 221974 268165 222026 268171
rect 221974 268107 222026 268113
rect 222178 267875 222206 271733
rect 222274 267949 222302 272103
rect 223042 270983 223070 278018
rect 223030 270977 223082 270983
rect 223030 270919 223082 270925
rect 224290 270909 224318 278018
rect 224278 270903 224330 270909
rect 224278 270845 224330 270851
rect 225442 270835 225470 278018
rect 225430 270829 225482 270835
rect 225430 270771 225482 270777
rect 226594 270761 226622 278018
rect 227842 273499 227870 278018
rect 227830 273493 227882 273499
rect 227830 273435 227882 273441
rect 228994 272167 229022 278018
rect 230146 273573 230174 278018
rect 230134 273567 230186 273573
rect 230134 273509 230186 273515
rect 228982 272161 229034 272167
rect 228982 272103 229034 272109
rect 231394 271945 231422 278018
rect 232546 272019 232574 278018
rect 233698 272759 233726 278018
rect 233686 272753 233738 272759
rect 233686 272695 233738 272701
rect 234550 272531 234602 272537
rect 234550 272473 234602 272479
rect 232630 272457 232682 272463
rect 232630 272399 232682 272405
rect 232534 272013 232586 272019
rect 232534 271955 232586 271961
rect 231382 271939 231434 271945
rect 231382 271881 231434 271887
rect 227158 271865 227210 271871
rect 227158 271807 227210 271813
rect 226582 270755 226634 270761
rect 226582 270697 226634 270703
rect 225526 270311 225578 270317
rect 225526 270253 225578 270259
rect 222838 270163 222890 270169
rect 222838 270105 222890 270111
rect 222358 269719 222410 269725
rect 222358 269661 222410 269667
rect 222262 267943 222314 267949
rect 222262 267885 222314 267891
rect 222166 267869 222218 267875
rect 222166 267811 222218 267817
rect 221218 263796 221472 263824
rect 221794 263796 221952 263824
rect 222370 263810 222398 269661
rect 222850 263810 222878 270105
rect 224758 270089 224810 270095
rect 224758 270031 224810 270037
rect 224086 269941 224138 269947
rect 224086 269883 224138 269889
rect 223414 268461 223466 268467
rect 223414 268403 223466 268409
rect 223426 263810 223454 268403
rect 223606 268313 223658 268319
rect 223606 268255 223658 268261
rect 223618 263824 223646 268255
rect 224098 263824 224126 269883
rect 223618 263796 223872 263824
rect 224098 263796 224352 263824
rect 224770 263810 224798 270031
rect 225238 269793 225290 269799
rect 225238 269735 225290 269741
rect 225250 263810 225278 269735
rect 225538 263824 225566 270253
rect 226678 270237 226730 270243
rect 226678 270179 226730 270185
rect 226006 269867 226058 269873
rect 226006 269809 226058 269815
rect 226018 263824 226046 269809
rect 225538 263796 225792 263824
rect 226018 263796 226272 263824
rect 226690 263810 226718 270179
rect 227170 263810 227198 271807
rect 232150 269497 232202 269503
rect 232150 269439 232202 269445
rect 231958 269423 232010 269429
rect 231958 269365 232010 269371
rect 230998 269349 231050 269355
rect 230998 269291 231050 269297
rect 229558 269275 229610 269281
rect 229558 269217 229610 269223
rect 227830 268313 227882 268319
rect 227830 268255 227882 268261
rect 227638 267869 227690 267875
rect 227638 267811 227690 267817
rect 227650 263810 227678 267811
rect 227842 263824 227870 268255
rect 229078 268017 229130 268023
rect 229078 267959 229130 267965
rect 228406 267943 228458 267949
rect 228406 267885 228458 267891
rect 228418 263824 228446 267885
rect 227842 263796 228096 263824
rect 228418 263796 228672 263824
rect 229090 263810 229118 267959
rect 229570 263810 229598 269217
rect 230038 268239 230090 268245
rect 230038 268181 230090 268187
rect 230050 263810 230078 268181
rect 230518 268091 230570 268097
rect 230518 268033 230570 268039
rect 230530 264120 230558 268033
rect 230482 264092 230558 264120
rect 230482 263810 230510 264092
rect 231010 263810 231038 269291
rect 231478 268165 231530 268171
rect 231478 268107 231530 268113
rect 231490 263810 231518 268107
rect 231970 263810 231998 269365
rect 232162 263824 232190 269439
rect 232642 263824 232670 272399
rect 233878 272383 233930 272389
rect 233878 272325 233930 272331
rect 233398 269571 233450 269577
rect 233398 269513 233450 269519
rect 232162 263796 232416 263824
rect 232642 263796 232896 263824
rect 233410 263810 233438 269513
rect 233890 263810 233918 272325
rect 234358 272309 234410 272315
rect 234358 272251 234410 272257
rect 234370 263810 234398 272251
rect 234562 263824 234590 272473
rect 234946 272315 234974 278018
rect 235030 272827 235082 272833
rect 235030 272769 235082 272775
rect 234934 272309 234986 272315
rect 234934 272251 234986 272257
rect 235042 263824 235070 272769
rect 236098 272537 236126 278018
rect 236950 272975 237002 272981
rect 236950 272917 237002 272923
rect 236278 272679 236330 272685
rect 236278 272621 236330 272627
rect 236086 272531 236138 272537
rect 236086 272473 236138 272479
rect 235702 271421 235754 271427
rect 235702 271363 235754 271369
rect 234562 263796 234816 263824
rect 235042 263796 235296 263824
rect 235714 263810 235742 271363
rect 236290 263810 236318 272621
rect 236470 272605 236522 272611
rect 236470 272547 236522 272553
rect 236482 263824 236510 272547
rect 236962 263824 236990 272917
rect 237250 271279 237278 278018
rect 237622 273123 237674 273129
rect 237622 273065 237674 273071
rect 237238 271273 237290 271279
rect 237238 271215 237290 271221
rect 236482 263796 236736 263824
rect 236962 263796 237216 263824
rect 237634 263810 237662 273065
rect 238102 273049 238154 273055
rect 238102 272991 238154 272997
rect 238114 263810 238142 272991
rect 238498 271205 238526 278018
rect 238678 273345 238730 273351
rect 238678 273287 238730 273293
rect 238486 271199 238538 271205
rect 238486 271141 238538 271147
rect 238690 263810 238718 273287
rect 239158 272901 239210 272907
rect 239158 272843 239210 272849
rect 239170 263824 239198 272843
rect 239350 271051 239402 271057
rect 239350 270993 239402 270999
rect 239542 271051 239594 271057
rect 239542 270993 239594 270999
rect 239136 263796 239198 263824
rect 239362 263824 239390 270993
rect 239554 270761 239582 270993
rect 239650 270761 239678 278018
rect 240802 271131 240830 278018
rect 240790 271125 240842 271131
rect 240790 271067 240842 271073
rect 241954 271057 241982 278018
rect 242902 273567 242954 273573
rect 242902 273509 242954 273515
rect 242134 273493 242186 273499
rect 242134 273435 242186 273441
rect 241270 271051 241322 271057
rect 241270 270993 241322 270999
rect 241942 271051 241994 271057
rect 241942 270993 241994 270999
rect 240022 270977 240074 270983
rect 240022 270919 240074 270925
rect 239542 270755 239594 270761
rect 239542 270697 239594 270703
rect 239638 270755 239690 270761
rect 239638 270697 239690 270703
rect 239362 263796 239616 263824
rect 240034 263810 240062 270919
rect 240502 270903 240554 270909
rect 240502 270845 240554 270851
rect 240514 263810 240542 270845
rect 241078 270829 241130 270835
rect 241078 270771 241130 270777
rect 241090 263810 241118 270771
rect 241282 263824 241310 270993
rect 242146 263824 242174 273435
rect 242422 272161 242474 272167
rect 242422 272103 242474 272109
rect 241282 263796 241536 263824
rect 242016 263796 242174 263824
rect 242434 263810 242462 272103
rect 242914 263810 242942 273509
rect 243094 271939 243146 271945
rect 243094 271881 243146 271887
rect 243106 263824 243134 271881
rect 243202 270983 243230 278018
rect 244054 272753 244106 272759
rect 244054 272695 244106 272701
rect 243670 272013 243722 272019
rect 243670 271955 243722 271961
rect 243190 270977 243242 270983
rect 243190 270919 243242 270925
rect 243682 263824 243710 271955
rect 244066 263824 244094 272695
rect 244354 270909 244382 278018
rect 245302 272531 245354 272537
rect 245302 272473 245354 272479
rect 244822 272309 244874 272315
rect 244822 272251 244874 272257
rect 244342 270903 244394 270909
rect 244342 270845 244394 270851
rect 243106 263796 243360 263824
rect 243682 263796 243936 263824
rect 244066 263796 244368 263824
rect 244834 263810 244862 272251
rect 245314 263810 245342 272473
rect 245506 270835 245534 278018
rect 245590 271273 245642 271279
rect 245590 271215 245642 271221
rect 245494 270829 245546 270835
rect 245494 270771 245546 270777
rect 245602 263824 245630 271215
rect 246070 271199 246122 271205
rect 246070 271141 246122 271147
rect 246082 263824 246110 271141
rect 246754 270761 246782 278018
rect 247222 271125 247274 271131
rect 247222 271067 247274 271073
rect 246454 270755 246506 270761
rect 246454 270697 246506 270703
rect 246742 270755 246794 270761
rect 246742 270697 246794 270703
rect 246466 263824 246494 270697
rect 245602 263796 245760 263824
rect 246082 263796 246336 263824
rect 246466 263796 246768 263824
rect 247234 263810 247262 271067
rect 247702 271051 247754 271057
rect 247702 270993 247754 270999
rect 247714 263810 247742 270993
rect 247906 268393 247934 278018
rect 247990 270977 248042 270983
rect 247990 270919 248042 270925
rect 247894 268387 247946 268393
rect 247894 268329 247946 268335
rect 248002 263824 248030 270919
rect 248662 270903 248714 270909
rect 248662 270845 248714 270851
rect 248002 263796 248160 263824
rect 248674 263810 248702 270845
rect 249058 269651 249086 278018
rect 250320 278004 250526 278032
rect 249142 270829 249194 270835
rect 249142 270771 249194 270777
rect 250498 270780 250526 278004
rect 249046 269645 249098 269651
rect 249046 269587 249098 269593
rect 249154 263810 249182 270771
rect 249622 270755 249674 270761
rect 250498 270752 250718 270780
rect 249622 270697 249674 270703
rect 249634 263810 249662 270697
rect 250294 269645 250346 269651
rect 250294 269587 250346 269593
rect 249814 268387 249866 268393
rect 249814 268329 249866 268335
rect 249826 263824 249854 268329
rect 250306 263824 250334 269587
rect 250690 263824 250718 270752
rect 251458 263824 251486 278018
rect 252322 278004 252624 278032
rect 252322 263824 252350 278004
rect 253366 269127 253418 269133
rect 253366 269069 253418 269075
rect 253174 268535 253226 268541
rect 253174 268477 253226 268483
rect 252694 268091 252746 268097
rect 252694 268033 252746 268039
rect 252706 263824 252734 268033
rect 253186 263824 253214 268477
rect 249826 263796 250080 263824
rect 250306 263796 250560 263824
rect 250690 263796 250992 263824
rect 251458 263796 251568 263824
rect 252048 263796 252350 263824
rect 252480 263796 252734 263824
rect 252960 263796 253214 263824
rect 253378 263810 253406 269069
rect 253762 268097 253790 278018
rect 253942 270459 253994 270465
rect 253942 270401 253994 270407
rect 253750 268091 253802 268097
rect 253750 268033 253802 268039
rect 253954 263810 253982 270401
rect 254614 268683 254666 268689
rect 254614 268625 254666 268631
rect 254626 263824 254654 268625
rect 255010 268541 255038 278018
rect 255286 270311 255338 270317
rect 255286 270253 255338 270259
rect 254998 268535 255050 268541
rect 254998 268477 255050 268483
rect 255094 268387 255146 268393
rect 255094 268329 255146 268335
rect 255106 263824 255134 268329
rect 254400 263796 254654 263824
rect 254880 263796 255134 263824
rect 255298 263810 255326 270253
rect 255766 269645 255818 269651
rect 255766 269587 255818 269593
rect 255778 263810 255806 269587
rect 256162 269133 256190 278018
rect 257314 270465 257342 278018
rect 257302 270459 257354 270465
rect 257302 270401 257354 270407
rect 256246 269941 256298 269947
rect 256246 269883 256298 269889
rect 256150 269127 256202 269133
rect 256150 269069 256202 269075
rect 256258 263810 256286 269883
rect 258166 269719 258218 269725
rect 258166 269661 258218 269667
rect 257686 269349 257738 269355
rect 257686 269291 257738 269297
rect 257494 268831 257546 268837
rect 257494 268773 257546 268779
rect 257014 268535 257066 268541
rect 257014 268477 257066 268483
rect 257026 263824 257054 268477
rect 257506 263824 257534 268773
rect 256800 263796 257054 263824
rect 257280 263796 257534 263824
rect 257698 263810 257726 269291
rect 258178 263810 258206 269661
rect 258562 268689 258590 278018
rect 258646 269571 258698 269577
rect 258646 269513 258698 269519
rect 258550 268683 258602 268689
rect 258550 268625 258602 268631
rect 258658 263810 258686 269513
rect 259414 268979 259466 268985
rect 259414 268921 259466 268927
rect 259426 263824 259454 268921
rect 259714 268393 259742 278018
rect 260866 270317 260894 278018
rect 260854 270311 260906 270317
rect 260854 270253 260906 270259
rect 261238 270237 261290 270243
rect 261238 270179 261290 270185
rect 260566 269867 260618 269873
rect 260566 269809 260618 269815
rect 259894 269793 259946 269799
rect 259894 269735 259946 269741
rect 259702 268387 259754 268393
rect 259702 268329 259754 268335
rect 259906 263824 259934 269735
rect 260086 269497 260138 269503
rect 260086 269439 260138 269445
rect 259200 263796 259454 263824
rect 259680 263796 259934 263824
rect 260098 263810 260126 269439
rect 260578 263810 260606 269809
rect 261250 263824 261278 270179
rect 261814 270015 261866 270021
rect 261814 269957 261866 269963
rect 261826 263824 261854 269957
rect 262114 269651 262142 278018
rect 262966 270459 263018 270465
rect 262966 270401 263018 270407
rect 262486 270385 262538 270391
rect 262486 270327 262538 270333
rect 262102 269645 262154 269651
rect 262102 269587 262154 269593
rect 262006 269201 262058 269207
rect 262006 269143 262058 269149
rect 261024 263796 261278 263824
rect 261600 263796 261854 263824
rect 262018 263810 262046 269143
rect 262498 263810 262526 270327
rect 262978 263810 263006 270401
rect 263266 269947 263294 278018
rect 263254 269941 263306 269947
rect 263254 269883 263306 269889
rect 263638 268905 263690 268911
rect 263638 268847 263690 268853
rect 263650 263824 263678 268847
rect 264418 268541 264446 278018
rect 265366 270163 265418 270169
rect 265366 270105 265418 270111
rect 264694 270089 264746 270095
rect 264694 270031 264746 270037
rect 264406 268535 264458 268541
rect 264406 268477 264458 268483
rect 264118 268091 264170 268097
rect 264118 268033 264170 268039
rect 264130 263824 264158 268033
rect 264706 263824 264734 270031
rect 264886 269941 264938 269947
rect 264886 269883 264938 269889
rect 263424 263796 263678 263824
rect 263904 263796 264158 263824
rect 264432 263796 264734 263824
rect 264898 263810 264926 269883
rect 265378 263810 265406 270105
rect 265666 268837 265694 278018
rect 266518 269423 266570 269429
rect 266518 269365 266570 269371
rect 266038 269127 266090 269133
rect 266038 269069 266090 269075
rect 265654 268831 265706 268837
rect 265654 268773 265706 268779
rect 266050 263824 266078 269069
rect 266530 263824 266558 269365
rect 266818 269355 266846 278018
rect 267970 269725 267998 278018
rect 267958 269719 268010 269725
rect 267958 269661 268010 269667
rect 268630 269719 268682 269725
rect 268630 269661 268682 269667
rect 267766 269645 267818 269651
rect 267766 269587 267818 269593
rect 266806 269349 266858 269355
rect 266806 269291 266858 269297
rect 266806 268609 266858 268615
rect 266806 268551 266858 268557
rect 265824 263796 266078 263824
rect 266304 263796 266558 263824
rect 266818 263810 266846 268551
rect 267286 268535 267338 268541
rect 267286 268477 267338 268483
rect 267298 263810 267326 268477
rect 267778 263824 267806 269587
rect 268438 268757 268490 268763
rect 268438 268699 268490 268705
rect 268450 263824 268478 268699
rect 267744 263796 267806 263824
rect 268224 263796 268478 263824
rect 268642 263810 268670 269661
rect 269122 269577 269150 278018
rect 270262 272605 270314 272611
rect 270262 272547 270314 272553
rect 269206 270681 269258 270687
rect 269206 270623 269258 270629
rect 269110 269571 269162 269577
rect 269110 269513 269162 269519
rect 269218 263810 269246 270623
rect 269686 269201 269738 269207
rect 269686 269143 269738 269149
rect 269698 263810 269726 269143
rect 270274 263824 270302 272547
rect 270370 268985 270398 278018
rect 270550 272457 270602 272463
rect 270550 272399 270602 272405
rect 270358 268979 270410 268985
rect 270358 268921 270410 268927
rect 270144 263796 270302 263824
rect 270562 263824 270590 272399
rect 271030 272013 271082 272019
rect 271030 271955 271082 271961
rect 270562 263796 270624 263824
rect 271042 263810 271070 271955
rect 271522 269799 271550 278018
rect 272278 272531 272330 272537
rect 272278 272473 272330 272479
rect 271510 269793 271562 269799
rect 271510 269735 271562 269741
rect 271702 269719 271754 269725
rect 271702 269661 271754 269667
rect 271510 269571 271562 269577
rect 271510 269513 271562 269519
rect 271522 263810 271550 269513
rect 271714 269429 271742 269661
rect 271702 269423 271754 269429
rect 271702 269365 271754 269371
rect 272290 263824 272318 272473
rect 272674 269503 272702 278018
rect 272758 272383 272810 272389
rect 272758 272325 272810 272331
rect 272662 269497 272714 269503
rect 272662 269439 272714 269445
rect 272770 263824 272798 272325
rect 273430 272309 273482 272315
rect 273430 272251 273482 272257
rect 272950 269497 273002 269503
rect 272950 269439 273002 269445
rect 272064 263796 272318 263824
rect 272544 263796 272798 263824
rect 272962 263810 272990 269439
rect 273442 263810 273470 272251
rect 273922 269873 273950 278018
rect 274198 272975 274250 272981
rect 274198 272917 274250 272923
rect 273910 269867 273962 269873
rect 273910 269809 273962 269815
rect 274210 263824 274238 272917
rect 275074 270243 275102 278018
rect 275158 273567 275210 273573
rect 275158 273509 275210 273515
rect 275062 270237 275114 270243
rect 275062 270179 275114 270185
rect 274678 269423 274730 269429
rect 274678 269365 274730 269371
rect 274690 263824 274718 269365
rect 275170 263824 275198 273509
rect 275350 273419 275402 273425
rect 275350 273361 275402 273367
rect 273936 263796 274238 263824
rect 274464 263796 274718 263824
rect 274944 263796 275198 263824
rect 275362 263810 275390 273361
rect 276226 270021 276254 278018
rect 276310 272235 276362 272241
rect 276310 272177 276362 272183
rect 276214 270015 276266 270021
rect 276214 269957 276266 269963
rect 275830 269349 275882 269355
rect 275830 269291 275882 269297
rect 275842 263810 275870 269291
rect 276322 263810 276350 272177
rect 277078 272161 277130 272167
rect 277078 272103 277130 272109
rect 277090 263824 277118 272103
rect 277474 269281 277502 278018
rect 277750 273493 277802 273499
rect 277750 273435 277802 273441
rect 277462 269275 277514 269281
rect 277462 269217 277514 269223
rect 277558 268683 277610 268689
rect 277558 268625 277610 268631
rect 277570 263824 277598 268625
rect 276864 263796 277118 263824
rect 277344 263796 277598 263824
rect 277762 263810 277790 273435
rect 278230 273345 278282 273351
rect 278230 273287 278282 273293
rect 278242 263810 278270 273287
rect 278626 270391 278654 278018
rect 279670 273271 279722 273277
rect 279670 273213 279722 273219
rect 279286 270607 279338 270613
rect 279286 270549 279338 270555
rect 278614 270385 278666 270391
rect 278614 270327 278666 270333
rect 278902 268831 278954 268837
rect 278902 268773 278954 268779
rect 278914 263824 278942 268773
rect 279298 263824 279326 270549
rect 278688 263796 278942 263824
rect 279168 263796 279326 263824
rect 279682 263810 279710 273213
rect 279778 270465 279806 278018
rect 280150 270533 280202 270539
rect 280150 270475 280202 270481
rect 279766 270459 279818 270465
rect 279766 270401 279818 270407
rect 280162 263810 280190 270475
rect 280630 270459 280682 270465
rect 280630 270401 280682 270407
rect 280642 263810 280670 270401
rect 281026 268985 281054 278018
rect 281782 274825 281834 274831
rect 281782 274767 281834 274773
rect 281302 269053 281354 269059
rect 281302 268995 281354 269001
rect 281014 268979 281066 268985
rect 281014 268921 281066 268927
rect 281314 263824 281342 268995
rect 281794 263824 281822 274767
rect 282070 268979 282122 268985
rect 282070 268921 282122 268927
rect 281088 263796 281342 263824
rect 281568 263796 281822 263824
rect 282082 263810 282110 268921
rect 282178 268097 282206 278018
rect 283030 274899 283082 274905
rect 283030 274841 283082 274847
rect 282166 268091 282218 268097
rect 282166 268033 282218 268039
rect 282550 267869 282602 267875
rect 282550 267811 282602 267817
rect 282562 263810 282590 267811
rect 283042 263810 283070 274841
rect 283330 270021 283358 278018
rect 284182 270385 284234 270391
rect 284182 270327 284234 270333
rect 283318 270015 283370 270021
rect 283318 269957 283370 269963
rect 283702 269275 283754 269281
rect 283702 269217 283754 269223
rect 283714 263824 283742 269217
rect 284194 263824 284222 270327
rect 284470 270237 284522 270243
rect 284470 270179 284522 270185
rect 284482 269799 284510 270179
rect 284578 269947 284606 278018
rect 284758 274973 284810 274979
rect 284758 274915 284810 274921
rect 284566 269941 284618 269947
rect 284566 269883 284618 269889
rect 284470 269793 284522 269799
rect 284470 269735 284522 269741
rect 284770 263824 284798 274915
rect 285622 273197 285674 273203
rect 285622 273139 285674 273145
rect 284950 273123 285002 273129
rect 284950 273065 285002 273071
rect 283488 263796 283742 263824
rect 283968 263796 284222 263824
rect 284496 263796 284798 263824
rect 284962 263810 284990 273065
rect 285634 263824 285662 273139
rect 285730 270169 285758 278018
rect 286102 276453 286154 276459
rect 286102 276395 286154 276401
rect 285718 270163 285770 270169
rect 285718 270105 285770 270111
rect 286114 263824 286142 276395
rect 286774 273049 286826 273055
rect 286774 272991 286826 272997
rect 286294 270311 286346 270317
rect 286294 270253 286346 270259
rect 285408 263796 285662 263824
rect 285888 263796 286142 263824
rect 286306 263810 286334 270253
rect 286486 270015 286538 270021
rect 286486 269957 286538 269963
rect 286498 269577 286526 269957
rect 286486 269571 286538 269577
rect 286486 269513 286538 269519
rect 286786 263810 286814 272991
rect 286882 269133 286910 278018
rect 287350 276379 287402 276385
rect 287350 276321 287402 276327
rect 286870 269127 286922 269133
rect 286870 269069 286922 269075
rect 287362 263810 287390 276321
rect 287926 270163 287978 270169
rect 287926 270105 287978 270111
rect 287938 263824 287966 270105
rect 288034 270095 288062 278018
rect 288694 276305 288746 276311
rect 288694 276247 288746 276253
rect 288022 270089 288074 270095
rect 288022 270031 288074 270037
rect 288502 269571 288554 269577
rect 288502 269513 288554 269519
rect 288514 263824 288542 269513
rect 287808 263796 287966 263824
rect 288288 263796 288542 263824
rect 288706 263810 288734 276247
rect 289174 268831 289226 268837
rect 289174 268773 289226 268779
rect 289186 263810 289214 268773
rect 289282 268615 289310 278018
rect 290326 276231 290378 276237
rect 290326 276173 290378 276179
rect 289942 272901 289994 272907
rect 289942 272843 289994 272849
rect 289270 268609 289322 268615
rect 289270 268551 289322 268557
rect 289954 263824 289982 272843
rect 290338 263824 290366 276173
rect 290434 268541 290462 278018
rect 290614 269941 290666 269947
rect 290614 269883 290666 269889
rect 290422 268535 290474 268541
rect 290422 268477 290474 268483
rect 289728 263796 289982 263824
rect 290208 263796 290366 263824
rect 290626 263810 290654 269883
rect 291094 269867 291146 269873
rect 291094 269809 291146 269815
rect 291106 263810 291134 269809
rect 291586 269651 291614 278018
rect 291862 276157 291914 276163
rect 291862 276099 291914 276105
rect 291574 269645 291626 269651
rect 291574 269587 291626 269593
rect 291874 263824 291902 276099
rect 292246 272827 292298 272833
rect 292246 272769 292298 272775
rect 292258 263824 292286 272769
rect 292726 272753 292778 272759
rect 292726 272695 292778 272701
rect 292738 263824 292766 272695
rect 292834 268763 292862 278018
rect 293014 276083 293066 276089
rect 293014 276025 293066 276031
rect 292822 268757 292874 268763
rect 292822 268699 292874 268705
rect 291600 263796 291902 263824
rect 292032 263796 292286 263824
rect 292608 263796 292766 263824
rect 293026 263810 293054 276025
rect 293986 270243 294014 278018
rect 294646 276009 294698 276015
rect 294646 275951 294698 275957
rect 293974 270237 294026 270243
rect 293974 270179 294026 270185
rect 293974 269793 294026 269799
rect 293974 269735 294026 269741
rect 293494 269719 293546 269725
rect 293494 269661 293546 269667
rect 293506 263810 293534 269661
rect 293986 263810 294014 269735
rect 294658 263824 294686 275951
rect 295138 270687 295166 278018
rect 295894 275935 295946 275941
rect 295894 275877 295946 275883
rect 295414 272679 295466 272685
rect 295414 272621 295466 272627
rect 295126 270681 295178 270687
rect 295126 270623 295178 270629
rect 295222 270681 295274 270687
rect 295222 270623 295274 270629
rect 295234 270021 295262 270623
rect 295222 270015 295274 270021
rect 295222 269957 295274 269963
rect 295222 268757 295274 268763
rect 295222 268699 295274 268705
rect 295234 263824 295262 268699
rect 294432 263796 294686 263824
rect 295008 263796 295262 263824
rect 295426 263810 295454 272621
rect 295906 263810 295934 275877
rect 296386 269207 296414 278018
rect 296470 275861 296522 275867
rect 296470 275803 296522 275809
rect 296374 269201 296426 269207
rect 296374 269143 296426 269149
rect 296482 263824 296510 275803
rect 297334 275787 297386 275793
rect 297334 275729 297386 275735
rect 297046 269645 297098 269651
rect 297046 269587 297098 269593
rect 297058 263824 297086 269587
rect 296352 263796 296510 263824
rect 296832 263796 297086 263824
rect 297346 263810 297374 275729
rect 297538 272611 297566 278018
rect 297814 275713 297866 275719
rect 297814 275655 297866 275661
rect 297526 272605 297578 272611
rect 297526 272547 297578 272553
rect 297826 263810 297854 275655
rect 298486 272605 298538 272611
rect 298486 272547 298538 272553
rect 298102 272087 298154 272093
rect 298102 272029 298154 272035
rect 298006 271865 298058 271871
rect 298006 271807 298058 271813
rect 298018 267875 298046 271807
rect 298114 268985 298142 272029
rect 298198 270607 298250 270613
rect 298198 270549 298250 270555
rect 298390 270607 298442 270613
rect 298390 270549 298442 270555
rect 298210 270391 298238 270549
rect 298198 270385 298250 270391
rect 298198 270327 298250 270333
rect 298294 270311 298346 270317
rect 298294 270253 298346 270259
rect 298198 270089 298250 270095
rect 298198 270031 298250 270037
rect 298210 269577 298238 270031
rect 298198 269571 298250 269577
rect 298198 269513 298250 269519
rect 298306 269281 298334 270253
rect 298294 269275 298346 269281
rect 298294 269217 298346 269223
rect 298102 268979 298154 268985
rect 298102 268921 298154 268927
rect 298402 268911 298430 270549
rect 298390 268905 298442 268911
rect 298390 268847 298442 268853
rect 298006 267869 298058 267875
rect 298498 267854 298526 272547
rect 298690 272463 298718 278018
rect 298966 275639 299018 275645
rect 298966 275581 299018 275587
rect 298678 272457 298730 272463
rect 298678 272399 298730 272405
rect 298006 267811 298058 267817
rect 298306 267826 298526 267854
rect 298306 263810 298334 267826
rect 298978 263824 299006 275581
rect 299446 275491 299498 275497
rect 299446 275433 299498 275439
rect 299458 263824 299486 275433
rect 299938 272019 299966 278018
rect 300214 275565 300266 275571
rect 300214 275507 300266 275513
rect 299926 272013 299978 272019
rect 299926 271955 299978 271961
rect 300118 271865 300170 271871
rect 300118 271807 300170 271813
rect 299638 269571 299690 269577
rect 299638 269513 299690 269519
rect 298752 263796 299006 263824
rect 299232 263796 299486 263824
rect 299650 263810 299678 269513
rect 300130 269059 300158 271807
rect 300118 269053 300170 269059
rect 300118 268995 300170 269001
rect 300226 263810 300254 275507
rect 301090 270687 301118 278018
rect 302242 272537 302270 278018
rect 303286 275417 303338 275423
rect 303286 275359 303338 275365
rect 302230 272531 302282 272537
rect 302230 272473 302282 272479
rect 301366 272457 301418 272463
rect 301366 272399 301418 272405
rect 301078 270681 301130 270687
rect 301078 270623 301130 270629
rect 300694 268979 300746 268985
rect 300694 268921 300746 268927
rect 300706 263810 300734 268921
rect 301378 263824 301406 272399
rect 302422 270681 302474 270687
rect 302422 270623 302474 270629
rect 302434 269503 302462 270623
rect 302422 269497 302474 269503
rect 302422 269439 302474 269445
rect 302614 269497 302666 269503
rect 302614 269439 302666 269445
rect 302038 269127 302090 269133
rect 302038 269069 302090 269075
rect 301846 266981 301898 266987
rect 301846 266923 301898 266929
rect 301858 263824 301886 266923
rect 301152 263796 301406 263824
rect 301632 263796 301886 263824
rect 302050 263810 302078 269069
rect 302626 263810 302654 269439
rect 303298 263824 303326 275359
rect 303490 272389 303518 278018
rect 304438 275343 304490 275349
rect 304438 275285 304490 275291
rect 303958 272457 304010 272463
rect 303958 272399 304010 272405
rect 303478 272383 303530 272389
rect 303478 272325 303530 272331
rect 303766 269201 303818 269207
rect 303766 269143 303818 269149
rect 303778 263824 303806 269143
rect 303072 263796 303326 263824
rect 303552 263796 303806 263824
rect 303970 263810 303998 272399
rect 304450 263810 304478 275285
rect 304642 270687 304670 278018
rect 305794 272315 305822 278018
rect 306946 272981 306974 278018
rect 307318 275269 307370 275275
rect 307318 275211 307370 275217
rect 306934 272975 306986 272981
rect 306934 272917 306986 272923
rect 307030 272975 307082 272981
rect 307030 272917 307082 272923
rect 305782 272309 305834 272315
rect 305782 272251 305834 272257
rect 304630 270681 304682 270687
rect 304630 270623 304682 270629
rect 306358 270681 306410 270687
rect 306358 270623 306410 270629
rect 305686 268165 305738 268171
rect 305686 268107 305738 268113
rect 305014 266907 305066 266913
rect 305014 266849 305066 266855
rect 305026 263810 305054 266849
rect 305698 263824 305726 268107
rect 306166 266833 306218 266839
rect 306166 266775 306218 266781
rect 306178 263824 306206 266775
rect 305472 263796 305726 263824
rect 305952 263796 306206 263824
rect 306370 263810 306398 270623
rect 307042 268763 307070 272917
rect 307126 272383 307178 272389
rect 307126 272325 307178 272331
rect 307030 268757 307082 268763
rect 307030 268699 307082 268705
rect 307138 263824 307166 272325
rect 306864 263796 307166 263824
rect 307330 263810 307358 275211
rect 308194 269429 308222 278018
rect 309346 273573 309374 278018
rect 310390 275195 310442 275201
rect 310390 275137 310442 275143
rect 309334 273567 309386 273573
rect 309334 273509 309386 273515
rect 309910 272309 309962 272315
rect 309910 272251 309962 272257
rect 308182 269423 308234 269429
rect 308182 269365 308234 269371
rect 308278 269423 308330 269429
rect 308278 269365 308330 269371
rect 308086 266685 308138 266691
rect 308086 266627 308138 266633
rect 308098 263824 308126 266627
rect 307872 263796 308126 263824
rect 308290 263810 308318 269365
rect 309238 268239 309290 268245
rect 309238 268181 309290 268187
rect 308758 266759 308810 266765
rect 308758 266701 308810 266707
rect 308770 263810 308798 266701
rect 309250 263810 309278 268181
rect 309922 263824 309950 272251
rect 310402 263824 310430 275137
rect 310498 273425 310526 278018
rect 311638 275047 311690 275053
rect 311638 274989 311690 274995
rect 310486 273419 310538 273425
rect 310486 273361 310538 273367
rect 310582 273419 310634 273425
rect 310582 273361 310634 273367
rect 310594 268837 310622 273361
rect 311158 269349 311210 269355
rect 311158 269291 311210 269297
rect 310582 268831 310634 268837
rect 310582 268773 310634 268779
rect 310678 266611 310730 266617
rect 310678 266553 310730 266559
rect 309696 263796 309950 263824
rect 310272 263796 310430 263824
rect 310690 263810 310718 266553
rect 311170 263810 311198 269291
rect 311650 263810 311678 274989
rect 311746 269281 311774 278018
rect 312898 272241 312926 278018
rect 312886 272235 312938 272241
rect 312886 272177 312938 272183
rect 312982 272235 313034 272241
rect 312982 272177 313034 272183
rect 311734 269275 311786 269281
rect 311734 269217 311786 269223
rect 312310 268313 312362 268319
rect 312310 268255 312362 268261
rect 312322 263824 312350 268255
rect 312994 263824 313022 272177
rect 314050 272167 314078 278018
rect 314710 275121 314762 275127
rect 314710 275063 314762 275069
rect 314038 272161 314090 272167
rect 314038 272103 314090 272109
rect 314230 269275 314282 269281
rect 314230 269217 314282 269223
rect 313558 266537 313610 266543
rect 313558 266479 313610 266485
rect 313078 266463 313130 266469
rect 313078 266405 313130 266411
rect 312096 263796 312350 263824
rect 312672 263796 313022 263824
rect 313090 263810 313118 266405
rect 313570 263810 313598 266479
rect 314242 263824 314270 269217
rect 314722 263824 314750 275063
rect 314016 263796 314270 263824
rect 314496 263796 314750 263824
rect 314914 263810 314942 278245
rect 319510 278229 319562 278235
rect 418966 278229 419018 278235
rect 319510 278171 319562 278177
rect 316630 278155 316682 278161
rect 316630 278097 316682 278103
rect 315298 268689 315326 278018
rect 315958 274233 316010 274239
rect 315958 274175 316010 274181
rect 315478 272161 315530 272167
rect 315478 272103 315530 272109
rect 315286 268683 315338 268689
rect 315286 268625 315338 268631
rect 315490 263810 315518 272103
rect 315970 263810 315998 274175
rect 316450 273499 316478 278018
rect 316438 273493 316490 273499
rect 316438 273435 316490 273441
rect 316642 263824 316670 278097
rect 317878 278081 317930 278087
rect 317878 278023 317930 278029
rect 317302 274159 317354 274165
rect 317302 274101 317354 274107
rect 317110 268387 317162 268393
rect 317110 268329 317162 268335
rect 317122 263824 317150 268329
rect 316416 263796 316670 263824
rect 316896 263796 317150 263824
rect 317314 263810 317342 274101
rect 317602 273351 317630 278018
rect 317590 273345 317642 273351
rect 317590 273287 317642 273293
rect 317890 263810 317918 278023
rect 318358 271273 318410 271279
rect 318358 271215 318410 271221
rect 318370 263810 318398 271215
rect 318850 270613 318878 278018
rect 318838 270607 318890 270613
rect 318838 270549 318890 270555
rect 319030 265501 319082 265507
rect 319030 265443 319082 265449
rect 319042 263824 319070 265443
rect 319522 263824 319550 278171
rect 411874 278161 412176 278180
rect 419018 278177 419280 278180
rect 418966 278171 419280 278177
rect 411862 278155 412176 278161
rect 411914 278152 412176 278155
rect 418978 278152 419280 278171
rect 411862 278097 411914 278103
rect 415414 278081 415466 278087
rect 320002 270391 320030 278018
rect 320950 276749 321002 276755
rect 320950 276691 321002 276697
rect 320182 274307 320234 274313
rect 320182 274249 320234 274255
rect 319990 270385 320042 270391
rect 319990 270327 320042 270333
rect 319702 268461 319754 268467
rect 319702 268403 319754 268409
rect 318816 263796 319070 263824
rect 319296 263796 319550 263824
rect 319714 263810 319742 268403
rect 320194 263810 320222 274249
rect 320962 263824 320990 276691
rect 321154 273277 321182 278018
rect 322102 278007 322154 278013
rect 322102 277949 322154 277955
rect 321142 273271 321194 273277
rect 321142 273213 321194 273219
rect 321430 271347 321482 271353
rect 321430 271289 321482 271295
rect 321442 263824 321470 271289
rect 321622 265649 321674 265655
rect 321622 265591 321674 265597
rect 320736 263796 320990 263824
rect 321216 263796 321470 263824
rect 321634 263810 321662 265591
rect 322114 263810 322142 277949
rect 322402 270539 322430 278018
rect 323350 274381 323402 274387
rect 323350 274323 323402 274329
rect 322390 270533 322442 270539
rect 322390 270475 322442 270481
rect 322582 268535 322634 268541
rect 322582 268477 322634 268483
rect 322594 263810 322622 268477
rect 323362 263824 323390 274323
rect 323554 270465 323582 278018
rect 323830 277785 323882 277791
rect 323830 277727 323882 277733
rect 323542 270459 323594 270465
rect 323542 270401 323594 270407
rect 323842 263824 323870 277727
rect 324706 271945 324734 278018
rect 325858 274831 325886 278018
rect 326422 277859 326474 277865
rect 326422 277801 326474 277807
rect 325846 274825 325898 274831
rect 325846 274767 325898 274773
rect 325942 274455 325994 274461
rect 325942 274397 325994 274403
rect 324694 271939 324746 271945
rect 324694 271881 324746 271887
rect 324022 271421 324074 271427
rect 324022 271363 324074 271369
rect 323136 263796 323390 263824
rect 323616 263796 323870 263824
rect 324034 263810 324062 271363
rect 325750 268609 325802 268615
rect 325750 268551 325802 268557
rect 324502 265723 324554 265729
rect 324502 265665 324554 265671
rect 324514 263810 324542 265665
rect 324982 264095 325034 264101
rect 324982 264037 325034 264043
rect 324994 263810 325022 264037
rect 325762 263824 325790 268551
rect 325536 263796 325790 263824
rect 325954 263810 325982 274397
rect 326134 273863 326186 273869
rect 326134 273805 326186 273811
rect 326146 268985 326174 273805
rect 326134 268979 326186 268985
rect 326134 268921 326186 268927
rect 326434 263810 326462 277801
rect 327106 272093 327134 278018
rect 327094 272087 327146 272093
rect 327094 272029 327146 272035
rect 328258 272019 328286 278018
rect 329302 277711 329354 277717
rect 329302 277653 329354 277659
rect 328822 274529 328874 274535
rect 328822 274471 328874 274477
rect 328246 272013 328298 272019
rect 328246 271955 328298 271961
rect 326902 271495 326954 271501
rect 326902 271437 326954 271443
rect 326914 263810 326942 271437
rect 328342 268683 328394 268689
rect 328342 268625 328394 268631
rect 327574 265797 327626 265803
rect 327574 265739 327626 265745
rect 327586 263824 327614 265739
rect 328054 264761 328106 264767
rect 328054 264703 328106 264709
rect 328066 263824 328094 264703
rect 327360 263796 327614 263824
rect 327840 263796 328094 263824
rect 328354 263810 328382 268625
rect 328834 263810 328862 274471
rect 329314 263810 329342 277653
rect 329410 274905 329438 278018
rect 329398 274899 329450 274905
rect 329398 274841 329450 274847
rect 330454 274603 330506 274609
rect 330454 274545 330506 274551
rect 329974 271569 330026 271575
rect 329974 271511 330026 271517
rect 329986 263824 330014 271511
rect 330466 263824 330494 274545
rect 330658 270317 330686 278018
rect 331222 273715 331274 273721
rect 331222 273657 331274 273663
rect 330646 270311 330698 270317
rect 330646 270253 330698 270259
rect 331234 269133 331262 273657
rect 331810 270243 331838 278018
rect 332374 277637 332426 277643
rect 332374 277579 332426 277585
rect 331798 270237 331850 270243
rect 331798 270179 331850 270185
rect 331222 269127 331274 269133
rect 331222 269069 331274 269075
rect 331222 268757 331274 268763
rect 331222 268699 331274 268705
rect 331126 264687 331178 264693
rect 331126 264629 331178 264635
rect 331138 263824 331166 264629
rect 329760 263796 330014 263824
rect 330240 263796 330494 263824
rect 330768 263796 331166 263824
rect 331234 263810 331262 268699
rect 331894 265871 331946 265877
rect 331894 265813 331946 265819
rect 331906 263824 331934 265813
rect 332386 263824 332414 277579
rect 332962 274979 332990 278018
rect 332950 274973 333002 274979
rect 332950 274915 333002 274921
rect 333142 274677 333194 274683
rect 333142 274619 333194 274625
rect 332566 271643 332618 271649
rect 332566 271585 332618 271591
rect 331680 263796 331934 263824
rect 332160 263796 332414 263824
rect 332578 263810 332606 271585
rect 333154 263810 333182 274619
rect 334210 273129 334238 278018
rect 334966 277563 335018 277569
rect 334966 277505 335018 277511
rect 334294 274011 334346 274017
rect 334294 273953 334346 273959
rect 334198 273123 334250 273129
rect 334198 273065 334250 273071
rect 334102 270755 334154 270761
rect 334102 270697 334154 270703
rect 334114 270169 334142 270697
rect 334102 270163 334154 270169
rect 334102 270105 334154 270111
rect 334306 269207 334334 273953
rect 334294 269201 334346 269207
rect 334294 269143 334346 269149
rect 334294 268831 334346 268837
rect 334294 268773 334346 268779
rect 333622 267943 333674 267949
rect 333622 267885 333674 267891
rect 333634 263810 333662 267885
rect 334306 263824 334334 268773
rect 334774 265945 334826 265951
rect 334774 265887 334826 265893
rect 334786 263824 334814 265887
rect 334080 263796 334334 263824
rect 334560 263796 334814 263824
rect 334978 263810 335006 277505
rect 335362 273203 335390 278018
rect 336514 276459 336542 278018
rect 336502 276453 336554 276459
rect 336502 276395 336554 276401
rect 336022 274751 336074 274757
rect 336022 274693 336074 274699
rect 335350 273197 335402 273203
rect 335350 273139 335402 273145
rect 335446 271717 335498 271723
rect 335446 271659 335498 271665
rect 335458 263810 335486 271659
rect 336034 263810 336062 274693
rect 337762 270761 337790 278018
rect 337846 277489 337898 277495
rect 337846 277431 337898 277437
rect 337750 270755 337802 270761
rect 337750 270697 337802 270703
rect 336886 268905 336938 268911
rect 336886 268847 336938 268853
rect 336694 268017 336746 268023
rect 336694 267959 336746 267965
rect 336706 263824 336734 267959
rect 336480 263796 336734 263824
rect 336898 263824 336926 268847
rect 337366 266019 337418 266025
rect 337366 265961 337418 265967
rect 336898 263796 336960 263824
rect 337378 263810 337406 265961
rect 337858 263810 337886 277431
rect 338914 273055 338942 278018
rect 340066 276385 340094 278018
rect 341014 277415 341066 277421
rect 341014 277357 341066 277363
rect 340054 276379 340106 276385
rect 340054 276321 340106 276327
rect 339094 274825 339146 274831
rect 339094 274767 339146 274773
rect 338902 273049 338954 273055
rect 338902 272991 338954 272997
rect 338614 271199 338666 271205
rect 338614 271141 338666 271147
rect 338134 270755 338186 270761
rect 338134 270697 338186 270703
rect 338146 270021 338174 270697
rect 338134 270015 338186 270021
rect 338134 269957 338186 269963
rect 338626 263824 338654 271141
rect 339106 263824 339134 274767
rect 339766 268979 339818 268985
rect 339766 268921 339818 268927
rect 339286 267869 339338 267875
rect 339286 267811 339338 267817
rect 338400 263796 338654 263824
rect 338880 263796 339134 263824
rect 339298 263810 339326 267811
rect 339778 263810 339806 268921
rect 340246 266093 340298 266099
rect 340246 266035 340298 266041
rect 340258 263810 340286 266035
rect 341026 263824 341054 277357
rect 341314 270761 341342 278018
rect 341684 274346 341740 274355
rect 341684 274281 341740 274290
rect 341494 271791 341546 271797
rect 341494 271733 341546 271739
rect 341302 270755 341354 270761
rect 341302 270697 341354 270703
rect 341506 263824 341534 271733
rect 340800 263796 341054 263824
rect 341280 263796 341534 263824
rect 341698 263810 341726 274281
rect 341974 273789 342026 273795
rect 341974 273731 342026 273737
rect 341986 270687 342014 273731
rect 341974 270681 342026 270687
rect 341974 270623 342026 270629
rect 342466 270095 342494 278018
rect 343618 276311 343646 278018
rect 343894 277341 343946 277347
rect 343894 277283 343946 277289
rect 343606 276305 343658 276311
rect 343606 276247 343658 276253
rect 342742 271939 342794 271945
rect 342742 271881 342794 271887
rect 342454 270089 342506 270095
rect 342454 270031 342506 270037
rect 342754 269947 342782 271881
rect 342742 269941 342794 269947
rect 342742 269883 342794 269889
rect 342646 269127 342698 269133
rect 342646 269069 342698 269075
rect 342166 268091 342218 268097
rect 342166 268033 342218 268039
rect 342178 263810 342206 268033
rect 342658 263810 342686 269069
rect 343318 266167 343370 266173
rect 343318 266109 343370 266115
rect 343330 263824 343358 266109
rect 343906 263824 343934 277283
rect 344566 274899 344618 274905
rect 344566 274841 344618 274847
rect 344086 271865 344138 271871
rect 344086 271807 344138 271813
rect 343104 263796 343358 263824
rect 343632 263796 343934 263824
rect 344098 263810 344126 271807
rect 344578 263810 344606 274841
rect 344770 273425 344798 278018
rect 344758 273419 344810 273425
rect 344758 273361 344810 273367
rect 346018 272907 346046 278018
rect 347170 276237 347198 278018
rect 347158 276231 347210 276237
rect 347158 276173 347210 276179
rect 347636 274494 347692 274503
rect 347636 274429 347692 274438
rect 347062 273937 347114 273943
rect 347062 273879 347114 273885
rect 346006 272901 346058 272907
rect 346006 272843 346058 272849
rect 346966 272087 347018 272093
rect 346966 272029 347018 272035
rect 346486 272013 346538 272019
rect 346486 271955 346538 271961
rect 345430 270681 345482 270687
rect 345430 270623 345482 270629
rect 345238 269201 345290 269207
rect 345238 269143 345290 269149
rect 345250 263824 345278 269143
rect 345024 263796 345278 263824
rect 345442 263676 345470 270623
rect 346006 266241 346058 266247
rect 346006 266183 346058 266189
rect 346018 263810 346046 266183
rect 346498 263810 346526 271955
rect 346978 263810 347006 272029
rect 347074 268245 347102 273879
rect 347062 268239 347114 268245
rect 347062 268181 347114 268187
rect 347650 263824 347678 274429
rect 348322 271945 348350 278018
rect 348502 274085 348554 274091
rect 348502 274027 348554 274033
rect 348310 271939 348362 271945
rect 348310 271881 348362 271887
rect 348118 270607 348170 270613
rect 348118 270549 348170 270555
rect 348130 263824 348158 270549
rect 348406 270533 348458 270539
rect 348406 270475 348458 270481
rect 347424 263796 347678 263824
rect 347904 263796 348158 263824
rect 348418 263810 348446 270475
rect 348514 268319 348542 274027
rect 349462 273493 349514 273499
rect 349462 273435 349514 273441
rect 348598 271791 348650 271797
rect 348598 271733 348650 271739
rect 348610 271205 348638 271733
rect 348598 271199 348650 271205
rect 348598 271141 348650 271147
rect 348502 268313 348554 268319
rect 348502 268255 348554 268261
rect 348886 266315 348938 266321
rect 348886 266257 348938 266263
rect 348898 263810 348926 266257
rect 349474 263824 349502 273435
rect 349570 269873 349598 278018
rect 350722 276163 350750 278018
rect 350710 276157 350762 276163
rect 350710 276099 350762 276105
rect 350228 274642 350284 274651
rect 350228 274577 350284 274586
rect 350038 273567 350090 273573
rect 350038 273509 350090 273515
rect 349558 269867 349610 269873
rect 349558 269809 349610 269815
rect 350050 263824 350078 273509
rect 349344 263796 349502 263824
rect 349824 263796 350078 263824
rect 350242 263810 350270 274577
rect 351874 272833 351902 278018
rect 352438 273419 352490 273425
rect 352438 273361 352490 273367
rect 351862 272827 351914 272833
rect 351862 272769 351914 272775
rect 351382 270903 351434 270909
rect 351382 270845 351434 270851
rect 350710 270459 350762 270465
rect 350710 270401 350762 270407
rect 350722 263810 350750 270401
rect 351286 270385 351338 270391
rect 351286 270327 351338 270333
rect 351298 263810 351326 270327
rect 351394 269725 351422 270845
rect 351382 269719 351434 269725
rect 351382 269661 351434 269667
rect 351382 267943 351434 267949
rect 351382 267885 351434 267891
rect 351394 264471 351422 267885
rect 351958 267795 352010 267801
rect 351958 267737 352010 267743
rect 351382 264465 351434 264471
rect 351382 264407 351434 264413
rect 351970 263824 351998 267737
rect 352450 263824 352478 273361
rect 352630 273345 352682 273351
rect 352630 273287 352682 273293
rect 351744 263796 351998 263824
rect 352224 263796 352478 263824
rect 352642 263810 352670 273287
rect 353122 272759 353150 278018
rect 354274 276089 354302 278018
rect 354262 276083 354314 276089
rect 354262 276025 354314 276031
rect 353396 274790 353452 274799
rect 353396 274725 353452 274734
rect 353110 272753 353162 272759
rect 353110 272695 353162 272701
rect 353410 263824 353438 274725
rect 355030 273197 355082 273203
rect 355030 273139 355082 273145
rect 354070 270311 354122 270317
rect 354070 270253 354122 270259
rect 353686 270237 353738 270243
rect 353686 270179 353738 270185
rect 353136 263796 353438 263824
rect 353698 263810 353726 270179
rect 354082 264120 354110 270253
rect 354262 268017 354314 268023
rect 354262 267959 354314 267965
rect 354274 264619 354302 267959
rect 354838 267721 354890 267727
rect 354838 267663 354890 267669
rect 354262 264613 354314 264619
rect 354262 264555 354314 264561
rect 354082 264092 354158 264120
rect 354130 263810 354158 264092
rect 354850 263824 354878 267663
rect 354624 263796 354878 263824
rect 355042 263810 355070 273139
rect 355426 270909 355454 278018
rect 356182 274973 356234 274979
rect 356182 274915 356234 274921
rect 355510 273271 355562 273277
rect 355510 273213 355562 273219
rect 355414 270903 355466 270909
rect 355414 270845 355466 270851
rect 355522 263810 355550 273213
rect 356194 263824 356222 274915
rect 356674 269799 356702 278018
rect 357826 276015 357854 278018
rect 357814 276009 357866 276015
rect 357814 275951 357866 275957
rect 358582 273123 358634 273129
rect 358582 273065 358634 273071
rect 357910 271199 357962 271205
rect 357910 271141 357962 271147
rect 356758 270163 356810 270169
rect 356758 270105 356810 270111
rect 356662 269793 356714 269799
rect 356662 269735 356714 269741
rect 356770 263824 356798 270105
rect 356950 270089 357002 270095
rect 356950 270031 357002 270037
rect 355968 263796 356222 263824
rect 356544 263796 356798 263824
rect 356962 263810 356990 270031
rect 357430 267647 357482 267653
rect 357430 267589 357482 267595
rect 357442 263810 357470 267589
rect 357922 263810 357950 271141
rect 358594 263824 358622 273065
rect 358978 272981 359006 278018
rect 359158 276453 359210 276459
rect 359158 276395 359210 276401
rect 358966 272975 359018 272981
rect 358966 272917 359018 272923
rect 359170 263824 359198 276395
rect 360226 272685 360254 278018
rect 361378 275941 361406 278018
rect 361750 276379 361802 276385
rect 361750 276321 361802 276327
rect 361366 275935 361418 275941
rect 361366 275877 361418 275883
rect 360982 273049 361034 273055
rect 360982 272991 361034 272997
rect 360214 272679 360266 272685
rect 360214 272621 360266 272627
rect 359350 270015 359402 270021
rect 359350 269957 359402 269963
rect 358368 263796 358622 263824
rect 358944 263796 359198 263824
rect 359362 263810 359390 269957
rect 359830 269941 359882 269947
rect 359830 269883 359882 269889
rect 359446 268091 359498 268097
rect 359446 268033 359498 268039
rect 359458 264841 359486 268033
rect 359446 264835 359498 264841
rect 359446 264777 359498 264783
rect 359842 263810 359870 269883
rect 360406 267869 360458 267875
rect 360406 267811 360458 267817
rect 360310 267573 360362 267579
rect 360310 267515 360362 267521
rect 360322 263810 360350 267515
rect 360418 264545 360446 267811
rect 360406 264539 360458 264545
rect 360406 264481 360458 264487
rect 360994 263824 361022 272991
rect 361270 272975 361322 272981
rect 361270 272917 361322 272923
rect 360768 263796 361022 263824
rect 361282 263810 361310 272917
rect 361762 263810 361790 276321
rect 362530 275867 362558 278018
rect 362518 275861 362570 275867
rect 362518 275803 362570 275809
rect 363574 272901 363626 272907
rect 363574 272843 363626 272849
rect 362230 269867 362282 269873
rect 362230 269809 362282 269815
rect 362242 263810 362270 269809
rect 362806 269793 362858 269799
rect 362806 269735 362858 269741
rect 362818 263824 362846 269735
rect 363382 267499 363434 267505
rect 363382 267441 363434 267447
rect 363394 263824 363422 267441
rect 362688 263796 362846 263824
rect 363168 263796 363422 263824
rect 363586 263810 363614 272843
rect 363682 269651 363710 278018
rect 364630 276305 364682 276311
rect 364630 276247 364682 276253
rect 364150 272827 364202 272833
rect 364150 272769 364202 272775
rect 363670 269645 363722 269651
rect 363670 269587 363722 269593
rect 364162 263810 364190 272769
rect 364642 263810 364670 276247
rect 364930 275793 364958 278018
rect 364918 275787 364970 275793
rect 364918 275729 364970 275735
rect 366082 275719 366110 278018
rect 366070 275713 366122 275719
rect 366070 275655 366122 275661
rect 366550 272753 366602 272759
rect 366550 272695 366602 272701
rect 365302 269719 365354 269725
rect 365302 269661 365354 269667
rect 365314 263824 365342 269661
rect 365686 268091 365738 268097
rect 365686 268033 365738 268039
rect 365698 263824 365726 268033
rect 365974 267425 366026 267431
rect 365974 267367 366026 267373
rect 365088 263796 365342 263824
rect 365568 263796 365726 263824
rect 365986 263810 366014 267367
rect 366562 263810 366590 272695
rect 367126 272679 367178 272685
rect 367126 272621 367178 272627
rect 367138 263824 367166 272621
rect 367234 272611 367262 278018
rect 367702 276231 367754 276237
rect 367702 276173 367754 276179
rect 367222 272605 367274 272611
rect 367222 272547 367274 272553
rect 367714 263824 367742 276173
rect 368482 275645 368510 278018
rect 368470 275639 368522 275645
rect 368470 275581 368522 275587
rect 369634 275497 369662 278018
rect 370294 276157 370346 276163
rect 370294 276099 370346 276105
rect 369622 275491 369674 275497
rect 369622 275433 369674 275439
rect 370100 271978 370156 271987
rect 370100 271913 370156 271922
rect 369620 271830 369676 271839
rect 369620 271765 369676 271774
rect 367892 269166 367948 269175
rect 367892 269101 367948 269110
rect 367008 263796 367166 263824
rect 367488 263796 367742 263824
rect 367906 263810 367934 269101
rect 368372 269018 368428 269027
rect 368372 268953 368428 268962
rect 368386 263810 368414 268953
rect 368950 267351 369002 267357
rect 368950 267293 369002 267299
rect 368962 263810 368990 267293
rect 369634 263824 369662 271765
rect 370114 263824 370142 271913
rect 369408 263796 369662 263824
rect 369888 263796 370142 263824
rect 370306 263810 370334 276099
rect 370786 269577 370814 278018
rect 371926 276083 371978 276089
rect 371926 276025 371978 276031
rect 371062 276009 371114 276015
rect 371062 275951 371114 275957
rect 370774 269571 370826 269577
rect 370774 269513 370826 269519
rect 371074 263824 371102 275951
rect 371254 269571 371306 269577
rect 371254 269513 371306 269519
rect 370800 263796 371102 263824
rect 371266 263810 371294 269513
rect 371938 263824 371966 276025
rect 372034 275571 372062 278018
rect 372022 275565 372074 275571
rect 372022 275507 372074 275513
rect 373186 273869 373214 278018
rect 373846 277267 373898 277273
rect 373846 277209 373898 277215
rect 373462 275935 373514 275941
rect 373462 275877 373514 275883
rect 373174 273863 373226 273869
rect 373174 273805 373226 273811
rect 372694 272605 372746 272611
rect 372694 272547 372746 272553
rect 372502 267277 372554 267283
rect 372502 267219 372554 267225
rect 372514 263824 372542 267219
rect 371808 263796 371966 263824
rect 372288 263796 372542 263824
rect 372706 263810 372734 272547
rect 373474 263824 373502 275877
rect 373858 263824 373886 277209
rect 374338 272537 374366 278018
rect 375298 278004 375600 278032
rect 375094 277193 375146 277199
rect 375094 277135 375146 277141
rect 374614 275861 374666 275867
rect 374614 275803 374666 275809
rect 374326 272531 374378 272537
rect 374326 272473 374378 272479
rect 374324 270498 374380 270507
rect 374324 270433 374380 270442
rect 374338 263824 374366 270433
rect 373200 263796 373502 263824
rect 373632 263796 373886 263824
rect 374208 263796 374366 263824
rect 374626 263810 374654 275803
rect 375106 263810 375134 277135
rect 375190 273123 375242 273129
rect 375190 273065 375242 273071
rect 375202 271205 375230 273065
rect 375190 271199 375242 271205
rect 375190 271141 375242 271147
rect 375298 266987 375326 278004
rect 376246 275713 376298 275719
rect 376246 275655 376298 275661
rect 375572 273458 375628 273467
rect 375572 273393 375628 273402
rect 375286 266981 375338 266987
rect 375286 266923 375338 266929
rect 375586 263810 375614 273393
rect 376258 263824 376286 275655
rect 376738 273721 376766 278018
rect 376822 277119 376874 277125
rect 376822 277061 376874 277067
rect 376726 273715 376778 273721
rect 376726 273657 376778 273663
rect 376834 263824 376862 277061
rect 377494 275787 377546 275793
rect 377494 275729 377546 275735
rect 377012 270350 377068 270359
rect 377012 270285 377068 270294
rect 376032 263796 376286 263824
rect 376608 263796 376862 263824
rect 377026 263810 377054 270285
rect 377506 263810 377534 275729
rect 377890 269503 377918 278018
rect 377974 277045 378026 277051
rect 377974 276987 378026 276993
rect 377878 269497 377930 269503
rect 377878 269439 377930 269445
rect 377986 263810 378014 276987
rect 379138 275423 379166 278018
rect 379414 276971 379466 276977
rect 379414 276913 379466 276919
rect 379126 275417 379178 275423
rect 379126 275359 379178 275365
rect 379124 274938 379180 274947
rect 379124 274873 379180 274882
rect 378644 273310 378700 273319
rect 378644 273245 378700 273254
rect 378658 263824 378686 273245
rect 379138 263824 379166 274873
rect 378432 263796 378686 263824
rect 378912 263796 379166 263824
rect 379426 263810 379454 276913
rect 380290 274017 380318 278018
rect 381046 276897 381098 276903
rect 381046 276839 381098 276845
rect 380566 275639 380618 275645
rect 380566 275581 380618 275587
rect 380278 274011 380330 274017
rect 380278 273953 380330 273959
rect 379894 269497 379946 269503
rect 379894 269439 379946 269445
rect 379906 263810 379934 269439
rect 380578 263824 380606 275581
rect 381058 263824 381086 276839
rect 381442 272463 381470 278018
rect 382294 277933 382346 277939
rect 382294 277875 382346 277881
rect 381814 275565 381866 275571
rect 381814 275507 381866 275513
rect 381430 272457 381482 272463
rect 381430 272399 381482 272405
rect 381526 272457 381578 272463
rect 381526 272399 381578 272405
rect 381538 263824 381566 272399
rect 380352 263796 380606 263824
rect 380832 263796 381086 263824
rect 381264 263796 381566 263824
rect 381826 263810 381854 275507
rect 382306 263810 382334 277875
rect 382594 275349 382622 278018
rect 383638 276823 383690 276829
rect 383638 276765 383690 276771
rect 383444 275974 383500 275983
rect 383444 275909 383500 275918
rect 382582 275343 382634 275349
rect 382582 275285 382634 275291
rect 382964 273162 383020 273171
rect 382964 273097 383020 273106
rect 382978 263824 383006 273097
rect 383458 263824 383486 275909
rect 382752 263796 383006 263824
rect 383232 263796 383486 263824
rect 383650 263810 383678 276765
rect 383842 266913 383870 278018
rect 384118 269053 384170 269059
rect 384118 268995 384170 269001
rect 383830 266907 383882 266913
rect 383830 266849 383882 266855
rect 384130 263810 384158 268995
rect 384994 268171 385022 278018
rect 385366 276601 385418 276607
rect 385366 276543 385418 276549
rect 384982 268165 385034 268171
rect 384982 268107 385034 268113
rect 384886 267203 384938 267209
rect 384886 267145 384938 267151
rect 384898 263824 384926 267145
rect 385378 263824 385406 276543
rect 385556 270202 385612 270211
rect 385556 270137 385612 270146
rect 384672 263796 384926 263824
rect 385152 263796 385406 263824
rect 385570 263810 385598 270137
rect 386038 267129 386090 267135
rect 386038 267071 386090 267077
rect 386050 263810 386078 267071
rect 386146 266839 386174 278018
rect 386518 276675 386570 276681
rect 386518 276617 386570 276623
rect 386134 266833 386186 266839
rect 386134 266775 386186 266781
rect 386530 263810 386558 276617
rect 387394 273795 387422 278018
rect 387382 273789 387434 273795
rect 387382 273731 387434 273737
rect 388546 272389 388574 278018
rect 388918 275491 388970 275497
rect 388918 275433 388970 275439
rect 388534 272383 388586 272389
rect 388534 272325 388586 272331
rect 387286 271199 387338 271205
rect 387286 271141 387338 271147
rect 387298 263824 387326 271141
rect 388436 270054 388492 270063
rect 388436 269989 388492 269998
rect 387766 267055 387818 267061
rect 387766 266997 387818 267003
rect 387778 263824 387806 266997
rect 387958 264021 388010 264027
rect 387958 263963 388010 263969
rect 387072 263796 387326 263824
rect 387552 263796 387806 263824
rect 387970 263810 387998 263963
rect 388450 263810 388478 269989
rect 388930 263810 388958 275433
rect 389590 275417 389642 275423
rect 389590 275359 389642 275365
rect 389602 263824 389630 275359
rect 389698 275275 389726 278018
rect 390356 275826 390412 275835
rect 390356 275761 390412 275770
rect 389686 275269 389738 275275
rect 389686 275211 389738 275217
rect 390164 273014 390220 273023
rect 390164 272949 390220 272958
rect 390178 263824 390206 272949
rect 389472 263796 389630 263824
rect 389952 263796 390206 263824
rect 390370 263810 390398 275761
rect 390946 266691 390974 278018
rect 391990 275343 392042 275349
rect 391990 275285 392042 275291
rect 391508 269906 391564 269915
rect 391508 269841 391564 269850
rect 390934 266685 390986 266691
rect 390934 266627 390986 266633
rect 390838 263947 390890 263953
rect 390838 263889 390890 263895
rect 390850 263810 390878 263889
rect 391522 263824 391550 269841
rect 392002 263824 392030 275285
rect 392098 269429 392126 278018
rect 392962 278004 393264 278032
rect 415466 278029 415728 278032
rect 415414 278023 415728 278029
rect 392278 276527 392330 276533
rect 392278 276469 392330 276475
rect 392086 269423 392138 269429
rect 392086 269365 392138 269371
rect 391296 263796 391550 263824
rect 391776 263796 392030 263824
rect 392290 263810 392318 276469
rect 392756 272866 392812 272875
rect 392756 272801 392812 272810
rect 392770 263810 392798 272801
rect 392962 266765 392990 278004
rect 394498 273943 394526 278018
rect 395156 276566 395212 276575
rect 395156 276501 395212 276510
rect 394486 273937 394538 273943
rect 394486 273879 394538 273885
rect 394390 269423 394442 269429
rect 394390 269365 394442 269371
rect 393238 266907 393290 266913
rect 393238 266849 393290 266855
rect 392950 266759 393002 266765
rect 392950 266701 393002 266707
rect 393250 263810 393278 266849
rect 393910 263873 393962 263879
rect 393696 263821 393910 263824
rect 394402 263824 394430 269365
rect 394678 266981 394730 266987
rect 394678 266923 394730 266929
rect 393696 263815 393962 263821
rect 393696 263796 393950 263815
rect 394176 263796 394430 263824
rect 394690 263810 394718 266923
rect 395170 263810 395198 276501
rect 395650 272315 395678 278018
rect 396310 275269 396362 275275
rect 396310 275211 396362 275217
rect 395638 272309 395690 272315
rect 395638 272251 395690 272257
rect 395926 272309 395978 272315
rect 395926 272251 395978 272257
rect 395938 263824 395966 272251
rect 396322 263824 396350 275211
rect 396802 275201 396830 278018
rect 396790 275195 396842 275201
rect 396790 275137 396842 275143
rect 397076 268870 397132 268879
rect 397076 268805 397132 268814
rect 395664 263796 395966 263824
rect 396096 263796 396350 263824
rect 396576 263805 396830 263824
rect 397090 263810 397118 268805
rect 397558 266833 397610 266839
rect 397558 266775 397610 266781
rect 397570 263810 397598 266775
rect 398050 266617 398078 278018
rect 398900 275678 398956 275687
rect 398900 275613 398956 275622
rect 398708 272718 398764 272727
rect 398708 272653 398764 272662
rect 398230 266759 398282 266765
rect 398230 266701 398282 266707
rect 398038 266611 398090 266617
rect 398038 266553 398090 266559
rect 398242 263824 398270 266701
rect 398722 263824 398750 272653
rect 396576 263799 396842 263805
rect 396576 263796 396790 263799
rect 398016 263796 398270 263824
rect 398496 263796 398750 263824
rect 398914 263810 398942 275613
rect 399202 269355 399230 278018
rect 400354 275053 400382 278018
rect 400342 275047 400394 275053
rect 400342 274989 400394 274995
rect 401506 274091 401534 278018
rect 402548 276714 402604 276723
rect 402548 276649 402604 276658
rect 401494 274085 401546 274091
rect 401494 274027 401546 274033
rect 401782 274085 401834 274091
rect 401782 274027 401834 274033
rect 399190 269349 399242 269355
rect 399190 269291 399242 269297
rect 399958 269349 400010 269355
rect 399958 269291 400010 269297
rect 399382 264169 399434 264175
rect 399382 264111 399434 264117
rect 399394 263810 399422 264111
rect 399970 263810 399998 269291
rect 401302 267869 401354 267875
rect 401302 267811 401354 267817
rect 400630 266685 400682 266691
rect 400630 266627 400682 266633
rect 400642 263824 400670 266627
rect 400416 263796 400670 263824
rect 401314 263810 401342 267811
rect 401794 263810 401822 274027
rect 402562 263824 402590 276649
rect 402754 272241 402782 278018
rect 402742 272235 402794 272241
rect 402742 272177 402794 272183
rect 402838 272235 402890 272241
rect 402838 272177 402890 272183
rect 402850 267875 402878 272177
rect 403028 269758 403084 269767
rect 403028 269693 403084 269702
rect 402838 267869 402890 267875
rect 402838 267811 402890 267817
rect 403042 263824 403070 269693
rect 403222 266611 403274 266617
rect 403222 266553 403274 266559
rect 402336 263796 402590 263824
rect 402816 263796 403070 263824
rect 403234 263810 403262 266553
rect 403906 266469 403934 278018
rect 404950 275195 405002 275201
rect 404950 275137 405002 275143
rect 404180 272570 404236 272579
rect 404180 272505 404236 272514
rect 403894 266463 403946 266469
rect 403894 266405 403946 266411
rect 404194 263810 404222 272505
rect 404962 263824 404990 275137
rect 405058 266543 405086 278018
rect 405428 276862 405484 276871
rect 405428 276797 405484 276806
rect 405046 266537 405098 266543
rect 405046 266479 405098 266485
rect 405442 263824 405470 276797
rect 405620 269610 405676 269619
rect 405620 269545 405676 269554
rect 404736 263796 404990 263824
rect 405216 263796 405470 263824
rect 405634 263810 405662 269545
rect 406306 269281 406334 278018
rect 407458 275127 407486 278018
rect 407828 275530 407884 275539
rect 407828 275465 407884 275474
rect 407734 275195 407786 275201
rect 407734 275137 407786 275143
rect 407446 275121 407498 275127
rect 407446 275063 407498 275069
rect 407746 274091 407774 275137
rect 407734 274085 407786 274091
rect 407734 274027 407786 274033
rect 407252 272422 407308 272431
rect 407252 272357 407308 272366
rect 407446 272383 407498 272389
rect 406294 269275 406346 269281
rect 406294 269217 406346 269223
rect 406582 269275 406634 269281
rect 406582 269217 406634 269223
rect 406102 266537 406154 266543
rect 406102 266479 406154 266485
rect 406114 263810 406142 266479
rect 406594 263810 406622 269217
rect 407266 263824 407294 272357
rect 407446 272325 407498 272331
rect 407458 271205 407486 272325
rect 407446 271199 407498 271205
rect 407446 271141 407498 271147
rect 407842 263824 407870 275465
rect 408598 275121 408650 275127
rect 408598 275063 408650 275069
rect 408610 269281 408638 275063
rect 409858 272167 409886 278018
rect 411010 274239 411038 278018
rect 410998 274233 411050 274239
rect 410998 274175 411050 274181
rect 410900 272274 410956 272283
rect 410900 272209 410956 272218
rect 409846 272161 409898 272167
rect 409846 272103 409898 272109
rect 408982 270755 409034 270761
rect 408982 270697 409034 270703
rect 408598 269275 408650 269281
rect 408598 269217 408650 269223
rect 408994 268393 409022 270697
rect 410420 269462 410476 269471
rect 410420 269397 410476 269406
rect 408982 268387 409034 268393
rect 408982 268329 409034 268335
rect 408502 268239 408554 268245
rect 408502 268181 408554 268187
rect 408022 265575 408074 265581
rect 408022 265517 408074 265523
rect 407040 263796 407294 263824
rect 407616 263796 407870 263824
rect 408034 263810 408062 265517
rect 408514 263810 408542 268181
rect 409942 267869 409994 267875
rect 409942 267811 409994 267817
rect 409174 266463 409226 266469
rect 409174 266405 409226 266411
rect 409186 263824 409214 266405
rect 408960 263796 409214 263824
rect 409954 263810 409982 267811
rect 410434 263810 410462 269397
rect 410914 263810 410942 272209
rect 411764 272126 411820 272135
rect 411764 272061 411820 272070
rect 411572 269314 411628 269323
rect 411572 269249 411628 269258
rect 410998 264169 411050 264175
rect 410998 264111 411050 264117
rect 396790 263741 396842 263747
rect 411010 263731 411038 264111
rect 411586 263824 411614 269249
rect 411360 263796 411614 263824
rect 411778 263824 411806 272061
rect 413410 270761 413438 278018
rect 414562 274165 414590 278018
rect 415426 278004 415728 278023
rect 414550 274159 414602 274165
rect 414550 274101 414602 274107
rect 413686 272161 413738 272167
rect 413686 272103 413738 272109
rect 413398 270755 413450 270761
rect 413398 270697 413450 270703
rect 413698 267875 413726 272103
rect 416962 271279 416990 278018
rect 416950 271273 417002 271279
rect 416950 271215 417002 271221
rect 413686 267869 413738 267875
rect 413686 267811 413738 267817
rect 418114 265507 418142 278018
rect 420514 268467 420542 278018
rect 421666 274313 421694 278018
rect 422818 276755 422846 278018
rect 422806 276749 422858 276755
rect 422806 276691 422858 276697
rect 421654 274307 421706 274313
rect 421654 274249 421706 274255
rect 423970 271353 423998 278018
rect 423958 271347 424010 271353
rect 423958 271289 424010 271295
rect 420502 268461 420554 268467
rect 420502 268403 420554 268409
rect 425218 265655 425246 278018
rect 426274 278013 426384 278032
rect 426262 278007 426384 278013
rect 426314 278004 426384 278007
rect 426262 277949 426314 277955
rect 427522 268541 427550 278018
rect 428770 274387 428798 278018
rect 429922 277791 429950 278018
rect 429910 277785 429962 277791
rect 429910 277727 429962 277733
rect 428758 274381 428810 274387
rect 428758 274323 428810 274329
rect 431074 271427 431102 278018
rect 431062 271421 431114 271427
rect 431062 271363 431114 271369
rect 427510 268535 427562 268541
rect 427510 268477 427562 268483
rect 432322 265729 432350 278018
rect 432310 265723 432362 265729
rect 432310 265665 432362 265671
rect 425206 265649 425258 265655
rect 425206 265591 425258 265597
rect 418102 265501 418154 265507
rect 418102 265443 418154 265449
rect 433474 264101 433502 278018
rect 434626 268615 434654 278018
rect 435874 274461 435902 278018
rect 437026 277865 437054 278018
rect 437014 277859 437066 277865
rect 437014 277801 437066 277807
rect 435862 274455 435914 274461
rect 435862 274397 435914 274403
rect 438178 271501 438206 278018
rect 438166 271495 438218 271501
rect 438166 271437 438218 271443
rect 434614 268609 434666 268615
rect 434614 268551 434666 268557
rect 439330 265803 439358 278018
rect 439318 265797 439370 265803
rect 439318 265739 439370 265745
rect 440578 264767 440606 278018
rect 441730 268689 441758 278018
rect 442882 274535 442910 278018
rect 444130 277717 444158 278018
rect 444118 277711 444170 277717
rect 444118 277653 444170 277659
rect 442870 274529 442922 274535
rect 442870 274471 442922 274477
rect 445282 271575 445310 278018
rect 446434 274609 446462 278018
rect 446422 274603 446474 274609
rect 446422 274545 446474 274551
rect 445270 271569 445322 271575
rect 445270 271511 445322 271517
rect 441718 268683 441770 268689
rect 441718 268625 441770 268631
rect 440566 264761 440618 264767
rect 440566 264703 440618 264709
rect 447682 264693 447710 278018
rect 448834 268763 448862 278018
rect 448822 268757 448874 268763
rect 448822 268699 448874 268705
rect 449986 265877 450014 278018
rect 451234 277643 451262 278018
rect 451222 277637 451274 277643
rect 451222 277579 451274 277585
rect 452386 271649 452414 278018
rect 453538 274683 453566 278018
rect 453526 274677 453578 274683
rect 453526 274619 453578 274625
rect 452374 271643 452426 271649
rect 452374 271585 452426 271591
rect 449974 265871 450026 265877
rect 449974 265813 450026 265819
rect 447670 264687 447722 264693
rect 447670 264629 447722 264635
rect 454786 264471 454814 278018
rect 455938 268837 455966 278018
rect 455926 268831 455978 268837
rect 455926 268773 455978 268779
rect 457090 265951 457118 278018
rect 458242 277569 458270 278018
rect 458230 277563 458282 277569
rect 458230 277505 458282 277511
rect 459490 271723 459518 278018
rect 460642 274757 460670 278018
rect 460630 274751 460682 274757
rect 460630 274693 460682 274699
rect 459478 271717 459530 271723
rect 459478 271659 459530 271665
rect 457078 265945 457130 265951
rect 457078 265887 457130 265893
rect 461794 264619 461822 278018
rect 463042 268911 463070 278018
rect 463030 268905 463082 268911
rect 463030 268847 463082 268853
rect 464194 266025 464222 278018
rect 465346 277495 465374 278018
rect 465334 277489 465386 277495
rect 465334 277431 465386 277437
rect 466594 271797 466622 278018
rect 467746 274831 467774 278018
rect 467734 274825 467786 274831
rect 467734 274767 467786 274773
rect 466582 271791 466634 271797
rect 466582 271733 466634 271739
rect 464182 266019 464234 266025
rect 464182 265961 464234 265967
rect 461782 264613 461834 264619
rect 461782 264555 461834 264561
rect 468898 264545 468926 278018
rect 470146 268985 470174 278018
rect 470134 268979 470186 268985
rect 470134 268921 470186 268927
rect 471298 266099 471326 278018
rect 472450 277421 472478 278018
rect 472438 277415 472490 277421
rect 472438 277357 472490 277363
rect 473698 271871 473726 278018
rect 474850 274355 474878 278018
rect 474836 274346 474892 274355
rect 474836 274281 474892 274290
rect 473686 271865 473738 271871
rect 473686 271807 473738 271813
rect 471286 266093 471338 266099
rect 471286 266035 471338 266041
rect 476002 264841 476030 278018
rect 477154 269133 477182 278018
rect 477142 269127 477194 269133
rect 477142 269069 477194 269075
rect 478402 266173 478430 278018
rect 479554 277347 479582 278018
rect 479542 277341 479594 277347
rect 479542 277283 479594 277289
rect 480706 271945 480734 278018
rect 481954 274905 481982 278018
rect 481942 274899 481994 274905
rect 481942 274841 481994 274847
rect 480694 271939 480746 271945
rect 480694 271881 480746 271887
rect 483106 269207 483134 278018
rect 484258 270687 484286 278018
rect 484246 270681 484298 270687
rect 484246 270623 484298 270629
rect 483094 269201 483146 269207
rect 483094 269143 483146 269149
rect 485506 266247 485534 278018
rect 486658 272019 486686 278018
rect 487810 272093 487838 278018
rect 489058 274503 489086 278018
rect 489044 274494 489100 274503
rect 489044 274429 489100 274438
rect 487798 272087 487850 272093
rect 487798 272029 487850 272035
rect 486646 272013 486698 272019
rect 486646 271955 486698 271961
rect 490210 270613 490238 278018
rect 490198 270607 490250 270613
rect 490198 270549 490250 270555
rect 491362 270539 491390 278018
rect 491350 270533 491402 270539
rect 491350 270475 491402 270481
rect 492610 266321 492638 278018
rect 493762 273499 493790 278018
rect 494914 273573 494942 278018
rect 496066 274651 496094 278018
rect 496052 274642 496108 274651
rect 496052 274577 496108 274586
rect 494902 273567 494954 273573
rect 494902 273509 494954 273515
rect 493750 273493 493802 273499
rect 493750 273435 493802 273441
rect 497314 270465 497342 278018
rect 497302 270459 497354 270465
rect 497302 270401 497354 270407
rect 498466 270391 498494 278018
rect 498454 270385 498506 270391
rect 498454 270327 498506 270333
rect 499618 267801 499646 278018
rect 500866 273425 500894 278018
rect 500854 273419 500906 273425
rect 500854 273361 500906 273367
rect 502018 273351 502046 278018
rect 503170 274799 503198 278018
rect 503156 274790 503212 274799
rect 503156 274725 503212 274734
rect 502006 273345 502058 273351
rect 502006 273287 502058 273293
rect 504418 270243 504446 278018
rect 505570 270317 505598 278018
rect 505558 270311 505610 270317
rect 505558 270253 505610 270259
rect 504406 270237 504458 270243
rect 504406 270179 504458 270185
rect 499606 267795 499658 267801
rect 499606 267737 499658 267743
rect 506722 267727 506750 278018
rect 507970 273203 507998 278018
rect 509122 273277 509150 278018
rect 510274 274979 510302 278018
rect 510262 274973 510314 274979
rect 510262 274915 510314 274921
rect 509110 273271 509162 273277
rect 509110 273213 509162 273219
rect 507958 273197 508010 273203
rect 507958 273139 508010 273145
rect 508246 273197 508298 273203
rect 508246 273139 508298 273145
rect 506710 267721 506762 267727
rect 506710 267663 506762 267669
rect 492598 266315 492650 266321
rect 492598 266257 492650 266263
rect 485494 266241 485546 266247
rect 485494 266183 485546 266189
rect 478390 266167 478442 266173
rect 478390 266109 478442 266115
rect 508258 265581 508286 273139
rect 511522 270169 511550 278018
rect 511510 270163 511562 270169
rect 511510 270105 511562 270111
rect 512674 270095 512702 278018
rect 512662 270089 512714 270095
rect 512662 270031 512714 270037
rect 513826 267653 513854 278018
rect 514978 273129 515006 278018
rect 514966 273123 515018 273129
rect 514966 273065 515018 273071
rect 516226 273055 516254 278018
rect 517378 276459 517406 278018
rect 517366 276453 517418 276459
rect 517366 276395 517418 276401
rect 516214 273049 516266 273055
rect 516214 272991 516266 272997
rect 516310 273049 516362 273055
rect 516310 272991 516362 272997
rect 516322 269059 516350 272991
rect 518530 270021 518558 278018
rect 518518 270015 518570 270021
rect 518518 269957 518570 269963
rect 519778 269947 519806 278018
rect 519766 269941 519818 269947
rect 519766 269883 519818 269889
rect 516310 269053 516362 269059
rect 516310 268995 516362 269001
rect 513814 267647 513866 267653
rect 513814 267589 513866 267595
rect 520930 267579 520958 278018
rect 522082 272981 522110 278018
rect 522548 276862 522604 276871
rect 522548 276797 522604 276806
rect 522562 273573 522590 276797
rect 522550 273567 522602 273573
rect 522550 273509 522602 273515
rect 522070 272975 522122 272981
rect 522070 272917 522122 272923
rect 523330 272907 523358 278018
rect 524482 276385 524510 278018
rect 524470 276379 524522 276385
rect 524470 276321 524522 276327
rect 523318 272901 523370 272907
rect 523318 272843 523370 272849
rect 523798 272901 523850 272907
rect 523798 272843 523850 272849
rect 523810 268879 523838 272843
rect 525634 269873 525662 278018
rect 525622 269867 525674 269873
rect 525622 269809 525674 269815
rect 526882 269799 526910 278018
rect 526870 269793 526922 269799
rect 526870 269735 526922 269741
rect 523796 268870 523852 268879
rect 523796 268805 523852 268814
rect 520918 267573 520970 267579
rect 520918 267515 520970 267521
rect 528034 267505 528062 278018
rect 529186 272833 529214 278018
rect 529844 276714 529900 276723
rect 529844 276649 529900 276658
rect 529858 273499 529886 276649
rect 529846 273493 529898 273499
rect 529846 273435 529898 273441
rect 529174 272827 529226 272833
rect 529174 272769 529226 272775
rect 530434 272759 530462 278018
rect 531586 276311 531614 278018
rect 531574 276305 531626 276311
rect 531574 276247 531626 276253
rect 530422 272753 530474 272759
rect 530422 272695 530474 272701
rect 532738 269725 532766 278018
rect 532726 269719 532778 269725
rect 532726 269661 532778 269667
rect 533890 268097 533918 278018
rect 533878 268091 533930 268097
rect 533878 268033 533930 268039
rect 528022 267499 528074 267505
rect 528022 267441 528074 267447
rect 535138 267431 535166 278018
rect 536290 272685 536318 278018
rect 536278 272679 536330 272685
rect 536278 272621 536330 272627
rect 537442 272611 537470 278018
rect 538690 276237 538718 278018
rect 538678 276231 538730 276237
rect 538678 276173 538730 276179
rect 537430 272605 537482 272611
rect 537430 272547 537482 272553
rect 539842 269175 539870 278018
rect 539828 269166 539884 269175
rect 539828 269101 539884 269110
rect 540994 269027 541022 278018
rect 540980 269018 541036 269027
rect 540980 268953 541036 268962
rect 535126 267425 535178 267431
rect 535126 267367 535178 267373
rect 542242 267357 542270 278018
rect 543394 271839 543422 278018
rect 544546 271987 544574 278018
rect 545794 276163 545822 278018
rect 545782 276157 545834 276163
rect 545782 276099 545834 276105
rect 546946 276015 546974 278018
rect 546934 276009 546986 276015
rect 546934 275951 546986 275957
rect 544532 271978 544588 271987
rect 544532 271913 544588 271922
rect 543380 271830 543436 271839
rect 543380 271765 543436 271774
rect 548098 269577 548126 278018
rect 549346 276089 549374 278018
rect 549334 276083 549386 276089
rect 549334 276025 549386 276031
rect 548086 269571 548138 269577
rect 548086 269513 548138 269519
rect 542230 267351 542282 267357
rect 542230 267293 542282 267299
rect 550498 267283 550526 278018
rect 551650 272537 551678 278018
rect 552802 275941 552830 278018
rect 554050 277273 554078 278018
rect 554038 277267 554090 277273
rect 554038 277209 554090 277215
rect 552790 275935 552842 275941
rect 552790 275877 552842 275883
rect 551638 272531 551690 272537
rect 551638 272473 551690 272479
rect 555202 270507 555230 278018
rect 556354 275867 556382 278018
rect 557602 277199 557630 278018
rect 557590 277193 557642 277199
rect 557590 277135 557642 277141
rect 556342 275861 556394 275867
rect 556342 275803 556394 275809
rect 558754 273467 558782 278018
rect 559906 275719 559934 278018
rect 561154 277125 561182 278018
rect 561142 277119 561194 277125
rect 561142 277061 561194 277067
rect 559894 275713 559946 275719
rect 559894 275655 559946 275661
rect 558740 273458 558796 273467
rect 558740 273393 558796 273402
rect 555188 270498 555244 270507
rect 555188 270433 555244 270442
rect 562306 270359 562334 278018
rect 563458 275793 563486 278018
rect 564706 277051 564734 278018
rect 564694 277045 564746 277051
rect 564694 276987 564746 276993
rect 563446 275787 563498 275793
rect 563446 275729 563498 275735
rect 565858 273319 565886 278018
rect 567010 274947 567038 278018
rect 568258 276977 568286 278018
rect 568246 276971 568298 276977
rect 568246 276913 568298 276919
rect 566996 274938 567052 274947
rect 566996 274873 567052 274882
rect 565844 273310 565900 273319
rect 565844 273245 565900 273254
rect 562292 270350 562348 270359
rect 562292 270285 562348 270294
rect 569410 269503 569438 278018
rect 570562 275645 570590 278018
rect 571714 276903 571742 278018
rect 571702 276897 571754 276903
rect 571702 276839 571754 276845
rect 570550 275639 570602 275645
rect 570550 275581 570602 275587
rect 572962 272463 572990 278018
rect 574114 275571 574142 278018
rect 574978 278004 575280 278032
rect 574978 277939 575006 278004
rect 574966 277933 575018 277939
rect 574966 277875 575018 277881
rect 574102 275565 574154 275571
rect 574102 275507 574154 275513
rect 576514 273171 576542 278018
rect 577666 275983 577694 278018
rect 578818 276829 578846 278018
rect 578806 276823 578858 276829
rect 578806 276765 578858 276771
rect 577652 275974 577708 275983
rect 577652 275909 577708 275918
rect 576500 273162 576556 273171
rect 576500 273097 576556 273106
rect 580066 273055 580094 278018
rect 580054 273049 580106 273055
rect 580054 272991 580106 272997
rect 572950 272457 573002 272463
rect 572950 272399 573002 272405
rect 569398 269497 569450 269503
rect 569398 269439 569450 269445
rect 550486 267277 550538 267283
rect 550486 267219 550538 267225
rect 581218 267209 581246 278018
rect 582370 276607 582398 278018
rect 582358 276601 582410 276607
rect 582358 276543 582410 276549
rect 583618 270211 583646 278018
rect 583604 270202 583660 270211
rect 583604 270137 583660 270146
rect 581206 267203 581258 267209
rect 581206 267145 581258 267151
rect 584770 267135 584798 278018
rect 585922 276681 585950 278018
rect 585910 276675 585962 276681
rect 585910 276617 585962 276623
rect 587170 272389 587198 278018
rect 587158 272383 587210 272389
rect 587158 272325 587210 272331
rect 584758 267129 584810 267135
rect 584758 267071 584810 267077
rect 588322 267061 588350 278018
rect 588310 267055 588362 267061
rect 588310 266997 588362 267003
rect 508246 265575 508298 265581
rect 508246 265517 508298 265523
rect 475990 264835 476042 264841
rect 475990 264777 476042 264783
rect 468886 264539 468938 264545
rect 468886 264481 468938 264487
rect 454774 264465 454826 264471
rect 454774 264407 454826 264413
rect 433462 264095 433514 264101
rect 433462 264037 433514 264043
rect 589474 264027 589502 278018
rect 590626 270063 590654 278018
rect 591874 275497 591902 278018
rect 591862 275491 591914 275497
rect 591862 275433 591914 275439
rect 593026 275423 593054 278018
rect 593014 275417 593066 275423
rect 593014 275359 593066 275365
rect 594178 273023 594206 278018
rect 595426 275835 595454 278018
rect 595412 275826 595468 275835
rect 595412 275761 595468 275770
rect 594164 273014 594220 273023
rect 594164 272949 594220 272958
rect 590612 270054 590668 270063
rect 590612 269989 590668 269998
rect 589462 264021 589514 264027
rect 589462 263963 589514 263969
rect 596578 263953 596606 278018
rect 597730 269915 597758 278018
rect 598978 275349 599006 278018
rect 600130 276533 600158 278018
rect 600118 276527 600170 276533
rect 600118 276469 600170 276475
rect 598966 275343 599018 275349
rect 598966 275285 599018 275291
rect 601282 272875 601310 278018
rect 601268 272866 601324 272875
rect 601268 272801 601324 272810
rect 597716 269906 597772 269915
rect 597716 269841 597772 269850
rect 602530 266913 602558 278018
rect 602518 266907 602570 266913
rect 602518 266849 602570 266855
rect 596566 263947 596618 263953
rect 596566 263889 596618 263895
rect 603682 263879 603710 278018
rect 604834 269429 604862 278018
rect 604822 269423 604874 269429
rect 604822 269365 604874 269371
rect 606082 266987 606110 278018
rect 607234 276575 607262 278018
rect 607220 276566 607276 276575
rect 607220 276501 607276 276510
rect 608386 272315 608414 278018
rect 609538 275275 609566 278018
rect 609526 275269 609578 275275
rect 609526 275211 609578 275217
rect 608374 272309 608426 272315
rect 608374 272251 608426 272257
rect 606070 266981 606122 266987
rect 606070 266923 606122 266929
rect 603670 263873 603722 263879
rect 411778 263796 411840 263824
rect 603670 263815 603722 263821
rect 610786 263805 610814 278018
rect 611938 272907 611966 278018
rect 611926 272901 611978 272907
rect 611926 272843 611978 272849
rect 613090 266839 613118 278018
rect 613078 266833 613130 266839
rect 613078 266775 613130 266781
rect 614338 266765 614366 278018
rect 615490 272727 615518 278018
rect 616642 275687 616670 278018
rect 616628 275678 616684 275687
rect 616628 275613 616684 275622
rect 615476 272718 615532 272727
rect 615476 272653 615532 272662
rect 614326 266759 614378 266765
rect 614326 266701 614378 266707
rect 610774 263799 610826 263805
rect 610774 263741 610826 263747
rect 617890 263731 617918 278018
rect 619042 269355 619070 278018
rect 619030 269349 619082 269355
rect 619030 269291 619082 269297
rect 620194 266691 620222 278018
rect 620182 266685 620234 266691
rect 620182 266627 620234 266633
rect 401110 263725 401162 263731
rect 345442 263648 345504 263676
rect 400896 263673 401110 263676
rect 410998 263725 411050 263731
rect 400896 263667 401162 263673
rect 400896 263648 401150 263667
rect 403728 263657 404030 263676
rect 410998 263667 411050 263673
rect 617878 263725 617930 263731
rect 617878 263667 617930 263673
rect 621442 263657 621470 278018
rect 622594 272241 622622 278018
rect 623746 275201 623774 278018
rect 623734 275195 623786 275201
rect 623734 275137 623786 275143
rect 624994 273499 625022 278018
rect 624982 273493 625034 273499
rect 624982 273435 625034 273441
rect 622582 272235 622634 272241
rect 622582 272177 622634 272183
rect 626146 269767 626174 278018
rect 626132 269758 626188 269767
rect 626132 269693 626188 269702
rect 627298 266617 627326 278018
rect 627286 266611 627338 266617
rect 627286 266553 627338 266559
rect 403728 263651 404042 263657
rect 403728 263648 403990 263651
rect 403990 263593 404042 263599
rect 621430 263651 621482 263657
rect 621430 263593 621482 263599
rect 628450 263583 628478 278018
rect 629698 272579 629726 278018
rect 630850 275053 630878 278018
rect 630838 275047 630890 275053
rect 630838 274989 630890 274995
rect 632002 273573 632030 278018
rect 631990 273567 632042 273573
rect 631990 273509 632042 273515
rect 629684 272570 629740 272579
rect 629684 272505 629740 272514
rect 633250 269619 633278 278018
rect 633236 269610 633292 269619
rect 633236 269545 633292 269554
rect 634402 266543 634430 278018
rect 635554 275127 635582 278018
rect 635542 275121 635594 275127
rect 635542 275063 635594 275069
rect 636802 272431 636830 278018
rect 637954 275539 637982 278018
rect 637940 275530 637996 275539
rect 637940 275465 637996 275474
rect 639106 273203 639134 278018
rect 639094 273197 639146 273203
rect 639094 273139 639146 273145
rect 636788 272422 636844 272431
rect 636788 272357 636844 272366
rect 640354 268245 640382 278018
rect 640342 268239 640394 268245
rect 640342 268181 640394 268187
rect 634390 266537 634442 266543
rect 634390 266479 634442 266485
rect 641506 266469 641534 278018
rect 641494 266463 641546 266469
rect 641494 266405 641546 266411
rect 409654 263577 409706 263583
rect 409440 263525 409654 263528
rect 409440 263519 409706 263525
rect 628438 263577 628490 263583
rect 628438 263519 628490 263525
rect 409440 263500 409694 263519
rect 642658 263509 642686 278018
rect 643906 272167 643934 278018
rect 643894 272161 643946 272167
rect 643894 272103 643946 272109
rect 645058 269471 645086 278018
rect 646210 272283 646238 278018
rect 646484 275382 646540 275391
rect 646484 275317 646540 275326
rect 646196 272274 646252 272283
rect 646196 272209 646252 272218
rect 645044 269462 645100 269471
rect 645044 269397 645100 269406
rect 642646 263503 642698 263509
rect 642646 263445 642698 263451
rect 420404 262210 420460 262219
rect 420404 262145 420406 262154
rect 420458 262145 420460 262154
rect 606166 262171 606218 262177
rect 420406 262113 420458 262119
rect 606166 262113 606218 262119
rect 420404 259842 420460 259851
rect 420404 259777 420460 259786
rect 191540 259398 191596 259407
rect 191540 259333 191596 259342
rect 190196 251702 190252 251711
rect 190196 251637 190252 251646
rect 190210 228581 190238 251637
rect 190198 228575 190250 228581
rect 190198 228517 190250 228523
rect 190774 227539 190826 227545
rect 190774 227481 190826 227487
rect 190786 221792 190814 227481
rect 190786 221764 190862 221792
rect 190834 221482 190862 221764
rect 191554 221482 191582 259333
rect 420418 259291 420446 259777
rect 420406 259285 420458 259291
rect 420406 259227 420458 259233
rect 420404 257030 420460 257039
rect 420404 256965 420460 256974
rect 420418 256405 420446 256965
rect 420406 256399 420458 256405
rect 420406 256341 420458 256347
rect 420404 255254 420460 255263
rect 420404 255189 420460 255198
rect 420418 253519 420446 255189
rect 420406 253513 420458 253519
rect 420406 253455 420458 253461
rect 603286 253513 603338 253519
rect 603286 253455 603338 253461
rect 420404 252886 420460 252895
rect 420404 252821 420460 252830
rect 420418 250633 420446 252821
rect 420406 250627 420458 250633
rect 420406 250569 420458 250575
rect 420308 250518 420364 250527
rect 420308 250453 420364 250462
rect 420322 247821 420350 250453
rect 420404 248150 420460 248159
rect 420404 248085 420460 248094
rect 420310 247815 420362 247821
rect 420310 247757 420362 247763
rect 420418 247747 420446 248085
rect 420406 247741 420458 247747
rect 420406 247683 420458 247689
rect 420404 245338 420460 245347
rect 420404 245273 420460 245282
rect 420418 244861 420446 245273
rect 420406 244855 420458 244861
rect 420406 244797 420458 244803
rect 420308 243562 420364 243571
rect 420308 243497 420364 243506
rect 420322 241975 420350 243497
rect 420310 241969 420362 241975
rect 420310 241911 420362 241917
rect 600406 241969 600458 241975
rect 600406 241911 600458 241917
rect 420308 241194 420364 241203
rect 420308 241129 420364 241138
rect 412244 240306 412300 240315
rect 412244 240241 412300 240250
rect 412148 240158 412204 240167
rect 412148 240093 412204 240102
rect 412052 240010 412108 240019
rect 380640 239977 380894 239996
rect 380640 239971 380906 239977
rect 380640 239968 380854 239971
rect 412052 239945 412054 239954
rect 380854 239913 380906 239919
rect 412106 239945 412108 239954
rect 412054 239913 412106 239919
rect 412162 239903 412190 240093
rect 409558 239897 409610 239903
rect 409344 239845 409558 239848
rect 409344 239839 409610 239845
rect 412150 239897 412202 239903
rect 412150 239839 412202 239845
rect 360022 239823 360074 239829
rect 409344 239820 409598 239839
rect 360022 239765 360074 239771
rect 192418 233391 192446 239686
rect 192768 239672 192926 239700
rect 192898 233613 192926 239672
rect 193090 239672 193152 239700
rect 192886 233607 192938 233613
rect 192886 233549 192938 233555
rect 192406 233385 192458 233391
rect 192406 233327 192458 233333
rect 192310 228575 192362 228581
rect 192310 228517 192362 228523
rect 192322 221482 192350 228517
rect 193090 221792 193118 239672
rect 193474 233317 193502 239686
rect 193858 233391 193886 239686
rect 194242 233539 194270 239686
rect 194230 233533 194282 233539
rect 194230 233475 194282 233481
rect 194626 233465 194654 239686
rect 194976 239672 195230 239700
rect 195360 239672 195614 239700
rect 194614 233459 194666 233465
rect 194614 233401 194666 233407
rect 193750 233385 193802 233391
rect 193750 233327 193802 233333
rect 193846 233385 193898 233391
rect 193846 233327 193898 233333
rect 193462 233311 193514 233317
rect 193462 233253 193514 233259
rect 193042 221764 193118 221792
rect 193042 221482 193070 221764
rect 193762 221482 193790 233327
rect 195202 233317 195230 239672
rect 195586 233613 195614 239672
rect 195682 233687 195710 239686
rect 195670 233681 195722 233687
rect 195670 233623 195722 233629
rect 195286 233607 195338 233613
rect 195286 233549 195338 233555
rect 195574 233607 195626 233613
rect 195574 233549 195626 233555
rect 194614 233311 194666 233317
rect 194614 233253 194666 233259
rect 195190 233311 195242 233317
rect 195190 233253 195242 233259
rect 194626 221482 194654 233253
rect 195298 221792 195326 233549
rect 196162 233465 196190 239686
rect 196546 233761 196574 239686
rect 196930 233835 196958 239686
rect 197280 239672 197534 239700
rect 197664 239672 197918 239700
rect 197506 233983 197534 239672
rect 197494 233977 197546 233983
rect 197494 233919 197546 233925
rect 196918 233829 196970 233835
rect 196918 233771 196970 233777
rect 196534 233755 196586 233761
rect 196534 233697 196586 233703
rect 196054 233459 196106 233465
rect 196054 233401 196106 233407
rect 196150 233459 196202 233465
rect 196150 233401 196202 233407
rect 195298 221764 195374 221792
rect 195346 221482 195374 221764
rect 196066 221482 196094 233401
rect 196822 233385 196874 233391
rect 196822 233327 196874 233333
rect 196834 221482 196862 233327
rect 197890 233317 197918 239672
rect 197986 233391 198014 239686
rect 198370 234057 198398 239686
rect 198754 234131 198782 239686
rect 198742 234125 198794 234131
rect 198742 234067 198794 234073
rect 198358 234051 198410 234057
rect 198358 233993 198410 233999
rect 199138 233909 199166 239686
rect 199488 239672 199742 239700
rect 199968 239672 200222 239700
rect 199126 233903 199178 233909
rect 199126 233845 199178 233851
rect 198358 233533 198410 233539
rect 198358 233475 198410 233481
rect 197974 233385 198026 233391
rect 197974 233327 198026 233333
rect 197494 233311 197546 233317
rect 197494 233253 197546 233259
rect 197878 233311 197930 233317
rect 197878 233253 197930 233259
rect 197506 221792 197534 233253
rect 197506 221764 197582 221792
rect 197554 221482 197582 221764
rect 198370 221482 198398 233475
rect 199714 233465 199742 239672
rect 200194 234205 200222 239672
rect 200290 234279 200318 239686
rect 200278 234273 200330 234279
rect 200278 234215 200330 234221
rect 200182 234199 200234 234205
rect 200182 234141 200234 234147
rect 200566 233755 200618 233761
rect 200566 233697 200618 233703
rect 199798 233607 199850 233613
rect 199798 233549 199850 233555
rect 199126 233459 199178 233465
rect 199126 233401 199178 233407
rect 199702 233459 199754 233465
rect 199702 233401 199754 233407
rect 199138 221482 199166 233401
rect 199810 221792 199838 233549
rect 199810 221764 199886 221792
rect 199858 221482 199886 221764
rect 200578 221482 200606 233697
rect 200674 233539 200702 239686
rect 201058 233613 201086 239686
rect 201408 239672 201566 239700
rect 201792 239672 202046 239700
rect 202176 239672 202430 239700
rect 201538 233761 201566 239672
rect 202018 234501 202046 239672
rect 202006 234495 202058 234501
rect 202006 234437 202058 234443
rect 201526 233755 201578 233761
rect 201526 233697 201578 233703
rect 201334 233681 201386 233687
rect 201334 233623 201386 233629
rect 201046 233607 201098 233613
rect 201046 233549 201098 233555
rect 200662 233533 200714 233539
rect 200662 233475 200714 233481
rect 201346 221482 201374 233623
rect 202402 233317 202430 239672
rect 202498 233687 202526 239686
rect 202882 234575 202910 239686
rect 203266 234797 203294 239686
rect 203712 239672 203966 239700
rect 204096 239672 204254 239700
rect 203254 234791 203306 234797
rect 203254 234733 203306 234739
rect 202870 234569 202922 234575
rect 202870 234511 202922 234517
rect 202870 233829 202922 233835
rect 202870 233771 202922 233777
rect 202486 233681 202538 233687
rect 202486 233623 202538 233629
rect 202102 233311 202154 233317
rect 202102 233253 202154 233259
rect 202390 233311 202442 233317
rect 202390 233253 202442 233259
rect 202114 221792 202142 233253
rect 202114 221764 202190 221792
rect 202162 221482 202190 221764
rect 202882 221482 202910 233771
rect 203938 233391 203966 239672
rect 204226 233835 204254 239672
rect 204418 239672 204480 239700
rect 204418 233983 204446 239672
rect 204802 234649 204830 239686
rect 204790 234643 204842 234649
rect 204790 234585 204842 234591
rect 204310 233977 204362 233983
rect 204310 233919 204362 233925
rect 204406 233977 204458 233983
rect 204406 233919 204458 233925
rect 204214 233829 204266 233835
rect 204214 233771 204266 233777
rect 203638 233385 203690 233391
rect 203638 233327 203690 233333
rect 203926 233385 203978 233391
rect 203926 233327 203978 233333
rect 203650 221482 203678 233327
rect 204322 221792 204350 233919
rect 205186 233909 205214 239686
rect 205570 234723 205598 239686
rect 205920 239672 206174 239700
rect 206304 239672 206558 239700
rect 206688 239672 206942 239700
rect 205558 234717 205610 234723
rect 205558 234659 205610 234665
rect 206146 234427 206174 239672
rect 206530 234871 206558 239672
rect 206518 234865 206570 234871
rect 206518 234807 206570 234813
rect 206134 234421 206186 234427
rect 206134 234363 206186 234369
rect 205942 234051 205994 234057
rect 205942 233993 205994 233999
rect 205078 233903 205130 233909
rect 205078 233845 205130 233851
rect 205174 233903 205226 233909
rect 205174 233845 205226 233851
rect 204322 221764 204398 221792
rect 204370 221482 204398 221764
rect 205090 221482 205118 233845
rect 205954 221496 205982 233993
rect 206914 233983 206942 239672
rect 207010 235315 207038 239686
rect 207490 235981 207518 239686
rect 207478 235975 207530 235981
rect 207478 235917 207530 235923
rect 206998 235309 207050 235315
rect 206998 235251 207050 235257
rect 207286 234717 207338 234723
rect 207286 234659 207338 234665
rect 206902 233977 206954 233983
rect 206902 233919 206954 233925
rect 207298 233465 207326 234659
rect 207874 234353 207902 239686
rect 208224 239672 208478 239700
rect 208608 239672 208862 239700
rect 208450 236055 208478 239672
rect 208438 236049 208490 236055
rect 208438 235991 208490 235997
rect 208834 234945 208862 239672
rect 208930 235833 208958 239686
rect 208918 235827 208970 235833
rect 208918 235769 208970 235775
rect 208822 234939 208874 234945
rect 208822 234881 208874 234887
rect 209314 234797 209342 239686
rect 209698 235907 209726 239686
rect 209686 235901 209738 235907
rect 209686 235843 209738 235849
rect 210082 235611 210110 239686
rect 210432 239672 210686 239700
rect 210816 239672 211070 239700
rect 210658 235685 210686 239672
rect 210646 235679 210698 235685
rect 210646 235621 210698 235627
rect 210070 235605 210122 235611
rect 210070 235547 210122 235553
rect 211042 235019 211070 239672
rect 211234 235759 211262 239686
rect 211222 235753 211274 235759
rect 211222 235695 211274 235701
rect 211618 235167 211646 239686
rect 212002 235463 212030 239686
rect 211990 235457 212042 235463
rect 211990 235399 212042 235405
rect 211606 235161 211658 235167
rect 211606 235103 211658 235109
rect 211030 235013 211082 235019
rect 211030 234955 211082 234961
rect 209302 234791 209354 234797
rect 209302 234733 209354 234739
rect 211990 234643 212042 234649
rect 211990 234585 212042 234591
rect 207862 234347 207914 234353
rect 207862 234289 207914 234295
rect 212002 234279 212030 234585
rect 210358 234273 210410 234279
rect 210358 234215 210410 234221
rect 211990 234273 212042 234279
rect 211990 234215 212042 234221
rect 208822 234199 208874 234205
rect 208822 234141 208874 234147
rect 207382 234125 207434 234131
rect 207382 234067 207434 234073
rect 206614 233459 206666 233465
rect 206614 233401 206666 233407
rect 207286 233459 207338 233465
rect 207286 233401 207338 233407
rect 205920 221468 205982 221496
rect 206626 221496 206654 233401
rect 206626 221468 206688 221496
rect 207394 221482 207422 234067
rect 208150 233533 208202 233539
rect 208150 233475 208202 233481
rect 208162 221496 208190 233475
rect 208128 221468 208190 221496
rect 208834 221496 208862 234141
rect 209686 233607 209738 233613
rect 209686 233549 209738 233555
rect 208834 221468 208896 221496
rect 209698 221482 209726 233549
rect 210370 221792 210398 234215
rect 211894 233755 211946 233761
rect 211894 233697 211946 233703
rect 211126 233311 211178 233317
rect 211126 233253 211178 233259
rect 210370 221764 210446 221792
rect 210418 221482 210446 221764
rect 211138 221482 211166 233253
rect 211906 221482 211934 233697
rect 212386 226361 212414 239686
rect 212736 239672 212990 239700
rect 212962 235537 212990 239672
rect 213058 239672 213120 239700
rect 212950 235531 213002 235537
rect 212950 235473 213002 235479
rect 212566 233681 212618 233687
rect 212566 233623 212618 233629
rect 212374 226355 212426 226361
rect 212374 226297 212426 226303
rect 212578 221792 212606 233623
rect 213058 225991 213086 239672
rect 213442 235093 213470 239686
rect 213430 235087 213482 235093
rect 213430 235029 213482 235035
rect 213430 234495 213482 234501
rect 213430 234437 213482 234443
rect 213046 225985 213098 225991
rect 213046 225927 213098 225933
rect 212578 221764 212654 221792
rect 212626 221482 212654 221764
rect 213442 221482 213470 234437
rect 213826 227027 213854 239686
rect 214210 235389 214238 239686
rect 214198 235383 214250 235389
rect 214198 235325 214250 235331
rect 214198 233385 214250 233391
rect 214198 233327 214250 233333
rect 213814 227021 213866 227027
rect 213814 226963 213866 226969
rect 214210 221482 214238 233327
rect 214594 226065 214622 239686
rect 215040 239672 215294 239700
rect 215424 239672 215678 239700
rect 214870 234569 214922 234575
rect 214870 234511 214922 234517
rect 214582 226059 214634 226065
rect 214582 226001 214634 226007
rect 214882 221792 214910 234511
rect 215266 229691 215294 239672
rect 215542 233829 215594 233835
rect 215542 233771 215594 233777
rect 215254 229685 215306 229691
rect 215254 229627 215306 229633
rect 215554 226084 215582 233771
rect 215650 226213 215678 239672
rect 215746 227175 215774 239686
rect 215830 234717 215882 234723
rect 215830 234659 215882 234665
rect 215842 233909 215870 234659
rect 215830 233903 215882 233909
rect 215830 233845 215882 233851
rect 216130 227545 216158 239686
rect 216514 236174 216542 239686
rect 216864 239672 217118 239700
rect 217248 239672 217502 239700
rect 217632 239672 217886 239700
rect 216514 236146 216638 236174
rect 216502 233903 216554 233909
rect 216502 233845 216554 233851
rect 216118 227539 216170 227545
rect 216118 227481 216170 227487
rect 215734 227169 215786 227175
rect 215734 227111 215786 227117
rect 215638 226207 215690 226213
rect 215638 226149 215690 226155
rect 215554 226056 215678 226084
rect 214882 221764 214958 221792
rect 214930 221482 214958 221764
rect 215650 221482 215678 226056
rect 216514 221482 216542 233845
rect 216610 232725 216638 236146
rect 216598 232719 216650 232725
rect 216598 232661 216650 232667
rect 217090 227397 217118 239672
rect 217174 233755 217226 233761
rect 217174 233697 217226 233703
rect 217078 227391 217130 227397
rect 217078 227333 217130 227339
rect 217186 221792 217214 233697
rect 217474 225917 217502 239672
rect 217858 227249 217886 239672
rect 217954 236174 217982 239686
rect 217954 236146 218078 236174
rect 217942 234051 217994 234057
rect 217942 233993 217994 233999
rect 217846 227243 217898 227249
rect 217846 227185 217898 227191
rect 217462 225911 217514 225917
rect 217462 225853 217514 225859
rect 217186 221764 217262 221792
rect 217234 221482 217262 221764
rect 217954 221482 217982 233993
rect 218050 232651 218078 236146
rect 218038 232645 218090 232651
rect 218038 232587 218090 232593
rect 218338 225769 218366 239686
rect 218710 233607 218762 233613
rect 218710 233549 218762 233555
rect 218326 225763 218378 225769
rect 218326 225705 218378 225711
rect 218722 221482 218750 233549
rect 218818 225843 218846 239686
rect 219168 239672 219422 239700
rect 219552 239672 219806 239700
rect 219936 239672 220190 239700
rect 219394 236174 219422 239672
rect 219394 236146 219518 236174
rect 219382 234273 219434 234279
rect 219382 234215 219434 234221
rect 218806 225837 218858 225843
rect 218806 225779 218858 225785
rect 219394 221792 219422 234215
rect 219490 227101 219518 236146
rect 219778 232577 219806 239672
rect 219766 232571 219818 232577
rect 219766 232513 219818 232519
rect 220162 229617 220190 239672
rect 220258 236174 220286 239686
rect 220258 236146 220382 236174
rect 220246 233977 220298 233983
rect 220246 233919 220298 233925
rect 220150 229611 220202 229617
rect 220150 229553 220202 229559
rect 219478 227095 219530 227101
rect 219478 227037 219530 227043
rect 219394 221764 219470 221792
rect 219442 221482 219470 221764
rect 220258 221482 220286 233919
rect 220354 226287 220382 236146
rect 220642 235241 220670 239686
rect 221026 236174 221054 239686
rect 221376 239672 221630 239700
rect 221026 236146 221150 236174
rect 220630 235235 220682 235241
rect 220630 235177 220682 235183
rect 221014 234421 221066 234427
rect 221014 234363 221066 234369
rect 220342 226281 220394 226287
rect 220342 226223 220394 226229
rect 221026 221482 221054 234363
rect 221122 232503 221150 236146
rect 221110 232497 221162 232503
rect 221110 232439 221162 232445
rect 221602 229543 221630 239672
rect 221746 239404 221774 239686
rect 222144 239672 222398 239700
rect 221698 239376 221774 239404
rect 221590 229537 221642 229543
rect 221590 229479 221642 229485
rect 221698 226953 221726 239376
rect 222370 236129 222398 239672
rect 222358 236123 222410 236129
rect 222358 236065 222410 236071
rect 221782 235309 221834 235315
rect 221782 235251 221834 235257
rect 221686 226947 221738 226953
rect 221686 226889 221738 226895
rect 221794 221755 221822 235251
rect 222454 234865 222506 234871
rect 222454 234807 222506 234813
rect 221746 221727 221822 221755
rect 221746 221482 221774 221727
rect 222466 221482 222494 234807
rect 222562 232429 222590 239686
rect 222550 232423 222602 232429
rect 222550 232365 222602 232371
rect 222946 232355 222974 239686
rect 223222 236049 223274 236055
rect 223222 235991 223274 235997
rect 222934 232349 222986 232355
rect 222934 232291 222986 232297
rect 223234 221482 223262 235991
rect 223330 226879 223358 239686
rect 223680 239672 223934 239700
rect 224064 239672 224318 239700
rect 223906 235315 223934 239672
rect 223990 235975 224042 235981
rect 223990 235917 224042 235923
rect 223894 235309 223946 235315
rect 223894 235251 223946 235257
rect 223318 226873 223370 226879
rect 223318 226815 223370 226821
rect 224002 221792 224030 235917
rect 224290 232281 224318 239672
rect 224278 232275 224330 232281
rect 224278 232217 224330 232223
rect 224386 228507 224414 239686
rect 224784 239672 224990 239700
rect 224758 234939 224810 234945
rect 224758 234881 224810 234887
rect 224374 228501 224426 228507
rect 224374 228443 224426 228449
rect 224002 221764 224078 221792
rect 224050 221482 224078 221764
rect 224770 221482 224798 234881
rect 224962 226805 224990 239672
rect 225154 234723 225182 239686
rect 225538 234945 225566 239686
rect 225984 239672 226238 239700
rect 226368 239672 226622 239700
rect 226210 236174 226238 239672
rect 226210 236146 226334 236174
rect 226198 235901 226250 235907
rect 226198 235843 226250 235849
rect 225526 234939 225578 234945
rect 225526 234881 225578 234887
rect 225142 234717 225194 234723
rect 225142 234659 225194 234665
rect 225526 234199 225578 234205
rect 225526 234141 225578 234147
rect 224950 226799 225002 226805
rect 224950 226741 225002 226747
rect 225538 221482 225566 234141
rect 226210 221755 226238 235843
rect 226306 232207 226334 236146
rect 226294 232201 226346 232207
rect 226294 232143 226346 232149
rect 226594 226657 226622 239672
rect 226690 233465 226718 239686
rect 226966 235827 227018 235833
rect 226966 235769 227018 235775
rect 226678 233459 226730 233465
rect 226678 233401 226730 233407
rect 226582 226651 226634 226657
rect 226582 226593 226634 226599
rect 226210 221727 226286 221755
rect 226258 221482 226286 221727
rect 226978 221482 227006 235769
rect 227074 232133 227102 239686
rect 227062 232127 227114 232133
rect 227062 232069 227114 232075
rect 227458 230061 227486 239686
rect 227842 236174 227870 239686
rect 228192 239672 228446 239700
rect 228576 239672 228830 239700
rect 227842 236146 227966 236174
rect 227830 235605 227882 235611
rect 227830 235547 227882 235553
rect 227446 230055 227498 230061
rect 227446 229997 227498 230003
rect 227842 221482 227870 235547
rect 227938 226731 227966 236146
rect 228418 233391 228446 239672
rect 228502 234791 228554 234797
rect 228502 234733 228554 234739
rect 228406 233385 228458 233391
rect 228406 233327 228458 233333
rect 227926 226725 227978 226731
rect 227926 226667 227978 226673
rect 228514 221792 228542 234733
rect 228802 228581 228830 239672
rect 228898 230209 228926 239686
rect 229296 239672 229598 239700
rect 229270 235753 229322 235759
rect 229270 235695 229322 235701
rect 228886 230203 228938 230209
rect 228886 230145 228938 230151
rect 228790 228575 228842 228581
rect 228790 228517 228842 228523
rect 228514 221764 228590 221792
rect 228562 221482 228590 221764
rect 229282 221482 229310 235695
rect 229570 226583 229598 239672
rect 229762 234797 229790 239686
rect 230112 239672 230366 239700
rect 230496 239672 230654 239700
rect 230880 239672 231134 239700
rect 230038 235679 230090 235685
rect 230038 235621 230090 235627
rect 229750 234791 229802 234797
rect 229750 234733 229802 234739
rect 229558 226577 229610 226583
rect 229558 226519 229610 226525
rect 230050 221482 230078 235621
rect 230338 229321 230366 239672
rect 230626 229395 230654 239672
rect 230710 235161 230762 235167
rect 230710 235103 230762 235109
rect 230614 229389 230666 229395
rect 230614 229331 230666 229337
rect 230326 229315 230378 229321
rect 230326 229257 230378 229263
rect 230722 221792 230750 235103
rect 231106 226509 231134 239672
rect 231202 235759 231230 239686
rect 231600 239672 231902 239700
rect 231190 235753 231242 235759
rect 231190 235695 231242 235701
rect 231574 235013 231626 235019
rect 231574 234955 231626 234961
rect 231094 226503 231146 226509
rect 231094 226445 231146 226451
rect 230722 221764 230798 221792
rect 230770 221482 230798 221764
rect 231586 221482 231614 234955
rect 231874 228655 231902 239672
rect 231970 229173 231998 239686
rect 232320 239672 232574 239700
rect 232704 239672 232958 239700
rect 233088 239672 233246 239700
rect 232342 235531 232394 235537
rect 232342 235473 232394 235479
rect 231958 229167 232010 229173
rect 231958 229109 232010 229115
rect 231862 228649 231914 228655
rect 231862 228591 231914 228597
rect 232354 221482 232382 235473
rect 232546 226435 232574 239672
rect 232930 235167 232958 239672
rect 233014 235457 233066 235463
rect 233014 235399 233066 235405
rect 232918 235161 232970 235167
rect 232918 235103 232970 235109
rect 232534 226429 232586 226435
rect 232534 226371 232586 226377
rect 233026 221792 233054 235399
rect 233218 231985 233246 239672
rect 233206 231979 233258 231985
rect 233206 231921 233258 231927
rect 233506 229247 233534 239686
rect 233890 232059 233918 239686
rect 234274 235907 234302 239686
rect 234624 239672 234878 239700
rect 235008 239672 235262 239700
rect 235392 239672 235646 239700
rect 234262 235901 234314 235907
rect 234262 235843 234314 235849
rect 233878 232053 233930 232059
rect 233878 231995 233930 232001
rect 234850 231911 234878 239672
rect 234838 231905 234890 231911
rect 234838 231847 234890 231853
rect 233494 229241 233546 229247
rect 233494 229183 233546 229189
rect 235234 229099 235262 239672
rect 235318 235383 235370 235389
rect 235318 235325 235370 235331
rect 235222 229093 235274 229099
rect 235222 229035 235274 229041
rect 234550 226355 234602 226361
rect 234550 226297 234602 226303
rect 233782 225985 233834 225991
rect 233782 225927 233834 225933
rect 233026 221764 233102 221792
rect 233074 221482 233102 221764
rect 233794 221482 233822 225927
rect 234562 221482 234590 226297
rect 235330 221496 235358 235325
rect 235618 234575 235646 239672
rect 235714 235093 235742 239686
rect 235702 235087 235754 235093
rect 235702 235029 235754 235035
rect 235990 235013 236042 235019
rect 235990 234955 236042 234961
rect 235606 234569 235658 234575
rect 235606 234511 235658 234517
rect 236002 227534 236030 234955
rect 236098 231837 236126 239686
rect 236482 235685 236510 239686
rect 236832 239672 237086 239700
rect 237312 239672 237566 239700
rect 236470 235679 236522 235685
rect 236470 235621 236522 235627
rect 237058 234353 237086 239672
rect 237538 235833 237566 239672
rect 237526 235827 237578 235833
rect 237526 235769 237578 235775
rect 237046 234347 237098 234353
rect 237046 234289 237098 234295
rect 236758 233459 236810 233465
rect 236758 233401 236810 233407
rect 236086 231831 236138 231837
rect 236086 231773 236138 231779
rect 236002 227506 236126 227534
rect 235330 221468 235392 221496
rect 236098 221482 236126 227506
rect 236770 227323 236798 233401
rect 237634 232799 237662 239686
rect 238018 235463 238046 239686
rect 238006 235457 238058 235463
rect 238006 235399 238058 235405
rect 237622 232793 237674 232799
rect 237622 232735 237674 232741
rect 238402 229025 238430 239686
rect 238390 229019 238442 229025
rect 238390 228961 238442 228967
rect 238786 227471 238814 239686
rect 239136 239672 239390 239700
rect 239520 239672 239774 239700
rect 239362 235611 239390 239672
rect 239350 235605 239402 235611
rect 239350 235547 239402 235553
rect 238966 233385 239018 233391
rect 238966 233327 239018 233333
rect 238774 227465 238826 227471
rect 238774 227407 238826 227413
rect 236758 227317 236810 227323
rect 236758 227259 236810 227265
rect 238978 227175 239006 233327
rect 239062 229685 239114 229691
rect 239062 229627 239114 229633
rect 238390 227169 238442 227175
rect 238390 227111 238442 227117
rect 238966 227169 239018 227175
rect 238966 227111 239018 227117
rect 237526 227021 237578 227027
rect 237526 226963 237578 226969
rect 236854 226059 236906 226065
rect 236854 226001 236906 226007
rect 236866 221496 236894 226001
rect 236832 221468 236894 221496
rect 237538 221496 237566 226963
rect 237538 221468 237600 221496
rect 238402 221482 238430 227111
rect 239074 221792 239102 229627
rect 239746 228729 239774 239672
rect 239842 234501 239870 239686
rect 240226 234649 240254 239686
rect 240610 235241 240638 239686
rect 240502 235235 240554 235241
rect 240502 235177 240554 235183
rect 240598 235235 240650 235241
rect 240598 235177 240650 235183
rect 240214 234643 240266 234649
rect 240214 234585 240266 234591
rect 239830 234495 239882 234501
rect 239830 234437 239882 234443
rect 239734 228723 239786 228729
rect 239734 228665 239786 228671
rect 239830 227539 239882 227545
rect 239830 227481 239882 227487
rect 239074 221764 239150 221792
rect 239122 221482 239150 221764
rect 239842 221482 239870 227481
rect 240514 227027 240542 235177
rect 241090 230431 241118 239686
rect 241440 239672 241694 239700
rect 241078 230425 241130 230431
rect 241078 230367 241130 230373
rect 241666 228803 241694 239672
rect 241810 239404 241838 239686
rect 241810 239376 241886 239404
rect 241654 228797 241706 228803
rect 241654 228739 241706 228745
rect 240502 227021 240554 227027
rect 240502 226963 240554 226969
rect 240598 226207 240650 226213
rect 240598 226149 240650 226155
rect 240610 221482 240638 226149
rect 241858 226065 241886 239376
rect 242146 235389 242174 239686
rect 242134 235383 242186 235389
rect 242134 235325 242186 235331
rect 242134 232719 242186 232725
rect 242134 232661 242186 232667
rect 241846 226059 241898 226065
rect 241846 226001 241898 226007
rect 241270 225911 241322 225917
rect 241270 225853 241322 225859
rect 241282 221792 241310 225853
rect 241282 221764 241358 221792
rect 241330 221482 241358 221764
rect 242146 221482 242174 232661
rect 242530 228877 242558 239686
rect 242914 233317 242942 239686
rect 243298 235981 243326 239686
rect 243648 239672 243902 239700
rect 244032 239672 244286 239700
rect 243286 235975 243338 235981
rect 243286 235917 243338 235923
rect 243874 235019 243902 239672
rect 243958 236123 244010 236129
rect 243958 236065 244010 236071
rect 243862 235013 243914 235019
rect 243862 234955 243914 234961
rect 242902 233311 242954 233317
rect 242902 233253 242954 233259
rect 242518 228871 242570 228877
rect 242518 228813 242570 228819
rect 243574 227391 243626 227397
rect 243574 227333 243626 227339
rect 242902 227243 242954 227249
rect 242902 227185 242954 227191
rect 242914 221482 242942 227185
rect 243586 221792 243614 227333
rect 243970 226361 243998 236065
rect 244258 229765 244286 239672
rect 244354 234205 244382 239686
rect 244848 239672 245054 239700
rect 244726 235309 244778 235315
rect 244726 235251 244778 235257
rect 244342 234199 244394 234205
rect 244342 234141 244394 234147
rect 244246 229759 244298 229765
rect 244246 229701 244298 229707
rect 243958 226355 244010 226361
rect 243958 226297 244010 226303
rect 244342 225837 244394 225843
rect 244342 225779 244394 225785
rect 243586 221764 243662 221792
rect 243634 221482 243662 221764
rect 244354 221482 244382 225779
rect 244738 225621 244766 235251
rect 245026 226213 245054 239672
rect 245110 232645 245162 232651
rect 245110 232587 245162 232593
rect 245014 226207 245066 226213
rect 245014 226149 245066 226155
rect 244726 225615 244778 225621
rect 244726 225557 244778 225563
rect 245122 221482 245150 232587
rect 245218 231023 245246 239686
rect 245568 239672 245822 239700
rect 245952 239672 246206 239700
rect 246336 239672 246590 239700
rect 245206 231017 245258 231023
rect 245206 230959 245258 230965
rect 245794 230357 245822 239672
rect 245782 230351 245834 230357
rect 245782 230293 245834 230299
rect 246178 228951 246206 239672
rect 246166 228945 246218 228951
rect 246166 228887 246218 228893
rect 245878 227095 245930 227101
rect 245878 227037 245930 227043
rect 245890 221792 245918 227037
rect 246562 225991 246590 239672
rect 246658 235315 246686 239686
rect 246646 235309 246698 235315
rect 246646 235251 246698 235257
rect 247042 227915 247070 239686
rect 247426 234131 247454 239686
rect 247776 239672 248030 239700
rect 248160 239672 248414 239700
rect 248640 239672 248798 239700
rect 248002 236055 248030 239672
rect 247990 236049 248042 236055
rect 247990 235991 248042 235997
rect 247702 234717 247754 234723
rect 247702 234659 247754 234665
rect 247414 234125 247466 234131
rect 247414 234067 247466 234073
rect 247030 227909 247082 227915
rect 247030 227851 247082 227857
rect 247414 226281 247466 226287
rect 247414 226223 247466 226229
rect 246550 225985 246602 225991
rect 246550 225927 246602 225933
rect 246646 225763 246698 225769
rect 246646 225705 246698 225711
rect 245890 221764 245966 221792
rect 245938 221482 245966 221764
rect 246658 221482 246686 225705
rect 247426 221482 247454 226223
rect 247714 225769 247742 234659
rect 248086 232571 248138 232577
rect 248086 232513 248138 232519
rect 247702 225763 247754 225769
rect 247702 225705 247754 225711
rect 248098 221792 248126 232513
rect 248386 231541 248414 239672
rect 248374 231535 248426 231541
rect 248374 231477 248426 231483
rect 248770 230135 248798 239672
rect 248962 230283 248990 239686
rect 248950 230277 249002 230283
rect 248950 230219 249002 230225
rect 248758 230129 248810 230135
rect 248758 230071 248810 230077
rect 249346 227545 249374 239686
rect 249730 235537 249758 239686
rect 250080 239672 250334 239700
rect 249718 235531 249770 235537
rect 249718 235473 249770 235479
rect 250306 229913 250334 239672
rect 250450 239404 250478 239686
rect 250848 239672 251102 239700
rect 250450 239376 250526 239404
rect 250498 234427 250526 239376
rect 251074 236129 251102 239672
rect 251062 236123 251114 236129
rect 251062 236065 251114 236071
rect 251170 234723 251198 239686
rect 251158 234717 251210 234723
rect 251158 234659 251210 234665
rect 250582 234569 250634 234575
rect 250582 234511 250634 234517
rect 250486 234421 250538 234427
rect 250486 234363 250538 234369
rect 250294 229907 250346 229913
rect 250294 229849 250346 229855
rect 249718 229611 249770 229617
rect 249718 229553 249770 229559
rect 249334 227539 249386 227545
rect 249334 227481 249386 227487
rect 248854 227021 248906 227027
rect 248854 226963 248906 226969
rect 248098 221764 248174 221792
rect 248146 221482 248174 221764
rect 248866 221482 248894 226963
rect 249730 221482 249758 229553
rect 250594 228433 250622 234511
rect 251158 232497 251210 232503
rect 251158 232439 251210 232445
rect 250582 228427 250634 228433
rect 250582 228369 250634 228375
rect 250390 226947 250442 226953
rect 250390 226889 250442 226895
rect 250402 221792 250430 226889
rect 250402 221764 250478 221792
rect 250450 221482 250478 221764
rect 251170 221482 251198 232439
rect 251554 229839 251582 239686
rect 251938 229987 251966 239686
rect 252384 239672 252638 239700
rect 252768 239672 253022 239700
rect 252610 236174 252638 239672
rect 252610 236146 252734 236174
rect 251926 229981 251978 229987
rect 251926 229923 251978 229929
rect 251542 229833 251594 229839
rect 251542 229775 251594 229781
rect 252598 229537 252650 229543
rect 252598 229479 252650 229485
rect 252022 227465 252074 227471
rect 252022 227407 252074 227413
rect 252034 226361 252062 227407
rect 251926 226355 251978 226361
rect 251926 226297 251978 226303
rect 252022 226355 252074 226361
rect 252022 226297 252074 226303
rect 251938 221482 251966 226297
rect 252610 221792 252638 229479
rect 252706 225103 252734 236146
rect 252994 231097 253022 239672
rect 252982 231091 253034 231097
rect 252982 231033 253034 231039
rect 253090 229691 253118 239686
rect 253474 233909 253502 239686
rect 253558 234791 253610 234797
rect 253558 234733 253610 234739
rect 253462 233903 253514 233909
rect 253462 233845 253514 233851
rect 253078 229685 253130 229691
rect 253078 229627 253130 229633
rect 253570 227249 253598 234733
rect 253858 227471 253886 239686
rect 254242 234871 254270 239686
rect 254592 239672 254846 239700
rect 254976 239672 255230 239700
rect 254230 234865 254282 234871
rect 254230 234807 254282 234813
rect 254230 232423 254282 232429
rect 254230 232365 254282 232371
rect 253846 227465 253898 227471
rect 253846 227407 253898 227413
rect 253558 227243 253610 227249
rect 253558 227185 253610 227191
rect 253462 226873 253514 226879
rect 253462 226815 253514 226821
rect 252694 225097 252746 225103
rect 252694 225039 252746 225045
rect 252610 221764 252686 221792
rect 252658 221482 252686 221764
rect 253474 221482 253502 226815
rect 254242 221482 254270 232365
rect 254818 229543 254846 239672
rect 255202 229617 255230 239672
rect 255298 234575 255326 239686
rect 255286 234569 255338 234575
rect 255286 234511 255338 234517
rect 255670 232349 255722 232355
rect 255670 232291 255722 232297
rect 255190 229611 255242 229617
rect 255190 229553 255242 229559
rect 254806 229537 254858 229543
rect 254806 229479 254858 229485
rect 254902 225615 254954 225621
rect 254902 225557 254954 225563
rect 254914 221792 254942 225557
rect 254914 221764 254990 221792
rect 254962 221482 254990 221764
rect 255682 221482 255710 232291
rect 255778 231245 255806 239686
rect 256162 231615 256190 239686
rect 256546 234279 256574 239686
rect 256896 239672 257150 239700
rect 257280 239672 257534 239700
rect 256534 234273 256586 234279
rect 256534 234215 256586 234221
rect 256150 231609 256202 231615
rect 256150 231551 256202 231557
rect 255766 231239 255818 231245
rect 255766 231181 255818 231187
rect 257122 226805 257150 239672
rect 257506 234797 257534 239672
rect 257494 234791 257546 234797
rect 257494 234733 257546 234739
rect 257206 232275 257258 232281
rect 257206 232217 257258 232223
rect 256438 226799 256490 226805
rect 256438 226741 256490 226747
rect 257110 226799 257162 226805
rect 257110 226741 257162 226747
rect 256450 221482 256478 226741
rect 257218 221792 257246 232217
rect 257602 231689 257630 239686
rect 257986 233391 258014 239686
rect 258370 233983 258398 239686
rect 258454 234347 258506 234353
rect 258454 234289 258506 234295
rect 258358 233977 258410 233983
rect 258358 233919 258410 233925
rect 257974 233385 258026 233391
rect 257974 233327 258026 233333
rect 257590 231683 257642 231689
rect 257590 231625 257642 231631
rect 258466 228063 258494 234289
rect 258754 233243 258782 239686
rect 259104 239672 259166 239700
rect 259584 239672 259838 239700
rect 259030 235753 259082 235759
rect 259030 235695 259082 235701
rect 258742 233237 258794 233243
rect 258742 233179 258794 233185
rect 258742 228501 258794 228507
rect 258742 228443 258794 228449
rect 258454 228057 258506 228063
rect 258454 227999 258506 228005
rect 257974 225763 258026 225769
rect 257974 225705 258026 225711
rect 257218 221764 257294 221792
rect 257266 221482 257294 221764
rect 257986 221482 258014 225705
rect 258754 221482 258782 228443
rect 259042 225621 259070 235695
rect 259138 231763 259166 239672
rect 259810 234057 259838 239672
rect 259798 234051 259850 234057
rect 259798 233993 259850 233999
rect 259906 233539 259934 239686
rect 260290 234945 260318 239686
rect 260182 234939 260234 234945
rect 260182 234881 260234 234887
rect 260278 234939 260330 234945
rect 260278 234881 260330 234887
rect 259894 233533 259946 233539
rect 259894 233475 259946 233481
rect 259510 233311 259562 233317
rect 259510 233253 259562 233259
rect 259126 231757 259178 231763
rect 259126 231699 259178 231705
rect 259522 228359 259550 233253
rect 259510 228353 259562 228359
rect 259510 228295 259562 228301
rect 259414 226651 259466 226657
rect 259414 226593 259466 226599
rect 259030 225615 259082 225621
rect 259030 225557 259082 225563
rect 259426 221792 259454 226593
rect 259426 221764 259502 221792
rect 259474 221482 259502 221764
rect 260194 221482 260222 234881
rect 260470 234495 260522 234501
rect 260470 234437 260522 234443
rect 260482 228507 260510 234437
rect 260674 233095 260702 239686
rect 261024 239672 261278 239700
rect 261408 239672 261662 239700
rect 261792 239672 262046 239700
rect 261250 234353 261278 239672
rect 261238 234347 261290 234353
rect 261238 234289 261290 234295
rect 261634 233317 261662 239672
rect 262018 236174 262046 239672
rect 261922 236146 262046 236174
rect 261622 233311 261674 233317
rect 261622 233253 261674 233259
rect 260662 233089 260714 233095
rect 260662 233031 260714 233037
rect 261718 232201 261770 232207
rect 261718 232143 261770 232149
rect 260470 228501 260522 228507
rect 260470 228443 260522 228449
rect 261046 227317 261098 227323
rect 261046 227259 261098 227265
rect 261058 221482 261086 227259
rect 261730 221792 261758 232143
rect 261922 223845 261950 236146
rect 262006 235161 262058 235167
rect 262006 235103 262058 235109
rect 262018 225917 262046 235103
rect 262114 233169 262142 239686
rect 262498 234501 262526 239686
rect 262882 235759 262910 239686
rect 263328 239672 263582 239700
rect 263712 239672 263966 239700
rect 264096 239672 264350 239700
rect 262870 235753 262922 235759
rect 262870 235695 262922 235701
rect 262486 234495 262538 234501
rect 262486 234437 262538 234443
rect 262102 233163 262154 233169
rect 262102 233105 262154 233111
rect 263254 232127 263306 232133
rect 263254 232069 263306 232075
rect 262486 226725 262538 226731
rect 262486 226667 262538 226673
rect 262006 225911 262058 225917
rect 262006 225853 262058 225859
rect 261910 223839 261962 223845
rect 261910 223781 261962 223787
rect 261730 221764 261806 221792
rect 261778 221482 261806 221764
rect 262498 221482 262526 226667
rect 263266 221482 263294 232069
rect 263554 223771 263582 239672
rect 263638 234199 263690 234205
rect 263638 234141 263690 234147
rect 263650 227841 263678 234141
rect 263938 232873 263966 239672
rect 263926 232867 263978 232873
rect 263926 232809 263978 232815
rect 264322 229469 264350 239672
rect 264418 233465 264446 239686
rect 264610 239672 264816 239700
rect 264406 233459 264458 233465
rect 264406 233401 264458 233407
rect 264310 229463 264362 229469
rect 264310 229405 264362 229411
rect 263638 227835 263690 227841
rect 263638 227777 263690 227783
rect 264022 227169 264074 227175
rect 264022 227111 264074 227117
rect 263542 223765 263594 223771
rect 263542 223707 263594 223713
rect 264034 221496 264062 227111
rect 264610 223623 264638 239672
rect 264886 235901 264938 235907
rect 264886 235843 264938 235849
rect 264694 234643 264746 234649
rect 264694 234585 264746 234591
rect 264706 227175 264734 234585
rect 264790 230055 264842 230061
rect 264790 229997 264842 230003
rect 264694 227169 264746 227175
rect 264694 227111 264746 227117
rect 264598 223617 264650 223623
rect 264598 223559 264650 223565
rect 264034 221468 264096 221496
rect 264802 221482 264830 229997
rect 264898 226065 264926 235843
rect 265186 232725 265214 239686
rect 265536 239672 265790 239700
rect 265920 239672 266174 239700
rect 266304 239672 266558 239700
rect 265762 233021 265790 239672
rect 266146 235167 266174 239672
rect 266134 235161 266186 235167
rect 266134 235103 266186 235109
rect 266422 235087 266474 235093
rect 266422 235029 266474 235035
rect 266326 234125 266378 234131
rect 266326 234067 266378 234073
rect 265750 233015 265802 233021
rect 265750 232957 265802 232963
rect 265174 232719 265226 232725
rect 265174 232661 265226 232667
rect 266338 228581 266366 234067
rect 266230 228575 266282 228581
rect 266230 228517 266282 228523
rect 266326 228575 266378 228581
rect 266326 228517 266378 228523
rect 265558 226577 265610 226583
rect 265558 226519 265610 226525
rect 264886 226059 264938 226065
rect 264886 226001 264938 226007
rect 265570 221496 265598 226519
rect 265536 221468 265598 221496
rect 266242 221496 266270 228517
rect 266434 225769 266462 235029
rect 266422 225763 266474 225769
rect 266422 225705 266474 225711
rect 266530 223697 266558 239672
rect 266626 232577 266654 239686
rect 267106 234131 267134 239686
rect 267490 234649 267518 239686
rect 267840 239672 268094 239700
rect 268224 239672 268478 239700
rect 267478 234643 267530 234649
rect 267478 234585 267530 234591
rect 267958 234421 268010 234427
rect 267958 234363 268010 234369
rect 267094 234125 267146 234131
rect 267094 234067 267146 234073
rect 267766 233533 267818 233539
rect 267766 233475 267818 233481
rect 266614 232571 266666 232577
rect 266614 232513 266666 232519
rect 266998 227243 267050 227249
rect 266998 227185 267050 227191
rect 266518 223691 266570 223697
rect 266518 223633 266570 223639
rect 266242 221468 266304 221496
rect 267010 221482 267038 227185
rect 267778 225991 267806 233475
rect 267862 230203 267914 230209
rect 267862 230145 267914 230151
rect 267766 225985 267818 225991
rect 267766 225927 267818 225933
rect 267874 221755 267902 230145
rect 267970 228211 267998 234363
rect 267958 228205 268010 228211
rect 267958 228147 268010 228153
rect 268066 223549 268094 239672
rect 268150 235827 268202 235833
rect 268150 235769 268202 235775
rect 268162 226657 268190 235769
rect 268450 232651 268478 239672
rect 268546 234205 268574 239686
rect 268930 235093 268958 239686
rect 269314 236174 269342 239686
rect 269314 236146 269438 236174
rect 268918 235087 268970 235093
rect 268918 235029 268970 235035
rect 268534 234199 268586 234205
rect 268534 234141 268586 234147
rect 268438 232645 268490 232651
rect 268438 232587 268490 232593
rect 269302 229315 269354 229321
rect 269302 229257 269354 229263
rect 268150 226651 268202 226657
rect 268150 226593 268202 226599
rect 268534 226503 268586 226509
rect 268534 226445 268586 226451
rect 268054 223543 268106 223549
rect 268054 223485 268106 223491
rect 267826 221727 267902 221755
rect 267826 221482 267854 221727
rect 268546 221482 268574 226445
rect 269314 221482 269342 229257
rect 269410 223401 269438 236146
rect 269590 233311 269642 233317
rect 269590 233253 269642 233259
rect 269602 225843 269630 233253
rect 269698 232429 269726 239686
rect 270048 239672 270302 239700
rect 270432 239672 270590 239700
rect 269878 233385 269930 233391
rect 269878 233327 269930 233333
rect 269686 232423 269738 232429
rect 269686 232365 269738 232371
rect 269890 230209 269918 233327
rect 270274 233317 270302 239672
rect 270562 233391 270590 239672
rect 270850 236174 270878 239686
rect 270850 236146 270974 236174
rect 270838 233903 270890 233909
rect 270838 233845 270890 233851
rect 270550 233385 270602 233391
rect 270550 233327 270602 233333
rect 270262 233311 270314 233317
rect 270262 233253 270314 233259
rect 269878 230203 269930 230209
rect 269878 230145 269930 230151
rect 270742 229389 270794 229395
rect 270742 229331 270794 229337
rect 269590 225837 269642 225843
rect 269590 225779 269642 225785
rect 269974 225615 270026 225621
rect 269974 225557 270026 225563
rect 269398 223395 269450 223401
rect 269398 223337 269450 223343
rect 269986 221792 270014 225557
rect 269986 221764 270062 221792
rect 270034 221482 270062 221764
rect 270754 221482 270782 229331
rect 270850 228285 270878 233845
rect 270838 228279 270890 228285
rect 270838 228221 270890 228227
rect 270946 223475 270974 236146
rect 271030 235975 271082 235981
rect 271030 235917 271082 235923
rect 271042 226583 271070 235917
rect 271234 232503 271262 239686
rect 271618 234427 271646 239686
rect 271606 234421 271658 234427
rect 271606 234363 271658 234369
rect 271222 232497 271274 232503
rect 271222 232439 271274 232445
rect 272002 227249 272030 239686
rect 272352 239672 272606 239700
rect 272736 239672 272990 239700
rect 272374 233459 272426 233465
rect 272374 233401 272426 233407
rect 272278 228649 272330 228655
rect 272278 228591 272330 228597
rect 271990 227243 272042 227249
rect 271990 227185 272042 227191
rect 271030 226577 271082 226583
rect 271030 226519 271082 226525
rect 271606 226429 271658 226435
rect 271606 226371 271658 226377
rect 270934 223469 270986 223475
rect 270934 223411 270986 223417
rect 271618 221482 271646 226371
rect 272290 221792 272318 228591
rect 272386 225029 272414 233401
rect 272374 225023 272426 225029
rect 272374 224965 272426 224971
rect 272578 222439 272606 239672
rect 272962 232281 272990 239672
rect 273058 235907 273086 239686
rect 273046 235901 273098 235907
rect 273046 235843 273098 235849
rect 273334 233311 273386 233317
rect 273334 233253 273386 233259
rect 272950 232275 273002 232281
rect 272950 232217 273002 232223
rect 273346 229395 273374 233253
rect 273334 229389 273386 229395
rect 273334 229331 273386 229337
rect 273442 226953 273470 239686
rect 273840 239672 274142 239700
rect 273718 236123 273770 236129
rect 273718 236065 273770 236071
rect 273622 236049 273674 236055
rect 273622 235991 273674 235997
rect 273430 226947 273482 226953
rect 273430 226889 273482 226895
rect 273238 226799 273290 226805
rect 273238 226741 273290 226747
rect 273250 225991 273278 226741
rect 273238 225985 273290 225991
rect 273238 225927 273290 225933
rect 273046 225911 273098 225917
rect 273046 225853 273098 225859
rect 272566 222433 272618 222439
rect 272566 222375 272618 222381
rect 272290 221764 272366 221792
rect 272338 221482 272366 221764
rect 273058 221482 273086 225853
rect 273634 225547 273662 235991
rect 273730 225621 273758 236065
rect 273814 229167 273866 229173
rect 273814 229109 273866 229115
rect 273718 225615 273770 225621
rect 273718 225557 273770 225563
rect 273622 225541 273674 225547
rect 273622 225483 273674 225489
rect 273826 221482 273854 229109
rect 274114 222217 274142 239672
rect 274210 232207 274238 239686
rect 274656 239672 274910 239700
rect 275040 239672 275294 239700
rect 274678 233385 274730 233391
rect 274678 233327 274730 233333
rect 274198 232201 274250 232207
rect 274198 232143 274250 232149
rect 274486 232053 274538 232059
rect 274486 231995 274538 232001
rect 274102 222211 274154 222217
rect 274102 222153 274154 222159
rect 274498 221792 274526 231995
rect 274690 227323 274718 233327
rect 274882 232355 274910 239672
rect 274870 232349 274922 232355
rect 274870 232291 274922 232297
rect 274678 227317 274730 227323
rect 274678 227259 274730 227265
rect 275266 227027 275294 239672
rect 275362 237683 275390 239686
rect 275350 237677 275402 237683
rect 275350 237619 275402 237625
rect 275746 232133 275774 239686
rect 276130 235833 276158 239686
rect 276480 239672 276734 239700
rect 276864 239672 277118 239700
rect 277248 239672 277502 239700
rect 276118 235827 276170 235833
rect 276118 235769 276170 235775
rect 275734 232127 275786 232133
rect 275734 232069 275786 232075
rect 275350 231979 275402 231985
rect 275350 231921 275402 231927
rect 275254 227021 275306 227027
rect 275254 226963 275306 226969
rect 274498 221764 274574 221792
rect 274546 221482 274574 221764
rect 275362 221482 275390 231921
rect 276502 228427 276554 228433
rect 276502 228369 276554 228375
rect 276118 226059 276170 226065
rect 276118 226001 276170 226007
rect 276130 221482 276158 226001
rect 276406 221767 276458 221773
rect 276514 221755 276542 228369
rect 276706 227101 276734 239672
rect 277090 237609 277118 239672
rect 277078 237603 277130 237609
rect 277078 237545 277130 237551
rect 277078 233977 277130 233983
rect 277078 233919 277130 233925
rect 276790 229241 276842 229247
rect 276790 229183 276842 229189
rect 276694 227095 276746 227101
rect 276694 227037 276746 227043
rect 276802 221792 276830 229183
rect 277090 225251 277118 233919
rect 277474 232059 277502 239672
rect 277570 236129 277598 239686
rect 277558 236123 277610 236129
rect 277558 236065 277610 236071
rect 277462 232053 277514 232059
rect 277462 231995 277514 232001
rect 277078 225245 277130 225251
rect 277078 225187 277130 225193
rect 277954 224733 277982 239686
rect 278434 236869 278462 239686
rect 278784 239672 279038 239700
rect 279168 239672 279326 239700
rect 279552 239672 279806 239700
rect 278422 236863 278474 236869
rect 278422 236805 278474 236811
rect 278230 234569 278282 234575
rect 278230 234511 278282 234517
rect 278134 234273 278186 234279
rect 278134 234215 278186 234221
rect 278146 227619 278174 234215
rect 278134 227613 278186 227619
rect 278134 227555 278186 227561
rect 278242 225695 278270 234511
rect 279010 231911 279038 239672
rect 279298 235981 279326 239672
rect 279286 235975 279338 235981
rect 279286 235917 279338 235923
rect 278326 231905 278378 231911
rect 278326 231847 278378 231853
rect 278998 231905 279050 231911
rect 278998 231847 279050 231853
rect 278230 225689 278282 225695
rect 278230 225631 278282 225637
rect 277942 224727 277994 224733
rect 277942 224669 277994 224675
rect 276802 221764 276878 221792
rect 276458 221727 276542 221755
rect 276406 221709 276458 221715
rect 276850 221482 276878 221764
rect 277558 221767 277610 221773
rect 277558 221709 277610 221715
rect 277570 221482 277598 221709
rect 278338 221482 278366 231847
rect 279778 226805 279806 239672
rect 279874 236943 279902 239686
rect 279862 236937 279914 236943
rect 279862 236879 279914 236885
rect 280258 231985 280286 239686
rect 280642 236055 280670 239686
rect 280992 239672 281246 239700
rect 281376 239672 281630 239700
rect 281760 239672 282014 239700
rect 280630 236049 280682 236055
rect 280630 235991 280682 235997
rect 280246 231979 280298 231985
rect 280246 231921 280298 231927
rect 281218 231467 281246 239672
rect 281302 231831 281354 231837
rect 281302 231773 281354 231779
rect 281206 231461 281258 231467
rect 281206 231403 281258 231409
rect 279862 229093 279914 229099
rect 279862 229035 279914 229041
rect 279766 226799 279818 226805
rect 279766 226741 279818 226747
rect 279094 225763 279146 225769
rect 279094 225705 279146 225711
rect 279106 221792 279134 225705
rect 279106 221764 279182 221792
rect 279154 221482 279182 221764
rect 279874 221482 279902 229035
rect 280630 228057 280682 228063
rect 280630 227999 280682 228005
rect 280642 221482 280670 227999
rect 281314 221792 281342 231773
rect 281602 222291 281630 239672
rect 281986 231837 282014 239672
rect 282070 234051 282122 234057
rect 282070 233993 282122 233999
rect 281974 231831 282026 231837
rect 281974 231773 282026 231779
rect 282082 227693 282110 233993
rect 282178 229247 282206 239686
rect 282562 233391 282590 239686
rect 282960 239672 283166 239700
rect 283296 239672 283550 239700
rect 283680 239672 283934 239700
rect 282934 235679 282986 235685
rect 282934 235621 282986 235627
rect 282550 233385 282602 233391
rect 282550 233327 282602 233333
rect 282166 229241 282218 229247
rect 282166 229183 282218 229189
rect 282070 227687 282122 227693
rect 282070 227629 282122 227635
rect 282070 226651 282122 226657
rect 282070 226593 282122 226599
rect 281590 222285 281642 222291
rect 281590 222227 281642 222233
rect 281314 221764 281390 221792
rect 281362 221482 281390 221764
rect 282082 221482 282110 226593
rect 282946 221482 282974 235621
rect 283138 222365 283166 239672
rect 283522 229321 283550 239672
rect 283906 234575 283934 239672
rect 283894 234569 283946 234575
rect 283894 234511 283946 234517
rect 284002 233613 284030 239686
rect 284400 239672 284702 239700
rect 283990 233607 284042 233613
rect 283990 233549 284042 233555
rect 284374 232793 284426 232799
rect 284374 232735 284426 232741
rect 283510 229315 283562 229321
rect 283510 229257 283562 229263
rect 283606 229019 283658 229025
rect 283606 228961 283658 228967
rect 283126 222359 283178 222365
rect 283126 222301 283178 222307
rect 283618 221792 283646 228961
rect 283618 221764 283694 221792
rect 283666 221482 283694 221764
rect 284386 221482 284414 232735
rect 284674 226731 284702 239672
rect 284770 229173 284798 239686
rect 285154 235685 285182 239686
rect 285504 239672 285758 239700
rect 285984 239672 286238 239700
rect 285142 235679 285194 235685
rect 285142 235621 285194 235627
rect 285334 235605 285386 235611
rect 285334 235547 285386 235553
rect 285046 234643 285098 234649
rect 285046 234585 285098 234591
rect 284758 229167 284810 229173
rect 284758 229109 284810 229115
rect 284662 226725 284714 226731
rect 284662 226667 284714 226673
rect 285058 225769 285086 234585
rect 285346 233317 285374 235547
rect 285334 233311 285386 233317
rect 285334 233253 285386 233259
rect 285730 226657 285758 239672
rect 285910 235457 285962 235463
rect 285910 235399 285962 235405
rect 285718 226651 285770 226657
rect 285718 226593 285770 226599
rect 285142 226355 285194 226361
rect 285142 226297 285194 226303
rect 285046 225763 285098 225769
rect 285046 225705 285098 225711
rect 285154 221482 285182 226297
rect 285922 221792 285950 235399
rect 286210 222513 286238 239672
rect 286306 229099 286334 239686
rect 286690 235611 286718 239686
rect 286678 235605 286730 235611
rect 286678 235547 286730 235553
rect 287074 234649 287102 239686
rect 287062 234643 287114 234649
rect 287062 234585 287114 234591
rect 287458 233539 287486 239686
rect 287808 239672 287966 239700
rect 288192 239672 288446 239700
rect 287446 233533 287498 233539
rect 287446 233475 287498 233481
rect 287446 233311 287498 233317
rect 287446 233253 287498 233259
rect 286294 229093 286346 229099
rect 286294 229035 286346 229041
rect 286678 228501 286730 228507
rect 286678 228443 286730 228449
rect 286198 222507 286250 222513
rect 286198 222449 286250 222455
rect 285922 221764 285998 221792
rect 285970 221482 285998 221764
rect 286690 221482 286718 228443
rect 287458 221482 287486 233253
rect 287938 229025 287966 239672
rect 288022 234347 288074 234353
rect 288022 234289 288074 234295
rect 287926 229019 287978 229025
rect 287926 228961 287978 228967
rect 288034 228433 288062 234289
rect 288418 233465 288446 239672
rect 288406 233459 288458 233465
rect 288406 233401 288458 233407
rect 288022 228427 288074 228433
rect 288022 228369 288074 228375
rect 288118 227169 288170 227175
rect 288118 227111 288170 227117
rect 288130 221792 288158 227111
rect 288514 226509 288542 239686
rect 288898 233317 288926 239686
rect 288886 233311 288938 233317
rect 288886 233253 288938 233259
rect 288886 228723 288938 228729
rect 288886 228665 288938 228671
rect 288502 226503 288554 226509
rect 288502 226445 288554 226451
rect 288130 221764 288206 221792
rect 288178 221482 288206 221764
rect 288898 221482 288926 228665
rect 289378 228507 289406 239686
rect 289728 239672 289982 239700
rect 290112 239672 290366 239700
rect 290496 239672 290654 239700
rect 289954 232947 289982 239672
rect 290338 234279 290366 239672
rect 290422 235235 290474 235241
rect 290422 235177 290474 235183
rect 290326 234273 290378 234279
rect 290326 234215 290378 234221
rect 289942 232941 289994 232947
rect 289942 232883 289994 232889
rect 289654 231461 289706 231467
rect 289654 231403 289706 231409
rect 289366 228501 289418 228507
rect 289366 228443 289418 228449
rect 289666 227175 289694 231403
rect 289750 228797 289802 228803
rect 289750 228739 289802 228745
rect 289654 227169 289706 227175
rect 289654 227111 289706 227117
rect 289762 221482 289790 228739
rect 290434 221792 290462 235177
rect 290626 230653 290654 239672
rect 290818 231393 290846 239686
rect 290902 234495 290954 234501
rect 290902 234437 290954 234443
rect 290806 231387 290858 231393
rect 290806 231329 290858 231335
rect 290614 230647 290666 230653
rect 290614 230589 290666 230595
rect 290914 230061 290942 234437
rect 290998 234125 291050 234131
rect 290998 234067 291050 234073
rect 290902 230055 290954 230061
rect 290902 229997 290954 230003
rect 291010 227989 291038 234067
rect 291202 228655 291230 239686
rect 291190 228649 291242 228655
rect 291190 228591 291242 228597
rect 290998 227983 291050 227989
rect 290998 227925 291050 227931
rect 291586 226361 291614 239686
rect 291936 239672 292190 239700
rect 292320 239672 292574 239700
rect 292704 239672 292958 239700
rect 291958 230425 292010 230431
rect 291958 230367 292010 230373
rect 291574 226355 291626 226361
rect 291574 226297 291626 226303
rect 291190 226207 291242 226213
rect 291190 226149 291242 226155
rect 290434 221764 290510 221792
rect 290482 221482 290510 221764
rect 291202 221482 291230 226149
rect 291970 221482 291998 230367
rect 292162 228919 292190 239672
rect 292546 231467 292574 239672
rect 292930 234353 292958 239672
rect 292918 234347 292970 234353
rect 292918 234289 292970 234295
rect 292534 231461 292586 231467
rect 292534 231403 292586 231409
rect 293122 231319 293150 239686
rect 293398 235383 293450 235389
rect 293398 235325 293450 235331
rect 293110 231313 293162 231319
rect 293110 231255 293162 231261
rect 292148 228910 292204 228919
rect 292148 228845 292204 228854
rect 292630 228353 292682 228359
rect 292630 228295 292682 228301
rect 292642 221792 292670 228295
rect 293410 228156 293438 235325
rect 293506 231171 293534 239686
rect 293782 234199 293834 234205
rect 293782 234141 293834 234147
rect 293494 231165 293546 231171
rect 293494 231107 293546 231113
rect 293410 228128 293534 228156
rect 293794 228137 293822 234141
rect 293890 228359 293918 239686
rect 294240 239672 294494 239700
rect 294624 239672 294878 239700
rect 295008 239672 295262 239700
rect 294466 234131 294494 239672
rect 294454 234125 294506 234131
rect 294454 234067 294506 234073
rect 294850 233983 294878 239672
rect 295234 235463 295262 239672
rect 295222 235457 295274 235463
rect 295222 235399 295274 235405
rect 294838 233977 294890 233983
rect 294838 233919 294890 233925
rect 295330 232799 295358 239686
rect 295714 234205 295742 239686
rect 295702 234199 295754 234205
rect 295702 234141 295754 234147
rect 296098 233909 296126 239686
rect 296448 239672 296606 239700
rect 296928 239672 297182 239700
rect 296578 235019 296606 239672
rect 296470 235013 296522 235019
rect 296470 234955 296522 234961
rect 296566 235013 296618 235019
rect 296566 234955 296618 234961
rect 296086 233903 296138 233909
rect 296086 233845 296138 233851
rect 295318 232793 295370 232799
rect 295318 232735 295370 232741
rect 294934 228871 294986 228877
rect 294934 228813 294986 228819
rect 293878 228353 293930 228359
rect 293878 228295 293930 228301
rect 292642 221764 292718 221792
rect 292690 221482 292718 221764
rect 293506 221482 293534 228128
rect 293782 228131 293834 228137
rect 293782 228073 293834 228079
rect 294262 226577 294314 226583
rect 294262 226519 294314 226525
rect 294274 221496 294302 226519
rect 294240 221468 294302 221496
rect 294946 221496 294974 228813
rect 295702 227835 295754 227841
rect 295702 227777 295754 227783
rect 294946 221468 295008 221496
rect 295714 221482 295742 227777
rect 296482 221496 296510 234955
rect 297154 234501 297182 239672
rect 297142 234495 297194 234501
rect 297142 234437 297194 234443
rect 297250 233761 297278 239686
rect 297238 233755 297290 233761
rect 297238 233697 297290 233703
rect 297334 230647 297386 230653
rect 297334 230589 297386 230595
rect 297346 226583 297374 230589
rect 297334 226577 297386 226583
rect 297334 226519 297386 226525
rect 297634 226287 297662 239686
rect 298018 236174 298046 239686
rect 298416 239672 298622 239700
rect 298752 239672 299006 239700
rect 299136 239672 299390 239700
rect 298018 236146 298142 236174
rect 298006 229759 298058 229765
rect 298006 229701 298058 229707
rect 297238 226281 297290 226287
rect 297238 226223 297290 226229
rect 297622 226281 297674 226287
rect 297622 226223 297674 226229
rect 296448 221468 296510 221496
rect 297250 221482 297278 226223
rect 298018 221482 298046 229701
rect 298114 228063 298142 236146
rect 298594 229765 298622 239672
rect 298978 231879 299006 239672
rect 299254 235309 299306 235315
rect 299254 235251 299306 235257
rect 299158 233385 299210 233391
rect 299158 233327 299210 233333
rect 298964 231870 299020 231879
rect 298964 231805 299020 231814
rect 298582 229759 298634 229765
rect 298582 229701 298634 229707
rect 298678 228945 298730 228951
rect 298678 228887 298730 228893
rect 298102 228057 298154 228063
rect 298102 227999 298154 228005
rect 298210 226805 298430 226824
rect 298198 226799 298442 226805
rect 298250 226796 298390 226799
rect 298198 226741 298250 226747
rect 298390 226741 298442 226747
rect 298102 226725 298154 226731
rect 298102 226667 298154 226673
rect 298114 226435 298142 226667
rect 298102 226429 298154 226435
rect 298102 226371 298154 226377
rect 298690 221792 298718 228887
rect 299170 226731 299198 233327
rect 299266 230505 299294 235251
rect 299362 234691 299390 239672
rect 299458 234987 299486 239686
rect 299842 235389 299870 239686
rect 300226 237017 300254 239686
rect 300214 237011 300266 237017
rect 300214 236953 300266 236959
rect 299830 235383 299882 235389
rect 299830 235325 299882 235331
rect 299444 234978 299500 234987
rect 299444 234913 299500 234922
rect 299348 234682 299404 234691
rect 299348 234617 299404 234626
rect 299446 231017 299498 231023
rect 299446 230959 299498 230965
rect 299254 230499 299306 230505
rect 299254 230441 299306 230447
rect 299158 226725 299210 226731
rect 299158 226667 299210 226673
rect 298690 221764 298766 221792
rect 298738 221482 298766 221764
rect 299458 221482 299486 230959
rect 300706 226213 300734 239686
rect 301056 239672 301310 239700
rect 301440 239672 301694 239700
rect 300982 230351 301034 230357
rect 300982 230293 301034 230299
rect 300694 226207 300746 226213
rect 300694 226149 300746 226155
rect 300214 226133 300266 226139
rect 300214 226075 300266 226081
rect 300226 221482 300254 226075
rect 300994 221792 301022 230293
rect 301282 226139 301310 239672
rect 301666 234839 301694 239672
rect 301762 235315 301790 239686
rect 301750 235309 301802 235315
rect 301750 235251 301802 235257
rect 301652 234830 301708 234839
rect 301652 234765 301708 234774
rect 301750 228575 301802 228581
rect 301750 228517 301802 228523
rect 301270 226133 301322 226139
rect 301270 226075 301322 226081
rect 300994 221764 301070 221792
rect 301042 221482 301070 221764
rect 301762 221482 301790 228517
rect 302146 225325 302174 239686
rect 302544 239672 302846 239700
rect 302326 235531 302378 235537
rect 302326 235473 302378 235479
rect 302230 234421 302282 234427
rect 302230 234363 302282 234369
rect 302242 227841 302270 234363
rect 302338 230653 302366 235473
rect 302326 230647 302378 230653
rect 302326 230589 302378 230595
rect 302518 230499 302570 230505
rect 302518 230441 302570 230447
rect 302230 227835 302282 227841
rect 302230 227777 302282 227783
rect 302134 225319 302186 225325
rect 302134 225261 302186 225267
rect 302530 221482 302558 230441
rect 302818 222661 302846 239672
rect 302914 233687 302942 239686
rect 303264 239672 303518 239700
rect 303648 239672 303902 239700
rect 303984 239672 304286 239700
rect 302902 233681 302954 233687
rect 302902 233623 302954 233629
rect 303490 228581 303518 239672
rect 303478 228575 303530 228581
rect 303478 228517 303530 228523
rect 303190 225541 303242 225547
rect 303190 225483 303242 225489
rect 302806 222655 302858 222661
rect 302806 222597 302858 222603
rect 303202 221792 303230 225483
rect 303874 225399 303902 239672
rect 304150 234717 304202 234723
rect 304150 234659 304202 234665
rect 304162 230505 304190 234659
rect 304150 230499 304202 230505
rect 304150 230441 304202 230447
rect 303958 227909 304010 227915
rect 303958 227851 304010 227857
rect 303862 225393 303914 225399
rect 303862 225335 303914 225341
rect 303202 221764 303278 221792
rect 303250 221482 303278 221764
rect 303970 221482 303998 227851
rect 304258 222735 304286 239672
rect 304450 228803 304478 239686
rect 304834 236174 304862 239686
rect 305184 239672 305246 239700
rect 305568 239672 305822 239700
rect 305952 239672 306206 239700
rect 304834 236146 304958 236174
rect 304822 230277 304874 230283
rect 304822 230219 304874 230225
rect 304438 228797 304490 228803
rect 304438 228739 304490 228745
rect 304246 222729 304298 222735
rect 304246 222671 304298 222677
rect 304834 221482 304862 230219
rect 304930 222587 304958 236146
rect 305014 235901 305066 235907
rect 305014 235843 305066 235849
rect 305026 230283 305054 235843
rect 305110 235753 305162 235759
rect 305110 235695 305162 235701
rect 305014 230277 305066 230283
rect 305014 230219 305066 230225
rect 305122 225177 305150 235695
rect 305218 234057 305246 239672
rect 305794 237091 305822 239672
rect 305782 237085 305834 237091
rect 305782 237027 305834 237033
rect 305206 234051 305258 234057
rect 305206 233993 305258 233999
rect 305494 231535 305546 231541
rect 305494 231477 305546 231483
rect 305110 225171 305162 225177
rect 305110 225113 305162 225119
rect 304918 222581 304970 222587
rect 304918 222523 304970 222529
rect 305506 221792 305534 231477
rect 306178 228729 306206 239672
rect 306274 233835 306302 239686
rect 306658 236174 306686 239686
rect 307056 239672 307262 239700
rect 307392 239672 307646 239700
rect 307776 239672 308030 239700
rect 308256 239672 308510 239700
rect 306658 236146 306782 236174
rect 306646 234865 306698 234871
rect 306646 234807 306698 234813
rect 306262 233829 306314 233835
rect 306262 233771 306314 233777
rect 306658 230579 306686 234807
rect 306646 230573 306698 230579
rect 306646 230515 306698 230521
rect 306166 228723 306218 228729
rect 306166 228665 306218 228671
rect 306262 227539 306314 227545
rect 306262 227481 306314 227487
rect 305506 221764 305582 221792
rect 305554 221482 305582 221764
rect 306274 221482 306302 227481
rect 306754 225473 306782 236146
rect 307030 230129 307082 230135
rect 307030 230071 307082 230077
rect 306742 225467 306794 225473
rect 306742 225409 306794 225415
rect 307042 221482 307070 230071
rect 307234 222809 307262 239672
rect 307618 231139 307646 239672
rect 307604 231130 307660 231139
rect 307604 231065 307660 231074
rect 307702 228205 307754 228211
rect 307702 228147 307754 228153
rect 307222 222803 307274 222809
rect 307222 222745 307274 222751
rect 307714 221792 307742 228147
rect 308002 222957 308030 239672
rect 308278 235827 308330 235833
rect 308278 235769 308330 235775
rect 308182 234791 308234 234797
rect 308182 234733 308234 234739
rect 308194 231023 308222 234733
rect 308182 231017 308234 231023
rect 308182 230959 308234 230965
rect 308290 227915 308318 235769
rect 308482 234723 308510 239672
rect 308578 237239 308606 239686
rect 308566 237233 308618 237239
rect 308566 237175 308618 237181
rect 308470 234717 308522 234723
rect 308470 234659 308522 234665
rect 308566 230647 308618 230653
rect 308566 230589 308618 230595
rect 308278 227909 308330 227915
rect 308278 227851 308330 227857
rect 307990 222951 308042 222957
rect 307990 222893 308042 222899
rect 307714 221764 307790 221792
rect 307762 221482 307790 221764
rect 308578 221482 308606 230589
rect 308962 228951 308990 239686
rect 309346 235537 309374 239686
rect 309696 239672 309950 239700
rect 310080 239672 310334 239700
rect 310464 239672 310718 239700
rect 309334 235531 309386 235537
rect 309334 235473 309386 235479
rect 308950 228945 309002 228951
rect 308950 228887 309002 228893
rect 309334 225615 309386 225621
rect 309334 225557 309386 225563
rect 309346 221482 309374 225557
rect 309922 225547 309950 239672
rect 310006 229907 310058 229913
rect 310006 229849 310058 229855
rect 309910 225541 309962 225547
rect 309910 225483 309962 225489
rect 310018 221792 310046 229849
rect 310306 223031 310334 239672
rect 310690 228877 310718 239672
rect 310786 237165 310814 239686
rect 310774 237159 310826 237165
rect 310774 237101 310826 237107
rect 311062 233459 311114 233465
rect 311062 233401 311114 233407
rect 310774 229981 310826 229987
rect 310774 229923 310826 229929
rect 310678 228871 310730 228877
rect 310678 228813 310730 228819
rect 310294 223025 310346 223031
rect 310294 222967 310346 222973
rect 310018 221764 310094 221792
rect 310066 221482 310094 221764
rect 310786 221482 310814 229923
rect 311074 228211 311102 233401
rect 311170 233391 311198 239686
rect 311554 237313 311582 239686
rect 312000 239672 312254 239700
rect 312384 239672 312638 239700
rect 311542 237307 311594 237313
rect 311542 237249 311594 237255
rect 311254 233607 311306 233613
rect 311254 233549 311306 233555
rect 311158 233385 311210 233391
rect 311158 233327 311210 233333
rect 311062 228205 311114 228211
rect 311062 228147 311114 228153
rect 311266 227545 311294 233549
rect 311350 233533 311402 233539
rect 311350 233475 311402 233481
rect 311254 227539 311306 227545
rect 311254 227481 311306 227487
rect 311362 227397 311390 233475
rect 312226 231541 312254 239672
rect 312214 231535 312266 231541
rect 312214 231477 312266 231483
rect 311638 230499 311690 230505
rect 311638 230441 311690 230447
rect 311350 227391 311402 227397
rect 311350 227333 311402 227339
rect 311650 221482 311678 230441
rect 312310 225097 312362 225103
rect 312310 225039 312362 225045
rect 312322 221792 312350 225039
rect 312610 222883 312638 239672
rect 312706 234353 312734 239686
rect 313104 239672 313406 239700
rect 312694 234347 312746 234353
rect 312694 234289 312746 234295
rect 313078 229833 313130 229839
rect 313078 229775 313130 229781
rect 312598 222877 312650 222883
rect 312598 222819 312650 222825
rect 312322 221764 312398 221792
rect 312370 221482 312398 221764
rect 313090 221482 313118 229775
rect 313378 223105 313406 239672
rect 313474 228179 313502 239686
rect 313858 235759 313886 239686
rect 314208 239672 314462 239700
rect 314592 239672 314846 239700
rect 313942 236123 313994 236129
rect 313942 236065 313994 236071
rect 313846 235753 313898 235759
rect 313846 235695 313898 235701
rect 313846 234421 313898 234427
rect 313846 234363 313898 234369
rect 313858 228452 313886 234363
rect 313954 230653 313982 236065
rect 314434 234427 314462 239672
rect 314818 237387 314846 239672
rect 314806 237381 314858 237387
rect 314806 237323 314858 237329
rect 314422 234421 314474 234427
rect 314422 234363 314474 234369
rect 314518 231091 314570 231097
rect 314518 231033 314570 231039
rect 313942 230647 313994 230653
rect 313942 230589 313994 230595
rect 313858 228424 313982 228452
rect 313954 228285 313982 228424
rect 313846 228279 313898 228285
rect 313846 228221 313898 228227
rect 313942 228279 313994 228285
rect 313942 228221 313994 228227
rect 313460 228170 313516 228179
rect 313460 228105 313516 228114
rect 313366 223099 313418 223105
rect 313366 223041 313418 223047
rect 313858 221482 313886 228221
rect 314530 221792 314558 231033
rect 314914 230431 314942 239686
rect 315298 234797 315326 239686
rect 315286 234791 315338 234797
rect 315286 234733 315338 234739
rect 314902 230425 314954 230431
rect 314902 230367 314954 230373
rect 315382 227465 315434 227471
rect 315382 227407 315434 227413
rect 314530 221764 314606 221792
rect 314578 221482 314606 221764
rect 315394 221482 315422 227407
rect 315778 225621 315806 239686
rect 316176 239672 316382 239700
rect 316512 239672 316766 239700
rect 316896 239672 317150 239700
rect 316150 229685 316202 229691
rect 316150 229627 316202 229633
rect 315766 225615 315818 225621
rect 315766 225557 315818 225563
rect 316162 221482 316190 229627
rect 316354 224659 316382 239672
rect 316738 231287 316766 239672
rect 317122 237461 317150 239672
rect 317110 237455 317162 237461
rect 317110 237397 317162 237403
rect 317218 233465 317246 239686
rect 317602 237535 317630 239686
rect 317590 237529 317642 237535
rect 317590 237471 317642 237477
rect 317206 233459 317258 233465
rect 317206 233401 317258 233407
rect 316724 231278 316780 231287
rect 316724 231213 316780 231222
rect 317590 230573 317642 230579
rect 317590 230515 317642 230521
rect 316822 229611 316874 229617
rect 316822 229553 316874 229559
rect 316342 224653 316394 224659
rect 316342 224595 316394 224601
rect 316834 221792 316862 229553
rect 316834 221764 316910 221792
rect 316882 221482 316910 221764
rect 317602 221482 317630 230515
rect 317986 229987 318014 239686
rect 318384 239672 318590 239700
rect 318720 239672 318974 239700
rect 319200 239672 319454 239700
rect 318358 234643 318410 234649
rect 318358 234585 318410 234591
rect 317974 229981 318026 229987
rect 317974 229923 318026 229929
rect 318370 227471 318398 234585
rect 318358 227465 318410 227471
rect 318358 227407 318410 227413
rect 318358 225689 318410 225695
rect 318358 225631 318410 225637
rect 318370 221482 318398 225631
rect 318562 223179 318590 239672
rect 318946 225219 318974 239672
rect 319426 236174 319454 239672
rect 319330 236146 319454 236174
rect 319126 229537 319178 229543
rect 319126 229479 319178 229485
rect 318932 225210 318988 225219
rect 318932 225145 318988 225154
rect 318550 223173 318602 223179
rect 318550 223115 318602 223121
rect 319138 221792 319166 229479
rect 319330 224511 319358 236146
rect 319414 234495 319466 234501
rect 319414 234437 319466 234443
rect 319426 227767 319454 234437
rect 319522 233613 319550 239686
rect 319906 236129 319934 239686
rect 319894 236123 319946 236129
rect 319894 236065 319946 236071
rect 319606 235975 319658 235981
rect 319606 235917 319658 235923
rect 319510 233607 319562 233613
rect 319510 233549 319562 233555
rect 319618 230801 319646 235917
rect 320290 234649 320318 239686
rect 320640 239672 320894 239700
rect 321024 239672 321278 239700
rect 321408 239672 321662 239700
rect 320866 236795 320894 239672
rect 320854 236789 320906 236795
rect 320854 236731 320906 236737
rect 320278 234643 320330 234649
rect 320278 234585 320330 234591
rect 320854 234569 320906 234575
rect 320854 234511 320906 234517
rect 320662 231239 320714 231245
rect 320662 231181 320714 231187
rect 319606 230795 319658 230801
rect 319606 230737 319658 230743
rect 319414 227761 319466 227767
rect 319414 227703 319466 227709
rect 319894 227613 319946 227619
rect 319894 227555 319946 227561
rect 319318 224505 319370 224511
rect 319318 224447 319370 224453
rect 319138 221764 319214 221792
rect 319186 221482 319214 221764
rect 319906 221482 319934 227555
rect 320674 221482 320702 231181
rect 320866 230727 320894 234511
rect 320854 230721 320906 230727
rect 320854 230663 320906 230669
rect 321250 230357 321278 239672
rect 321634 234871 321662 239672
rect 321622 234865 321674 234871
rect 321622 234807 321674 234813
rect 321238 230351 321290 230357
rect 321238 230293 321290 230299
rect 321334 225985 321386 225991
rect 321334 225927 321386 225933
rect 321346 221792 321374 225927
rect 321730 225695 321758 239686
rect 322128 239672 322334 239700
rect 322006 236049 322058 236055
rect 322006 235991 322058 235997
rect 322018 230505 322046 235991
rect 322102 231609 322154 231615
rect 322102 231551 322154 231557
rect 322006 230499 322058 230505
rect 322006 230441 322058 230447
rect 321718 225689 321770 225695
rect 321718 225631 321770 225637
rect 321346 221764 321422 221792
rect 321394 221482 321422 221764
rect 322114 221482 322142 231551
rect 322306 224437 322334 239672
rect 322498 231435 322526 239686
rect 322944 239672 323198 239700
rect 323328 239672 323582 239700
rect 323712 239672 323966 239700
rect 322484 231426 322540 231435
rect 322484 231361 322540 231370
rect 322966 230203 323018 230209
rect 322966 230145 323018 230151
rect 322294 224431 322346 224437
rect 322294 224373 322346 224379
rect 322978 221496 323006 230145
rect 323170 224585 323198 239672
rect 323554 234501 323582 239672
rect 323938 238867 323966 239672
rect 323926 238861 323978 238867
rect 323926 238803 323978 238809
rect 323830 235679 323882 235685
rect 323830 235621 323882 235627
rect 323542 234495 323594 234501
rect 323542 234437 323594 234443
rect 323638 231017 323690 231023
rect 323638 230959 323690 230965
rect 323158 224579 323210 224585
rect 323158 224521 323210 224527
rect 322944 221468 323006 221496
rect 323650 221496 323678 230959
rect 323842 230579 323870 235621
rect 323830 230573 323882 230579
rect 323830 230515 323882 230521
rect 324034 230135 324062 239686
rect 324418 238941 324446 239686
rect 324406 238935 324458 238941
rect 324406 238877 324458 238883
rect 324118 235161 324170 235167
rect 324118 235103 324170 235109
rect 324022 230129 324074 230135
rect 324022 230071 324074 230077
rect 324130 226879 324158 235103
rect 324802 233539 324830 239686
rect 325152 239672 325214 239700
rect 325536 239672 325790 239700
rect 325920 239672 326174 239700
rect 325186 236174 325214 239672
rect 325186 236146 325406 236174
rect 325270 234939 325322 234945
rect 325270 234881 325322 234887
rect 324790 233533 324842 233539
rect 324790 233475 324842 233481
rect 325174 231683 325226 231689
rect 325174 231625 325226 231631
rect 324118 226873 324170 226879
rect 324118 226815 324170 226821
rect 324406 225245 324458 225251
rect 324406 225187 324458 225193
rect 323650 221468 323712 221496
rect 324418 221482 324446 225187
rect 325186 221496 325214 231625
rect 325282 230949 325310 234881
rect 325270 230943 325322 230949
rect 325270 230885 325322 230891
rect 325378 224363 325406 236146
rect 325762 230209 325790 239672
rect 326146 235685 326174 239672
rect 326134 235679 326186 235685
rect 326134 235621 326186 235627
rect 326242 233539 326270 239686
rect 326722 238793 326750 239686
rect 326710 238787 326762 238793
rect 326710 238729 326762 238735
rect 326710 235605 326762 235611
rect 326710 235547 326762 235553
rect 325942 233533 325994 233539
rect 325942 233475 325994 233481
rect 326230 233533 326282 233539
rect 326230 233475 326282 233481
rect 325750 230203 325802 230209
rect 325750 230145 325802 230151
rect 325846 227687 325898 227693
rect 325846 227629 325898 227635
rect 325366 224357 325418 224363
rect 325366 224299 325418 224305
rect 325152 221468 325214 221496
rect 325858 221496 325886 227629
rect 325954 225367 325982 233475
rect 326614 233237 326666 233243
rect 326614 233179 326666 233185
rect 326626 227120 326654 233179
rect 326722 230875 326750 235547
rect 327106 231583 327134 239686
rect 327456 239672 327710 239700
rect 327840 239672 327998 239700
rect 327682 234945 327710 239672
rect 327670 234939 327722 234945
rect 327670 234881 327722 234887
rect 327092 231574 327148 231583
rect 327092 231509 327148 231518
rect 326710 230869 326762 230875
rect 326710 230811 326762 230817
rect 326806 230277 326858 230283
rect 326806 230219 326858 230225
rect 326818 227767 326846 230219
rect 326806 227761 326858 227767
rect 326806 227703 326858 227709
rect 326626 227092 326750 227120
rect 325940 225358 325996 225367
rect 325940 225293 325996 225302
rect 325858 221468 325920 221496
rect 326722 221482 326750 227092
rect 327382 225911 327434 225917
rect 327382 225853 327434 225859
rect 327394 221792 327422 225853
rect 327970 225663 327998 239672
rect 328162 236174 328190 239686
rect 328162 236146 328286 236174
rect 328150 233607 328202 233613
rect 328150 233549 328202 233555
rect 328054 231757 328106 231763
rect 328054 231699 328106 231705
rect 328066 226380 328094 231699
rect 328162 231615 328190 233549
rect 328150 231609 328202 231615
rect 328150 231551 328202 231557
rect 328066 226352 328190 226380
rect 327956 225654 328012 225663
rect 327956 225589 328012 225598
rect 327394 221764 327470 221792
rect 327442 221482 327470 221764
rect 328162 221482 328190 226352
rect 328258 224289 328286 236146
rect 328342 233755 328394 233761
rect 328342 233697 328394 233703
rect 328354 231023 328382 233697
rect 328342 231017 328394 231023
rect 328342 230959 328394 230965
rect 328546 229839 328574 239686
rect 328930 238719 328958 239686
rect 328918 238713 328970 238719
rect 328918 238655 328970 238661
rect 329314 234575 329342 239686
rect 329664 239672 329918 239700
rect 330048 239672 330302 239700
rect 330480 239672 330782 239700
rect 330864 239672 331166 239700
rect 331248 239672 331550 239700
rect 329890 238645 329918 239672
rect 329878 238639 329930 238645
rect 329878 238581 329930 238587
rect 329302 234569 329354 234575
rect 329302 234511 329354 234517
rect 330274 231731 330302 239672
rect 330754 233761 330782 239672
rect 331138 236174 331166 239672
rect 331042 236146 331166 236174
rect 330742 233755 330794 233761
rect 330742 233697 330794 233703
rect 330260 231722 330316 231731
rect 330260 231657 330316 231666
rect 329590 230943 329642 230949
rect 329590 230885 329642 230891
rect 329206 230351 329258 230357
rect 329206 230293 329258 230299
rect 329218 229987 329246 230293
rect 329206 229981 329258 229987
rect 329206 229923 329258 229929
rect 328534 229833 328586 229839
rect 328534 229775 328586 229781
rect 328918 228427 328970 228433
rect 328918 228369 328970 228375
rect 328246 224283 328298 224289
rect 328246 224225 328298 224231
rect 328930 221482 328958 228369
rect 329602 221792 329630 230885
rect 330454 225837 330506 225843
rect 331042 225811 331070 236146
rect 331414 235087 331466 235093
rect 331414 235029 331466 235035
rect 331222 234125 331274 234131
rect 331222 234067 331274 234073
rect 331234 230949 331262 234067
rect 331318 233089 331370 233095
rect 331318 233031 331370 233037
rect 331222 230943 331274 230949
rect 331222 230885 331274 230891
rect 331126 229833 331178 229839
rect 331126 229775 331178 229781
rect 331138 228433 331166 229775
rect 331126 228427 331178 228433
rect 331126 228369 331178 228375
rect 331330 226972 331358 233031
rect 331234 226944 331358 226972
rect 330454 225779 330506 225785
rect 331028 225802 331084 225811
rect 329602 221764 329678 221792
rect 329650 221482 329678 221764
rect 330466 221482 330494 225779
rect 331028 225737 331084 225746
rect 331234 221482 331262 226944
rect 331426 225917 331454 235029
rect 331414 225911 331466 225917
rect 331414 225853 331466 225859
rect 331522 224215 331550 239672
rect 331618 229987 331646 239686
rect 331968 239672 332222 239700
rect 332352 239672 332606 239700
rect 332194 235611 332222 239672
rect 332578 235981 332606 239672
rect 332674 238571 332702 239686
rect 332662 238565 332714 238571
rect 332662 238507 332714 238513
rect 332566 235975 332618 235981
rect 332566 235917 332618 235923
rect 332182 235605 332234 235611
rect 332182 235547 332234 235553
rect 331894 230055 331946 230061
rect 331894 229997 331946 230003
rect 331606 229981 331658 229987
rect 331606 229923 331658 229929
rect 331510 224209 331562 224215
rect 331510 224151 331562 224157
rect 331906 221792 331934 229997
rect 333058 228327 333086 239686
rect 333442 235093 333470 239686
rect 333430 235087 333482 235093
rect 333430 235029 333482 235035
rect 333044 228318 333100 228327
rect 333044 228253 333100 228262
rect 333826 225959 333854 239686
rect 334272 239672 334526 239700
rect 334656 239672 334910 239700
rect 334294 234273 334346 234279
rect 334294 234215 334346 234221
rect 334102 233681 334154 233687
rect 334102 233623 334154 233629
rect 334114 231245 334142 233623
rect 334198 233163 334250 233169
rect 334198 233105 334250 233111
rect 334102 231239 334154 231245
rect 334102 231181 334154 231187
rect 333812 225950 333868 225959
rect 333812 225885 333868 225894
rect 333526 225171 333578 225177
rect 333526 225113 333578 225119
rect 332662 223839 332714 223845
rect 332662 223781 332714 223787
rect 331906 221764 331982 221792
rect 331954 221482 331982 221764
rect 332674 221482 332702 223781
rect 333538 221482 333566 225113
rect 334210 221792 334238 233105
rect 334306 226065 334334 234215
rect 334294 226059 334346 226065
rect 334294 226001 334346 226007
rect 334498 224141 334526 239672
rect 334882 233211 334910 239672
rect 334978 235167 335006 239686
rect 334966 235161 335018 235167
rect 334966 235103 335018 235109
rect 335362 233613 335390 239686
rect 335746 238497 335774 239686
rect 336096 239672 336350 239700
rect 336480 239672 336734 239700
rect 335734 238491 335786 238497
rect 335734 238433 335786 238439
rect 335350 233607 335402 233613
rect 335350 233549 335402 233555
rect 334868 233202 334924 233211
rect 334868 233137 334924 233146
rect 336322 229913 336350 239672
rect 336706 238423 336734 239672
rect 336850 239404 336878 239686
rect 336850 239376 336926 239404
rect 336694 238417 336746 238423
rect 336694 238359 336746 238365
rect 336310 229907 336362 229913
rect 336310 229849 336362 229855
rect 334966 229463 335018 229469
rect 334966 229405 335018 229411
rect 334486 224135 334538 224141
rect 334486 224077 334538 224083
rect 334210 221764 334286 221792
rect 334258 221482 334286 221764
rect 334978 221482 335006 229405
rect 336898 227439 336926 239376
rect 336884 227430 336940 227439
rect 336884 227365 336940 227374
rect 336406 225023 336458 225029
rect 336406 224965 336458 224971
rect 335734 223765 335786 223771
rect 335734 223707 335786 223713
rect 335746 221482 335774 223707
rect 336418 221792 336446 224965
rect 337186 224067 337214 239686
rect 337270 232867 337322 232873
rect 337270 232809 337322 232815
rect 337174 224061 337226 224067
rect 337174 224003 337226 224009
rect 336418 221764 336494 221792
rect 336466 221482 336494 221764
rect 337282 221482 337310 232809
rect 337570 231689 337598 239686
rect 338050 234131 338078 239686
rect 338400 239672 338654 239700
rect 338784 239672 339038 239700
rect 339168 239672 339422 239700
rect 338626 234247 338654 239672
rect 339010 238349 339038 239672
rect 338998 238343 339050 238349
rect 338998 238285 339050 238291
rect 338612 234238 338668 234247
rect 338612 234173 338668 234182
rect 338038 234125 338090 234131
rect 338038 234067 338090 234073
rect 339094 233903 339146 233909
rect 339094 233845 339146 233851
rect 338038 233015 338090 233021
rect 338038 232957 338090 232963
rect 337558 231683 337610 231689
rect 337558 231625 337610 231631
rect 338050 221482 338078 232957
rect 339106 225177 339134 233845
rect 339190 232867 339242 232873
rect 339190 232809 339242 232815
rect 339202 232355 339230 232809
rect 339286 232497 339338 232503
rect 339286 232439 339338 232445
rect 339298 232355 339326 232439
rect 339190 232349 339242 232355
rect 339190 232291 339242 232297
rect 339286 232349 339338 232355
rect 339286 232291 339338 232297
rect 339394 228475 339422 239672
rect 339490 234279 339518 239686
rect 339478 234273 339530 234279
rect 339478 234215 339530 234221
rect 339766 233977 339818 233983
rect 339766 233919 339818 233925
rect 339478 232571 339530 232577
rect 339478 232513 339530 232519
rect 339490 232133 339518 232513
rect 339478 232127 339530 232133
rect 339478 232069 339530 232075
rect 339380 228466 339436 228475
rect 339380 228401 339436 228410
rect 339478 226873 339530 226879
rect 339478 226815 339530 226821
rect 339094 225171 339146 225177
rect 339094 225113 339146 225119
rect 338710 223617 338762 223623
rect 338710 223559 338762 223565
rect 338722 221792 338750 223559
rect 338722 221764 338798 221792
rect 338770 221482 338798 221764
rect 339490 221482 339518 226815
rect 339778 225103 339806 233919
rect 339874 230399 339902 239686
rect 340272 239672 340478 239700
rect 340608 239672 340862 239700
rect 340992 239672 341246 239700
rect 341376 239672 341630 239700
rect 340246 232719 340298 232725
rect 340246 232661 340298 232667
rect 339860 230390 339916 230399
rect 339860 230325 339916 230334
rect 339766 225097 339818 225103
rect 339766 225039 339818 225045
rect 340258 221482 340286 232661
rect 340450 223993 340478 239672
rect 340834 233243 340862 239672
rect 341218 239237 341246 239672
rect 341206 239231 341258 239237
rect 341206 239173 341258 239179
rect 341602 234395 341630 239672
rect 341794 238275 341822 239686
rect 341782 238269 341834 238275
rect 341782 238211 341834 238217
rect 341588 234386 341644 234395
rect 341588 234321 341644 234330
rect 340822 233237 340874 233243
rect 340822 233179 340874 233185
rect 342178 228771 342206 239686
rect 342562 235241 342590 239686
rect 342912 239672 343166 239700
rect 343296 239672 343550 239700
rect 342550 235235 342602 235241
rect 342550 235177 342602 235183
rect 342358 234199 342410 234205
rect 342358 234141 342410 234147
rect 342164 228762 342220 228771
rect 342164 228697 342220 228706
rect 342370 227989 342398 234141
rect 341014 227983 341066 227989
rect 341014 227925 341066 227931
rect 342358 227983 342410 227989
rect 342358 227925 342410 227931
rect 340438 223987 340490 223993
rect 340438 223929 340490 223935
rect 341026 221792 341054 227925
rect 343138 227291 343166 239672
rect 343522 235907 343550 239672
rect 343510 235901 343562 235907
rect 343510 235843 343562 235849
rect 343222 232497 343274 232503
rect 343222 232439 343274 232445
rect 343124 227282 343180 227291
rect 343124 227217 343180 227226
rect 342550 225763 342602 225769
rect 342550 225705 342602 225711
rect 341782 223691 341834 223697
rect 341782 223633 341834 223639
rect 341026 221764 341102 221792
rect 341074 221482 341102 221764
rect 341794 221482 341822 223633
rect 342562 221482 342590 225705
rect 343234 221792 343262 232439
rect 343618 223919 343646 239686
rect 344016 239672 344318 239700
rect 344182 232497 344234 232503
rect 344182 232439 344234 232445
rect 344194 232281 344222 232439
rect 344290 232281 344318 239672
rect 344386 235135 344414 239686
rect 344372 235126 344428 235135
rect 344372 235061 344428 235070
rect 344182 232275 344234 232281
rect 344182 232217 344234 232223
rect 344278 232275 344330 232281
rect 344278 232217 344330 232223
rect 343990 228131 344042 228137
rect 343990 228073 344042 228079
rect 343606 223913 343658 223919
rect 343606 223855 343658 223861
rect 343234 221764 343310 221792
rect 343282 221482 343310 221764
rect 344002 221482 344030 228073
rect 344770 227143 344798 239686
rect 345120 239672 345374 239700
rect 345346 238201 345374 239672
rect 345538 239672 345600 239700
rect 345334 238195 345386 238201
rect 345334 238137 345386 238143
rect 345538 236174 345566 239672
rect 345442 236146 345566 236174
rect 345332 234830 345388 234839
rect 345332 234765 345388 234774
rect 345346 228137 345374 234765
rect 345442 228623 345470 236146
rect 345922 234205 345950 239686
rect 346320 239672 346622 239700
rect 345910 234199 345962 234205
rect 345910 234141 345962 234147
rect 345526 233829 345578 233835
rect 345526 233771 345578 233777
rect 345538 231097 345566 233771
rect 346294 232645 346346 232651
rect 346294 232587 346346 232593
rect 345526 231091 345578 231097
rect 345526 231033 345578 231039
rect 345428 228614 345484 228623
rect 345428 228549 345484 228558
rect 345334 228131 345386 228137
rect 345334 228073 345386 228079
rect 344756 227134 344812 227143
rect 344756 227069 344812 227078
rect 345526 225911 345578 225917
rect 345526 225853 345578 225859
rect 344854 223543 344906 223549
rect 344854 223485 344906 223491
rect 344866 221482 344894 223485
rect 345538 221792 345566 225853
rect 345538 221764 345614 221792
rect 345586 221482 345614 221764
rect 346306 221482 346334 232587
rect 346594 223845 346622 239672
rect 346690 238127 346718 239686
rect 346678 238121 346730 238127
rect 346678 238063 346730 238069
rect 346966 233311 347018 233317
rect 346966 233253 347018 233259
rect 346978 225917 347006 233253
rect 347074 233169 347102 239686
rect 347424 239672 347678 239700
rect 347808 239672 348062 239700
rect 347650 234839 347678 239672
rect 347636 234830 347692 234839
rect 347636 234765 347692 234774
rect 347062 233163 347114 233169
rect 347062 233105 347114 233111
rect 347062 229389 347114 229395
rect 347062 229331 347114 229337
rect 346966 225911 347018 225917
rect 346966 225853 347018 225859
rect 346582 223839 346634 223845
rect 346582 223781 346634 223787
rect 347074 221482 347102 229331
rect 348034 223549 348062 239672
rect 348130 223771 348158 239686
rect 348514 229839 348542 239686
rect 348898 235833 348926 239686
rect 349344 239672 349598 239700
rect 349728 239672 349982 239700
rect 350112 239672 350366 239700
rect 348886 235827 348938 235833
rect 348886 235769 348938 235775
rect 348694 235457 348746 235463
rect 348694 235399 348746 235405
rect 348502 229833 348554 229839
rect 348502 229775 348554 229781
rect 348598 227317 348650 227323
rect 348598 227259 348650 227265
rect 348118 223765 348170 223771
rect 348118 223707 348170 223713
rect 348022 223543 348074 223549
rect 348022 223485 348074 223491
rect 347734 223395 347786 223401
rect 347734 223337 347786 223343
rect 347746 221792 347774 223337
rect 347746 221764 347822 221792
rect 347794 221482 347822 221764
rect 348610 221482 348638 227259
rect 348706 224955 348734 235399
rect 349366 232423 349418 232429
rect 349366 232365 349418 232371
rect 348694 224949 348746 224955
rect 348694 224891 348746 224897
rect 349378 221482 349406 232365
rect 349570 223697 349598 239672
rect 349954 238053 349982 239672
rect 349942 238047 349994 238053
rect 349942 237989 349994 237995
rect 350338 233095 350366 239672
rect 350434 239163 350462 239686
rect 350832 239672 351134 239700
rect 350422 239157 350474 239163
rect 350422 239099 350474 239105
rect 350326 233089 350378 233095
rect 350326 233031 350378 233037
rect 350038 227835 350090 227841
rect 350038 227777 350090 227783
rect 349558 223691 349610 223697
rect 349558 223633 349610 223639
rect 350050 221792 350078 227777
rect 351106 223475 351134 239672
rect 351202 223623 351230 239686
rect 351552 239672 351806 239700
rect 351936 239672 352190 239700
rect 352320 239672 352574 239700
rect 351382 234051 351434 234057
rect 351382 233993 351434 233999
rect 351394 225251 351422 233993
rect 351778 229691 351806 239672
rect 352162 233909 352190 239672
rect 352150 233903 352202 233909
rect 352150 233845 352202 233851
rect 352342 232349 352394 232355
rect 352342 232291 352394 232297
rect 351766 229685 351818 229691
rect 351766 229627 351818 229633
rect 351574 227243 351626 227249
rect 351574 227185 351626 227191
rect 351382 225245 351434 225251
rect 351382 225187 351434 225193
rect 351190 223617 351242 223623
rect 351190 223559 351242 223565
rect 350806 223469 350858 223475
rect 350806 223411 350858 223417
rect 351094 223469 351146 223475
rect 351094 223411 351146 223417
rect 350050 221764 350126 221792
rect 350098 221482 350126 221764
rect 350818 221482 350846 223411
rect 351586 221482 351614 227185
rect 352354 221496 352382 232291
rect 352546 223401 352574 239672
rect 352738 237905 352766 239686
rect 352726 237899 352778 237905
rect 352726 237841 352778 237847
rect 353122 233021 353150 239686
rect 353506 237979 353534 239686
rect 353856 239672 354110 239700
rect 353494 237973 353546 237979
rect 353494 237915 353546 237921
rect 353110 233015 353162 233021
rect 353110 232957 353162 232963
rect 352726 230869 352778 230875
rect 352724 230834 352726 230843
rect 352778 230834 352780 230843
rect 352724 230769 352780 230778
rect 353110 227761 353162 227767
rect 353110 227703 353162 227709
rect 352534 223395 352586 223401
rect 352534 223337 352586 223343
rect 352354 221468 352416 221496
rect 353122 221482 353150 227703
rect 354082 223253 354110 239672
rect 354226 239404 354254 239686
rect 354624 239672 354878 239700
rect 354178 239376 354254 239404
rect 354178 224479 354206 239376
rect 354356 234978 354412 234987
rect 354356 234913 354412 234922
rect 354260 230390 354316 230399
rect 354260 230325 354316 230334
rect 354274 225515 354302 230325
rect 354260 225506 354316 225515
rect 354260 225441 354316 225450
rect 354370 225029 354398 234913
rect 354850 229617 354878 239672
rect 354946 233835 354974 239686
rect 355344 239672 355646 239700
rect 354934 233829 354986 233835
rect 354934 233771 354986 233777
rect 355318 232497 355370 232503
rect 355318 232439 355370 232445
rect 354838 229611 354890 229617
rect 354838 229553 354890 229559
rect 354550 226947 354602 226953
rect 354550 226889 354602 226895
rect 354358 225023 354410 225029
rect 354358 224965 354410 224971
rect 354164 224470 354220 224479
rect 354164 224405 354220 224414
rect 354070 223247 354122 223253
rect 354070 223189 354122 223195
rect 353878 222433 353930 222439
rect 353878 222375 353930 222381
rect 353890 221496 353918 222375
rect 353856 221468 353918 221496
rect 354562 221496 354590 226889
rect 354562 221468 354624 221496
rect 355330 221482 355358 232439
rect 355618 223327 355646 239672
rect 355714 237831 355742 239686
rect 356064 239672 356318 239700
rect 356544 239672 356798 239700
rect 355702 237825 355754 237831
rect 355702 237767 355754 237773
rect 356290 232873 356318 239672
rect 356470 235383 356522 235389
rect 356470 235325 356522 235331
rect 356086 232867 356138 232873
rect 356086 232809 356138 232815
rect 356278 232867 356330 232873
rect 356278 232809 356330 232815
rect 355606 223321 355658 223327
rect 355606 223263 355658 223269
rect 356098 221792 356126 232809
rect 356482 232207 356510 235325
rect 356770 235283 356798 239672
rect 356756 235274 356812 235283
rect 356756 235209 356812 235218
rect 356866 234987 356894 239686
rect 357264 239672 357470 239700
rect 356852 234978 356908 234987
rect 356852 234913 356908 234922
rect 356470 232201 356522 232207
rect 356470 232143 356522 232149
rect 357442 222999 357470 239672
rect 357634 229543 357662 239686
rect 358018 234057 358046 239686
rect 358368 239672 358622 239700
rect 358752 239672 359006 239700
rect 358594 237757 358622 239672
rect 358582 237751 358634 237757
rect 358582 237693 358634 237699
rect 358582 235309 358634 235315
rect 358582 235251 358634 235257
rect 358006 234051 358058 234057
rect 358006 233993 358058 233999
rect 358486 232275 358538 232281
rect 358486 232217 358538 232223
rect 358198 232127 358250 232133
rect 358198 232069 358250 232075
rect 357622 229537 357674 229543
rect 357622 229479 357674 229485
rect 358210 227534 358238 232069
rect 358498 231763 358526 232217
rect 358594 232133 358622 235251
rect 358582 232127 358634 232133
rect 358582 232069 358634 232075
rect 358486 231757 358538 231763
rect 358486 231699 358538 231705
rect 358594 230940 358910 230968
rect 358594 230801 358622 230940
rect 358774 230869 358826 230875
rect 358774 230811 358826 230817
rect 358582 230795 358634 230801
rect 358582 230737 358634 230743
rect 358786 230672 358814 230811
rect 358882 230801 358910 230940
rect 358870 230795 358922 230801
rect 358870 230737 358922 230743
rect 358402 230653 358622 230672
rect 358390 230647 358634 230653
rect 358442 230644 358582 230647
rect 358390 230589 358442 230595
rect 358582 230589 358634 230595
rect 358690 230644 358814 230672
rect 358690 230505 358718 230644
rect 358294 230499 358346 230505
rect 358294 230441 358346 230447
rect 358678 230499 358730 230505
rect 358678 230441 358730 230447
rect 358774 230499 358826 230505
rect 358774 230441 358826 230447
rect 358306 230376 358334 230441
rect 358786 230376 358814 230441
rect 358306 230348 358814 230376
rect 358978 229955 359006 239672
rect 359074 233063 359102 239686
rect 359060 233054 359116 233063
rect 359060 232989 359116 232998
rect 359060 230834 359116 230843
rect 359060 230769 359116 230778
rect 359074 230727 359102 230769
rect 359062 230721 359114 230727
rect 359062 230663 359114 230669
rect 358964 229946 359020 229955
rect 358964 229881 359020 229890
rect 359158 227909 359210 227915
rect 359158 227851 359210 227857
rect 358210 227506 358334 227534
rect 357622 227021 357674 227027
rect 357622 226963 357674 226969
rect 357428 222990 357484 222999
rect 357428 222925 357484 222934
rect 356854 222211 356906 222217
rect 356854 222153 356906 222159
rect 356098 221764 356174 221792
rect 356146 221482 356174 221764
rect 356866 221482 356894 222153
rect 357634 221482 357662 226963
rect 358306 221792 358334 227506
rect 358306 221764 358382 221792
rect 358354 221482 358382 221764
rect 359170 221482 359198 227851
rect 359458 224627 359486 239686
rect 359746 239672 359856 239700
rect 359444 224618 359500 224627
rect 359444 224553 359500 224562
rect 359746 224183 359774 239672
rect 359926 237677 359978 237683
rect 359926 237619 359978 237625
rect 359828 228910 359884 228919
rect 359828 228845 359884 228854
rect 359842 226953 359870 228845
rect 359830 226947 359882 226953
rect 359830 226889 359882 226895
rect 359732 224174 359788 224183
rect 359732 224109 359788 224118
rect 359938 221482 359966 237619
rect 360034 235759 360062 239765
rect 371446 239749 371498 239755
rect 360022 235753 360074 235759
rect 360022 235695 360074 235701
rect 360214 235013 360266 235019
rect 360214 234955 360266 234961
rect 360226 227534 360254 234955
rect 360322 233687 360350 239686
rect 360672 239672 360926 239700
rect 361056 239672 361310 239700
rect 360310 233681 360362 233687
rect 360310 233623 360362 233629
rect 360898 230399 360926 239672
rect 361282 233983 361310 239672
rect 361378 235315 361406 239686
rect 361762 237059 361790 239686
rect 361748 237050 361804 237059
rect 361748 236985 361804 236994
rect 361366 235309 361418 235315
rect 361366 235251 361418 235257
rect 361270 233977 361322 233983
rect 361270 233919 361322 233925
rect 361078 233903 361130 233909
rect 361078 233845 361130 233851
rect 361090 233687 361118 233845
rect 360982 233681 361034 233687
rect 360982 233623 361034 233629
rect 361078 233681 361130 233687
rect 361078 233623 361130 233629
rect 360884 230390 360940 230399
rect 360884 230325 360940 230334
rect 360226 227506 360350 227534
rect 360322 224807 360350 227506
rect 360598 227095 360650 227101
rect 360598 227037 360650 227043
rect 360310 224801 360362 224807
rect 360310 224743 360362 224749
rect 360610 221792 360638 227037
rect 360994 224331 361022 233623
rect 362146 232725 362174 239686
rect 362530 233317 362558 239686
rect 362880 239672 363134 239700
rect 363264 239672 363518 239700
rect 363106 237683 363134 239672
rect 363094 237677 363146 237683
rect 363094 237619 363146 237625
rect 362806 235531 362858 235537
rect 362806 235473 362858 235479
rect 362518 233311 362570 233317
rect 362518 233253 362570 233259
rect 362134 232719 362186 232725
rect 362134 232661 362186 232667
rect 361366 232571 361418 232577
rect 361366 232513 361418 232519
rect 360980 224322 361036 224331
rect 360980 224257 361036 224266
rect 360610 221764 360686 221792
rect 360658 221482 360686 221764
rect 361378 221482 361406 232513
rect 362230 232127 362282 232133
rect 362230 232069 362282 232075
rect 362242 230653 362270 232069
rect 362134 230647 362186 230653
rect 362134 230589 362186 230595
rect 362230 230647 362282 230653
rect 362230 230589 362282 230595
rect 362146 221482 362174 230589
rect 362818 228156 362846 235473
rect 362818 228128 362942 228156
rect 362914 228063 362942 228128
rect 362806 228057 362858 228063
rect 362806 227999 362858 228005
rect 362902 228057 362954 228063
rect 362902 227999 362954 228005
rect 362818 224881 362846 227999
rect 362806 224875 362858 224881
rect 362806 224817 362858 224823
rect 363490 224035 363518 239672
rect 363586 230103 363614 239686
rect 363670 237603 363722 237609
rect 363670 237545 363722 237551
rect 363572 230094 363628 230103
rect 363572 230029 363628 230038
rect 363476 224026 363532 224035
rect 363476 223961 363532 223970
rect 363682 221940 363710 237545
rect 364066 234543 364094 239686
rect 364450 237609 364478 239686
rect 364800 239672 365054 239700
rect 365184 239672 365438 239700
rect 365568 239672 365726 239700
rect 365904 239672 366206 239700
rect 364438 237603 364490 237609
rect 364438 237545 364490 237551
rect 364052 234534 364108 234543
rect 364052 234469 364108 234478
rect 365026 232503 365054 239672
rect 365410 232651 365438 239672
rect 365698 233359 365726 239672
rect 365684 233350 365740 233359
rect 365684 233285 365740 233294
rect 365398 232645 365450 232651
rect 365398 232587 365450 232593
rect 365014 232497 365066 232503
rect 365014 232439 365066 232445
rect 365206 232201 365258 232207
rect 365206 232143 365258 232149
rect 364438 232053 364490 232059
rect 364438 231995 364490 232001
rect 364054 231165 364106 231171
rect 364054 231107 364106 231113
rect 364066 226879 364094 231107
rect 364054 226873 364106 226879
rect 364054 226815 364106 226821
rect 363766 224727 363818 224733
rect 363766 224669 363818 224675
rect 363010 221912 363710 221940
rect 363010 221792 363038 221912
rect 362962 221764 363038 221792
rect 362962 221482 362990 221764
rect 363778 221755 363806 224669
rect 363682 221727 363806 221755
rect 363682 221482 363710 221727
rect 364450 221482 364478 231995
rect 365218 230801 365246 232143
rect 365110 230795 365162 230801
rect 365110 230737 365162 230743
rect 365206 230795 365258 230801
rect 365206 230737 365258 230743
rect 365122 221792 365150 230737
rect 366178 223887 366206 239672
rect 366274 232429 366302 239686
rect 366262 232423 366314 232429
rect 366262 232365 366314 232371
rect 366658 229469 366686 239686
rect 367008 239672 367262 239700
rect 367392 239672 367646 239700
rect 367872 239672 368126 239700
rect 366742 236863 366794 236869
rect 366742 236805 366794 236811
rect 366646 229463 366698 229469
rect 366646 229405 366698 229411
rect 366754 226972 366782 236805
rect 367234 236023 367262 239672
rect 367220 236014 367276 236023
rect 367220 235949 367276 235958
rect 367414 231905 367466 231911
rect 367414 231847 367466 231853
rect 367030 229389 367082 229395
rect 367030 229331 367082 229337
rect 366274 226944 366782 226972
rect 366164 223878 366220 223887
rect 366164 223813 366220 223822
rect 366274 223716 366302 226944
rect 366742 226799 366794 226805
rect 366742 226741 366794 226747
rect 365890 223688 366302 223716
rect 365122 221764 365198 221792
rect 365170 221482 365198 221764
rect 365890 221482 365918 223688
rect 366754 221482 366782 226741
rect 367042 224807 367070 229331
rect 367030 224801 367082 224807
rect 367030 224743 367082 224749
rect 367426 221792 367454 231847
rect 367618 223739 367646 239672
rect 368098 232207 368126 239672
rect 368194 232577 368222 239686
rect 368578 239089 368606 239686
rect 368566 239083 368618 239089
rect 368566 239025 368618 239031
rect 368962 237059 368990 239686
rect 369312 239672 369566 239700
rect 369696 239672 369950 239700
rect 370080 239672 370334 239700
rect 371446 239691 371498 239697
rect 368948 237050 369004 237059
rect 368948 236985 369004 236994
rect 368950 236937 369002 236943
rect 368950 236879 369002 236885
rect 368182 232571 368234 232577
rect 368182 232513 368234 232519
rect 368086 232201 368138 232207
rect 368086 232143 368138 232149
rect 368182 230499 368234 230505
rect 368182 230441 368234 230447
rect 367604 223730 367660 223739
rect 367604 223665 367660 223674
rect 367426 221764 367502 221792
rect 367474 221482 367502 221764
rect 368194 221482 368222 230441
rect 368962 221482 368990 236879
rect 369538 232281 369566 239672
rect 369526 232275 369578 232281
rect 369526 232217 369578 232223
rect 369922 229469 369950 239672
rect 370198 235309 370250 235315
rect 370198 235251 370250 235257
rect 370210 234871 370238 235251
rect 370306 234871 370334 239672
rect 370402 236911 370430 239686
rect 370388 236902 370444 236911
rect 370388 236837 370444 236846
rect 370198 234865 370250 234871
rect 370198 234807 370250 234813
rect 370294 234865 370346 234871
rect 370294 234807 370346 234813
rect 370786 232915 370814 239686
rect 370772 232906 370828 232915
rect 370772 232841 370828 232850
rect 371170 232355 371198 239686
rect 371458 236129 371486 239691
rect 371616 239672 371870 239700
rect 372000 239672 372254 239700
rect 371842 236129 371870 239672
rect 372226 236319 372254 239672
rect 372212 236310 372268 236319
rect 372212 236245 372268 236254
rect 371446 236123 371498 236129
rect 371446 236065 371498 236071
rect 371830 236123 371882 236129
rect 371830 236065 371882 236071
rect 371638 233755 371690 233761
rect 371638 233697 371690 233703
rect 371158 232349 371210 232355
rect 371158 232291 371210 232297
rect 370390 232127 370442 232133
rect 370390 232069 370442 232075
rect 369910 229463 369962 229469
rect 369910 229405 369962 229411
rect 370402 227534 370430 232069
rect 371446 229463 371498 229469
rect 371446 229405 371498 229411
rect 371458 229321 371486 229405
rect 371254 229315 371306 229321
rect 371254 229257 371306 229263
rect 371446 229315 371498 229321
rect 371446 229257 371498 229263
rect 370402 227506 370526 227534
rect 369622 227169 369674 227175
rect 369622 227111 369674 227117
rect 369634 221792 369662 227111
rect 369634 221764 369710 221792
rect 369682 221482 369710 221764
rect 370498 221482 370526 227506
rect 371266 221482 371294 229257
rect 371542 229241 371594 229247
rect 371542 229183 371594 229189
rect 371554 225769 371582 229183
rect 371542 225763 371594 225769
rect 371542 225705 371594 225711
rect 371650 222439 371678 233697
rect 372322 231985 372350 239686
rect 372706 232133 372734 239686
rect 372694 232127 372746 232133
rect 372694 232069 372746 232075
rect 372310 231979 372362 231985
rect 372310 231921 372362 231927
rect 372790 231313 372842 231319
rect 372790 231255 372842 231261
rect 372802 226731 372830 231255
rect 373090 229807 373118 239686
rect 373474 236615 373502 239686
rect 373824 239672 374078 239700
rect 374208 239672 374366 239700
rect 373460 236606 373516 236615
rect 373460 236541 373516 236550
rect 373462 232053 373514 232059
rect 373462 231995 373514 232001
rect 373076 229798 373132 229807
rect 373076 229733 373132 229742
rect 372694 226725 372746 226731
rect 372694 226667 372746 226673
rect 372790 226725 372842 226731
rect 372790 226667 372842 226673
rect 371638 222433 371690 222439
rect 371638 222375 371690 222381
rect 371926 222285 371978 222291
rect 371926 222227 371978 222233
rect 371938 221792 371966 222227
rect 371938 221764 372014 221792
rect 371986 221482 372014 221764
rect 372706 221482 372734 226667
rect 373474 221482 373502 231995
rect 374050 231837 374078 239672
rect 374038 231831 374090 231837
rect 374038 231773 374090 231779
rect 374230 230573 374282 230579
rect 374230 230515 374282 230521
rect 374242 221792 374270 230515
rect 374338 229247 374366 239672
rect 374530 231911 374558 239686
rect 374914 236763 374942 239686
rect 374900 236754 374956 236763
rect 374900 236689 374956 236698
rect 375394 232767 375422 239686
rect 375380 232758 375436 232767
rect 375380 232693 375436 232702
rect 375778 231985 375806 239686
rect 376128 239672 376382 239700
rect 376512 239672 376766 239700
rect 376354 233655 376382 239672
rect 376534 236493 376586 236499
rect 376534 236435 376586 236441
rect 376546 236319 376574 236435
rect 376738 236319 376766 239672
rect 376532 236310 376588 236319
rect 376532 236245 376588 236254
rect 376724 236310 376780 236319
rect 376724 236245 376780 236254
rect 376340 233646 376396 233655
rect 376340 233581 376396 233590
rect 375766 231979 375818 231985
rect 375766 231921 375818 231927
rect 374518 231905 374570 231911
rect 374518 231847 374570 231853
rect 374614 231387 374666 231393
rect 374614 231329 374666 231335
rect 374326 229241 374378 229247
rect 374326 229183 374378 229189
rect 374518 229167 374570 229173
rect 374518 229109 374570 229115
rect 374422 229019 374474 229025
rect 374422 228961 374474 228967
rect 374434 225917 374462 228961
rect 374422 225911 374474 225917
rect 374422 225853 374474 225859
rect 374530 225843 374558 229109
rect 374626 226805 374654 231329
rect 376834 229659 376862 239686
rect 377026 239672 377232 239700
rect 376820 229650 376876 229659
rect 376820 229585 376876 229594
rect 377026 229173 377054 239672
rect 377204 233350 377260 233359
rect 377204 233285 377260 233294
rect 377110 230869 377162 230875
rect 377110 230811 377162 230817
rect 377014 229167 377066 229173
rect 377014 229109 377066 229115
rect 375766 227539 375818 227545
rect 377122 227534 377150 230811
rect 377218 229469 377246 233285
rect 377206 229463 377258 229469
rect 377206 229405 377258 229411
rect 377122 227506 377246 227534
rect 375766 227481 375818 227487
rect 374614 226799 374666 226805
rect 374614 226741 374666 226747
rect 374518 225837 374570 225843
rect 374518 225779 374570 225785
rect 374998 222359 375050 222365
rect 374998 222301 375050 222307
rect 374242 221764 374318 221792
rect 374290 221482 374318 221764
rect 375010 221482 375038 222301
rect 375778 221482 375806 227481
rect 376438 224801 376490 224807
rect 376438 224743 376490 224749
rect 376450 221792 376478 224743
rect 376450 221764 376526 221792
rect 376498 221482 376526 221764
rect 377218 221482 377246 227506
rect 377602 223591 377630 239686
rect 377986 237059 378014 239686
rect 378336 239672 378494 239700
rect 377780 237050 377836 237059
rect 377780 236985 377836 236994
rect 377972 237050 378028 237059
rect 377972 236985 378028 236994
rect 377794 236721 377822 236985
rect 377782 236715 377834 236721
rect 377782 236657 377834 236663
rect 378466 235019 378494 239672
rect 378706 239404 378734 239686
rect 378838 239675 378890 239681
rect 378838 239617 378890 239623
rect 378706 239376 378782 239404
rect 378646 238417 378698 238423
rect 378646 238359 378698 238365
rect 378658 237979 378686 238359
rect 378550 237973 378602 237979
rect 378550 237915 378602 237921
rect 378646 237973 378698 237979
rect 378646 237915 378698 237921
rect 378562 236869 378590 237915
rect 378550 236863 378602 236869
rect 378550 236805 378602 236811
rect 378454 235013 378506 235019
rect 378454 234955 378506 234961
rect 378646 234273 378698 234279
rect 378646 234215 378698 234221
rect 378658 234131 378686 234215
rect 378550 234125 378602 234131
rect 378550 234067 378602 234073
rect 378646 234125 378698 234131
rect 378646 234067 378698 234073
rect 378562 233909 378590 234067
rect 378550 233903 378602 233909
rect 378550 233845 378602 233851
rect 378754 232619 378782 239376
rect 378850 235685 378878 239617
rect 378838 235679 378890 235685
rect 378838 235621 378890 235627
rect 378838 234273 378890 234279
rect 378838 234215 378890 234221
rect 378850 234057 378878 234215
rect 378838 234051 378890 234057
rect 378838 233993 378890 233999
rect 379138 233951 379166 239686
rect 379536 239672 379838 239700
rect 379124 233942 379180 233951
rect 379124 233877 379180 233886
rect 378740 232610 378796 232619
rect 378740 232545 378796 232554
rect 378742 226651 378794 226657
rect 378742 226593 378794 226599
rect 378070 226429 378122 226435
rect 378070 226371 378122 226377
rect 377588 223582 377644 223591
rect 377588 223517 377644 223526
rect 378082 221482 378110 226371
rect 378754 221792 378782 226593
rect 379510 225763 379562 225769
rect 379510 225705 379562 225711
rect 378754 221764 378830 221792
rect 378802 221482 378830 221764
rect 379522 221482 379550 225705
rect 379810 223443 379838 239672
rect 379906 229025 379934 239686
rect 380256 239672 380510 239700
rect 381024 239672 381278 239700
rect 379990 231461 380042 231467
rect 379990 231403 380042 231409
rect 379894 229019 379946 229025
rect 379894 228961 379946 228967
rect 380002 226657 380030 231403
rect 380278 230721 380330 230727
rect 380278 230663 380330 230669
rect 380086 228501 380138 228507
rect 380086 228443 380138 228449
rect 379990 226651 380042 226657
rect 379990 226593 380042 226599
rect 380098 225769 380126 228443
rect 380086 225763 380138 225769
rect 380086 225705 380138 225711
rect 379796 223434 379852 223443
rect 379796 223369 379852 223378
rect 380290 221482 380318 230663
rect 380482 229099 380510 239672
rect 380470 229093 380522 229099
rect 380470 229035 380522 229041
rect 380758 228353 380810 228359
rect 380758 228295 380810 228301
rect 380566 226503 380618 226509
rect 380566 226445 380618 226451
rect 380578 226065 380606 226445
rect 380566 226059 380618 226065
rect 380566 226001 380618 226007
rect 380770 225991 380798 228295
rect 380758 225985 380810 225991
rect 380758 225927 380810 225933
rect 381250 223295 381278 239672
rect 381346 229511 381374 239686
rect 381730 232471 381758 239686
rect 382114 233803 382142 239686
rect 382560 239672 382814 239700
rect 382786 239015 382814 239672
rect 382930 239404 382958 239686
rect 383328 239672 383582 239700
rect 383062 239601 383114 239607
rect 383062 239543 383114 239549
rect 382930 239376 383006 239404
rect 382774 239009 382826 239015
rect 382774 238951 382826 238957
rect 382100 233794 382156 233803
rect 382100 233729 382156 233738
rect 382198 232941 382250 232947
rect 382198 232883 382250 232889
rect 381716 232462 381772 232471
rect 381716 232397 381772 232406
rect 381332 229502 381388 229511
rect 381332 229437 381388 229446
rect 381814 227465 381866 227471
rect 381814 227407 381866 227413
rect 381236 223286 381292 223295
rect 381236 223221 381292 223230
rect 381046 222507 381098 222513
rect 381046 222449 381098 222455
rect 381058 221496 381086 222449
rect 381058 221468 381120 221496
rect 381826 221482 381854 227407
rect 382210 224733 382238 232883
rect 382978 232027 383006 239376
rect 383074 235611 383102 239543
rect 383062 235605 383114 235611
rect 383062 235547 383114 235553
rect 382964 232018 383020 232027
rect 382964 231953 383020 231962
rect 383554 229363 383582 239672
rect 383650 233761 383678 239686
rect 384048 239672 384350 239700
rect 383638 233755 383690 233761
rect 383638 233697 383690 233703
rect 383540 229354 383596 229363
rect 383540 229289 383596 229298
rect 382966 228649 383018 228655
rect 382966 228591 383018 228597
rect 382978 225843 383006 228591
rect 383254 228205 383306 228211
rect 383254 228147 383306 228153
rect 382582 225837 382634 225843
rect 382582 225779 382634 225785
rect 382966 225837 383018 225843
rect 382966 225779 383018 225785
rect 382198 224727 382250 224733
rect 382198 224669 382250 224675
rect 382594 221496 382622 225779
rect 382560 221468 382622 221496
rect 383266 221496 383294 228147
rect 384022 227391 384074 227397
rect 384022 227333 384074 227339
rect 383266 221468 383328 221496
rect 384034 221482 384062 227333
rect 384322 223147 384350 239672
rect 384418 229215 384446 239686
rect 384768 239672 385022 239700
rect 385152 239672 385406 239700
rect 385536 239672 385694 239700
rect 384994 232323 385022 239672
rect 384980 232314 385036 232323
rect 384980 232249 385036 232258
rect 385378 232175 385406 239672
rect 385364 232166 385420 232175
rect 385364 232101 385420 232110
rect 384404 229206 384460 229215
rect 384404 229141 384460 229150
rect 385666 227175 385694 239672
rect 385858 235685 385886 239686
rect 386352 239672 386654 239700
rect 385846 235679 385898 235685
rect 385846 235621 385898 235627
rect 385750 235383 385802 235389
rect 385750 235325 385802 235331
rect 385654 227169 385706 227175
rect 385654 227111 385706 227117
rect 384790 226429 384842 226435
rect 384790 226371 384842 226377
rect 384308 223138 384364 223147
rect 384308 223073 384364 223082
rect 384802 221792 384830 226371
rect 385558 225911 385610 225917
rect 385558 225853 385610 225859
rect 384802 221764 384878 221792
rect 384850 221482 384878 221764
rect 385570 221482 385598 225853
rect 385762 222851 385790 235325
rect 385942 235309 385994 235315
rect 385942 235251 385994 235257
rect 385844 231870 385900 231879
rect 385844 231805 385900 231814
rect 385858 226435 385886 231805
rect 385954 230875 385982 235251
rect 385942 230869 385994 230875
rect 385942 230811 385994 230817
rect 385846 226429 385898 226435
rect 385846 226371 385898 226377
rect 386626 225991 386654 239672
rect 386722 236055 386750 239686
rect 387072 239672 387326 239700
rect 387456 239672 387710 239700
rect 386710 236049 386762 236055
rect 386710 235991 386762 235997
rect 386902 234865 386954 234871
rect 386902 234807 386954 234813
rect 386914 233909 386942 234807
rect 386806 233903 386858 233909
rect 386806 233845 386858 233851
rect 386902 233903 386954 233909
rect 386902 233845 386954 233851
rect 386422 225985 386474 225991
rect 386422 225927 386474 225933
rect 386614 225985 386666 225991
rect 386614 225927 386666 225933
rect 386434 224733 386462 225927
rect 386326 224727 386378 224733
rect 386326 224669 386378 224675
rect 386422 224727 386474 224733
rect 386422 224669 386474 224675
rect 385748 222842 385804 222851
rect 385748 222777 385804 222786
rect 386338 221482 386366 224669
rect 386818 222365 386846 233845
rect 386998 226059 387050 226065
rect 386998 226001 387050 226007
rect 386806 222359 386858 222365
rect 386806 222301 386858 222307
rect 387010 221792 387038 226001
rect 387298 225917 387326 239672
rect 387682 235537 387710 239672
rect 387670 235531 387722 235537
rect 387670 235473 387722 235479
rect 387778 227693 387806 239686
rect 387766 227687 387818 227693
rect 387766 227629 387818 227635
rect 388162 226509 388190 239686
rect 388436 237050 388492 237059
rect 388436 236985 388492 236994
rect 388450 236943 388478 236985
rect 388438 236937 388490 236943
rect 388438 236879 388490 236885
rect 388546 227249 388574 239686
rect 388724 237050 388780 237059
rect 388724 236985 388780 236994
rect 388738 236721 388766 236985
rect 388726 236715 388778 236721
rect 388726 236657 388778 236663
rect 388930 227534 388958 239686
rect 389280 239672 389534 239700
rect 389664 239672 389918 239700
rect 389506 227545 389534 239672
rect 389890 235463 389918 239672
rect 389878 235457 389930 235463
rect 389878 235399 389930 235405
rect 389494 227539 389546 227545
rect 388930 227506 389054 227534
rect 388534 227243 388586 227249
rect 388534 227185 388586 227191
rect 387766 226503 387818 226509
rect 387766 226445 387818 226451
rect 388150 226503 388202 226509
rect 388150 226445 388202 226451
rect 387286 225911 387338 225917
rect 387286 225853 387338 225859
rect 387010 221764 387086 221792
rect 387058 221482 387086 221764
rect 387778 221482 387806 226445
rect 388822 226429 388874 226435
rect 388822 226371 388874 226377
rect 388918 226429 388970 226435
rect 388918 226371 388970 226377
rect 388834 226065 388862 226371
rect 388930 226287 388958 226371
rect 389026 226287 389054 227506
rect 389494 227481 389546 227487
rect 390082 227471 390110 239686
rect 390070 227465 390122 227471
rect 390070 227407 390122 227413
rect 390466 227101 390494 239686
rect 390850 227323 390878 239686
rect 390838 227317 390890 227323
rect 390838 227259 390890 227265
rect 390454 227095 390506 227101
rect 390454 227037 390506 227043
rect 391234 226995 391262 239686
rect 391570 239404 391598 239686
rect 391968 239672 392222 239700
rect 391522 239376 391598 239404
rect 391522 231560 391550 239376
rect 391606 236345 391658 236351
rect 391606 236287 391658 236293
rect 391618 235241 391646 236287
rect 392194 235611 392222 239672
rect 392182 235605 392234 235611
rect 392182 235547 392234 235553
rect 391606 235235 391658 235241
rect 391606 235177 391658 235183
rect 391702 235161 391754 235167
rect 391702 235103 391754 235109
rect 391522 231532 391646 231560
rect 391220 226986 391276 226995
rect 391220 226921 391276 226930
rect 391618 226847 391646 231532
rect 391714 228359 391742 235103
rect 391702 228353 391754 228359
rect 391702 228295 391754 228301
rect 392290 227397 392318 239686
rect 392470 234939 392522 234945
rect 392470 234881 392522 234887
rect 392482 228285 392510 234881
rect 392374 228279 392426 228285
rect 392374 228221 392426 228227
rect 392470 228279 392522 228285
rect 392470 228221 392522 228227
rect 392278 227391 392330 227397
rect 392278 227333 392330 227339
rect 391604 226838 391660 226847
rect 391510 226799 391562 226805
rect 391604 226773 391660 226782
rect 391510 226741 391562 226747
rect 390070 226577 390122 226583
rect 390070 226519 390122 226525
rect 388918 226281 388970 226287
rect 388918 226223 388970 226229
rect 389014 226281 389066 226287
rect 389014 226223 389066 226229
rect 388822 226059 388874 226065
rect 388822 226001 388874 226007
rect 389302 225837 389354 225843
rect 389302 225779 389354 225785
rect 388630 225763 388682 225769
rect 388630 225705 388682 225711
rect 388642 221482 388670 225705
rect 389314 221792 389342 225779
rect 389314 221764 389390 221792
rect 389362 221482 389390 221764
rect 390082 221482 390110 226519
rect 390838 226355 390890 226361
rect 390838 226297 390890 226303
rect 390850 221482 390878 226297
rect 391522 221792 391550 226741
rect 391522 221764 391598 221792
rect 391570 221482 391598 221764
rect 392386 221482 392414 228221
rect 392674 227027 392702 239686
rect 393058 235875 393086 239686
rect 393044 235866 393100 235875
rect 393044 235801 393100 235810
rect 393442 235759 393470 239686
rect 393888 239672 394142 239700
rect 394272 239672 394526 239700
rect 394608 239672 394910 239700
rect 393430 235753 393482 235759
rect 393430 235695 393482 235701
rect 392662 227021 392714 227027
rect 392662 226963 392714 226969
rect 393142 226947 393194 226953
rect 393142 226889 393194 226895
rect 393154 221482 393182 226889
rect 393814 226725 393866 226731
rect 393814 226667 393866 226673
rect 393826 221792 393854 226667
rect 394114 226551 394142 239672
rect 394498 226699 394526 239672
rect 394774 239527 394826 239533
rect 394774 239469 394826 239475
rect 394582 236271 394634 236277
rect 394582 236213 394634 236219
rect 394594 235833 394622 236213
rect 394582 235827 394634 235833
rect 394582 235769 394634 235775
rect 394678 235087 394730 235093
rect 394678 235029 394730 235035
rect 394582 234125 394634 234131
rect 394582 234067 394634 234073
rect 394594 231319 394622 234067
rect 394582 231313 394634 231319
rect 394582 231255 394634 231261
rect 394690 231171 394718 235029
rect 394786 233317 394814 239469
rect 394882 235389 394910 239672
rect 394870 235383 394922 235389
rect 394870 235325 394922 235331
rect 394978 235315 395006 239686
rect 395376 239672 395582 239700
rect 395712 239672 395966 239700
rect 396096 239672 396350 239700
rect 396480 239672 396734 239700
rect 394966 235309 395018 235315
rect 394966 235251 395018 235257
rect 394870 234791 394922 234797
rect 394870 234733 394922 234739
rect 394774 233311 394826 233317
rect 394774 233253 394826 233259
rect 394678 231165 394730 231171
rect 394678 231107 394730 231113
rect 394882 228211 394910 234733
rect 395350 230943 395402 230949
rect 395350 230885 395402 230891
rect 394870 228205 394922 228211
rect 394870 228147 394922 228153
rect 394484 226690 394540 226699
rect 394484 226625 394540 226634
rect 394582 226651 394634 226657
rect 394582 226593 394634 226599
rect 394100 226542 394156 226551
rect 394100 226477 394156 226486
rect 394390 224949 394442 224955
rect 394390 224891 394442 224897
rect 394402 222291 394430 224891
rect 394390 222285 394442 222291
rect 394390 222227 394442 222233
rect 393826 221764 393902 221792
rect 393874 221482 393902 221764
rect 394594 221482 394622 226593
rect 395362 221482 395390 230885
rect 395554 226953 395582 239672
rect 395938 234057 395966 239672
rect 396322 235241 396350 239672
rect 396310 235235 396362 235241
rect 396310 235177 396362 235183
rect 396706 234131 396734 239672
rect 396802 235727 396830 239686
rect 397078 238417 397130 238423
rect 397078 238359 397130 238365
rect 397090 236467 397118 238359
rect 397076 236458 397132 236467
rect 397076 236393 397132 236402
rect 396788 235718 396844 235727
rect 396788 235653 396844 235662
rect 396980 235126 397036 235135
rect 396980 235061 397036 235070
rect 396694 234125 396746 234131
rect 396694 234067 396746 234073
rect 395926 234051 395978 234057
rect 395926 233993 395978 233999
rect 396406 227687 396458 227693
rect 396406 227629 396458 227635
rect 395542 226947 395594 226953
rect 395542 226889 395594 226895
rect 396118 226873 396170 226879
rect 396118 226815 396170 226821
rect 396130 221792 396158 226815
rect 396418 225769 396446 227629
rect 396406 225763 396458 225769
rect 396406 225705 396458 225711
rect 396790 225097 396842 225103
rect 396790 225039 396842 225045
rect 396802 222976 396830 225039
rect 396802 222948 396926 222976
rect 396130 221764 396206 221792
rect 396178 221482 396206 221764
rect 396898 221482 396926 222948
rect 396994 222513 397022 235061
rect 397186 226805 397214 239686
rect 397460 237050 397516 237059
rect 397460 236985 397516 236994
rect 397474 236721 397502 236985
rect 397556 236902 397612 236911
rect 397556 236837 397612 236846
rect 397462 236715 397514 236721
rect 397462 236657 397514 236663
rect 397570 236573 397598 236837
rect 397558 236567 397610 236573
rect 397558 236509 397610 236515
rect 397366 236493 397418 236499
rect 397364 236458 397366 236467
rect 397418 236458 397420 236467
rect 397364 236393 397420 236402
rect 397366 232793 397418 232799
rect 397366 232735 397418 232741
rect 397378 232596 397406 232735
rect 397378 232568 397502 232596
rect 397174 226799 397226 226805
rect 397174 226741 397226 226747
rect 397474 224733 397502 232568
rect 397666 226657 397694 239686
rect 398016 239672 398270 239700
rect 398400 239672 398654 239700
rect 398784 239672 399038 239700
rect 399120 239672 399422 239700
rect 397750 238417 397802 238423
rect 397750 238359 397802 238365
rect 397762 237059 397790 238359
rect 397748 237050 397804 237059
rect 397748 236985 397804 236994
rect 397750 236937 397802 236943
rect 397748 236902 397750 236911
rect 397802 236902 397804 236911
rect 397748 236837 397804 236846
rect 398242 234057 398270 239672
rect 398626 235093 398654 239672
rect 399010 235167 399038 239672
rect 398998 235161 399050 235167
rect 398998 235103 399050 235109
rect 398614 235087 398666 235093
rect 398614 235029 398666 235035
rect 398134 234051 398186 234057
rect 398134 233993 398186 233999
rect 398230 234051 398282 234057
rect 398230 233993 398282 233999
rect 398146 229067 398174 233993
rect 398132 229058 398188 229067
rect 398132 228993 398188 229002
rect 398326 227983 398378 227989
rect 398326 227925 398378 227931
rect 397654 226651 397706 226657
rect 397654 226593 397706 226599
rect 397654 224801 397706 224807
rect 397654 224743 397706 224749
rect 397462 224727 397514 224733
rect 397462 224669 397514 224675
rect 396982 222507 397034 222513
rect 396982 222449 397034 222455
rect 397666 221482 397694 224743
rect 398338 221792 398366 227925
rect 398806 227169 398858 227175
rect 398806 227111 398858 227117
rect 398902 227169 398954 227175
rect 398902 227111 398954 227117
rect 398710 226355 398762 226361
rect 398710 226297 398762 226303
rect 398722 226065 398750 226297
rect 398818 226065 398846 227111
rect 398914 226509 398942 227111
rect 399394 226879 399422 239672
rect 399490 228919 399518 239686
rect 399874 235579 399902 239686
rect 400224 239672 400286 239700
rect 400608 239672 400862 239700
rect 400992 239672 401246 239700
rect 399860 235570 399916 235579
rect 399860 235505 399916 235514
rect 399574 235013 399626 235019
rect 399574 234955 399626 234961
rect 399586 232799 399614 234955
rect 400054 234273 400106 234279
rect 400054 234215 400106 234221
rect 399574 232793 399626 232799
rect 399574 232735 399626 232741
rect 399476 228910 399532 228919
rect 399476 228845 399532 228854
rect 399382 226873 399434 226879
rect 399382 226815 399434 226821
rect 398902 226503 398954 226509
rect 398902 226445 398954 226451
rect 398998 226281 399050 226287
rect 398998 226223 399050 226229
rect 399010 226065 399038 226223
rect 398710 226059 398762 226065
rect 398710 226001 398762 226007
rect 398806 226059 398858 226065
rect 398806 226001 398858 226007
rect 398998 226059 399050 226065
rect 398998 226001 399050 226007
rect 398626 225917 398942 225936
rect 398614 225911 398954 225917
rect 398666 225908 398902 225911
rect 398614 225853 398666 225859
rect 398902 225853 398954 225859
rect 399958 225171 400010 225177
rect 399958 225113 400010 225119
rect 399094 222285 399146 222291
rect 399094 222227 399146 222233
rect 398338 221764 398414 221792
rect 398386 221482 398414 221764
rect 399106 221482 399134 222227
rect 399970 221482 399998 225113
rect 400066 222703 400094 234215
rect 400150 234199 400202 234205
rect 400150 234141 400202 234147
rect 400162 231393 400190 234141
rect 400258 233317 400286 239672
rect 400438 239305 400490 239311
rect 400438 239247 400490 239253
rect 400342 236641 400394 236647
rect 400342 236583 400394 236589
rect 400354 233687 400382 236583
rect 400450 236023 400478 239247
rect 400436 236014 400492 236023
rect 400436 235949 400492 235958
rect 400342 233681 400394 233687
rect 400342 233623 400394 233629
rect 400246 233311 400298 233317
rect 400246 233253 400298 233259
rect 400150 231387 400202 231393
rect 400150 231329 400202 231335
rect 400834 226731 400862 239672
rect 400822 226725 400874 226731
rect 400822 226667 400874 226673
rect 401218 226583 401246 239672
rect 401410 235431 401438 239686
rect 401396 235422 401452 235431
rect 401396 235357 401452 235366
rect 401794 234205 401822 239686
rect 401782 234199 401834 234205
rect 401782 234141 401834 234147
rect 401398 231017 401450 231023
rect 401398 230959 401450 230965
rect 401206 226577 401258 226583
rect 401206 226519 401258 226525
rect 400630 224727 400682 224733
rect 400630 224669 400682 224675
rect 400052 222694 400108 222703
rect 400052 222629 400108 222638
rect 400642 221792 400670 224669
rect 400642 221764 400718 221792
rect 400690 221482 400718 221764
rect 401410 221482 401438 230959
rect 402178 226509 402206 239686
rect 402528 239672 402686 239700
rect 402548 235274 402604 235283
rect 402548 235209 402604 235218
rect 402562 231467 402590 235209
rect 402550 231461 402602 231467
rect 402550 231403 402602 231409
rect 402166 226503 402218 226509
rect 402166 226445 402218 226451
rect 402658 226403 402686 239672
rect 402754 239672 402912 239700
rect 403248 239672 403550 239700
rect 402754 235283 402782 239672
rect 403414 238417 403466 238423
rect 403414 238359 403466 238365
rect 403426 237979 403454 238359
rect 403522 237979 403550 239672
rect 403414 237973 403466 237979
rect 403414 237915 403466 237921
rect 403510 237973 403562 237979
rect 403510 237915 403562 237921
rect 403618 235833 403646 239686
rect 403702 237973 403754 237979
rect 403702 237915 403754 237921
rect 403606 235827 403658 235833
rect 403606 235769 403658 235775
rect 402740 235274 402796 235283
rect 402740 235209 402796 235218
rect 403412 234978 403468 234987
rect 403412 234913 403468 234922
rect 402838 226429 402890 226435
rect 402644 226394 402700 226403
rect 402838 226371 402890 226377
rect 402644 226329 402700 226338
rect 402166 224875 402218 224881
rect 402166 224817 402218 224823
rect 402178 221482 402206 224817
rect 402850 221792 402878 226371
rect 403426 222555 403454 234913
rect 403714 234279 403742 237915
rect 404002 236171 404030 239686
rect 403988 236162 404044 236171
rect 403988 236097 404044 236106
rect 403702 234273 403754 234279
rect 403702 234215 403754 234221
rect 403702 227613 403754 227619
rect 403702 227555 403754 227561
rect 403412 222546 403468 222555
rect 403412 222481 403468 222490
rect 402850 221764 402926 221792
rect 402898 221482 402926 221764
rect 403714 221482 403742 227555
rect 404386 226361 404414 239686
rect 404736 239672 404990 239700
rect 405216 239672 405470 239700
rect 404662 233829 404714 233835
rect 404662 233771 404714 233777
rect 404674 228655 404702 233771
rect 404662 228649 404714 228655
rect 404662 228591 404714 228597
rect 404962 226435 404990 239672
rect 405442 236023 405470 239672
rect 405428 236014 405484 236023
rect 405428 235949 405484 235958
rect 405538 234691 405566 239686
rect 405826 239672 405936 239700
rect 405332 234682 405388 234691
rect 405524 234682 405580 234691
rect 405388 234640 405470 234668
rect 405332 234617 405388 234626
rect 405238 234051 405290 234057
rect 405238 233993 405290 233999
rect 405250 231879 405278 233993
rect 405236 231870 405292 231879
rect 405236 231805 405292 231814
rect 405442 227534 405470 234640
rect 405524 234617 405580 234626
rect 405442 227506 405758 227534
rect 404950 226429 405002 226435
rect 404950 226371 405002 226377
rect 404374 226355 404426 226361
rect 404374 226297 404426 226303
rect 404470 226281 404522 226287
rect 404470 226223 404522 226229
rect 404482 221482 404510 226223
rect 405142 225023 405194 225029
rect 405142 224965 405194 224971
rect 405154 221792 405182 224965
rect 405730 224160 405758 227506
rect 405826 226107 405854 239672
rect 406198 239379 406250 239385
rect 406198 239321 406250 239327
rect 405910 236937 405962 236943
rect 405910 236879 405962 236885
rect 405922 234543 405950 236879
rect 406210 236129 406238 239321
rect 406306 236129 406334 239686
rect 406198 236123 406250 236129
rect 406198 236065 406250 236071
rect 406294 236123 406346 236129
rect 406294 236065 406346 236071
rect 406690 235019 406718 239686
rect 407040 239672 407294 239700
rect 407424 239672 407678 239700
rect 406774 237011 406826 237017
rect 406774 236953 406826 236959
rect 406786 236174 406814 236953
rect 406786 236146 407198 236174
rect 406678 235013 406730 235019
rect 406678 234955 406730 234961
rect 405908 234534 405964 234543
rect 405908 234469 405964 234478
rect 406774 229759 406826 229765
rect 406774 229701 406826 229707
rect 405812 226098 405868 226107
rect 405812 226033 405868 226042
rect 405730 224132 405950 224160
rect 405154 221764 405230 221792
rect 405202 221482 405230 221764
rect 405922 221482 405950 224132
rect 406786 221482 406814 229701
rect 407170 227534 407198 236146
rect 407266 234099 407294 239672
rect 407446 237973 407498 237979
rect 407446 237915 407498 237921
rect 407458 236869 407486 237915
rect 407446 236863 407498 236869
rect 407446 236805 407498 236811
rect 407650 236174 407678 239672
rect 407554 236146 407678 236174
rect 407444 234830 407500 234839
rect 407444 234765 407500 234774
rect 407252 234090 407308 234099
rect 407252 234025 407308 234034
rect 407458 228507 407486 234765
rect 407446 228501 407498 228507
rect 407446 228443 407498 228449
rect 407170 227506 407486 227534
rect 407458 221792 407486 227506
rect 407554 226255 407582 236146
rect 407638 233755 407690 233761
rect 407638 233697 407690 233703
rect 407650 230251 407678 233697
rect 407636 230242 407692 230251
rect 407636 230177 407692 230186
rect 407746 226287 407774 239686
rect 408130 235135 408158 239686
rect 408116 235126 408172 235135
rect 408116 235061 408172 235070
rect 408514 234987 408542 239686
rect 408960 239672 409214 239700
rect 409728 239672 409982 239700
rect 408790 237011 408842 237017
rect 408790 236953 408842 236959
rect 408500 234978 408556 234987
rect 408500 234913 408556 234922
rect 408802 233655 408830 236953
rect 409186 234945 409214 239672
rect 409174 234939 409226 234945
rect 409174 234881 409226 234887
rect 409954 234839 409982 239672
rect 409940 234830 409996 234839
rect 410050 234797 410078 239686
rect 409940 234765 409996 234774
rect 410038 234791 410090 234797
rect 410038 234733 410090 234739
rect 408788 233646 408844 233655
rect 408788 233581 408844 233590
rect 409654 230795 409706 230801
rect 409654 230737 409706 230743
rect 407734 226281 407786 226287
rect 407540 226246 407596 226255
rect 407734 226223 407786 226229
rect 407540 226181 407596 226190
rect 408982 226207 409034 226213
rect 408982 226149 409034 226155
rect 408214 225097 408266 225103
rect 408214 225039 408266 225045
rect 407458 221764 407534 221792
rect 407506 221482 407534 221764
rect 408226 221482 408254 225039
rect 408994 221482 409022 226149
rect 409666 221792 409694 230737
rect 410434 225177 410462 239686
rect 410818 234871 410846 239686
rect 411168 239672 411326 239700
rect 411552 239672 411710 239700
rect 411936 239672 412190 239700
rect 411190 237159 411242 237165
rect 411190 237101 411242 237107
rect 411202 236869 411230 237101
rect 411190 236863 411242 236869
rect 411190 236805 411242 236811
rect 410806 234865 410858 234871
rect 410806 234807 410858 234813
rect 411298 234691 411326 239672
rect 411574 239453 411626 239459
rect 411394 239401 411574 239404
rect 411394 239395 411626 239401
rect 411394 239376 411614 239395
rect 411394 239311 411422 239376
rect 411382 239305 411434 239311
rect 411382 239247 411434 239253
rect 411478 239305 411530 239311
rect 411478 239247 411530 239253
rect 411382 237085 411434 237091
rect 411380 237050 411382 237059
rect 411434 237050 411436 237059
rect 411380 236985 411436 236994
rect 411490 236055 411518 239247
rect 411572 237050 411628 237059
rect 411572 236985 411628 236994
rect 411586 236319 411614 236985
rect 411572 236310 411628 236319
rect 411572 236245 411628 236254
rect 411478 236049 411530 236055
rect 411478 235991 411530 235997
rect 411574 234717 411626 234723
rect 411284 234682 411340 234691
rect 411574 234659 411626 234665
rect 411284 234617 411340 234626
rect 411476 233942 411532 233951
rect 411476 233877 411532 233886
rect 410518 230647 410570 230653
rect 410518 230589 410570 230595
rect 410422 225171 410474 225177
rect 410422 225113 410474 225119
rect 409666 221764 409742 221792
rect 409714 221482 409742 221764
rect 410530 221482 410558 230589
rect 411490 229765 411518 233877
rect 411586 231023 411614 234659
rect 411574 231017 411626 231023
rect 411574 230959 411626 230965
rect 411478 229759 411530 229765
rect 411478 229701 411530 229707
rect 411682 226139 411710 239672
rect 412054 236493 412106 236499
rect 412054 236435 412106 236441
rect 411764 236310 411820 236319
rect 411764 236245 411820 236254
rect 411778 236129 411806 236245
rect 411766 236123 411818 236129
rect 411766 236065 411818 236071
rect 411764 233794 411820 233803
rect 411764 233729 411820 233738
rect 411778 232947 411806 233729
rect 412066 233391 412094 236435
rect 412162 234723 412190 239672
rect 412258 239311 412286 240241
rect 420322 239311 420350 241129
rect 581780 240306 581836 240315
rect 581780 240241 581836 240250
rect 567380 240010 567436 240019
rect 567380 239945 567436 239954
rect 434614 239823 434666 239829
rect 434614 239765 434666 239771
rect 412246 239305 412298 239311
rect 412246 239247 412298 239253
rect 420310 239305 420362 239311
rect 420310 239247 420362 239253
rect 414646 239009 414698 239015
rect 413396 238974 413452 238983
rect 414646 238951 414698 238957
rect 413396 238909 413452 238918
rect 413410 236573 413438 238909
rect 414658 238835 414686 238951
rect 414644 238826 414700 238835
rect 414644 238761 414700 238770
rect 413684 238678 413740 238687
rect 413684 238613 413740 238622
rect 413698 236721 413726 238613
rect 413972 238382 414028 238391
rect 413972 238317 414028 238326
rect 413986 237091 414014 238317
rect 414260 238234 414316 238243
rect 414260 238169 414316 238178
rect 413974 237085 414026 237091
rect 413974 237027 414026 237033
rect 414274 237017 414302 238169
rect 414452 238086 414508 238095
rect 414452 238021 414508 238030
rect 414262 237011 414314 237017
rect 414262 236953 414314 236959
rect 414466 236943 414494 238021
rect 432406 237307 432458 237313
rect 432406 237249 432458 237255
rect 426358 237233 426410 237239
rect 419156 237198 419212 237207
rect 426358 237175 426410 237181
rect 419156 237133 419212 237142
rect 420310 237159 420362 237165
rect 414454 236937 414506 236943
rect 419170 236911 419198 237133
rect 420310 237101 420362 237107
rect 414454 236879 414506 236885
rect 419156 236902 419212 236911
rect 419156 236837 419212 236846
rect 413686 236715 413738 236721
rect 413686 236657 413738 236663
rect 413398 236567 413450 236573
rect 413398 236509 413450 236515
rect 412726 236419 412778 236425
rect 412726 236361 412778 236367
rect 412150 234717 412202 234723
rect 412150 234659 412202 234665
rect 412738 233465 412766 236361
rect 418294 234347 418346 234353
rect 418294 234289 418346 234295
rect 412726 233459 412778 233465
rect 412726 233401 412778 233407
rect 412054 233385 412106 233391
rect 412054 233327 412106 233333
rect 411766 232941 411818 232947
rect 411766 232883 411818 232889
rect 415702 231239 415754 231245
rect 415702 231181 415754 231187
rect 413494 228575 413546 228581
rect 413494 228517 413546 228523
rect 412726 228131 412778 228137
rect 412726 228073 412778 228079
rect 411286 226133 411338 226139
rect 411286 226075 411338 226081
rect 411670 226133 411722 226139
rect 411670 226075 411722 226081
rect 411298 221496 411326 226075
rect 411958 225319 412010 225325
rect 411958 225261 412010 225267
rect 411264 221468 411326 221496
rect 411970 221496 411998 225261
rect 411970 221468 412032 221496
rect 412738 221482 412766 228073
rect 413506 221496 413534 228517
rect 415030 225393 415082 225399
rect 415030 225335 415082 225341
rect 414262 222655 414314 222661
rect 414262 222597 414314 222603
rect 413472 221468 413534 221496
rect 414274 221482 414302 222597
rect 415042 221482 415070 225335
rect 415714 221792 415742 231181
rect 418306 227619 418334 234289
rect 419254 231091 419306 231097
rect 419254 231033 419306 231039
rect 418774 228797 418826 228803
rect 418774 228739 418826 228745
rect 418294 227613 418346 227619
rect 418294 227555 418346 227561
rect 418678 226651 418730 226657
rect 418678 226593 418730 226599
rect 418690 226213 418718 226593
rect 418678 226207 418730 226213
rect 418678 226149 418730 226155
rect 418006 225245 418058 225251
rect 418006 225187 418058 225193
rect 417238 222729 417290 222735
rect 417238 222671 417290 222677
rect 416470 222581 416522 222587
rect 416470 222523 416522 222529
rect 415714 221764 415790 221792
rect 415762 221482 415790 221764
rect 416482 221482 416510 222523
rect 417250 221482 417278 222671
rect 418018 221792 418046 225187
rect 418018 221764 418094 221792
rect 418066 221482 418094 221764
rect 418786 221482 418814 228739
rect 419266 221774 419294 231033
rect 419362 226944 419678 226972
rect 419362 226879 419390 226944
rect 419350 226873 419402 226879
rect 419350 226815 419402 226821
rect 419446 226873 419498 226879
rect 419446 226815 419498 226821
rect 419458 226213 419486 226815
rect 419650 226731 419678 226944
rect 419638 226725 419690 226731
rect 419638 226667 419690 226673
rect 419446 226207 419498 226213
rect 419446 226149 419498 226155
rect 420322 221792 420350 237101
rect 423382 234421 423434 234427
rect 423382 234363 423434 234369
rect 423394 230505 423422 234363
rect 424724 231130 424780 231139
rect 424724 231065 424780 231074
rect 424054 231017 424106 231023
rect 424054 230959 424106 230965
rect 423382 230499 423434 230505
rect 423382 230441 423434 230447
rect 421846 228723 421898 228729
rect 421846 228665 421898 228671
rect 420982 225467 421034 225473
rect 420982 225409 421034 225415
rect 419266 221746 419582 221774
rect 419554 221482 419582 221746
rect 420274 221764 420350 221792
rect 420274 221482 420302 221764
rect 420994 221482 421022 225409
rect 421858 221482 421886 228665
rect 422518 222951 422570 222957
rect 422518 222893 422570 222899
rect 422530 221792 422558 222893
rect 423286 222803 423338 222809
rect 423286 222745 423338 222751
rect 422530 221764 422606 221792
rect 422578 221482 422606 221764
rect 423298 221482 423326 222745
rect 424066 221482 424094 230959
rect 424738 221792 424766 231065
rect 425590 228057 425642 228063
rect 425590 227999 425642 228005
rect 424738 221764 424814 221792
rect 424786 221482 424814 221764
rect 425602 221482 425630 227999
rect 426370 221482 426398 237175
rect 428662 236863 428714 236869
rect 428662 236805 428714 236811
rect 427894 233903 427946 233909
rect 427894 233845 427946 233851
rect 427906 228951 427934 233845
rect 427798 228945 427850 228951
rect 427798 228887 427850 228893
rect 427894 228945 427946 228951
rect 427894 228887 427946 228893
rect 427030 225541 427082 225547
rect 427030 225483 427082 225489
rect 427042 221792 427070 225483
rect 427042 221764 427118 221792
rect 427090 221482 427118 221764
rect 427810 221482 427838 228887
rect 428674 221482 428702 236805
rect 430102 236493 430154 236499
rect 430102 236435 430154 236441
rect 429334 223025 429386 223031
rect 429334 222967 429386 222973
rect 429346 221792 429374 222967
rect 429346 221764 429422 221792
rect 429394 221482 429422 221764
rect 430114 221482 430142 236435
rect 432022 233977 432074 233983
rect 432022 233919 432074 233925
rect 432034 228877 432062 233919
rect 430870 228871 430922 228877
rect 430870 228813 430922 228819
rect 432022 228871 432074 228877
rect 432022 228813 432074 228819
rect 430882 221482 430910 228813
rect 431542 222877 431594 222883
rect 431542 222819 431594 222825
rect 431554 221792 431582 222819
rect 431554 221764 431630 221792
rect 431602 221482 431630 221764
rect 432418 221482 432446 237249
rect 433846 231535 433898 231541
rect 433846 231477 433898 231483
rect 433174 227613 433226 227619
rect 433174 227555 433226 227561
rect 433186 221482 433214 227555
rect 433858 221792 433886 231477
rect 433858 221764 433934 221792
rect 433906 221482 433934 221764
rect 434626 221482 434654 239765
rect 446710 239749 446762 239755
rect 446710 239691 446762 239697
rect 444502 237529 444554 237535
rect 444502 237471 444554 237477
rect 441430 237455 441482 237461
rect 441430 237397 441482 237403
rect 438358 237381 438410 237387
rect 438358 237323 438410 237329
rect 434902 234495 434954 234501
rect 434902 234437 434954 234443
rect 434914 228803 434942 234437
rect 436150 230499 436202 230505
rect 436150 230441 436202 230447
rect 434902 228797 434954 228803
rect 434902 228739 434954 228745
rect 435382 223099 435434 223105
rect 435382 223041 435434 223047
rect 435394 221482 435422 223041
rect 436162 221792 436190 230441
rect 437686 228205 437738 228211
rect 436916 228170 436972 228179
rect 437686 228147 437738 228153
rect 436916 228105 436972 228114
rect 436162 221764 436238 221792
rect 436210 221482 436238 221764
rect 436930 221482 436958 228105
rect 437698 221482 437726 228147
rect 438370 221792 438398 237323
rect 441442 236174 441470 237397
rect 442198 236419 442250 236425
rect 442198 236361 442250 236367
rect 440770 236146 441470 236174
rect 439990 230425 440042 230431
rect 439990 230367 440042 230373
rect 439126 225615 439178 225621
rect 439126 225557 439178 225563
rect 438370 221764 438446 221792
rect 438418 221482 438446 221764
rect 439138 221482 439166 225557
rect 440002 221496 440030 230367
rect 440770 221792 440798 236146
rect 441430 224653 441482 224659
rect 441430 224595 441482 224601
rect 439968 221468 440030 221496
rect 440722 221764 440798 221792
rect 440722 221482 440750 221764
rect 441442 221482 441470 224595
rect 442210 221496 442238 236361
rect 442868 231278 442924 231287
rect 442868 231213 442924 231222
rect 442176 221468 442238 221496
rect 442882 221496 442910 231213
rect 443734 223173 443786 223179
rect 443734 223115 443786 223121
rect 442882 221468 442944 221496
rect 443746 221482 443774 223115
rect 444514 221792 444542 237471
rect 445942 230351 445994 230357
rect 445942 230293 445994 230299
rect 445172 225210 445228 225219
rect 445172 225145 445228 225154
rect 444466 221764 444542 221792
rect 444466 221482 444494 221764
rect 445186 221482 445214 225145
rect 445954 221482 445982 230293
rect 446722 221792 446750 239691
rect 458806 239675 458858 239681
rect 458806 239617 458858 239623
rect 455158 238935 455210 238941
rect 455158 238877 455210 238883
rect 455062 238861 455114 238867
rect 455062 238803 455114 238809
rect 450454 236789 450506 236795
rect 450454 236731 450506 236737
rect 448246 234643 448298 234649
rect 448246 234585 448298 234591
rect 447478 224505 447530 224511
rect 447478 224447 447530 224453
rect 446674 221764 446750 221792
rect 446674 221482 446702 221764
rect 447490 221482 447518 224447
rect 448258 221482 448286 234585
rect 449302 234569 449354 234575
rect 449302 234511 449354 234517
rect 448918 231609 448970 231615
rect 448918 231551 448970 231557
rect 448930 221792 448958 231551
rect 449314 230357 449342 234511
rect 449686 230869 449738 230875
rect 449686 230811 449738 230817
rect 449302 230351 449354 230357
rect 449302 230293 449354 230299
rect 448930 221764 449006 221792
rect 448978 221482 449006 221764
rect 449698 221482 449726 230811
rect 450466 221482 450494 236731
rect 451990 230277 452042 230283
rect 451990 230219 452042 230225
rect 451222 225689 451274 225695
rect 451222 225631 451274 225637
rect 451234 221792 451262 225631
rect 451234 221764 451310 221792
rect 451282 221482 451310 221764
rect 452002 221482 452030 230219
rect 454294 228797 454346 228803
rect 454294 228739 454346 228745
rect 452758 224579 452810 224585
rect 452758 224521 452810 224527
rect 452770 221482 452798 224521
rect 453430 224431 453482 224437
rect 453430 224373 453482 224379
rect 453442 221792 453470 224373
rect 453442 221764 453518 221792
rect 453490 221482 453518 221764
rect 454306 221482 454334 228739
rect 455074 228581 455102 238803
rect 455170 236174 455198 238877
rect 455170 236146 455774 236174
rect 455156 231426 455212 231435
rect 455156 231361 455212 231370
rect 455062 228575 455114 228581
rect 455062 228517 455114 228523
rect 455170 226084 455198 231361
rect 455074 226056 455198 226084
rect 455074 221482 455102 226056
rect 455746 221792 455774 236146
rect 458038 230129 458090 230135
rect 458038 230071 458090 230077
rect 456502 228575 456554 228581
rect 456502 228517 456554 228523
rect 455746 221764 455822 221792
rect 455794 221482 455822 221764
rect 456514 221482 456542 228517
rect 457268 225358 457324 225367
rect 457268 225293 457324 225302
rect 457282 221482 457310 225293
rect 458050 221792 458078 230071
rect 458050 221764 458126 221792
rect 458098 221482 458126 221764
rect 458818 221482 458846 239617
rect 470902 239601 470954 239607
rect 470902 239543 470954 239549
rect 462550 238787 462602 238793
rect 462550 238729 462602 238735
rect 460246 233533 460298 233539
rect 460246 233475 460298 233481
rect 459574 224357 459626 224363
rect 459574 224299 459626 224305
rect 459586 221482 459614 224299
rect 460258 221792 460286 233475
rect 461014 230203 461066 230209
rect 461014 230145 461066 230151
rect 460258 221764 460334 221792
rect 460306 221482 460334 221764
rect 461026 221482 461054 230145
rect 461878 228279 461930 228285
rect 461878 228221 461930 228227
rect 461890 221482 461918 228221
rect 462562 221792 462590 238729
rect 464758 238713 464810 238719
rect 464758 238655 464810 238661
rect 463606 233607 463658 233613
rect 463606 233549 463658 233555
rect 463618 230209 463646 233549
rect 464084 231574 464140 231583
rect 464084 231509 464140 231518
rect 463606 230203 463658 230209
rect 463606 230145 463658 230151
rect 463316 225654 463372 225663
rect 463316 225589 463372 225598
rect 462562 221764 462638 221792
rect 462610 221482 462638 221764
rect 463330 221482 463358 225589
rect 464098 221482 464126 231509
rect 464770 221792 464798 238655
rect 468598 238639 468650 238645
rect 468598 238581 468650 238587
rect 466484 234238 466540 234247
rect 466484 234173 466540 234182
rect 466390 230351 466442 230357
rect 466390 230293 466442 230299
rect 465622 224283 465674 224289
rect 465622 224225 465674 224231
rect 464770 221764 464846 221792
rect 464818 221482 464846 221764
rect 465634 221482 465662 224225
rect 466402 221482 466430 230293
rect 466498 230135 466526 234173
rect 466486 230129 466538 230135
rect 466486 230071 466538 230077
rect 467062 228427 467114 228433
rect 467062 228369 467114 228375
rect 467074 221792 467102 228369
rect 467830 222433 467882 222439
rect 467830 222375 467882 222381
rect 467074 221764 467150 221792
rect 467122 221482 467150 221764
rect 467842 221482 467870 222375
rect 468610 221482 468638 238581
rect 470132 231722 470188 231731
rect 470132 231657 470188 231666
rect 469364 225802 469420 225811
rect 469364 225737 469420 225746
rect 469378 221496 469406 225737
rect 469378 221468 469440 221496
rect 470146 221482 470174 231657
rect 470914 221496 470942 239543
rect 532822 239527 532874 239533
rect 532822 239469 532874 239475
rect 488278 239231 488330 239237
rect 488278 239173 488330 239179
rect 474646 238565 474698 238571
rect 474646 238507 474698 238513
rect 472342 235975 472394 235981
rect 472342 235917 472394 235923
rect 471574 224209 471626 224215
rect 471574 224151 471626 224157
rect 470880 221468 470942 221496
rect 471586 221496 471614 224151
rect 471586 221468 471648 221496
rect 472354 221482 472382 235917
rect 473878 231165 473930 231171
rect 473878 231107 473930 231113
rect 473110 229981 473162 229987
rect 473110 229923 473162 229929
rect 473122 221792 473150 229923
rect 473122 221764 473198 221792
rect 473170 221482 473198 221764
rect 473890 221482 473918 231107
rect 474658 221482 474686 238507
rect 478198 238491 478250 238497
rect 478198 238433 478250 238439
rect 475222 234125 475274 234131
rect 475222 234067 475274 234073
rect 475234 230061 475262 234067
rect 475222 230055 475274 230061
rect 475222 229997 475274 230003
rect 478210 228581 478238 238433
rect 478390 238417 478442 238423
rect 478390 238359 478442 238365
rect 478294 230203 478346 230209
rect 478294 230145 478346 230151
rect 478198 228575 478250 228581
rect 478198 228517 478250 228523
rect 476950 228353 477002 228359
rect 476180 228318 476236 228327
rect 476950 228295 477002 228301
rect 476180 228253 476236 228262
rect 475316 225950 475372 225959
rect 475316 225885 475372 225894
rect 475330 221792 475358 225885
rect 475330 221764 475406 221792
rect 475378 221482 475406 221764
rect 476194 221482 476222 228253
rect 476962 221482 476990 228295
rect 477622 224135 477674 224141
rect 477622 224077 477674 224083
rect 477634 221792 477662 224077
rect 478306 223568 478334 230145
rect 478402 227534 478430 238359
rect 486742 238343 486794 238349
rect 486742 238285 486794 238291
rect 484630 234199 484682 234205
rect 484630 234141 484682 234147
rect 479158 233311 479210 233317
rect 479158 233253 479210 233259
rect 479060 233202 479116 233211
rect 479060 233137 479116 233146
rect 479074 227534 479102 233137
rect 479170 229987 479198 233253
rect 484438 230129 484490 230135
rect 484438 230071 484490 230077
rect 479158 229981 479210 229987
rect 479158 229923 479210 229929
rect 482134 229907 482186 229913
rect 482134 229849 482186 229855
rect 480694 228575 480746 228581
rect 480694 228517 480746 228523
rect 478402 227506 478526 227534
rect 479074 227506 479198 227534
rect 478306 223540 478430 223568
rect 477634 221764 477710 221792
rect 477682 221482 477710 221764
rect 478402 221482 478430 223540
rect 478498 221773 478526 227506
rect 478486 221767 478538 221773
rect 478486 221709 478538 221715
rect 479170 221482 479198 227506
rect 479974 221767 480026 221773
rect 479974 221709 480026 221715
rect 479986 221482 480014 221709
rect 480706 221482 480734 228517
rect 481460 227430 481516 227439
rect 481460 227365 481516 227374
rect 481474 221482 481502 227365
rect 482146 221792 482174 229849
rect 483766 224061 483818 224067
rect 483766 224003 483818 224009
rect 482902 222359 482954 222365
rect 482902 222301 482954 222307
rect 482146 221764 482222 221792
rect 482194 221482 482222 221764
rect 482914 221482 482942 222301
rect 483778 221482 483806 224003
rect 484450 221792 484478 230071
rect 484642 229913 484670 234141
rect 485206 231683 485258 231689
rect 485206 231625 485258 231631
rect 484630 229907 484682 229913
rect 484630 229849 484682 229855
rect 484450 221764 484526 221792
rect 484498 221482 484526 221764
rect 485218 221482 485246 231625
rect 485974 231313 486026 231319
rect 485974 231255 486026 231261
rect 485986 221482 486014 231255
rect 486754 221792 486782 238285
rect 488290 236174 488318 239173
rect 508630 239157 508682 239163
rect 508630 239099 508682 239105
rect 492790 238269 492842 238275
rect 492790 238211 492842 238217
rect 492022 236345 492074 236351
rect 492022 236287 492074 236293
rect 488290 236146 488990 236174
rect 488276 228466 488332 228475
rect 488276 228401 488332 228410
rect 487508 225506 487564 225515
rect 487508 225441 487564 225450
rect 486706 221764 486782 221792
rect 486706 221482 486734 221764
rect 487522 221482 487550 225441
rect 488290 221482 488318 228401
rect 488962 221792 488990 236146
rect 490484 234386 490540 234395
rect 490484 234321 490540 234330
rect 489718 223987 489770 223993
rect 489718 223929 489770 223935
rect 488962 221764 489038 221792
rect 489010 221482 489038 221764
rect 489730 221482 489758 223929
rect 490498 221482 490526 234321
rect 491254 233237 491306 233243
rect 491254 233179 491306 233185
rect 491266 221792 491294 233179
rect 491266 221764 491342 221792
rect 491314 221482 491342 221764
rect 492034 221482 492062 236287
rect 492802 221482 492830 238211
rect 500278 238195 500330 238201
rect 500278 238137 500330 238143
rect 495766 235901 495818 235907
rect 495766 235843 495818 235849
rect 495094 231757 495146 231763
rect 495094 231699 495146 231705
rect 494228 228762 494284 228771
rect 494228 228697 494284 228706
rect 493460 227282 493516 227291
rect 493460 227217 493516 227226
rect 493474 221792 493502 227217
rect 493474 221764 493550 221792
rect 493522 221482 493550 221764
rect 494242 221482 494270 228697
rect 495106 221482 495134 231699
rect 495778 221792 495806 235843
rect 499606 231387 499658 231393
rect 499606 231329 499658 231335
rect 497972 228614 498028 228623
rect 497972 228549 498028 228558
rect 497302 223913 497354 223919
rect 497302 223855 497354 223861
rect 496534 222507 496586 222513
rect 496534 222449 496586 222455
rect 495778 221764 495854 221792
rect 495826 221482 495854 221764
rect 496546 221482 496574 222449
rect 497314 221482 497342 223855
rect 497986 221792 498014 228549
rect 498836 227134 498892 227143
rect 498836 227069 498892 227078
rect 497986 221764 498062 221792
rect 498034 221482 498062 221764
rect 498850 221482 498878 227069
rect 499618 221496 499646 231329
rect 499584 221468 499646 221496
rect 500290 221496 500318 238137
rect 503350 238121 503402 238127
rect 503350 238063 503402 238069
rect 501046 234273 501098 234279
rect 501046 234215 501098 234221
rect 501058 233243 501086 234215
rect 501046 233237 501098 233243
rect 501046 233179 501098 233185
rect 501046 233089 501098 233095
rect 501046 233031 501098 233037
rect 500854 233015 500906 233021
rect 500854 232957 500906 232963
rect 500866 231763 500894 232957
rect 500854 231757 500906 231763
rect 500854 231699 500906 231705
rect 500290 221468 500352 221496
rect 501058 221482 501086 233031
rect 502582 228501 502634 228507
rect 502582 228443 502634 228449
rect 501814 223839 501866 223845
rect 501814 223781 501866 223787
rect 501826 221792 501854 223781
rect 501826 221764 501902 221792
rect 501874 221482 501902 221764
rect 502594 221482 502622 228443
rect 503362 221482 503390 238063
rect 505654 236271 505706 236277
rect 505654 236213 505706 236219
rect 504022 229833 504074 229839
rect 504022 229775 504074 229781
rect 504034 221792 504062 229775
rect 504790 223543 504842 223549
rect 504790 223485 504842 223491
rect 504034 221764 504110 221792
rect 504082 221482 504110 221764
rect 504802 221482 504830 223485
rect 505666 221482 505694 236213
rect 506804 234090 506860 234099
rect 506804 234025 506860 234034
rect 506818 229839 506846 234025
rect 507094 233015 507146 233021
rect 507094 232957 507146 232963
rect 506806 229833 506858 229839
rect 506806 229775 506858 229781
rect 506326 223765 506378 223771
rect 506326 223707 506378 223713
rect 506338 221792 506366 223707
rect 506338 221764 506414 221792
rect 506386 221482 506414 221764
rect 507106 221482 507134 232957
rect 507862 223691 507914 223697
rect 507862 223633 507914 223639
rect 507874 221482 507902 223633
rect 508642 221792 508670 239099
rect 509398 238047 509450 238053
rect 509398 237989 509450 237995
rect 508594 221764 508670 221792
rect 508594 221482 508622 221764
rect 509410 221482 509438 237989
rect 512758 237973 512810 237979
rect 512758 237915 512810 237921
rect 511606 236567 511658 236573
rect 511606 236509 511658 236515
rect 510166 229685 510218 229691
rect 510166 229627 510218 229633
rect 510178 221482 510206 229627
rect 510838 223469 510890 223475
rect 510838 223411 510890 223417
rect 510850 221792 510878 223411
rect 510850 221764 510926 221792
rect 510898 221482 510926 221764
rect 511618 221482 511646 236509
rect 512770 228581 512798 237915
rect 513910 237899 513962 237905
rect 513910 237841 513962 237847
rect 513142 231757 513194 231763
rect 513142 231699 513194 231705
rect 512758 228575 512810 228581
rect 512758 228517 512810 228523
rect 512374 223617 512426 223623
rect 512374 223559 512426 223565
rect 512386 221482 512414 223559
rect 513154 221792 513182 231699
rect 513154 221764 513230 221792
rect 513202 221482 513230 221764
rect 513814 221767 513866 221773
rect 513922 221755 513950 237841
rect 521494 237825 521546 237831
rect 521494 237767 521546 237773
rect 519190 232867 519242 232873
rect 519190 232809 519242 232815
rect 516118 229611 516170 229617
rect 516118 229553 516170 229559
rect 514678 228575 514730 228581
rect 514678 228517 514730 228523
rect 514006 223395 514058 223401
rect 514006 223337 514058 223343
rect 514018 221797 514046 223337
rect 513866 221727 513950 221755
rect 514004 221788 514060 221797
rect 514004 221723 514060 221732
rect 513814 221709 513866 221715
rect 513908 221658 513964 221667
rect 513908 221593 513964 221602
rect 513922 221482 513950 221593
rect 514690 221482 514718 228517
rect 515398 221767 515450 221773
rect 515398 221709 515450 221715
rect 515410 221482 515438 221709
rect 516130 221482 516158 229553
rect 517654 228649 517706 228655
rect 517654 228591 517706 228597
rect 516982 223247 517034 223253
rect 516982 223189 517034 223195
rect 516994 221482 517022 223189
rect 517666 221792 517694 228591
rect 518420 224470 518476 224479
rect 518420 224405 518476 224414
rect 517666 221764 517742 221792
rect 517714 221482 517742 221764
rect 518434 221482 518462 224405
rect 519202 221482 519230 232809
rect 520726 231461 520778 231467
rect 520726 231403 520778 231409
rect 519862 223321 519914 223327
rect 519862 223263 519914 223269
rect 519874 221792 519902 223263
rect 519874 221764 519950 221792
rect 519922 221482 519950 221764
rect 520738 221482 520766 231403
rect 521506 221482 521534 237767
rect 526006 237751 526058 237757
rect 526006 237693 526058 237699
rect 525236 233054 525292 233063
rect 525236 232989 525292 232998
rect 522166 229537 522218 229543
rect 522166 229479 522218 229485
rect 522178 221792 522206 229479
rect 524468 222990 524524 222999
rect 524468 222925 524524 222934
rect 523796 222694 523852 222703
rect 523796 222629 523852 222638
rect 522932 222546 522988 222555
rect 522932 222481 522988 222490
rect 522178 221764 522254 221792
rect 522226 221482 522254 221764
rect 522946 221482 522974 222481
rect 523810 221482 523838 222629
rect 524482 221792 524510 222925
rect 524482 221764 524558 221792
rect 524530 221482 524558 221764
rect 525250 221482 525278 232989
rect 526018 221482 526046 237693
rect 531286 232719 531338 232725
rect 531286 232661 531338 232667
rect 528308 230390 528364 230399
rect 528308 230325 528364 230334
rect 527540 229946 527596 229955
rect 527540 229881 527596 229890
rect 526676 224618 526732 224627
rect 526676 224553 526732 224562
rect 526690 221792 526718 224553
rect 526690 221764 526766 221792
rect 526738 221482 526766 221764
rect 527554 221482 527582 229881
rect 528322 221496 528350 230325
rect 529750 228871 529802 228877
rect 529750 228813 529802 228819
rect 528980 224174 529036 224183
rect 528980 224109 529036 224118
rect 528288 221468 528350 221496
rect 528994 221496 529022 224109
rect 528994 221468 529056 221496
rect 529762 221482 529790 228813
rect 530516 224322 530572 224331
rect 530516 224257 530572 224266
rect 530530 221496 530558 224257
rect 530496 221468 530558 221496
rect 531298 221482 531326 232661
rect 532052 222842 532108 222851
rect 532052 222777 532108 222786
rect 532066 221482 532094 222777
rect 532834 221792 532862 239469
rect 541462 239453 541514 239459
rect 541462 239395 541514 239401
rect 533492 238382 533548 238391
rect 533492 238317 533548 238326
rect 532786 221764 532862 221792
rect 532786 221482 532814 221764
rect 533506 221482 533534 238317
rect 538004 238086 538060 238095
rect 538004 238021 538060 238030
rect 535126 237677 535178 237683
rect 535126 237619 535178 237625
rect 534260 230094 534316 230103
rect 534260 230029 534316 230038
rect 534274 221482 534302 230029
rect 535138 221792 535166 237619
rect 535798 237603 535850 237609
rect 535798 237545 535850 237551
rect 535810 228581 535838 237545
rect 538018 236174 538046 238021
rect 537922 236146 538046 236174
rect 541474 236174 541502 239395
rect 550870 239379 550922 239385
rect 550870 239321 550922 239327
rect 544822 239083 544874 239089
rect 544822 239025 544874 239031
rect 544340 238678 544396 238687
rect 544340 238613 544396 238622
rect 541474 236146 541790 236174
rect 537238 232645 537290 232651
rect 537238 232587 537290 232593
rect 535798 228575 535850 228581
rect 535798 228517 535850 228523
rect 535798 228427 535850 228433
rect 535798 228369 535850 228375
rect 535090 221764 535166 221792
rect 535090 221482 535118 221764
rect 535810 221482 535838 228369
rect 536564 224026 536620 224035
rect 536564 223961 536620 223970
rect 536578 221482 536606 223961
rect 537250 221792 537278 232587
rect 537922 228433 537950 236146
rect 539542 232497 539594 232503
rect 539542 232439 539594 232445
rect 538870 229463 538922 229469
rect 538870 229405 538922 229411
rect 538006 228575 538058 228581
rect 538006 228517 538058 228523
rect 537910 228427 537962 228433
rect 537910 228369 537962 228375
rect 537250 221764 537326 221792
rect 537298 221482 537326 221764
rect 538018 221482 538046 228517
rect 538882 221482 538910 229405
rect 539554 221792 539582 232439
rect 540310 229389 540362 229395
rect 540310 229331 540362 229337
rect 539554 221764 539630 221792
rect 539602 221482 539630 221764
rect 540322 221482 540350 229331
rect 541076 223878 541132 223887
rect 541076 223813 541132 223822
rect 541090 221482 541118 223813
rect 541762 221792 541790 236146
rect 543382 232571 543434 232577
rect 543382 232513 543434 232519
rect 542614 232423 542666 232429
rect 542614 232365 542666 232371
rect 541762 221764 541838 221792
rect 541810 221482 541838 221764
rect 542626 221482 542654 232365
rect 543394 221482 543422 232513
rect 544354 228581 544382 238613
rect 544342 228575 544394 228581
rect 544342 228517 544394 228523
rect 544052 223730 544108 223739
rect 544052 223665 544108 223674
rect 544066 221792 544094 223665
rect 544066 221764 544142 221792
rect 544114 221482 544142 221764
rect 544834 221482 544862 239025
rect 550196 238974 550252 238983
rect 550196 238909 550252 238918
rect 549430 232349 549482 232355
rect 549430 232291 549482 232297
rect 548566 232275 548618 232281
rect 548566 232217 548618 232223
rect 545590 232201 545642 232207
rect 545590 232143 545642 232149
rect 545602 221482 545630 232143
rect 546358 229315 546410 229321
rect 546358 229257 546410 229263
rect 546370 221792 546398 229257
rect 547894 228945 547946 228951
rect 547894 228887 547946 228893
rect 547126 228575 547178 228581
rect 547126 228517 547178 228523
rect 546370 221764 546446 221792
rect 546418 221482 546446 221764
rect 547138 221482 547166 228517
rect 547906 221482 547934 228887
rect 548578 221792 548606 232217
rect 548578 221764 548654 221792
rect 548626 221482 548654 221764
rect 549442 221482 549470 232291
rect 550210 221482 550238 238909
rect 550882 221792 550910 239321
rect 559892 238234 559948 238243
rect 559892 238169 559948 238178
rect 559220 236754 559276 236763
rect 559220 236689 559276 236698
rect 557012 236606 557068 236615
rect 557012 236541 557068 236550
rect 553940 236458 553996 236467
rect 553940 236393 553996 236402
rect 553954 236174 553982 236393
rect 557026 236174 557054 236541
rect 553282 236146 553982 236174
rect 556162 236146 557054 236174
rect 551636 232906 551692 232915
rect 551636 232841 551692 232850
rect 550882 221764 550958 221792
rect 550930 221482 550958 221764
rect 551650 221482 551678 232841
rect 552406 232127 552458 232133
rect 552406 232069 552458 232075
rect 552418 221482 552446 232069
rect 553282 221792 553310 236146
rect 554710 232053 554762 232059
rect 554710 231995 554762 232001
rect 553940 229798 553996 229807
rect 553940 229733 553996 229742
rect 553234 221764 553310 221792
rect 553234 221482 553262 221764
rect 553954 221482 553982 229733
rect 554722 221482 554750 231995
rect 555382 229241 555434 229247
rect 555382 229183 555434 229189
rect 555394 221792 555422 229183
rect 555394 221764 555470 221792
rect 555442 221482 555470 221764
rect 556162 221482 556190 236146
rect 558454 231979 558506 231985
rect 558454 231921 558506 231927
rect 557014 231905 557066 231911
rect 557014 231847 557066 231853
rect 557026 221496 557054 231847
rect 557686 231831 557738 231837
rect 557686 231773 557738 231779
rect 556992 221468 557054 221496
rect 557698 221496 557726 231773
rect 557698 221468 557760 221496
rect 558466 221482 558494 231921
rect 559234 221496 559262 236689
rect 559200 221468 559262 221496
rect 559906 221496 559934 238169
rect 565268 237050 565324 237059
rect 565268 236985 565324 236994
rect 562196 236902 562252 236911
rect 562196 236837 562252 236846
rect 560756 232758 560812 232767
rect 560756 232693 560812 232702
rect 559906 221468 559968 221496
rect 560770 221482 560798 232693
rect 561430 229167 561482 229173
rect 561430 229109 561482 229115
rect 561442 221792 561470 229109
rect 561442 221764 561518 221792
rect 561490 221482 561518 221764
rect 562210 221482 562238 236837
rect 564500 232610 564556 232619
rect 564500 232545 564556 232554
rect 563636 229650 563692 229659
rect 563636 229585 563692 229594
rect 562964 223582 563020 223591
rect 562964 223517 563020 223526
rect 562978 221482 563006 223517
rect 563650 221792 563678 229585
rect 563650 221764 563726 221792
rect 563698 221482 563726 221764
rect 564514 221482 564542 232545
rect 565282 221482 565310 236985
rect 566710 232793 566762 232799
rect 566710 232735 566762 232741
rect 565942 229759 565994 229765
rect 565942 229701 565994 229707
rect 565954 221792 565982 229701
rect 565954 221764 566030 221792
rect 566002 221482 566030 221764
rect 566722 221482 566750 232735
rect 567394 228581 567422 239945
rect 573140 238826 573196 238835
rect 573140 238761 573196 238770
rect 573154 236174 573182 238761
rect 573154 236146 574334 236174
rect 572086 232941 572138 232947
rect 572086 232883 572138 232889
rect 570452 232462 570508 232471
rect 570452 232397 570508 232406
rect 567478 229093 567530 229099
rect 567478 229035 567530 229041
rect 567382 228575 567434 228581
rect 567382 228517 567434 228523
rect 567490 221482 567518 229035
rect 569782 229019 569834 229025
rect 569782 228961 569834 228967
rect 569014 228575 569066 228581
rect 569014 228517 569066 228523
rect 568244 223434 568300 223443
rect 568244 223369 568300 223378
rect 568258 221792 568286 223369
rect 568258 221764 568334 221792
rect 568306 221482 568334 221764
rect 569026 221482 569054 228517
rect 569794 221482 569822 228961
rect 570466 221792 570494 232397
rect 571316 223286 571372 223295
rect 571316 223221 571372 223230
rect 570466 221764 570542 221792
rect 570514 221482 570542 221764
rect 571330 221482 571358 223221
rect 572098 221482 572126 232883
rect 572756 229502 572812 229511
rect 572756 229437 572812 229446
rect 572770 221792 572798 229437
rect 573524 229354 573580 229363
rect 573524 229289 573580 229298
rect 572770 221764 572846 221792
rect 572818 221482 572846 221764
rect 573538 221482 573566 229289
rect 574306 221482 574334 236146
rect 580342 235679 580394 235685
rect 580342 235621 580394 235627
rect 576596 232314 576652 232323
rect 576596 232249 576652 232258
rect 575828 232018 575884 232027
rect 575828 231953 575884 231962
rect 575060 230242 575116 230251
rect 575060 230177 575116 230186
rect 575074 221792 575102 230177
rect 575074 221764 575150 221792
rect 575122 221482 575150 221764
rect 575842 221482 575870 231953
rect 576610 221482 576638 232249
rect 578036 232166 578092 232175
rect 578036 232101 578092 232110
rect 577268 223138 577324 223147
rect 577268 223073 577324 223082
rect 577282 221792 577310 223073
rect 577282 221764 577358 221792
rect 577330 221482 577358 221764
rect 578050 221482 578078 232101
rect 578900 229206 578956 229215
rect 578900 229141 578956 229150
rect 578914 221482 578942 229141
rect 579574 225985 579626 225991
rect 579574 225927 579626 225933
rect 579586 221792 579614 225927
rect 579586 221764 579662 221792
rect 579634 221482 579662 221764
rect 580354 221482 580382 235621
rect 581110 225837 581162 225843
rect 581110 225779 581162 225785
rect 581122 221482 581150 225779
rect 581794 221792 581822 240241
rect 599062 239305 599114 239311
rect 599062 239247 599114 239253
rect 587348 236162 587404 236171
rect 587348 236097 587404 236106
rect 587062 235753 587114 235759
rect 587062 235695 587114 235701
rect 586294 235605 586346 235611
rect 586294 235547 586346 235553
rect 583414 235531 583466 235537
rect 583414 235473 583466 235479
rect 582646 225911 582698 225917
rect 582646 225853 582698 225859
rect 581794 221764 581870 221792
rect 581842 221482 581870 221764
rect 582658 221482 582686 225853
rect 583426 221482 583454 235473
rect 585622 227243 585674 227249
rect 585622 227185 585674 227191
rect 584854 227169 584906 227175
rect 584854 227111 584906 227117
rect 584086 225763 584138 225769
rect 584086 225705 584138 225711
rect 584098 221792 584126 225705
rect 584098 221764 584174 221792
rect 584146 221482 584174 221764
rect 584866 221482 584894 227111
rect 585634 221482 585662 227185
rect 586306 224807 586334 235547
rect 586390 226059 586442 226065
rect 586390 226001 586442 226007
rect 586294 224801 586346 224807
rect 586294 224743 586346 224749
rect 586402 221496 586430 226001
rect 587074 225991 587102 235695
rect 587158 227539 587210 227545
rect 587158 227481 587210 227487
rect 587062 225985 587114 225991
rect 587062 225927 587114 225933
rect 586402 221468 586464 221496
rect 587170 221482 587198 227481
rect 587362 227249 587390 236097
rect 588980 236014 589036 236023
rect 588980 235949 589036 235958
rect 587828 235866 587884 235875
rect 587828 235801 587884 235810
rect 588886 235827 588938 235833
rect 587444 234534 587500 234543
rect 587444 234469 587500 234478
rect 587350 227243 587402 227249
rect 587350 227185 587402 227191
rect 587458 227175 587486 234469
rect 587446 227169 587498 227175
rect 587446 227111 587498 227117
rect 587842 226065 587870 235801
rect 588886 235769 588938 235775
rect 587926 235457 587978 235463
rect 587926 235399 587978 235405
rect 587830 226059 587882 226065
rect 587830 226001 587882 226007
rect 587938 221496 587966 235399
rect 588898 227545 588926 235769
rect 588886 227539 588938 227545
rect 588886 227481 588938 227487
rect 588994 227471 589022 235949
rect 597718 235383 597770 235389
rect 597718 235325 597770 235331
rect 588598 227465 588650 227471
rect 588598 227407 588650 227413
rect 588982 227465 589034 227471
rect 588982 227407 589034 227413
rect 587904 221468 587966 221496
rect 588610 221496 588638 227407
rect 593110 227391 593162 227397
rect 593110 227333 593162 227339
rect 590134 227317 590186 227323
rect 590134 227259 590186 227265
rect 589366 227095 589418 227101
rect 589366 227037 589418 227043
rect 588610 221468 588672 221496
rect 589378 221482 589406 227037
rect 590146 221792 590174 227259
rect 590900 226986 590956 226995
rect 590900 226921 590956 226930
rect 590146 221764 590222 221792
rect 590194 221482 590222 221764
rect 590914 221482 590942 226921
rect 591668 226838 591724 226847
rect 591668 226773 591724 226782
rect 591682 221482 591710 226773
rect 592342 224801 592394 224807
rect 592342 224743 592394 224749
rect 592354 221792 592382 224743
rect 592354 221764 592430 221792
rect 592402 221482 592430 221764
rect 593122 221482 593150 227333
rect 593974 227021 594026 227027
rect 593974 226963 594026 226969
rect 593986 221482 594014 226963
rect 596948 226690 597004 226699
rect 596948 226625 597004 226634
rect 596180 226542 596236 226551
rect 596180 226477 596236 226486
rect 594646 226059 594698 226065
rect 594646 226001 594698 226007
rect 594658 221792 594686 226001
rect 595414 225985 595466 225991
rect 595414 225927 595466 225933
rect 594658 221764 594734 221792
rect 594706 221482 594734 221764
rect 595426 221482 595454 225927
rect 596194 221482 596222 226477
rect 596962 221792 596990 226625
rect 596962 221764 597038 221792
rect 597010 221482 597038 221764
rect 597730 221482 597758 235325
rect 598486 235309 598538 235315
rect 598486 235251 598538 235257
rect 598498 221482 598526 235251
rect 599074 227323 599102 239247
rect 599924 229058 599980 229067
rect 599924 228993 599980 229002
rect 599062 227317 599114 227323
rect 599062 227259 599114 227265
rect 599158 226947 599210 226953
rect 599158 226889 599210 226895
rect 599170 221792 599198 226889
rect 599170 221764 599246 221792
rect 599218 221482 599246 221764
rect 599938 221482 599966 228993
rect 600418 226953 600446 241911
rect 602228 235718 602284 235727
rect 602228 235653 602284 235662
rect 600790 235235 600842 235241
rect 600790 235177 600842 235183
rect 600406 226947 600458 226953
rect 600406 226889 600458 226895
rect 600802 221482 600830 235177
rect 601462 230055 601514 230061
rect 601462 229997 601514 230003
rect 601474 221792 601502 229997
rect 601474 221764 601550 221792
rect 601522 221482 601550 221764
rect 602242 221482 602270 235653
rect 602998 226799 603050 226805
rect 602998 226741 603050 226747
rect 603010 221482 603038 226741
rect 603298 226065 603326 253455
rect 603382 250627 603434 250633
rect 603382 250569 603434 250575
rect 603394 226805 603422 250569
rect 603478 247815 603530 247821
rect 603478 247757 603530 247763
rect 603490 227027 603518 247757
rect 605974 235161 606026 235167
rect 605974 235103 606026 235109
rect 605302 235087 605354 235093
rect 605302 235029 605354 235035
rect 604532 231870 604588 231879
rect 604532 231805 604588 231814
rect 603478 227021 603530 227027
rect 603478 226963 603530 226969
rect 603670 226873 603722 226879
rect 603670 226815 603722 226821
rect 603382 226799 603434 226805
rect 603382 226741 603434 226747
rect 603286 226059 603338 226065
rect 603286 226001 603338 226007
rect 603682 221792 603710 226815
rect 603682 221764 603758 221792
rect 603730 221482 603758 221764
rect 604546 221482 604574 231805
rect 605314 221482 605342 235029
rect 605986 221792 606014 235103
rect 606178 226879 606206 262113
rect 606262 259285 606314 259291
rect 606262 259227 606314 259233
rect 606274 227397 606302 259227
rect 606358 256399 606410 256405
rect 606358 256341 606410 256347
rect 606262 227391 606314 227397
rect 606262 227333 606314 227339
rect 606370 227101 606398 256341
rect 629206 247741 629258 247747
rect 629206 247683 629258 247689
rect 627188 240158 627244 240167
rect 627188 240093 627244 240102
rect 621140 236310 621196 236319
rect 621140 236245 621196 236254
rect 608276 235570 608332 235579
rect 608276 235505 608332 235514
rect 607508 228910 607564 228919
rect 607508 228845 607564 228854
rect 606358 227095 606410 227101
rect 606358 227037 606410 227043
rect 606166 226873 606218 226879
rect 606166 226815 606218 226821
rect 606742 226725 606794 226731
rect 606742 226667 606794 226673
rect 605986 221764 606062 221792
rect 606034 221482 606062 221764
rect 606754 221482 606782 226667
rect 607522 221482 607550 228845
rect 608290 221792 608318 235505
rect 611252 235422 611308 235431
rect 611252 235357 611308 235366
rect 609046 229981 609098 229987
rect 609046 229923 609098 229929
rect 608290 221764 608366 221792
rect 608338 221482 608366 221764
rect 609058 221482 609086 229923
rect 609814 226651 609866 226657
rect 609814 226593 609866 226599
rect 609826 221482 609854 226593
rect 610486 226577 610538 226583
rect 610486 226519 610538 226525
rect 610498 221792 610526 226519
rect 610498 221764 610574 221792
rect 610546 221482 610574 221764
rect 611266 221482 611294 235357
rect 614324 235274 614380 235283
rect 614324 235209 614380 235218
rect 612118 229907 612170 229913
rect 612118 229849 612170 229855
rect 612130 221482 612158 229849
rect 612790 226503 612842 226509
rect 612790 226445 612842 226451
rect 612802 221792 612830 226445
rect 613556 226394 613612 226403
rect 613556 226329 613612 226338
rect 612802 221764 612878 221792
rect 612850 221482 612878 221764
rect 613570 221482 613598 226329
rect 614338 221482 614366 235209
rect 614998 233237 615050 233243
rect 614998 233179 615050 233185
rect 615010 221792 615038 233179
rect 615862 227539 615914 227545
rect 615862 227481 615914 227487
rect 615010 221764 615086 221792
rect 615058 221482 615086 221764
rect 615874 221482 615902 227481
rect 618838 227465 618890 227471
rect 618838 227407 618890 227413
rect 616630 227243 616682 227249
rect 616630 227185 616682 227191
rect 616642 221496 616670 227185
rect 618070 226429 618122 226435
rect 618070 226371 618122 226377
rect 617302 226355 617354 226361
rect 617302 226297 617354 226303
rect 616608 221468 616670 221496
rect 617314 221496 617342 226297
rect 617314 221468 617376 221496
rect 618082 221482 618110 226371
rect 618850 221792 618878 227407
rect 619606 227169 619658 227175
rect 619606 227111 619658 227117
rect 618850 221764 618926 221792
rect 618898 221482 618926 221764
rect 619618 221482 619646 227111
rect 620372 226098 620428 226107
rect 620372 226033 620428 226042
rect 620386 221482 620414 226033
rect 621154 221792 621182 236245
rect 624884 235126 624940 235135
rect 624884 235061 624940 235070
rect 621814 235013 621866 235019
rect 621814 234955 621866 234961
rect 621106 221764 621182 221792
rect 621106 221482 621134 221764
rect 621826 221482 621854 234955
rect 622678 229833 622730 229839
rect 622678 229775 622730 229781
rect 622690 221482 622718 229775
rect 624118 226281 624170 226287
rect 623348 226246 623404 226255
rect 624118 226223 624170 226229
rect 623348 226181 623404 226190
rect 623362 221792 623390 226181
rect 623362 221764 623438 221792
rect 623410 221482 623438 221764
rect 624130 221482 624158 226223
rect 624898 221482 624926 235061
rect 625556 234978 625612 234987
rect 625556 234913 625612 234922
rect 626422 234939 626474 234945
rect 625570 221792 625598 234913
rect 626422 234881 626474 234887
rect 625570 221764 625646 221792
rect 625618 221482 625646 221764
rect 626434 221482 626462 234881
rect 627202 221482 627230 240093
rect 627860 234830 627916 234839
rect 627860 234765 627916 234774
rect 628630 234791 628682 234797
rect 627874 221792 627902 234765
rect 628630 234733 628682 234739
rect 627874 221764 627950 221792
rect 627922 221482 627950 221764
rect 628642 221482 628670 234733
rect 629218 225917 629246 247683
rect 629302 244855 629354 244861
rect 629302 244797 629354 244803
rect 629314 226657 629342 244797
rect 630166 234865 630218 234871
rect 630166 234807 630218 234813
rect 629302 226651 629354 226657
rect 629302 226593 629354 226599
rect 629206 225911 629258 225917
rect 629206 225853 629258 225859
rect 629398 225171 629450 225177
rect 629398 225113 629450 225119
rect 629410 221482 629438 225113
rect 630178 221792 630206 234807
rect 632374 234717 632426 234723
rect 630932 234682 630988 234691
rect 632374 234659 632426 234665
rect 630932 234617 630988 234626
rect 630178 221764 630254 221792
rect 630226 221482 630254 221764
rect 630946 221482 630974 234617
rect 631702 226133 631754 226139
rect 631702 226075 631754 226081
rect 631714 221482 631742 226075
rect 632386 221792 632414 234659
rect 639190 227391 639242 227397
rect 639190 227333 639242 227339
rect 633142 227317 633194 227323
rect 633142 227259 633194 227265
rect 632386 221764 632462 221792
rect 632434 221482 632462 221764
rect 633154 221482 633182 227259
rect 638518 227095 638570 227101
rect 638518 227037 638570 227043
rect 636214 227021 636266 227027
rect 636214 226963 636266 226969
rect 634678 226947 634730 226953
rect 634678 226889 634730 226895
rect 634006 226651 634058 226657
rect 634006 226593 634058 226599
rect 634018 221482 634046 226593
rect 634690 221792 634718 226889
rect 635446 225911 635498 225917
rect 635446 225853 635498 225859
rect 634690 221764 634766 221792
rect 634738 221482 634766 221764
rect 635458 221482 635486 225853
rect 636226 221482 636254 226963
rect 636886 226799 636938 226805
rect 636886 226741 636938 226747
rect 636898 221792 636926 226741
rect 637750 226059 637802 226065
rect 637750 226001 637802 226007
rect 636898 221764 636974 221792
rect 636946 221482 636974 221764
rect 637762 221482 637790 226001
rect 638530 221482 638558 227037
rect 639202 221792 639230 227333
rect 639958 226873 640010 226879
rect 639958 226815 640010 226821
rect 639202 221764 639278 221792
rect 639250 221482 639278 221764
rect 639970 221482 639998 226815
rect 640148 212334 640204 212343
rect 640148 212269 640204 212278
rect 640162 211603 640190 212269
rect 640148 211594 640204 211603
rect 640148 211529 640204 211538
rect 190292 201382 190348 201391
rect 190292 201317 190348 201326
rect 190306 200577 190334 201317
rect 640148 200938 640204 200947
rect 640148 200873 640204 200882
rect 190292 200568 190348 200577
rect 190292 200503 190348 200512
rect 640162 200207 640190 200873
rect 640148 200198 640204 200207
rect 640148 200133 640204 200142
rect 187220 199162 187276 199171
rect 187220 199097 187276 199106
rect 185890 195826 186398 195854
rect 185974 185803 186026 185809
rect 185974 185745 186026 185751
rect 185780 182438 185836 182447
rect 185780 182373 185836 182382
rect 185684 174742 185740 174751
rect 185684 174677 185740 174686
rect 185506 155506 185822 155534
rect 184534 155479 184586 155485
rect 184438 155389 184490 155395
rect 184438 155331 184490 155337
rect 184342 155315 184394 155321
rect 184342 155257 184394 155263
rect 184354 155067 184382 155257
rect 184340 155058 184396 155067
rect 184340 154993 184396 155002
rect 184450 154179 184478 155331
rect 184436 154170 184492 154179
rect 184436 154105 184492 154114
rect 184546 153587 184574 155479
rect 184630 155463 184682 155469
rect 184630 155405 184682 155411
rect 184532 153578 184588 153587
rect 184532 153513 184588 153522
rect 184642 152699 184670 155405
rect 184628 152690 184684 152699
rect 184534 152651 184586 152657
rect 184628 152625 184684 152634
rect 184534 152593 184586 152599
rect 184438 152577 184490 152583
rect 184438 152519 184490 152525
rect 184342 152503 184394 152509
rect 184342 152445 184394 152451
rect 184354 151959 184382 152445
rect 184340 151950 184396 151959
rect 184340 151885 184396 151894
rect 184450 151219 184478 152519
rect 184436 151210 184492 151219
rect 184436 151145 184492 151154
rect 184546 150479 184574 152593
rect 184532 150470 184588 150479
rect 184532 150405 184588 150414
rect 184726 149765 184778 149771
rect 184340 149730 184396 149739
rect 184726 149707 184778 149713
rect 184340 149665 184396 149674
rect 184438 149691 184490 149697
rect 184354 149549 184382 149665
rect 184438 149633 184490 149639
rect 184342 149543 184394 149549
rect 184342 149485 184394 149491
rect 184450 148999 184478 149633
rect 184534 149617 184586 149623
rect 184534 149559 184586 149565
rect 184436 148990 184492 148999
rect 184436 148925 184492 148934
rect 184546 147371 184574 149559
rect 184738 148111 184766 149707
rect 184724 148102 184780 148111
rect 184724 148037 184780 148046
rect 184532 147362 184588 147371
rect 184532 147297 184588 147306
rect 184534 146879 184586 146885
rect 184534 146821 184586 146827
rect 184438 146805 184490 146811
rect 184438 146747 184490 146753
rect 184342 146731 184394 146737
rect 184342 146673 184394 146679
rect 184354 145891 184382 146673
rect 184340 145882 184396 145891
rect 184340 145817 184396 145826
rect 184450 145151 184478 146747
rect 184436 145142 184492 145151
rect 184436 145077 184492 145086
rect 184546 144411 184574 146821
rect 184630 146657 184682 146663
rect 184628 146622 184630 146631
rect 184682 146622 184684 146631
rect 184628 146557 184684 146566
rect 184532 144402 184588 144411
rect 184532 144337 184588 144346
rect 183094 143993 183146 143999
rect 183094 143935 183146 143941
rect 184630 143993 184682 143999
rect 184630 143935 184682 143941
rect 184438 143919 184490 143925
rect 184438 143861 184490 143867
rect 184342 143845 184394 143851
rect 184342 143787 184394 143793
rect 184354 143671 184382 143787
rect 184340 143662 184396 143671
rect 184340 143597 184396 143606
rect 184450 142783 184478 143861
rect 184534 143771 184586 143777
rect 184534 143713 184586 143719
rect 184436 142774 184492 142783
rect 184436 142709 184492 142718
rect 184546 141303 184574 143713
rect 184642 142191 184670 143935
rect 184628 142182 184684 142191
rect 184628 142117 184684 142126
rect 184532 141294 184588 141303
rect 184532 141229 184588 141238
rect 184534 141107 184586 141113
rect 184534 141049 184586 141055
rect 184438 141033 184490 141039
rect 184438 140975 184490 140981
rect 184342 140959 184394 140965
rect 184342 140901 184394 140907
rect 184354 140563 184382 140901
rect 184340 140554 184396 140563
rect 184340 140489 184396 140498
rect 184450 139823 184478 140975
rect 184436 139814 184492 139823
rect 184436 139749 184492 139758
rect 184546 138935 184574 141049
rect 184532 138926 184588 138935
rect 184532 138861 184588 138870
rect 184438 135335 184490 135341
rect 184438 135277 184490 135283
rect 184342 135261 184394 135267
rect 184342 135203 184394 135209
rect 184354 134495 184382 135203
rect 184340 134486 184396 134495
rect 184340 134421 184396 134430
rect 184450 133015 184478 135277
rect 185794 135235 185822 155506
rect 185986 138343 186014 185745
rect 186262 182991 186314 182997
rect 186262 182933 186314 182939
rect 186070 182917 186122 182923
rect 186070 182859 186122 182865
rect 185972 138334 186028 138343
rect 185972 138269 186028 138278
rect 186082 137455 186110 182859
rect 186166 174259 186218 174265
rect 186166 174201 186218 174207
rect 186068 137446 186124 137455
rect 186068 137381 186124 137390
rect 185780 135226 185836 135235
rect 185780 135161 185836 135170
rect 186178 133755 186206 174201
rect 186274 136863 186302 182933
rect 186370 173271 186398 195826
rect 640244 185694 640300 185703
rect 640244 185629 640300 185638
rect 640258 184963 640286 185629
rect 640244 184954 640300 184963
rect 640244 184889 640300 184898
rect 186742 184175 186794 184181
rect 186742 184117 186794 184123
rect 186754 183187 186782 184117
rect 186740 183178 186796 183187
rect 186740 183113 186796 183122
rect 645142 183139 645194 183145
rect 645142 183081 645194 183087
rect 645154 183039 645182 183081
rect 645140 183030 645196 183039
rect 645140 182965 645196 182974
rect 186454 180031 186506 180037
rect 186454 179973 186506 179979
rect 186356 173262 186412 173271
rect 186356 173197 186412 173206
rect 186260 136854 186316 136863
rect 186260 136789 186316 136798
rect 186466 135975 186494 179973
rect 645142 179439 645194 179445
rect 645142 179381 645194 179387
rect 645154 179339 645182 179381
rect 645140 179330 645196 179339
rect 645140 179265 645196 179274
rect 645142 174925 645194 174931
rect 645140 174890 645142 174899
rect 645194 174890 645196 174899
rect 645140 174825 645196 174834
rect 645142 171077 645194 171083
rect 645140 171042 645142 171051
rect 645194 171042 645196 171051
rect 645140 170977 645196 170986
rect 645142 168265 645194 168271
rect 645142 168207 645194 168213
rect 645154 167795 645182 168207
rect 645140 167786 645196 167795
rect 645140 167721 645196 167730
rect 645142 163381 645194 163387
rect 645140 163346 645142 163355
rect 645194 163346 645196 163355
rect 645140 163281 645196 163290
rect 645142 159755 645194 159761
rect 645142 159697 645194 159703
rect 645154 159507 645182 159697
rect 645140 159498 645196 159507
rect 645140 159433 645196 159442
rect 645142 156055 645194 156061
rect 645142 155997 645194 156003
rect 645154 155511 645182 155997
rect 645140 155502 645196 155511
rect 645140 155437 645196 155446
rect 645142 152577 645194 152583
rect 645140 152542 645142 152551
rect 645194 152542 645196 152551
rect 645140 152477 645196 152486
rect 645142 148211 645194 148217
rect 645142 148153 645194 148159
rect 645154 148111 645182 148153
rect 645140 148102 645196 148111
rect 645140 148037 645196 148046
rect 186452 135966 186508 135975
rect 186452 135901 186508 135910
rect 186164 133746 186220 133755
rect 186164 133681 186220 133690
rect 184436 133006 184492 133015
rect 184436 132941 184492 132950
rect 184726 132597 184778 132603
rect 184726 132539 184778 132545
rect 182998 132523 183050 132529
rect 182998 132465 183050 132471
rect 182902 112247 182954 112253
rect 182902 112189 182954 112195
rect 183010 106555 183038 132465
rect 184630 132449 184682 132455
rect 184630 132391 184682 132397
rect 184534 132375 184586 132381
rect 184534 132317 184586 132323
rect 184438 132301 184490 132307
rect 184340 132266 184396 132275
rect 184438 132243 184490 132249
rect 184340 132201 184342 132210
rect 184394 132201 184396 132210
rect 184342 132169 184394 132175
rect 184450 131535 184478 132243
rect 184436 131526 184492 131535
rect 184436 131461 184492 131470
rect 184546 130647 184574 132317
rect 184532 130638 184588 130647
rect 184532 130573 184588 130582
rect 184642 129907 184670 132391
rect 184628 129898 184684 129907
rect 184628 129833 184684 129842
rect 184438 129489 184490 129495
rect 184438 129431 184490 129437
rect 184342 129341 184394 129347
rect 184342 129283 184394 129289
rect 184354 128427 184382 129283
rect 184340 128418 184396 128427
rect 184340 128353 184396 128362
rect 184450 127687 184478 129431
rect 184534 129415 184586 129421
rect 184534 129357 184586 129363
rect 184436 127678 184492 127687
rect 184436 127613 184492 127622
rect 184546 126947 184574 129357
rect 184532 126938 184588 126947
rect 184532 126873 184588 126882
rect 184534 126677 184586 126683
rect 184534 126619 184586 126625
rect 184438 126603 184490 126609
rect 184438 126545 184490 126551
rect 184342 126529 184394 126535
rect 184342 126471 184394 126477
rect 184354 126059 184382 126471
rect 184340 126050 184396 126059
rect 184340 125985 184396 125994
rect 184450 125467 184478 126545
rect 184436 125458 184492 125467
rect 184436 125393 184492 125402
rect 184546 124579 184574 126619
rect 184532 124570 184588 124579
rect 184532 124505 184588 124514
rect 184630 123865 184682 123871
rect 184436 123830 184492 123839
rect 184630 123807 184682 123813
rect 184436 123765 184492 123774
rect 184534 123791 184586 123797
rect 184450 123723 184478 123765
rect 184534 123733 184586 123739
rect 184438 123717 184490 123723
rect 184438 123659 184490 123665
rect 184342 123643 184394 123649
rect 184342 123585 184394 123591
rect 184354 123099 184382 123585
rect 184340 123090 184396 123099
rect 184340 123025 184396 123034
rect 184546 121619 184574 123733
rect 184642 122211 184670 123807
rect 184628 122202 184684 122211
rect 184628 122137 184684 122146
rect 184532 121610 184588 121619
rect 184532 121545 184588 121554
rect 184534 120979 184586 120985
rect 184534 120921 184586 120927
rect 184342 120905 184394 120911
rect 184342 120847 184394 120853
rect 184354 120731 184382 120847
rect 184438 120831 184490 120837
rect 184438 120773 184490 120779
rect 184340 120722 184396 120731
rect 184340 120657 184396 120666
rect 184450 119251 184478 120773
rect 184546 120139 184574 120921
rect 184532 120130 184588 120139
rect 184532 120065 184588 120074
rect 184436 119242 184492 119251
rect 184436 119177 184492 119186
rect 184738 118659 184766 132539
rect 185590 132079 185642 132085
rect 185590 132021 185642 132027
rect 184724 118650 184780 118659
rect 184724 118585 184780 118594
rect 184630 118093 184682 118099
rect 184630 118035 184682 118041
rect 184534 118019 184586 118025
rect 184534 117961 184586 117967
rect 184438 117945 184490 117951
rect 184438 117887 184490 117893
rect 184342 117871 184394 117877
rect 184342 117813 184394 117819
rect 184354 117771 184382 117813
rect 184340 117762 184396 117771
rect 184340 117697 184396 117706
rect 184450 117031 184478 117887
rect 184436 117022 184492 117031
rect 184436 116957 184492 116966
rect 184546 116291 184574 117961
rect 184532 116282 184588 116291
rect 184532 116217 184588 116226
rect 184642 115403 184670 118035
rect 184628 115394 184684 115403
rect 184628 115329 184684 115338
rect 184534 115207 184586 115213
rect 184534 115149 184586 115155
rect 184438 115133 184490 115139
rect 184438 115075 184490 115081
rect 184342 115059 184394 115065
rect 184342 115001 184394 115007
rect 184354 114811 184382 115001
rect 184340 114802 184396 114811
rect 184340 114737 184396 114746
rect 184450 113923 184478 115075
rect 184436 113914 184492 113923
rect 184436 113849 184492 113858
rect 184546 113183 184574 115149
rect 184630 114171 184682 114177
rect 184630 114113 184682 114119
rect 184532 113174 184588 113183
rect 184532 113109 184588 113118
rect 184642 112443 184670 114113
rect 184628 112434 184684 112443
rect 184628 112369 184684 112378
rect 184342 112321 184394 112327
rect 184342 112263 184394 112269
rect 184354 111703 184382 112263
rect 184534 112247 184586 112253
rect 184534 112189 184586 112195
rect 184438 112173 184490 112179
rect 184438 112115 184490 112121
rect 184340 111694 184396 111703
rect 184340 111629 184396 111638
rect 184450 110963 184478 112115
rect 184436 110954 184492 110963
rect 184436 110889 184492 110898
rect 184546 110223 184574 112189
rect 184532 110214 184588 110223
rect 184532 110149 184588 110158
rect 184438 109435 184490 109441
rect 184438 109377 184490 109383
rect 184342 109361 184394 109367
rect 184340 109326 184342 109335
rect 184394 109326 184396 109335
rect 184340 109261 184396 109270
rect 184450 107115 184478 109377
rect 185602 108743 185630 132021
rect 645718 129637 645770 129643
rect 645718 129579 645770 129585
rect 186742 129563 186794 129569
rect 186742 129505 186794 129511
rect 186754 129167 186782 129505
rect 186740 129158 186796 129167
rect 186740 129093 186796 129102
rect 645730 129019 645758 129579
rect 645716 129010 645772 129019
rect 645716 128945 645772 128954
rect 646498 126979 646526 275317
rect 647362 269323 647390 278018
rect 648610 272135 648638 278018
rect 648596 272126 648652 272135
rect 648596 272061 648652 272070
rect 647348 269314 647404 269323
rect 647348 269249 647404 269258
rect 646580 267094 646636 267103
rect 646580 267029 646636 267038
rect 646486 126973 646538 126979
rect 646486 126915 646538 126921
rect 186166 122459 186218 122465
rect 186166 122401 186218 122407
rect 185588 108734 185644 108743
rect 185588 108669 185644 108678
rect 186178 107855 186206 122401
rect 646498 122063 646526 126915
rect 646594 126831 646622 267029
rect 646678 253513 646730 253519
rect 646678 253455 646730 253461
rect 646690 144263 646718 253455
rect 646774 207411 646826 207417
rect 646774 207353 646826 207359
rect 646676 144254 646732 144263
rect 646676 144189 646732 144198
rect 646786 141007 646814 207353
rect 649378 183145 649406 861106
rect 655126 792085 655178 792091
rect 655126 792027 655178 792033
rect 654358 780541 654410 780547
rect 654358 780483 654410 780489
rect 654370 773559 654398 780483
rect 655138 775927 655166 792027
rect 656566 783501 656618 783507
rect 656566 783443 656618 783449
rect 655220 778286 655276 778295
rect 655220 778221 655276 778230
rect 655124 775918 655180 775927
rect 655124 775853 655180 775862
rect 654356 773550 654412 773559
rect 654356 773485 654412 773494
rect 654070 737473 654122 737479
rect 654070 737415 654122 737421
rect 654082 730195 654110 737415
rect 654166 737399 654218 737405
rect 654166 737341 654218 737347
rect 654068 730186 654124 730195
rect 654068 730121 654124 730130
rect 654178 728567 654206 737341
rect 655124 734478 655180 734487
rect 655124 734413 655180 734422
rect 654164 728558 654220 728567
rect 654164 728493 654220 728502
rect 653782 702841 653834 702847
rect 653782 702783 653834 702789
rect 649462 702767 649514 702773
rect 649462 702709 649514 702715
rect 649366 183139 649418 183145
rect 649366 183081 649418 183087
rect 649474 179445 649502 702709
rect 653794 686979 653822 702783
rect 654166 694183 654218 694189
rect 654166 694125 654218 694131
rect 654070 691371 654122 691377
rect 654070 691313 654122 691319
rect 653780 686970 653836 686979
rect 653780 686905 653836 686914
rect 654082 684611 654110 691313
rect 654178 685351 654206 694125
rect 654164 685342 654220 685351
rect 654164 685277 654220 685286
rect 654068 684602 654124 684611
rect 654068 684537 654124 684546
rect 655138 668215 655166 734413
rect 655234 714465 655262 778221
rect 655412 777694 655468 777703
rect 655412 777629 655468 777638
rect 655316 731666 655372 731675
rect 655316 731601 655372 731610
rect 655222 714459 655274 714465
rect 655222 714401 655274 714407
rect 655220 689486 655276 689495
rect 655220 689421 655276 689430
rect 655126 668209 655178 668215
rect 655126 668151 655178 668157
rect 652246 666803 652298 666809
rect 652246 666745 652298 666751
rect 649750 666729 649802 666735
rect 649750 666671 649802 666677
rect 649558 656739 649610 656745
rect 649558 656681 649610 656687
rect 649462 179439 649514 179445
rect 649462 179381 649514 179387
rect 649570 174931 649598 656681
rect 649654 610637 649706 610643
rect 649654 610579 649706 610585
rect 649558 174925 649610 174931
rect 649558 174867 649610 174873
rect 649666 171083 649694 610579
rect 649762 263551 649790 666671
rect 649846 564535 649898 564541
rect 649846 564477 649898 564483
rect 649748 263542 649804 263551
rect 649748 263477 649804 263486
rect 649654 171077 649706 171083
rect 649654 171019 649706 171025
rect 649858 168271 649886 564477
rect 649942 521319 649994 521325
rect 649942 521261 649994 521267
rect 649846 168265 649898 168271
rect 649846 168207 649898 168213
rect 646870 164417 646922 164423
rect 646870 164359 646922 164365
rect 646772 140998 646828 141007
rect 646772 140933 646828 140942
rect 646582 126825 646634 126831
rect 646582 126767 646634 126773
rect 646594 123839 646622 126767
rect 646882 125763 646910 164359
rect 647062 164343 647114 164349
rect 647062 164285 647114 164291
rect 646966 164269 647018 164275
rect 646966 164211 647018 164217
rect 646978 127687 647006 164211
rect 647074 134791 647102 164285
rect 649954 163387 649982 521261
rect 650038 478177 650090 478183
rect 650038 478119 650090 478125
rect 649942 163381 649994 163387
rect 649942 163323 649994 163329
rect 650050 159761 650078 478119
rect 650134 388859 650186 388865
rect 650134 388801 650186 388807
rect 650038 159755 650090 159761
rect 650038 159697 650090 159703
rect 650146 156061 650174 388801
rect 650230 345865 650282 345871
rect 650230 345807 650282 345813
rect 650134 156055 650186 156061
rect 650134 155997 650186 156003
rect 650242 152583 650270 345807
rect 650326 299763 650378 299769
rect 650326 299705 650378 299711
rect 650230 152577 650282 152583
rect 650230 152519 650282 152525
rect 650338 148217 650366 299705
rect 652258 266955 652286 666745
rect 654166 656813 654218 656819
rect 654166 656755 654218 656761
rect 654178 640655 654206 656755
rect 655124 642422 655180 642431
rect 655124 642357 655180 642366
rect 654164 640646 654220 640655
rect 654164 640581 654220 640590
rect 653974 602053 654026 602059
rect 653974 601995 654026 602001
rect 653986 594183 654014 601995
rect 653972 594174 654028 594183
rect 653972 594109 654028 594118
rect 655138 576233 655166 642357
rect 655234 622261 655262 689421
rect 655330 668437 655358 731601
rect 655426 714613 655454 777629
rect 655604 776066 655660 776075
rect 655604 776001 655660 776010
rect 655508 732702 655564 732711
rect 655508 732637 655564 732646
rect 655414 714607 655466 714613
rect 655414 714549 655466 714555
rect 655412 688450 655468 688459
rect 655412 688385 655468 688394
rect 655318 668431 655370 668437
rect 655318 668373 655370 668379
rect 655316 643014 655372 643023
rect 655316 642949 655372 642958
rect 655222 622255 655274 622261
rect 655222 622197 655274 622203
rect 655220 597874 655276 597883
rect 655220 597809 655276 597818
rect 655126 576227 655178 576233
rect 655126 576169 655178 576175
rect 654166 555951 654218 555957
rect 654166 555893 654218 555899
rect 654178 548599 654206 555893
rect 655124 553326 655180 553335
rect 655124 553261 655180 553270
rect 654164 548590 654220 548599
rect 654164 548525 654220 548534
rect 655138 489801 655166 553261
rect 655234 533017 655262 597809
rect 655330 576381 655358 642949
rect 655426 624999 655454 688385
rect 655522 668585 655550 732637
rect 655618 714761 655646 776001
rect 656578 774743 656606 783443
rect 656564 774734 656620 774743
rect 656564 774669 656620 774678
rect 655702 748869 655754 748875
rect 655702 748811 655754 748817
rect 655714 731379 655742 748811
rect 655700 731370 655756 731379
rect 655700 731305 655756 731314
rect 655606 714755 655658 714761
rect 655606 714697 655658 714703
rect 669718 713127 669770 713133
rect 669718 713069 669770 713075
rect 669526 711943 669578 711949
rect 669526 711885 669578 711891
rect 655604 687118 655660 687127
rect 655604 687053 655660 687062
rect 655510 668579 655562 668585
rect 655510 668521 655562 668527
rect 655508 640794 655564 640803
rect 655508 640729 655564 640738
rect 655414 624993 655466 624999
rect 655414 624935 655466 624941
rect 655412 596690 655468 596699
rect 655412 596625 655468 596634
rect 655318 576375 655370 576381
rect 655318 576317 655370 576323
rect 655316 550958 655372 550967
rect 655316 550893 655372 550902
rect 655222 533011 655274 533017
rect 655222 532953 655274 532959
rect 655330 489949 655358 550893
rect 655426 533165 655454 596625
rect 655522 576529 655550 640729
rect 655618 622409 655646 687053
rect 655798 648229 655850 648235
rect 655798 648171 655850 648177
rect 655810 639175 655838 648171
rect 655990 645195 656042 645201
rect 655990 645137 656042 645143
rect 655796 639166 655852 639175
rect 655796 639101 655852 639110
rect 656002 638287 656030 645137
rect 655988 638278 656044 638287
rect 655988 638213 656044 638222
rect 655606 622403 655658 622409
rect 655606 622345 655658 622351
rect 655798 613523 655850 613529
rect 655798 613465 655850 613471
rect 655604 595506 655660 595515
rect 655604 595441 655660 595450
rect 655510 576523 655562 576529
rect 655510 576465 655562 576471
rect 655508 552142 655564 552151
rect 655508 552077 655564 552086
rect 655414 533159 655466 533165
rect 655414 533101 655466 533107
rect 655522 490097 655550 552077
rect 655618 533313 655646 595441
rect 655810 595367 655838 613465
rect 656566 602201 656618 602207
rect 656566 602143 656618 602149
rect 655796 595358 655852 595367
rect 655796 595293 655852 595302
rect 656578 592999 656606 602143
rect 656564 592990 656620 592999
rect 656564 592925 656620 592934
rect 655702 567495 655754 567501
rect 655702 567437 655754 567443
rect 655714 550819 655742 567437
rect 656566 558837 656618 558843
rect 656566 558779 656618 558785
rect 655700 550810 655756 550819
rect 655700 550745 655756 550754
rect 656578 549783 656606 558779
rect 656564 549774 656620 549783
rect 656564 549709 656620 549718
rect 655606 533307 655658 533313
rect 655606 533249 655658 533255
rect 655510 490091 655562 490097
rect 655510 490033 655562 490039
rect 655318 489943 655370 489949
rect 655318 489885 655370 489891
rect 655126 489795 655178 489801
rect 655126 489737 655178 489743
rect 655126 400625 655178 400631
rect 655126 400567 655178 400573
rect 655138 373367 655166 400567
rect 655510 400551 655562 400557
rect 655510 400493 655562 400499
rect 655318 400477 655370 400483
rect 655318 400419 655370 400425
rect 655124 373358 655180 373367
rect 655124 373293 655180 373302
rect 655330 372183 655358 400419
rect 655522 374403 655550 400493
rect 656566 381607 656618 381613
rect 656566 381549 656618 381555
rect 655508 374394 655564 374403
rect 655508 374329 655564 374338
rect 655316 372174 655372 372183
rect 655316 372109 655372 372118
rect 656578 370999 656606 381549
rect 656564 370990 656620 370999
rect 656564 370925 656620 370934
rect 655318 357335 655370 357341
rect 655318 357277 655370 357283
rect 655222 357261 655274 357267
rect 655222 357203 655274 357209
rect 655126 357187 655178 357193
rect 655126 357129 655178 357135
rect 654166 328327 654218 328333
rect 654166 328269 654218 328275
rect 654178 326303 654206 328269
rect 655138 328079 655166 357129
rect 655234 329855 655262 357203
rect 655220 329846 655276 329855
rect 655220 329781 655276 329790
rect 655124 328070 655180 328079
rect 655124 328005 655180 328014
rect 655330 327487 655358 357277
rect 666742 340019 666794 340025
rect 666742 339961 666794 339967
rect 666754 328333 666782 339961
rect 666742 328327 666794 328333
rect 666742 328269 666794 328275
rect 655316 327478 655372 327487
rect 655316 327413 655372 327422
rect 654164 326294 654220 326303
rect 654164 326229 654220 326238
rect 654262 311233 654314 311239
rect 654262 311175 654314 311181
rect 654166 311159 654218 311165
rect 654166 311101 654218 311107
rect 654070 311085 654122 311091
rect 654070 311027 654122 311033
rect 654082 302179 654110 311027
rect 654178 303363 654206 311101
rect 654164 303354 654220 303363
rect 654164 303289 654220 303298
rect 654068 302170 654124 302179
rect 654068 302105 654124 302114
rect 654274 300995 654302 311175
rect 654260 300986 654316 300995
rect 654260 300921 654316 300930
rect 656564 298766 656620 298775
rect 656564 298701 656620 298710
rect 656084 297582 656140 297591
rect 656084 297517 656140 297526
rect 655892 294030 655948 294039
rect 655892 293965 655948 293974
rect 655796 292846 655852 292855
rect 655796 292781 655852 292790
rect 655604 289294 655660 289303
rect 655604 289229 655660 289238
rect 655412 288110 655468 288119
rect 655412 288045 655468 288054
rect 653780 284558 653836 284567
rect 653780 284493 653836 284502
rect 653794 284303 653822 284493
rect 653782 284297 653834 284303
rect 653782 284239 653834 284245
rect 655124 283374 655180 283383
rect 655124 283309 655180 283318
rect 654164 279822 654220 279831
rect 654164 279757 654220 279766
rect 654178 279493 654206 279757
rect 654166 279487 654218 279493
rect 654166 279429 654218 279435
rect 652244 266946 652300 266955
rect 652244 266881 652300 266890
rect 650326 148211 650378 148217
rect 650326 148153 650378 148159
rect 647060 134782 647116 134791
rect 647060 134717 647116 134726
rect 647828 130934 647884 130943
rect 647828 130869 647884 130878
rect 646964 127678 647020 127687
rect 646964 127613 647020 127622
rect 646868 125754 646924 125763
rect 646868 125689 646924 125698
rect 646580 123830 646636 123839
rect 646580 123765 646636 123774
rect 646484 122054 646540 122063
rect 646484 121989 646540 121998
rect 647842 118395 647870 130869
rect 655138 129865 655166 283309
rect 655316 282338 655372 282347
rect 655316 282273 655372 282282
rect 655220 281006 655276 281015
rect 655220 280941 655276 280950
rect 655234 130013 655262 280941
rect 655330 130161 655358 282273
rect 655426 175893 655454 288045
rect 655508 286926 655564 286935
rect 655508 286861 655564 286870
rect 655522 176041 655550 286861
rect 655618 201571 655646 289229
rect 655700 285742 655756 285751
rect 655700 285677 655756 285686
rect 655606 201565 655658 201571
rect 655606 201507 655658 201513
rect 655714 176189 655742 285677
rect 655810 219109 655838 292781
rect 655906 247673 655934 293965
rect 655988 290922 656044 290931
rect 655988 290857 656044 290866
rect 655894 247667 655946 247673
rect 655894 247609 655946 247615
rect 656002 219257 656030 290857
rect 656098 265137 656126 297517
rect 656276 296842 656332 296851
rect 656276 296777 656332 296786
rect 656180 291662 656236 291671
rect 656180 291597 656236 291606
rect 656086 265131 656138 265137
rect 656086 265073 656138 265079
rect 656194 221847 656222 291597
rect 656290 265285 656318 296777
rect 656372 295214 656428 295223
rect 656372 295149 656428 295158
rect 656386 290464 656414 295149
rect 656578 290889 656606 298701
rect 656566 290883 656618 290889
rect 656566 290825 656618 290831
rect 656386 290436 656606 290464
rect 656578 265433 656606 290436
rect 658006 284297 658058 284303
rect 658006 284239 658058 284245
rect 656566 265427 656618 265433
rect 656566 265369 656618 265375
rect 656278 265279 656330 265285
rect 656278 265221 656330 265227
rect 656182 221841 656234 221847
rect 656182 221783 656234 221789
rect 655990 219251 656042 219257
rect 655990 219193 656042 219199
rect 655798 219103 655850 219109
rect 655798 219045 655850 219051
rect 655702 176183 655754 176189
rect 655702 176125 655754 176131
rect 655510 176035 655562 176041
rect 655510 175977 655562 175983
rect 655414 175887 655466 175893
rect 655414 175829 655466 175835
rect 658018 155543 658046 284239
rect 663766 279487 663818 279493
rect 663766 279429 663818 279435
rect 658006 155537 658058 155543
rect 658006 155479 658058 155485
rect 655318 130155 655370 130161
rect 655318 130097 655370 130103
rect 655222 130007 655274 130013
rect 655222 129949 655274 129955
rect 655126 129859 655178 129865
rect 655126 129801 655178 129807
rect 647924 119538 647980 119547
rect 647924 119473 647980 119482
rect 647830 118389 647882 118395
rect 647830 118331 647882 118337
rect 647938 118247 647966 119473
rect 647926 118241 647978 118247
rect 647926 118183 647978 118189
rect 645238 118167 645290 118173
rect 645238 118109 645290 118115
rect 645250 117623 645278 118109
rect 645236 117614 645292 117623
rect 645236 117549 645292 117558
rect 647924 115690 647980 115699
rect 647924 115625 647980 115634
rect 647938 115287 647966 115625
rect 647926 115281 647978 115287
rect 647926 115223 647978 115229
rect 646580 113174 646636 113183
rect 646580 113109 646636 113118
rect 186164 107846 186220 107855
rect 186164 107781 186220 107790
rect 184436 107106 184492 107115
rect 184436 107041 184492 107050
rect 182998 106549 183050 106555
rect 182998 106491 183050 106497
rect 184534 106549 184586 106555
rect 184534 106491 184586 106497
rect 184342 106475 184394 106481
rect 184342 106417 184394 106423
rect 179926 106401 179978 106407
rect 179926 106343 179978 106349
rect 184354 105635 184382 106417
rect 184438 106327 184490 106333
rect 184438 106269 184490 106275
rect 184340 105626 184396 105635
rect 184340 105561 184396 105570
rect 184450 104007 184478 106269
rect 184546 104895 184574 106491
rect 185302 106401 185354 106407
rect 185300 106366 185302 106375
rect 185354 106366 185356 106375
rect 185300 106301 185356 106310
rect 645908 106070 645964 106079
rect 645908 106005 645964 106014
rect 184726 105143 184778 105149
rect 184726 105085 184778 105091
rect 184532 104886 184588 104895
rect 184532 104821 184588 104830
rect 184436 103998 184492 104007
rect 184436 103933 184492 103942
rect 184438 103663 184490 103669
rect 184438 103605 184490 103611
rect 184342 103441 184394 103447
rect 184450 103415 184478 103605
rect 184630 103589 184682 103595
rect 184630 103531 184682 103537
rect 184534 103515 184586 103521
rect 184534 103457 184586 103463
rect 184342 103383 184394 103389
rect 184436 103406 184492 103415
rect 184354 102527 184382 103383
rect 184436 103341 184492 103350
rect 184340 102518 184396 102527
rect 184340 102453 184396 102462
rect 184546 101935 184574 103457
rect 184532 101926 184588 101935
rect 184532 101861 184588 101870
rect 184642 101047 184670 103531
rect 184628 101038 184684 101047
rect 184628 100973 184684 100982
rect 184630 100777 184682 100783
rect 184630 100719 184682 100725
rect 184438 100703 184490 100709
rect 184438 100645 184490 100651
rect 184342 100555 184394 100561
rect 184342 100497 184394 100503
rect 184354 100307 184382 100497
rect 184340 100298 184396 100307
rect 184340 100233 184396 100242
rect 184450 99567 184478 100645
rect 184534 100629 184586 100635
rect 184534 100571 184586 100577
rect 184436 99558 184492 99567
rect 184436 99493 184492 99502
rect 184546 98087 184574 100571
rect 184642 98679 184670 100719
rect 184628 98670 184684 98679
rect 184628 98605 184684 98614
rect 184532 98078 184588 98087
rect 184246 98039 184298 98045
rect 184532 98013 184588 98022
rect 184246 97981 184298 97987
rect 179926 95079 179978 95085
rect 179926 95021 179978 95027
rect 177142 91897 177194 91903
rect 177142 91839 177194 91845
rect 171286 83461 171338 83467
rect 171286 83403 171338 83409
rect 165238 80501 165290 80507
rect 165238 80443 165290 80449
rect 179938 80433 179966 95021
rect 184258 81955 184286 97981
rect 184342 97891 184394 97897
rect 184342 97833 184394 97839
rect 184354 97199 184382 97833
rect 184438 97817 184490 97823
rect 184438 97759 184490 97765
rect 184340 97190 184396 97199
rect 184340 97125 184396 97134
rect 184450 96459 184478 97759
rect 184436 96450 184492 96459
rect 184436 96385 184492 96394
rect 184738 95719 184766 105085
rect 645922 103743 645950 106005
rect 645910 103737 645962 103743
rect 645910 103679 645962 103685
rect 645140 102222 645196 102231
rect 645140 102157 645196 102166
rect 645154 102115 645182 102157
rect 645142 102109 645194 102115
rect 645142 102051 645194 102057
rect 186166 97965 186218 97971
rect 186166 97907 186218 97913
rect 184724 95710 184780 95719
rect 184724 95645 184780 95654
rect 184630 95005 184682 95011
rect 184630 94947 184682 94953
rect 184534 94931 184586 94937
rect 184534 94873 184586 94879
rect 184438 94857 184490 94863
rect 184340 94822 184396 94831
rect 184438 94799 184490 94805
rect 184340 94757 184342 94766
rect 184394 94757 184396 94766
rect 184342 94725 184394 94731
rect 184450 94239 184478 94799
rect 184436 94230 184492 94239
rect 184436 94165 184492 94174
rect 184546 93499 184574 94873
rect 184532 93490 184588 93499
rect 184532 93425 184588 93434
rect 184642 92759 184670 94947
rect 184628 92750 184684 92759
rect 184628 92685 184684 92694
rect 184438 92119 184490 92125
rect 184438 92061 184490 92067
rect 184340 92010 184396 92019
rect 184340 91945 184342 91954
rect 184394 91945 184396 91954
rect 184342 91913 184394 91919
rect 184450 90391 184478 92061
rect 184534 92045 184586 92051
rect 184534 91987 184586 91993
rect 184436 90382 184492 90391
rect 184436 90317 184492 90326
rect 184546 89651 184574 91987
rect 184630 91897 184682 91903
rect 184630 91839 184682 91845
rect 184642 91131 184670 91839
rect 184628 91122 184684 91131
rect 184628 91057 184684 91066
rect 184532 89642 184588 89651
rect 184532 89577 184588 89586
rect 184534 89233 184586 89239
rect 184534 89175 184586 89181
rect 184438 89085 184490 89091
rect 184438 89027 184490 89033
rect 184342 89011 184394 89017
rect 184342 88953 184394 88959
rect 184354 88911 184382 88953
rect 184340 88902 184396 88911
rect 184340 88837 184396 88846
rect 184450 88171 184478 89027
rect 184436 88162 184492 88171
rect 184436 88097 184492 88106
rect 184546 87283 184574 89175
rect 184630 89159 184682 89165
rect 184630 89101 184682 89107
rect 184532 87274 184588 87283
rect 184532 87209 184588 87218
rect 184642 86691 184670 89101
rect 184628 86682 184684 86691
rect 184628 86617 184684 86626
rect 184342 86421 184394 86427
rect 184342 86363 184394 86369
rect 184354 85803 184382 86363
rect 184438 86347 184490 86353
rect 184438 86289 184490 86295
rect 184340 85794 184396 85803
rect 184340 85729 184396 85738
rect 184450 85211 184478 86289
rect 184534 86273 184586 86279
rect 184534 86215 184586 86221
rect 184436 85202 184492 85211
rect 184436 85137 184492 85146
rect 184546 84323 184574 86215
rect 184532 84314 184588 84323
rect 184532 84249 184588 84258
rect 184438 83535 184490 83541
rect 184438 83477 184490 83483
rect 184342 83461 184394 83467
rect 184340 83426 184342 83435
rect 184394 83426 184396 83435
rect 184340 83361 184396 83370
rect 184244 81946 184300 81955
rect 184244 81881 184300 81890
rect 184450 81363 184478 83477
rect 186178 82843 186206 97907
rect 642262 96485 642314 96491
rect 642262 96427 642314 96433
rect 642274 83541 642302 96427
rect 645428 96006 645484 96015
rect 645428 95941 645430 95950
rect 645482 95941 645484 95950
rect 645430 95909 645482 95915
rect 646486 92415 646538 92421
rect 646486 92357 646538 92363
rect 645526 92341 645578 92347
rect 645526 92283 645578 92289
rect 640726 83535 640778 83541
rect 640726 83477 640778 83483
rect 642262 83535 642314 83541
rect 642262 83477 642314 83483
rect 186164 82834 186220 82843
rect 186164 82769 186220 82778
rect 184436 81354 184492 81363
rect 184436 81289 184492 81298
rect 184438 80649 184490 80655
rect 184438 80591 184490 80597
rect 184342 80501 184394 80507
rect 184342 80443 184394 80449
rect 179926 80427 179978 80433
rect 179926 80369 179978 80375
rect 184354 78995 184382 80443
rect 184450 79883 184478 80591
rect 184534 80575 184586 80581
rect 184534 80517 184586 80523
rect 184436 79874 184492 79883
rect 184436 79809 184492 79818
rect 184340 78986 184396 78995
rect 184340 78921 184396 78930
rect 184546 78255 184574 80517
rect 184628 80466 184684 80475
rect 184628 80401 184630 80410
rect 184682 80401 184684 80410
rect 184630 80369 184682 80375
rect 184532 78246 184588 78255
rect 184532 78181 184588 78190
rect 184438 77763 184490 77769
rect 184438 77705 184490 77711
rect 159766 77541 159818 77547
rect 159766 77483 159818 77489
rect 184342 77541 184394 77547
rect 184450 77515 184478 77705
rect 184534 77689 184586 77695
rect 184534 77631 184586 77637
rect 184342 77483 184394 77489
rect 184436 77506 184492 77515
rect 184354 76775 184382 77483
rect 184436 77441 184492 77450
rect 184340 76766 184396 76775
rect 184340 76701 184396 76710
rect 184546 76035 184574 77631
rect 184630 77615 184682 77621
rect 184630 77557 184682 77563
rect 184532 76026 184588 76035
rect 184532 75961 184588 75970
rect 184642 75147 184670 77557
rect 184628 75138 184684 75147
rect 184628 75073 184684 75082
rect 184534 74877 184586 74883
rect 184534 74819 184586 74825
rect 184438 74729 184490 74735
rect 184438 74671 184490 74677
rect 154102 74655 154154 74661
rect 154102 74597 154154 74603
rect 184342 74655 184394 74661
rect 184342 74597 184394 74603
rect 184354 74407 184382 74597
rect 184340 74398 184396 74407
rect 184340 74333 184396 74342
rect 184450 72927 184478 74671
rect 184546 73667 184574 74819
rect 184630 74803 184682 74809
rect 184630 74745 184682 74751
rect 184532 73658 184588 73667
rect 184532 73593 184588 73602
rect 184436 72918 184492 72927
rect 184436 72853 184492 72862
rect 184642 72187 184670 74745
rect 184628 72178 184684 72187
rect 184628 72113 184684 72122
rect 184438 71991 184490 71997
rect 184438 71933 184490 71939
rect 149686 71917 149738 71923
rect 149686 71859 149738 71865
rect 149590 71843 149642 71849
rect 149590 71785 149642 71791
rect 184342 71843 184394 71849
rect 184342 71785 184394 71791
rect 149506 70952 149630 70980
rect 149492 70846 149548 70855
rect 149492 70781 149548 70790
rect 149396 69514 149452 69523
rect 149396 69449 149452 69458
rect 149302 68883 149354 68889
rect 149302 68825 149354 68831
rect 149204 68330 149260 68339
rect 149204 68265 149260 68274
rect 149110 66219 149162 66225
rect 149110 66161 149162 66167
rect 149014 65997 149066 66003
rect 149014 65939 149066 65945
rect 149218 63339 149246 68265
rect 149410 66151 149438 69449
rect 149398 66145 149450 66151
rect 149398 66087 149450 66093
rect 149506 66077 149534 70781
rect 149602 69111 149630 70952
rect 184354 70559 184382 71785
rect 184450 71447 184478 71933
rect 184534 71917 184586 71923
rect 184534 71859 184586 71865
rect 184436 71438 184492 71447
rect 184436 71373 184492 71382
rect 184340 70550 184396 70559
rect 184340 70485 184396 70494
rect 184546 69967 184574 71859
rect 184532 69958 184588 69967
rect 184532 69893 184588 69902
rect 149590 69105 149642 69111
rect 184534 69105 184586 69111
rect 149590 69047 149642 69053
rect 184340 69070 184396 69079
rect 184534 69047 184586 69053
rect 184340 69005 184342 69014
rect 184394 69005 184396 69014
rect 184342 68973 184394 68979
rect 184438 68957 184490 68963
rect 184438 68899 184490 68905
rect 184342 68883 184394 68889
rect 184342 68825 184394 68831
rect 149588 67146 149644 67155
rect 149588 67081 149644 67090
rect 149494 66071 149546 66077
rect 149494 66013 149546 66019
rect 149492 65370 149548 65379
rect 149492 65305 149548 65314
rect 149396 64630 149452 64639
rect 149396 64565 149452 64574
rect 149300 63446 149356 63455
rect 149300 63381 149356 63390
rect 149206 63333 149258 63339
rect 149206 63275 149258 63281
rect 149314 60453 149342 63381
rect 149410 63191 149438 64565
rect 149506 63265 149534 65305
rect 149494 63259 149546 63265
rect 149494 63201 149546 63207
rect 149398 63185 149450 63191
rect 149398 63127 149450 63133
rect 149602 63117 149630 67081
rect 184354 66859 184382 68825
rect 184450 67599 184478 68899
rect 184546 68487 184574 69047
rect 184532 68478 184588 68487
rect 184532 68413 184588 68422
rect 184436 67590 184492 67599
rect 184436 67525 184492 67534
rect 184340 66850 184396 66859
rect 184340 66785 184396 66794
rect 184534 66219 184586 66225
rect 184534 66161 184586 66167
rect 184340 66110 184396 66119
rect 184340 66045 184396 66054
rect 184438 66071 184490 66077
rect 184354 66003 184382 66045
rect 184438 66013 184490 66019
rect 184342 65997 184394 66003
rect 184342 65939 184394 65945
rect 184450 64639 184478 66013
rect 184546 65231 184574 66161
rect 184630 66145 184682 66151
rect 184630 66087 184682 66093
rect 184532 65222 184588 65231
rect 184532 65157 184588 65166
rect 184436 64630 184492 64639
rect 184436 64565 184492 64574
rect 184642 63751 184670 66087
rect 184628 63742 184684 63751
rect 184628 63677 184684 63686
rect 184438 63333 184490 63339
rect 184438 63275 184490 63281
rect 184450 63159 184478 63275
rect 184534 63259 184586 63265
rect 184534 63201 184586 63207
rect 184436 63150 184492 63159
rect 149590 63111 149642 63117
rect 149590 63053 149642 63059
rect 184342 63111 184394 63117
rect 184436 63085 184492 63094
rect 184342 63053 184394 63059
rect 184354 62271 184382 63053
rect 149396 62262 149452 62271
rect 149396 62197 149452 62206
rect 184340 62262 184396 62271
rect 184340 62197 184396 62206
rect 149302 60447 149354 60453
rect 149302 60389 149354 60395
rect 149410 60305 149438 62197
rect 184546 61531 184574 63201
rect 184630 63185 184682 63191
rect 184630 63127 184682 63133
rect 184532 61522 184588 61531
rect 184532 61457 184588 61466
rect 184642 60791 184670 63127
rect 184628 60782 184684 60791
rect 184628 60717 184684 60726
rect 149492 60634 149548 60643
rect 149492 60569 149548 60578
rect 149506 60379 149534 60569
rect 184438 60447 184490 60453
rect 184438 60389 184490 60395
rect 149494 60373 149546 60379
rect 149494 60315 149546 60321
rect 149398 60299 149450 60305
rect 149398 60241 149450 60247
rect 184342 60299 184394 60305
rect 184342 60241 184394 60247
rect 149396 59746 149452 59755
rect 149396 59681 149452 59690
rect 149410 59047 149438 59681
rect 184354 59311 184382 60241
rect 184450 60051 184478 60389
rect 184534 60373 184586 60379
rect 184534 60315 184586 60321
rect 184436 60042 184492 60051
rect 184436 59977 184492 59986
rect 184340 59302 184396 59311
rect 184340 59237 184396 59246
rect 149398 59041 149450 59047
rect 149398 58983 149450 58989
rect 184342 59041 184394 59047
rect 184342 58983 184394 58989
rect 149396 58562 149452 58571
rect 149396 58497 149452 58506
rect 149410 57567 149438 58497
rect 184354 57683 184382 58983
rect 184546 58423 184574 60315
rect 184532 58414 184588 58423
rect 184532 58349 184588 58358
rect 184340 57674 184396 57683
rect 184340 57609 184396 57618
rect 149398 57561 149450 57567
rect 149398 57503 149450 57509
rect 184342 57561 184394 57567
rect 184342 57503 184394 57509
rect 149492 57378 149548 57387
rect 149492 57313 149548 57322
rect 149398 56229 149450 56235
rect 149396 56194 149398 56203
rect 149450 56194 149452 56203
rect 149506 56161 149534 57313
rect 184354 56943 184382 57503
rect 184340 56934 184396 56943
rect 184340 56869 184396 56878
rect 184438 56229 184490 56235
rect 184340 56194 184396 56203
rect 149396 56129 149452 56138
rect 149494 56155 149546 56161
rect 184438 56171 184490 56177
rect 184340 56129 184342 56138
rect 149494 56097 149546 56103
rect 184394 56129 184396 56138
rect 184342 56097 184394 56103
rect 184450 55463 184478 56171
rect 184436 55454 184492 55463
rect 184436 55389 184492 55398
rect 149684 54862 149740 54871
rect 149684 54797 149740 54806
rect 149698 54681 149726 54797
rect 184340 54714 184396 54723
rect 149686 54675 149738 54681
rect 184340 54649 184342 54658
rect 149686 54617 149738 54623
rect 184394 54649 184396 54658
rect 184342 54617 184394 54623
rect 184340 53974 184396 53983
rect 184340 53909 184396 53918
rect 149396 53826 149452 53835
rect 149396 53761 149452 53770
rect 149410 53275 149438 53761
rect 184354 53275 184382 53909
rect 149398 53269 149450 53275
rect 149398 53211 149450 53217
rect 184342 53269 184394 53275
rect 184342 53211 184394 53217
rect 175606 53195 175658 53201
rect 175606 53137 175658 53143
rect 145104 49788 145406 49816
rect 145378 47133 145406 49788
rect 145366 47127 145418 47133
rect 145366 47069 145418 47075
rect 142114 46680 142416 46708
rect 142114 40219 142142 46680
rect 175618 44198 175646 53137
rect 199138 47133 199166 53650
rect 199126 47127 199178 47133
rect 199126 47069 199178 47075
rect 216418 46171 216446 53650
rect 233698 47725 233726 53650
rect 233686 47719 233738 47725
rect 233686 47661 233738 47667
rect 250978 47577 251006 53650
rect 268320 53636 268574 53664
rect 285600 53636 285854 53664
rect 268546 47651 268574 53636
rect 268534 47645 268586 47651
rect 268534 47587 268586 47593
rect 250966 47571 251018 47577
rect 250966 47513 251018 47519
rect 207382 46165 207434 46171
rect 207382 46107 207434 46113
rect 216406 46165 216458 46171
rect 216406 46107 216458 46113
rect 175606 44192 175658 44198
rect 175606 44134 175658 44140
rect 186262 42021 186314 42027
rect 186262 41963 186314 41969
rect 187030 42021 187082 42027
rect 194326 42021 194378 42027
rect 187082 41969 187344 41972
rect 187030 41963 187344 41969
rect 186274 41509 186302 41963
rect 187042 41944 187344 41963
rect 194064 41969 194326 41972
rect 194064 41963 194378 41969
rect 194064 41944 194366 41963
rect 207394 41509 207422 46107
rect 285826 43285 285854 53636
rect 302914 47873 302942 53650
rect 311062 47941 311114 47947
rect 311062 47883 311114 47889
rect 302902 47867 302954 47873
rect 302902 47809 302954 47815
rect 285814 43279 285866 43285
rect 285814 43221 285866 43227
rect 311074 42268 311102 47883
rect 320194 47799 320222 53650
rect 320182 47793 320234 47799
rect 320182 47735 320234 47741
rect 337474 46615 337502 53650
rect 331222 46609 331274 46615
rect 331222 46551 331274 46557
rect 337462 46609 337514 46615
rect 337462 46551 337514 46557
rect 310498 42240 311102 42268
rect 302902 42169 302954 42175
rect 302688 42117 302902 42120
rect 310498 42120 310526 42240
rect 302688 42111 302954 42117
rect 302688 42092 302942 42111
rect 307008 42101 307262 42120
rect 307008 42095 307274 42101
rect 307008 42092 307222 42095
rect 310128 42092 310526 42120
rect 311158 42169 311210 42175
rect 311158 42111 311210 42117
rect 311062 42095 311114 42101
rect 307222 42037 307274 42043
rect 311062 42037 311114 42043
rect 186262 41503 186314 41509
rect 186262 41445 186314 41451
rect 207382 41503 207434 41509
rect 207382 41445 207434 41451
rect 142100 40210 142156 40219
rect 142100 40145 142156 40154
rect 311074 37259 311102 42037
rect 311060 37250 311116 37259
rect 311060 37185 311116 37194
rect 311170 31635 311198 42111
rect 331234 37259 331262 46551
rect 354850 42101 354878 53650
rect 371938 53636 372192 53664
rect 389218 53636 389472 53664
rect 371938 47947 371966 53636
rect 371926 47941 371978 47947
rect 371926 47883 371978 47889
rect 365314 42240 365726 42268
rect 357718 42169 357770 42175
rect 357456 42117 357718 42120
rect 365314 42120 365342 42240
rect 357456 42111 357770 42117
rect 335446 42095 335498 42101
rect 335446 42037 335498 42043
rect 354838 42095 354890 42101
rect 357456 42092 357758 42111
rect 361776 42101 362078 42120
rect 361776 42095 362090 42101
rect 361776 42092 362038 42095
rect 354838 42037 354890 42043
rect 364944 42092 365342 42120
rect 362038 42037 362090 42043
rect 331220 37250 331276 37259
rect 331220 37185 331276 37194
rect 335458 31667 335486 42037
rect 365698 41824 365726 42240
rect 365974 42095 366026 42101
rect 365974 42037 366026 42043
rect 365698 41796 365918 41824
rect 365890 37439 365918 41796
rect 365878 37433 365930 37439
rect 365878 37375 365930 37381
rect 365986 37365 366014 42037
rect 389218 37365 389246 53636
rect 405526 47941 405578 47947
rect 405526 47883 405578 47889
rect 402166 46165 402218 46171
rect 402166 46107 402218 46113
rect 402178 42101 402206 46107
rect 403510 43205 403562 43211
rect 403510 43147 403562 43153
rect 402166 42095 402218 42101
rect 402166 42037 402218 42043
rect 403522 37513 403550 43147
rect 405538 42106 405566 47883
rect 406786 46171 406814 53650
rect 417526 48015 417578 48021
rect 417526 47957 417578 47963
rect 406774 46165 406826 46171
rect 406774 46107 406826 46113
rect 417538 44955 417566 47957
rect 424066 47503 424094 53650
rect 441346 47947 441374 53650
rect 441334 47941 441386 47947
rect 441334 47883 441386 47889
rect 418870 47497 418922 47503
rect 418870 47439 418922 47445
rect 424054 47497 424106 47503
rect 424054 47439 424106 47445
rect 417524 44946 417580 44955
rect 417524 44881 417580 44890
rect 418882 43211 418910 47439
rect 458626 43211 458654 53650
rect 475714 53636 475968 53664
rect 492994 53636 493248 53664
rect 510370 53636 510624 53664
rect 460342 48089 460394 48095
rect 460342 48031 460394 48037
rect 418870 43205 418922 43211
rect 418870 43147 418922 43153
rect 444886 43205 444938 43211
rect 444886 43147 444938 43153
rect 458614 43205 458666 43211
rect 458614 43147 458666 43153
rect 415220 41986 415276 41995
rect 415220 41921 415276 41930
rect 415234 41810 415262 41921
rect 416852 41838 416908 41847
rect 416592 41796 416852 41824
rect 416852 41773 416908 41782
rect 420788 40506 420844 40515
rect 420788 40441 420844 40450
rect 403510 37507 403562 37513
rect 403510 37449 403562 37455
rect 365974 37359 366026 37365
rect 365974 37301 366026 37307
rect 389206 37359 389258 37365
rect 389206 37301 389258 37307
rect 420802 34553 420830 40441
rect 444898 34553 444926 43147
rect 460354 42106 460382 48031
rect 472246 47941 472298 47947
rect 472246 47883 472298 47889
rect 464854 46461 464906 46467
rect 464854 46403 464906 46409
rect 464866 41847 464894 46403
rect 472258 44955 472286 47883
rect 475510 47719 475562 47725
rect 475510 47661 475562 47667
rect 472244 44946 472300 44955
rect 472244 44881 472300 44890
rect 471408 42101 471710 42120
rect 471408 42095 471722 42101
rect 471408 42092 471670 42095
rect 471670 42037 471722 42043
rect 464852 41838 464908 41847
rect 470324 41838 470380 41847
rect 470160 41796 470324 41824
rect 464852 41773 464908 41782
rect 470324 41773 470380 41782
rect 475522 37439 475550 47661
rect 475714 46467 475742 53636
rect 480982 48163 481034 48169
rect 480982 48105 481034 48111
rect 475702 46461 475754 46467
rect 475702 46403 475754 46409
rect 480994 42101 481022 48105
rect 492994 48021 493022 53636
rect 510370 48095 510398 53636
rect 527938 48169 527966 53650
rect 527926 48163 527978 48169
rect 527926 48105 527978 48111
rect 510358 48089 510410 48095
rect 510358 48031 510410 48037
rect 492982 48015 493034 48021
rect 492982 47957 493034 47963
rect 506806 47867 506858 47873
rect 506806 47809 506858 47815
rect 506818 44913 506846 47809
rect 529270 47793 529322 47799
rect 529270 47735 529322 47741
rect 520630 47645 520682 47651
rect 520630 47587 520682 47593
rect 506806 44907 506858 44913
rect 506806 44849 506858 44855
rect 512182 44907 512234 44913
rect 512182 44849 512234 44855
rect 480982 42095 481034 42101
rect 480982 42037 481034 42043
rect 512194 41847 512222 44849
rect 518722 43285 518834 43304
rect 518710 43279 518834 43285
rect 518762 43276 518834 43279
rect 518710 43221 518762 43227
rect 520642 42106 520670 47587
rect 521206 47571 521258 47577
rect 521206 47513 521258 47519
rect 521218 43304 521246 47513
rect 521218 43276 521534 43304
rect 521506 42120 521534 43276
rect 521506 42092 521856 42120
rect 529282 42106 529310 47735
rect 545218 46245 545246 53650
rect 562498 47947 562526 53650
rect 579796 53602 579852 54402
rect 597092 53602 597148 54402
rect 614388 53602 614444 54402
rect 631684 53602 631740 54402
rect 640738 49057 640766 83477
rect 645538 79439 645566 92283
rect 645908 88902 645964 88911
rect 645908 88837 645964 88846
rect 645922 87537 645950 88837
rect 645910 87531 645962 87537
rect 645910 87473 645962 87479
rect 645908 84462 645964 84471
rect 645908 84397 645964 84406
rect 645922 84207 645950 84397
rect 645910 84201 645962 84207
rect 645910 84143 645962 84149
rect 645524 79430 645580 79439
rect 645524 79365 645580 79374
rect 646006 76135 646058 76141
rect 646006 76077 646058 76083
rect 646018 75591 646046 76077
rect 646004 75582 646060 75591
rect 646004 75517 646060 75526
rect 646004 66258 646060 66267
rect 646004 66193 646006 66202
rect 646058 66193 646060 66202
rect 646006 66161 646058 66167
rect 646006 59115 646058 59121
rect 646006 59057 646058 59063
rect 646018 59015 646046 59057
rect 646004 59006 646060 59015
rect 646004 58941 646060 58950
rect 646498 54723 646526 92357
rect 646594 77695 646622 113109
rect 663778 112993 663806 279429
rect 669538 275243 669566 711885
rect 669622 622995 669674 623001
rect 669622 622937 669674 622943
rect 669524 275234 669580 275243
rect 669524 275169 669580 275178
rect 669634 264915 669662 622937
rect 669730 275095 669758 713069
rect 670678 712683 670730 712689
rect 670678 712625 670730 712631
rect 670690 668067 670718 712625
rect 670882 711949 670910 890373
rect 670978 713133 671006 891409
rect 673078 778765 673130 778771
rect 673078 778707 673130 778713
rect 672118 737621 672170 737627
rect 672118 737563 672170 737569
rect 670966 713127 671018 713133
rect 670966 713069 671018 713075
rect 670870 711943 670922 711949
rect 670870 711885 670922 711891
rect 670774 711573 670826 711579
rect 670774 711515 670826 711521
rect 670786 679694 670814 711515
rect 672022 689373 672074 689379
rect 672022 689315 672074 689321
rect 670786 679666 670910 679694
rect 670678 668061 670730 668067
rect 670678 668003 670730 668009
rect 670690 666735 670718 668003
rect 670774 667691 670826 667697
rect 670774 667633 670826 667639
rect 670678 666729 670730 666735
rect 670678 666671 670730 666677
rect 670678 642309 670730 642315
rect 670678 642251 670730 642257
rect 670582 622477 670634 622483
rect 670582 622419 670634 622425
rect 670486 621367 670538 621373
rect 670486 621309 670538 621315
rect 669814 619887 669866 619893
rect 669814 619829 669866 619835
rect 669716 275086 669772 275095
rect 669716 275021 669772 275030
rect 669826 264989 669854 619829
rect 670498 574975 670526 621309
rect 670594 575937 670622 622419
rect 670582 575931 670634 575937
rect 670582 575873 670634 575879
rect 670486 574969 670538 574975
rect 670486 574911 670538 574917
rect 670498 573273 670526 574911
rect 669910 573267 669962 573273
rect 669910 573209 669962 573215
rect 670486 573267 670538 573273
rect 670486 573209 670538 573215
rect 669922 277611 669950 573209
rect 670594 573199 670622 575873
rect 670102 573193 670154 573199
rect 670102 573135 670154 573141
rect 670582 573193 670634 573199
rect 670582 573135 670634 573141
rect 670006 487131 670058 487137
rect 670006 487073 670058 487079
rect 669908 277602 669964 277611
rect 669908 277537 669964 277546
rect 670018 273615 670046 487073
rect 670114 277759 670142 573135
rect 670690 569573 670718 642251
rect 670786 623001 670814 667633
rect 670882 666809 670910 679666
rect 670870 666803 670922 666809
rect 670870 666745 670922 666751
rect 670966 666359 671018 666365
rect 670966 666301 671018 666307
rect 670870 648969 670922 648975
rect 670870 648911 670922 648917
rect 670774 622995 670826 623001
rect 670774 622937 670826 622943
rect 670774 603903 670826 603909
rect 670774 603845 670826 603851
rect 670678 569567 670730 569573
rect 670678 569509 670730 569515
rect 670786 527467 670814 603845
rect 670882 570683 670910 648911
rect 670978 621965 671006 666301
rect 670966 621959 671018 621965
rect 670966 621901 671018 621907
rect 670978 619893 671006 621901
rect 670966 619887 671018 619893
rect 670966 619829 671018 619835
rect 672034 615971 672062 689315
rect 672130 662147 672158 737563
rect 672886 734809 672938 734815
rect 672886 734751 672938 734757
rect 672310 734439 672362 734445
rect 672310 734381 672362 734387
rect 672214 689151 672266 689157
rect 672214 689093 672266 689099
rect 672118 662141 672170 662147
rect 672118 662083 672170 662089
rect 672022 615965 672074 615971
rect 672022 615907 672074 615913
rect 672226 614491 672254 689093
rect 672322 661407 672350 734381
rect 672406 734217 672458 734223
rect 672406 734159 672458 734165
rect 672310 661401 672362 661407
rect 672310 661343 672362 661349
rect 672418 659927 672446 734159
rect 672790 732367 672842 732373
rect 672790 732309 672842 732315
rect 672694 713423 672746 713429
rect 672694 713365 672746 713371
rect 672598 693665 672650 693671
rect 672598 693607 672650 693613
rect 672502 687375 672554 687381
rect 672502 687317 672554 687323
rect 672406 659921 672458 659927
rect 672406 659863 672458 659869
rect 672406 648303 672458 648309
rect 672406 648245 672458 648251
rect 672310 623439 672362 623445
rect 672310 623381 672362 623387
rect 672214 614485 672266 614491
rect 672214 614427 672266 614433
rect 670966 606937 671018 606943
rect 670966 606879 671018 606885
rect 670870 570677 670922 570683
rect 670870 570619 670922 570625
rect 670978 528059 671006 606879
rect 672322 577047 672350 623381
rect 672310 577041 672362 577047
rect 672310 576983 672362 576989
rect 672214 575487 672266 575493
rect 672214 575429 672266 575435
rect 672226 532721 672254 575429
rect 672310 574377 672362 574383
rect 672310 574319 672362 574325
rect 672214 532715 672266 532721
rect 672214 532657 672266 532663
rect 672322 531537 672350 574319
rect 672418 569943 672446 648245
rect 672514 616563 672542 687317
rect 672610 617155 672638 693607
rect 672706 669251 672734 713365
rect 672694 669245 672746 669251
rect 672694 669187 672746 669193
rect 672802 661703 672830 732309
rect 672790 661697 672842 661703
rect 672790 661639 672842 661645
rect 672898 660223 672926 734751
rect 673090 704919 673118 778707
rect 673174 738287 673226 738293
rect 673174 738229 673226 738235
rect 673078 704913 673130 704919
rect 673078 704855 673130 704861
rect 673078 692925 673130 692931
rect 673078 692867 673130 692873
rect 672982 689817 673034 689823
rect 672982 689759 673034 689765
rect 672886 660217 672938 660223
rect 672886 660159 672938 660165
rect 672886 644825 672938 644831
rect 672886 644767 672938 644773
rect 672790 644085 672842 644091
rect 672790 644027 672842 644033
rect 672694 643641 672746 643647
rect 672694 643583 672746 643589
rect 672598 617149 672650 617155
rect 672598 617091 672650 617097
rect 672502 616557 672554 616563
rect 672502 616499 672554 616505
rect 672598 598945 672650 598951
rect 672598 598887 672650 598893
rect 672502 597169 672554 597175
rect 672502 597111 672554 597117
rect 672406 569937 672458 569943
rect 672406 569879 672458 569885
rect 672406 532715 672458 532721
rect 672406 532657 672458 532663
rect 672310 531531 672362 531537
rect 672310 531473 672362 531479
rect 670966 528053 671018 528059
rect 670966 527995 671018 528001
rect 670774 527461 670826 527467
rect 670774 527403 670826 527409
rect 670294 488167 670346 488173
rect 670294 488109 670346 488115
rect 670198 398923 670250 398929
rect 670198 398865 670250 398871
rect 670100 277750 670156 277759
rect 670100 277685 670156 277694
rect 670004 273606 670060 273615
rect 670004 273541 670060 273550
rect 670210 270655 670238 398865
rect 670306 277463 670334 488109
rect 670486 398479 670538 398485
rect 670486 398421 670538 398427
rect 670498 277907 670526 398421
rect 672322 278647 672350 531473
rect 672308 278638 672364 278647
rect 672308 278573 672364 278582
rect 672418 278055 672446 532657
rect 672514 526357 672542 597111
rect 672502 526351 672554 526357
rect 672502 526293 672554 526299
rect 672610 524507 672638 598887
rect 672706 567723 672734 643583
rect 672802 569203 672830 644027
rect 672790 569197 672842 569203
rect 672790 569139 672842 569145
rect 672898 568019 672926 644767
rect 672994 615231 673022 689759
rect 673090 615675 673118 692867
rect 673186 660667 673214 738229
rect 673378 714243 673406 892371
rect 676052 891506 676108 891515
rect 676052 891441 676054 891450
rect 676106 891441 676108 891450
rect 676054 891409 676106 891415
rect 676052 890470 676108 890479
rect 676052 890405 676054 890414
rect 676106 890405 676108 890414
rect 676054 890373 676106 890379
rect 680180 890174 680236 890183
rect 680180 890109 680236 890118
rect 676244 889286 676300 889295
rect 676244 889221 676300 889230
rect 676258 887921 676286 889221
rect 679988 888694 680044 888703
rect 679988 888629 680044 888638
rect 673942 887915 673994 887921
rect 673942 887857 673994 887863
rect 676246 887915 676298 887921
rect 676246 887857 676298 887863
rect 673954 875267 673982 887857
rect 676244 887806 676300 887815
rect 676244 887741 676300 887750
rect 676052 887436 676108 887445
rect 676052 887371 676108 887380
rect 676066 887181 676094 887371
rect 674134 887175 674186 887181
rect 674134 887117 674186 887123
rect 676054 887175 676106 887181
rect 676054 887117 676106 887123
rect 674038 885103 674090 885109
rect 674038 885045 674090 885051
rect 673942 875261 673994 875267
rect 673942 875203 673994 875209
rect 674050 867423 674078 885045
rect 674146 868163 674174 887117
rect 676258 887107 676286 887741
rect 674230 887101 674282 887107
rect 674230 887043 674282 887049
rect 676246 887101 676298 887107
rect 676246 887043 676298 887049
rect 674242 876155 674270 887043
rect 679700 886770 679756 886779
rect 679700 886705 679756 886714
rect 676052 885512 676108 885521
rect 676052 885447 676108 885456
rect 676066 885109 676094 885447
rect 676054 885103 676106 885109
rect 676054 885045 676106 885051
rect 676052 884994 676108 885003
rect 676052 884929 676108 884938
rect 675764 884402 675820 884411
rect 675764 884337 675820 884346
rect 674518 884289 674570 884295
rect 674518 884231 674570 884237
rect 674422 883623 674474 883629
rect 674422 883565 674474 883571
rect 674326 881255 674378 881261
rect 674326 881197 674378 881203
rect 674230 876149 674282 876155
rect 674230 876091 674282 876097
rect 674338 874971 674366 881197
rect 674434 875360 674462 883565
rect 674530 875489 674558 884231
rect 675286 883253 675338 883259
rect 675286 883195 675338 883201
rect 675094 883179 675146 883185
rect 675094 883121 675146 883127
rect 674998 883105 675050 883111
rect 674818 883053 674998 883056
rect 674818 883047 675050 883053
rect 674818 883028 675038 883047
rect 674614 880145 674666 880151
rect 674614 880087 674666 880093
rect 674518 875483 674570 875489
rect 674518 875425 674570 875431
rect 674434 875332 674558 875360
rect 674422 875261 674474 875267
rect 674422 875203 674474 875209
rect 674326 874965 674378 874971
rect 674326 874907 674378 874913
rect 674134 868157 674186 868163
rect 674134 868099 674186 868105
rect 674038 867417 674090 867423
rect 674038 867359 674090 867365
rect 674434 865795 674462 875203
rect 674530 869865 674558 875332
rect 674626 874305 674654 880087
rect 674614 874299 674666 874305
rect 674614 874241 674666 874247
rect 674614 872671 674666 872677
rect 674614 872613 674666 872619
rect 674518 869859 674570 869865
rect 674518 869801 674570 869807
rect 674626 868089 674654 872613
rect 674818 868256 674846 883028
rect 674998 882883 675050 882889
rect 674998 882825 675050 882831
rect 674902 878369 674954 878375
rect 674902 878311 674954 878317
rect 674914 872973 674942 878311
rect 675010 877265 675038 882825
rect 674998 877259 675050 877265
rect 674998 877201 675050 877207
rect 675106 876396 675134 883121
rect 675190 879553 675242 879559
rect 675190 879495 675242 879501
rect 675202 876673 675230 879495
rect 675298 877537 675326 883195
rect 675478 881403 675530 881409
rect 675478 881345 675530 881351
rect 675490 878084 675518 881345
rect 675778 878375 675806 884337
rect 676066 884295 676094 884929
rect 676054 884289 676106 884295
rect 676054 884231 676106 884237
rect 676052 884032 676108 884041
rect 676052 883967 676108 883976
rect 676066 883629 676094 883967
rect 676054 883623 676106 883629
rect 676054 883565 676106 883571
rect 676052 883514 676108 883523
rect 676052 883449 676108 883458
rect 676066 883111 676094 883449
rect 676054 883105 676106 883111
rect 676054 883047 676106 883053
rect 679714 882889 679742 886705
rect 679796 886178 679852 886187
rect 679796 886113 679852 886122
rect 679702 882883 679754 882889
rect 679702 882825 679754 882831
rect 679700 882774 679756 882783
rect 679700 882709 679756 882718
rect 679714 882191 679742 882709
rect 679700 882182 679756 882191
rect 679700 882117 679756 882126
rect 679714 881483 679742 882117
rect 679702 881477 679754 881483
rect 679702 881419 679754 881425
rect 679810 880151 679838 886113
rect 679892 885734 679948 885743
rect 679892 885669 679948 885678
rect 679798 880145 679850 880151
rect 679798 880087 679850 880093
rect 679906 879559 679934 885669
rect 680002 883259 680030 888629
rect 680084 888250 680140 888259
rect 680084 888185 680140 888194
rect 679990 883253 680042 883259
rect 679990 883195 680042 883201
rect 680098 881261 680126 888185
rect 680194 883185 680222 890109
rect 680182 883179 680234 883185
rect 680182 883121 680234 883127
rect 685460 882182 685516 882191
rect 685460 882117 685516 882126
rect 685474 881747 685502 882117
rect 685460 881738 685516 881747
rect 685460 881673 685516 881682
rect 680086 881255 680138 881261
rect 680086 881197 680138 881203
rect 679894 879553 679946 879559
rect 679894 879495 679946 879501
rect 675766 878369 675818 878375
rect 675766 878311 675818 878317
rect 675298 877509 675408 877537
rect 675478 877259 675530 877265
rect 675478 877201 675530 877207
rect 675490 876900 675518 877201
rect 675190 876667 675242 876673
rect 675190 876609 675242 876615
rect 675106 876368 675422 876396
rect 675394 876234 675422 876368
rect 675190 876223 675242 876229
rect 675190 876165 675242 876171
rect 675094 876149 675146 876155
rect 675094 876091 675146 876097
rect 674998 875483 675050 875489
rect 674998 875425 675050 875431
rect 674902 872967 674954 872973
rect 674902 872909 674954 872915
rect 675010 868889 675038 875425
rect 675106 872654 675134 876091
rect 675202 873565 675230 876165
rect 675478 874965 675530 874971
rect 675478 874907 675530 874913
rect 675490 874384 675518 874907
rect 675478 874299 675530 874305
rect 675478 874241 675530 874247
rect 675490 873866 675518 874241
rect 675190 873559 675242 873565
rect 675190 873501 675242 873507
rect 675382 873559 675434 873565
rect 675382 873501 675434 873507
rect 675394 873200 675422 873501
rect 675382 872967 675434 872973
rect 675382 872909 675434 872915
rect 675106 872626 675230 872654
rect 675202 870032 675230 872626
rect 675394 872534 675422 872909
rect 675394 870032 675422 870092
rect 675202 870004 675422 870032
rect 675382 869859 675434 869865
rect 675382 869801 675434 869807
rect 675394 869500 675422 869801
rect 675010 868861 675408 868889
rect 674818 868228 675408 868256
rect 674998 868157 675050 868163
rect 674998 868099 675050 868105
rect 674614 868083 674666 868089
rect 674614 868025 674666 868031
rect 674422 865789 674474 865795
rect 674422 865731 674474 865737
rect 675010 863372 675038 868099
rect 675094 868083 675146 868089
rect 675094 868025 675146 868031
rect 675106 867693 675134 868025
rect 675106 867665 675408 867693
rect 675478 867417 675530 867423
rect 675478 867359 675530 867365
rect 675490 867058 675518 867359
rect 675106 865825 675408 865853
rect 675106 864019 675134 865825
rect 675190 865789 675242 865795
rect 675190 865731 675242 865737
rect 675202 865222 675230 865731
rect 675202 865194 675408 865222
rect 675094 864013 675146 864019
rect 675094 863955 675146 863961
rect 675010 863344 675408 863372
rect 675382 792085 675434 792091
rect 675382 792027 675434 792033
rect 675394 788875 675422 792027
rect 675394 788063 675422 788322
rect 675380 788054 675436 788063
rect 675380 787989 675436 787998
rect 675778 787471 675806 787656
rect 675764 787462 675820 787471
rect 675764 787397 675820 787406
rect 675490 786731 675518 787035
rect 675476 786722 675532 786731
rect 675476 786657 675532 786666
rect 675394 784807 675422 785214
rect 675380 784798 675436 784807
rect 675380 784733 675436 784742
rect 675490 784215 675518 784622
rect 675476 784206 675532 784215
rect 675476 784141 675532 784150
rect 675298 783985 675408 784013
rect 674998 783501 675050 783507
rect 675298 783475 675326 783985
rect 674998 783443 675050 783449
rect 675284 783466 675340 783475
rect 675010 778919 675038 783443
rect 675284 783401 675340 783410
rect 675778 783031 675806 783364
rect 675764 783022 675820 783031
rect 675764 782957 675820 782966
rect 675682 780663 675710 780848
rect 675668 780654 675724 780663
rect 675668 780589 675724 780598
rect 675286 780541 675338 780547
rect 675286 780483 675338 780489
rect 674998 778913 675050 778919
rect 674998 778855 675050 778861
rect 675298 776644 675326 780483
rect 675778 779923 675806 780330
rect 675764 779914 675820 779923
rect 675764 779849 675820 779858
rect 675778 779183 675806 779664
rect 675764 779174 675820 779183
rect 675764 779109 675820 779118
rect 675382 778913 675434 778919
rect 675382 778855 675434 778861
rect 675394 778480 675422 778855
rect 675490 778771 675518 779031
rect 675478 778765 675530 778771
rect 675478 778707 675530 778713
rect 675490 777703 675518 777814
rect 675476 777694 675532 777703
rect 675476 777629 675532 777638
rect 675298 776616 675408 776644
rect 675778 775483 675806 775995
rect 675764 775474 675820 775483
rect 675764 775409 675820 775418
rect 675298 774141 675408 774169
rect 675298 773665 675326 774141
rect 674518 773659 674570 773665
rect 674518 773601 674570 773607
rect 675286 773659 675338 773665
rect 675286 773601 675338 773607
rect 674422 742135 674474 742141
rect 674422 742077 674474 742083
rect 674434 730639 674462 742077
rect 674420 730630 674476 730639
rect 674420 730565 674476 730574
rect 674422 730517 674474 730523
rect 674422 730459 674474 730465
rect 674230 728667 674282 728673
rect 674230 728609 674282 728615
rect 673366 714237 673418 714243
rect 673366 714179 673418 714185
rect 673270 668505 673322 668511
rect 673270 668447 673322 668453
rect 673174 660661 673226 660667
rect 673174 660603 673226 660609
rect 673282 624037 673310 668447
rect 674242 665255 674270 728609
rect 674326 685525 674378 685531
rect 674326 685467 674378 685473
rect 674230 665249 674282 665255
rect 674230 665191 674282 665197
rect 673366 648081 673418 648087
rect 673366 648023 673418 648029
rect 673270 624031 673322 624037
rect 673270 623973 673322 623979
rect 673078 615669 673130 615675
rect 673078 615611 673130 615617
rect 672982 615225 673034 615231
rect 672982 615167 673034 615173
rect 673270 603089 673322 603095
rect 673270 603031 673322 603037
rect 673174 601979 673226 601985
rect 673174 601921 673226 601927
rect 672982 599833 673034 599839
rect 672982 599775 673034 599781
rect 672886 568013 672938 568019
rect 672886 567955 672938 567961
rect 672694 567717 672746 567723
rect 672694 567659 672746 567665
rect 672790 556099 672842 556105
rect 672790 556041 672842 556047
rect 672694 553953 672746 553959
rect 672694 553895 672746 553901
rect 672598 524501 672650 524507
rect 672598 524443 672650 524449
rect 672706 481587 672734 553895
rect 672694 481581 672746 481587
rect 672694 481523 672746 481529
rect 672802 480847 672830 556041
rect 672886 551955 672938 551961
rect 672886 551897 672938 551903
rect 672898 481957 672926 551897
rect 672994 524877 673022 599775
rect 673078 599315 673130 599321
rect 673078 599257 673130 599263
rect 673090 525987 673118 599257
rect 673186 526727 673214 601921
rect 673174 526721 673226 526727
rect 673174 526663 673226 526669
rect 673078 525981 673130 525987
rect 673078 525923 673130 525929
rect 673282 525247 673310 603031
rect 673378 568463 673406 648023
rect 674338 622039 674366 685467
rect 674434 668141 674462 730459
rect 674530 711135 674558 773601
rect 674996 772070 675052 772079
rect 674996 772005 675052 772014
rect 674900 771922 674956 771931
rect 674900 771857 674956 771866
rect 674614 737399 674666 737405
rect 674614 737341 674666 737347
rect 674626 732077 674654 737341
rect 674614 732071 674666 732077
rect 674614 732013 674666 732019
rect 674914 711357 674942 771857
rect 674902 711351 674954 711357
rect 674902 711293 674954 711299
rect 674518 711129 674570 711135
rect 674518 711071 674570 711077
rect 675010 708471 675038 772005
rect 675382 748869 675434 748875
rect 675382 748811 675434 748817
rect 675394 743848 675422 748811
rect 675202 743316 675408 743344
rect 675202 742141 675230 743316
rect 675490 742479 675518 742664
rect 675476 742470 675532 742479
rect 675476 742405 675532 742414
rect 675190 742135 675242 742141
rect 675190 742077 675242 742083
rect 675202 742021 675408 742049
rect 675202 741147 675230 742021
rect 675188 741138 675244 741147
rect 675188 741073 675244 741082
rect 675476 740398 675532 740407
rect 675476 740333 675532 740342
rect 675490 740222 675518 740333
rect 675490 739223 675518 739630
rect 675476 739214 675532 739223
rect 675476 739149 675532 739158
rect 675298 738985 675408 739013
rect 675298 737627 675326 738985
rect 675394 738293 675422 738372
rect 675382 738287 675434 738293
rect 675382 738229 675434 738235
rect 675286 737621 675338 737627
rect 675286 737563 675338 737569
rect 675286 737473 675338 737479
rect 675286 737415 675338 737421
rect 675298 736832 675326 737415
rect 675202 736804 675326 736832
rect 675202 733927 675230 736804
rect 675778 735523 675806 735856
rect 675764 735514 675820 735523
rect 675764 735449 675820 735458
rect 675394 734815 675422 735338
rect 675382 734809 675434 734815
rect 675382 734751 675434 734757
rect 675394 734445 675422 734672
rect 675382 734439 675434 734445
rect 675382 734381 675434 734387
rect 675382 734217 675434 734223
rect 675382 734159 675434 734165
rect 675394 734006 675422 734159
rect 675190 733921 675242 733927
rect 675190 733863 675242 733869
rect 675478 733921 675530 733927
rect 675478 733863 675530 733869
rect 675490 733488 675518 733863
rect 675490 732373 675518 732822
rect 675478 732367 675530 732373
rect 675478 732309 675530 732315
rect 675382 732071 675434 732077
rect 675382 732013 675434 732019
rect 675394 731638 675422 732013
rect 675490 730523 675518 730972
rect 675478 730517 675530 730523
rect 675478 730459 675530 730465
rect 675490 728673 675518 729155
rect 675478 728667 675530 728673
rect 675478 728609 675530 728615
rect 676340 715534 676396 715543
rect 676340 715469 676396 715478
rect 676148 714942 676204 714951
rect 676148 714877 676204 714886
rect 676162 714465 676190 714877
rect 676244 714794 676300 714803
rect 676244 714729 676246 714738
rect 676298 714729 676300 714738
rect 676246 714697 676298 714703
rect 676354 714613 676382 715469
rect 676342 714607 676394 714613
rect 676342 714549 676394 714555
rect 676150 714459 676202 714465
rect 676150 714401 676202 714407
rect 676054 714237 676106 714243
rect 676052 714202 676054 714211
rect 676106 714202 676108 714211
rect 676052 714137 676108 714146
rect 676244 713462 676300 713471
rect 676244 713397 676246 713406
rect 676298 713397 676300 713406
rect 676246 713365 676298 713371
rect 676052 713166 676108 713175
rect 676052 713101 676054 713110
rect 676106 713101 676108 713110
rect 676054 713069 676106 713075
rect 676052 712722 676108 712731
rect 676052 712657 676054 712666
rect 676106 712657 676108 712666
rect 676054 712625 676106 712631
rect 676244 711982 676300 711991
rect 676244 711917 676246 711926
rect 676298 711917 676300 711926
rect 676246 711885 676298 711891
rect 676052 711612 676108 711621
rect 676052 711547 676054 711556
rect 676106 711547 676108 711556
rect 676054 711515 676106 711521
rect 676054 711351 676106 711357
rect 676054 711293 676106 711299
rect 676066 711251 676094 711293
rect 676052 711242 676108 711251
rect 676052 711177 676108 711186
rect 676054 711129 676106 711135
rect 676054 711071 676106 711077
rect 676066 708587 676094 711071
rect 676052 708578 676108 708587
rect 676052 708513 676108 708522
rect 674998 708465 675050 708471
rect 674998 708407 675050 708413
rect 676054 708465 676106 708471
rect 676054 708407 676106 708413
rect 676066 708217 676094 708407
rect 676052 708208 676108 708217
rect 676052 708143 676108 708152
rect 676246 704913 676298 704919
rect 676244 704878 676246 704887
rect 676298 704878 676300 704887
rect 676244 704813 676300 704822
rect 679988 704434 680044 704443
rect 679988 704369 680044 704378
rect 680002 703407 680030 704369
rect 679796 703398 679852 703407
rect 679796 703333 679852 703342
rect 679988 703398 680044 703407
rect 679988 703333 680044 703342
rect 679810 702963 679838 703333
rect 679796 702954 679852 702963
rect 679796 702889 679852 702898
rect 675382 702841 675434 702847
rect 675382 702783 675434 702789
rect 675394 698856 675422 702783
rect 680002 702773 680030 703333
rect 679990 702767 680042 702773
rect 679990 702709 680042 702715
rect 675394 697931 675422 698338
rect 675380 697922 675436 697931
rect 675380 697857 675436 697866
rect 675202 697658 675408 697686
rect 675202 697191 675230 697658
rect 675188 697182 675244 697191
rect 675188 697117 675244 697126
rect 675202 697043 675408 697049
rect 675188 697034 675408 697043
rect 675244 697021 675408 697034
rect 675188 696969 675244 696978
rect 675682 694971 675710 695195
rect 675668 694962 675724 694971
rect 675668 694897 675724 694906
rect 675284 694666 675340 694675
rect 675340 694624 675408 694652
rect 675284 694601 675340 694610
rect 674998 694183 675050 694189
rect 674998 694125 675050 694131
rect 674902 690483 674954 690489
rect 674902 690425 674954 690431
rect 674518 683675 674570 683681
rect 674518 683617 674570 683623
rect 674422 668135 674474 668141
rect 674422 668077 674474 668083
rect 674326 622033 674378 622039
rect 674326 621975 674378 621981
rect 674530 618931 674558 683617
rect 674914 659534 674942 690425
rect 675010 688935 675038 694125
rect 675490 693671 675518 693972
rect 675478 693665 675530 693671
rect 675478 693607 675530 693613
rect 675394 692931 675422 693380
rect 675382 692925 675434 692931
rect 675382 692867 675434 692873
rect 675190 691371 675242 691377
rect 675190 691313 675242 691319
rect 674998 688929 675050 688935
rect 674998 688871 675050 688877
rect 675202 687085 675230 691313
rect 675490 690489 675518 690864
rect 675478 690483 675530 690489
rect 675478 690425 675530 690431
rect 675394 689823 675422 690346
rect 675382 689817 675434 689823
rect 675382 689759 675434 689765
rect 675394 689379 675422 689680
rect 675382 689373 675434 689379
rect 675382 689315 675434 689321
rect 675382 689151 675434 689157
rect 675382 689093 675434 689099
rect 675394 689014 675422 689093
rect 675478 688929 675530 688935
rect 675478 688871 675530 688877
rect 675490 688496 675518 688871
rect 675490 687381 675518 687830
rect 675478 687375 675530 687381
rect 675478 687317 675530 687323
rect 675190 687079 675242 687085
rect 675190 687021 675242 687027
rect 675478 687079 675530 687085
rect 675478 687021 675530 687027
rect 675490 686646 675518 687021
rect 675490 685531 675518 685980
rect 675478 685525 675530 685531
rect 675478 685467 675530 685473
rect 675490 683681 675518 684130
rect 675478 683675 675530 683681
rect 675478 683617 675530 683623
rect 676148 670394 676204 670403
rect 676148 670329 676204 670338
rect 676054 669245 676106 669251
rect 676052 669210 676054 669219
rect 676106 669210 676108 669219
rect 676052 669145 676108 669154
rect 676052 668618 676108 668627
rect 676162 668585 676190 670329
rect 676340 669802 676396 669811
rect 676340 669737 676396 669746
rect 676244 669358 676300 669367
rect 676244 669293 676300 669302
rect 676052 668553 676108 668562
rect 676150 668579 676202 668585
rect 676066 668511 676094 668553
rect 676150 668521 676202 668527
rect 676054 668505 676106 668511
rect 676054 668447 676106 668453
rect 676258 668437 676286 669293
rect 676246 668431 676298 668437
rect 676246 668373 676298 668379
rect 676354 668215 676382 669737
rect 676342 668209 676394 668215
rect 676342 668151 676394 668157
rect 676054 668135 676106 668141
rect 675956 668100 676012 668109
rect 676054 668077 676106 668083
rect 675956 668035 675958 668044
rect 676010 668035 676012 668044
rect 675958 668003 676010 668009
rect 675956 667730 676012 667739
rect 675956 667665 675958 667674
rect 676010 667665 676012 667674
rect 675958 667633 676010 667639
rect 676066 665667 676094 668077
rect 676244 666990 676300 666999
rect 676244 666925 676300 666934
rect 676258 666809 676286 666925
rect 676246 666803 676298 666809
rect 676246 666745 676298 666751
rect 676244 666398 676300 666407
rect 676244 666333 676246 666342
rect 676298 666333 676300 666342
rect 676246 666301 676298 666307
rect 676052 665658 676108 665667
rect 676052 665593 676108 665602
rect 676054 665249 676106 665255
rect 676054 665191 676106 665197
rect 676066 663595 676094 665191
rect 676052 663586 676108 663595
rect 676052 663521 676108 663530
rect 676054 662141 676106 662147
rect 676052 662106 676054 662115
rect 676106 662106 676108 662115
rect 676052 662041 676108 662050
rect 676054 661697 676106 661703
rect 676052 661662 676054 661671
rect 676106 661662 676108 661671
rect 676052 661597 676108 661606
rect 676246 661401 676298 661407
rect 676244 661366 676246 661375
rect 676298 661366 676300 661375
rect 676244 661301 676300 661310
rect 676054 660661 676106 660667
rect 676052 660626 676054 660635
rect 676106 660626 676108 660635
rect 676052 660561 676108 660570
rect 676054 660217 676106 660223
rect 676052 660182 676054 660191
rect 676106 660182 676108 660191
rect 676052 660117 676108 660126
rect 676246 659921 676298 659927
rect 676244 659886 676246 659895
rect 676298 659886 676300 659895
rect 676244 659821 676300 659830
rect 674818 659506 674942 659534
rect 674818 639374 674846 659506
rect 679796 659294 679852 659303
rect 679796 659229 679852 659238
rect 679810 658415 679838 659229
rect 679796 658406 679852 658415
rect 679796 658341 679852 658350
rect 685460 658406 685516 658415
rect 685460 658341 685516 658350
rect 675382 656813 675434 656819
rect 675382 656755 675434 656761
rect 675394 653675 675422 656755
rect 679810 656745 679838 658341
rect 685474 657971 685502 658341
rect 685460 657962 685516 657971
rect 685460 657897 685516 657906
rect 679798 656739 679850 656745
rect 679798 656681 679850 656687
rect 675394 652791 675422 653124
rect 675380 652782 675436 652791
rect 675380 652717 675436 652726
rect 675490 652199 675518 652458
rect 675476 652190 675532 652199
rect 675476 652125 675532 652134
rect 675394 651459 675422 651835
rect 675380 651450 675436 651459
rect 675380 651385 675436 651394
rect 675394 649683 675422 650016
rect 675380 649674 675436 649683
rect 675380 649609 675436 649618
rect 675298 649484 675422 649512
rect 675298 649438 675326 649484
rect 675202 649410 675326 649438
rect 675394 649424 675422 649484
rect 675202 648975 675230 649410
rect 675190 648969 675242 648975
rect 675190 648911 675242 648917
rect 675202 648785 675408 648813
rect 675202 648309 675230 648785
rect 675190 648303 675242 648309
rect 675190 648245 675242 648251
rect 674998 648229 675050 648235
rect 674998 648171 675050 648177
rect 675010 643721 675038 648171
rect 675202 648152 675408 648180
rect 675202 648087 675230 648152
rect 675190 648081 675242 648087
rect 675190 648023 675242 648029
rect 675490 645391 675518 645650
rect 675476 645382 675532 645391
rect 675476 645317 675532 645326
rect 675286 645195 675338 645201
rect 675286 645137 675338 645143
rect 674998 643715 675050 643721
rect 674998 643657 675050 643663
rect 675298 641446 675326 645137
rect 675394 644831 675422 645132
rect 675382 644825 675434 644831
rect 675382 644767 675434 644773
rect 675490 644091 675518 644466
rect 675478 644085 675530 644091
rect 675478 644027 675530 644033
rect 675382 643715 675434 643721
rect 675382 643657 675434 643663
rect 675394 643282 675422 643657
rect 675490 643647 675518 643831
rect 675478 643641 675530 643647
rect 675478 643583 675530 643589
rect 675490 642315 675518 642616
rect 675478 642309 675530 642315
rect 675478 642251 675530 642257
rect 675298 641418 675408 641446
rect 675778 640359 675806 640795
rect 675764 640350 675820 640359
rect 675764 640285 675820 640294
rect 674818 639346 674942 639374
rect 674914 619079 674942 639346
rect 675778 638583 675806 638955
rect 675764 638574 675820 638583
rect 675764 638509 675820 638518
rect 676244 625106 676300 625115
rect 676244 625041 676300 625050
rect 676258 624999 676286 625041
rect 676246 624993 676298 624999
rect 676246 624935 676298 624941
rect 676148 624662 676204 624671
rect 676148 624597 676204 624606
rect 676054 624031 676106 624037
rect 676052 623996 676054 624005
rect 676106 623996 676108 624005
rect 676052 623931 676108 623940
rect 676052 623478 676108 623487
rect 676052 623413 676054 623422
rect 676106 623413 676108 623422
rect 676054 623381 676106 623387
rect 676054 622995 676106 623001
rect 676054 622937 676106 622943
rect 676066 622895 676094 622937
rect 676052 622886 676108 622895
rect 676052 622821 676108 622830
rect 676052 622516 676108 622525
rect 676052 622451 676054 622460
rect 676106 622451 676108 622460
rect 676054 622419 676106 622425
rect 676162 622261 676190 624597
rect 676244 624218 676300 624227
rect 676244 624153 676300 624162
rect 676258 622409 676286 624153
rect 676246 622403 676298 622409
rect 676246 622345 676298 622351
rect 676150 622255 676202 622261
rect 676150 622197 676202 622203
rect 676246 622033 676298 622039
rect 676052 621998 676108 622007
rect 676246 621975 676298 621981
rect 676052 621933 676054 621942
rect 676106 621933 676108 621942
rect 676054 621901 676106 621907
rect 676052 621406 676108 621415
rect 676052 621341 676054 621350
rect 676106 621341 676108 621350
rect 676054 621309 676106 621315
rect 676258 620675 676286 621975
rect 676244 620666 676300 620675
rect 676244 620601 676300 620610
rect 674902 619073 674954 619079
rect 674902 619015 674954 619021
rect 676054 619073 676106 619079
rect 676054 619015 676106 619021
rect 676066 618973 676094 619015
rect 676052 618964 676108 618973
rect 674518 618925 674570 618931
rect 676052 618899 676108 618908
rect 676246 618925 676298 618931
rect 674518 618867 674570 618873
rect 676246 618867 676298 618873
rect 676258 618603 676286 618867
rect 676244 618594 676300 618603
rect 676244 618529 676300 618538
rect 676246 617149 676298 617155
rect 676244 617114 676246 617123
rect 676298 617114 676300 617123
rect 676244 617049 676300 617058
rect 676054 616557 676106 616563
rect 676052 616522 676054 616531
rect 676106 616522 676108 616531
rect 676052 616457 676108 616466
rect 676054 615965 676106 615971
rect 676052 615930 676054 615939
rect 676106 615930 676108 615939
rect 676052 615865 676108 615874
rect 676246 615669 676298 615675
rect 676244 615634 676246 615643
rect 676298 615634 676300 615643
rect 676244 615569 676300 615578
rect 676246 615225 676298 615231
rect 676244 615190 676246 615199
rect 676298 615190 676300 615199
rect 676244 615125 676300 615134
rect 676054 614485 676106 614491
rect 676052 614450 676054 614459
rect 676106 614450 676108 614459
rect 676052 614385 676108 614394
rect 679988 613710 680044 613719
rect 679988 613645 680044 613654
rect 675382 613523 675434 613529
rect 675382 613465 675434 613471
rect 675394 608650 675422 613465
rect 680002 613275 680030 613645
rect 679796 613266 679852 613275
rect 679796 613201 679852 613210
rect 679988 613266 680044 613275
rect 679988 613201 680044 613210
rect 679810 612831 679838 613201
rect 679796 612822 679852 612831
rect 679796 612757 679852 612766
rect 680002 610643 680030 613201
rect 679990 610637 680042 610643
rect 679990 610579 680042 610585
rect 675202 608118 675408 608146
rect 675202 607799 675230 608118
rect 675188 607790 675244 607799
rect 675188 607725 675244 607734
rect 675202 607452 675408 607480
rect 675202 606943 675230 607452
rect 675190 606937 675242 606943
rect 675190 606879 675242 606885
rect 675202 606821 675408 606849
rect 675202 606023 675230 606821
rect 675188 606014 675244 606023
rect 675188 605949 675244 605958
rect 675298 604981 675408 605009
rect 675298 604839 675326 604981
rect 675284 604830 675340 604839
rect 675284 604765 675340 604774
rect 675298 604418 675408 604446
rect 675298 603909 675326 604418
rect 675286 603903 675338 603909
rect 675286 603845 675338 603851
rect 675298 603785 675408 603813
rect 674902 602201 674954 602207
rect 674902 602143 674954 602149
rect 674914 596879 674942 602143
rect 674998 602053 675050 602059
rect 674998 601995 675050 602001
rect 675010 598729 675038 601995
rect 675298 601985 675326 603785
rect 675394 603095 675422 603174
rect 675382 603089 675434 603095
rect 675382 603031 675434 603037
rect 675286 601979 675338 601985
rect 675286 601921 675338 601927
rect 675490 600251 675518 600658
rect 675476 600242 675532 600251
rect 675476 600177 675532 600186
rect 675394 599839 675422 600140
rect 675382 599833 675434 599839
rect 675382 599775 675434 599781
rect 675394 599321 675422 599474
rect 675382 599315 675434 599321
rect 675382 599257 675434 599263
rect 675382 598945 675434 598951
rect 675382 598887 675434 598893
rect 675394 598808 675422 598887
rect 674998 598723 675050 598729
rect 674998 598665 675050 598671
rect 675478 598723 675530 598729
rect 675478 598665 675530 598671
rect 675490 598290 675518 598665
rect 675490 597175 675518 597624
rect 675478 597169 675530 597175
rect 675478 597111 675530 597117
rect 674902 596873 674954 596879
rect 674902 596815 674954 596821
rect 675382 596873 675434 596879
rect 675382 596815 675434 596821
rect 675394 596440 675422 596815
rect 675778 595367 675806 595774
rect 675764 595358 675820 595367
rect 675764 595293 675820 595302
rect 675682 593443 675710 593955
rect 675668 593434 675724 593443
rect 675668 593369 675724 593378
rect 676340 578338 676396 578347
rect 676340 578273 676396 578282
rect 676148 577598 676204 577607
rect 676148 577533 676204 577542
rect 676054 577041 676106 577047
rect 676052 577006 676054 577015
rect 676106 577006 676108 577015
rect 676052 576941 676108 576950
rect 676162 576381 676190 577533
rect 676244 577154 676300 577163
rect 676244 577089 676300 577098
rect 676258 576529 676286 577089
rect 676246 576523 676298 576529
rect 676246 576465 676298 576471
rect 676150 576375 676202 576381
rect 676150 576317 676202 576323
rect 676244 576266 676300 576275
rect 676354 576233 676382 578273
rect 676244 576201 676300 576210
rect 676342 576227 676394 576233
rect 676258 576159 676286 576201
rect 676342 576169 676394 576175
rect 673846 576153 673898 576159
rect 673846 576095 673898 576101
rect 676246 576153 676298 576159
rect 676246 576095 676298 576101
rect 673366 568457 673418 568463
rect 673366 568399 673418 568405
rect 673366 554397 673418 554403
rect 673366 554339 673418 554345
rect 673270 525241 673322 525247
rect 673270 525183 673322 525189
rect 672982 524871 673034 524877
rect 672982 524813 673034 524819
rect 672886 481951 672938 481957
rect 672886 481893 672938 481899
rect 672790 480841 672842 480847
rect 672790 480783 672842 480789
rect 673378 480477 673406 554339
rect 673750 553361 673802 553367
rect 673750 553303 673802 553309
rect 673366 480471 673418 480477
rect 673366 480413 673418 480419
rect 673762 480107 673790 553303
rect 673858 533831 673886 576095
rect 676052 575970 676108 575979
rect 676052 575905 676054 575914
rect 676106 575905 676108 575914
rect 676054 575873 676106 575879
rect 676052 575526 676108 575535
rect 676052 575461 676054 575470
rect 676106 575461 676108 575470
rect 676054 575429 676106 575435
rect 676054 574969 676106 574975
rect 676052 574934 676054 574943
rect 676106 574934 676108 574943
rect 676052 574869 676108 574878
rect 676052 574416 676108 574425
rect 676052 574351 676054 574360
rect 676106 574351 676108 574360
rect 676054 574319 676106 574325
rect 676246 570677 676298 570683
rect 676244 570642 676246 570651
rect 676298 570642 676300 570651
rect 676244 570577 676300 570586
rect 676054 569937 676106 569943
rect 676052 569902 676054 569911
rect 676106 569902 676108 569911
rect 676052 569837 676108 569846
rect 676054 569567 676106 569573
rect 676052 569532 676054 569541
rect 676106 569532 676108 569541
rect 676052 569467 676108 569476
rect 676246 569197 676298 569203
rect 676244 569162 676246 569171
rect 676298 569162 676300 569171
rect 676244 569097 676300 569106
rect 676054 568457 676106 568463
rect 676052 568422 676054 568431
rect 676106 568422 676108 568431
rect 676052 568357 676108 568366
rect 676054 568013 676106 568019
rect 676052 567978 676054 567987
rect 676106 567978 676108 567987
rect 676052 567913 676108 567922
rect 676246 567717 676298 567723
rect 676244 567682 676246 567691
rect 676298 567682 676300 567691
rect 676244 567617 676300 567626
rect 675382 567495 675434 567501
rect 675382 567437 675434 567443
rect 675394 563475 675422 567437
rect 679796 567090 679852 567099
rect 679796 567025 679852 567034
rect 679810 566211 679838 567025
rect 679796 566202 679852 566211
rect 679796 566137 679852 566146
rect 685460 566202 685516 566211
rect 685460 566137 685516 566146
rect 679810 564541 679838 566137
rect 685474 565767 685502 566137
rect 685460 565758 685516 565767
rect 685460 565693 685516 565702
rect 679798 564535 679850 564541
rect 679798 564477 679850 564483
rect 675490 562511 675518 562918
rect 675476 562502 675532 562511
rect 675476 562437 675532 562446
rect 675298 562312 675422 562340
rect 675298 562266 675326 562312
rect 675202 562238 675326 562266
rect 675394 562252 675422 562312
rect 675202 561771 675230 562238
rect 675188 561762 675244 561771
rect 675188 561697 675244 561706
rect 675394 561475 675422 561660
rect 675380 561466 675436 561475
rect 675380 561401 675436 561410
rect 675394 559583 675422 559810
rect 674422 559577 674474 559583
rect 674422 559519 674474 559525
rect 675382 559577 675434 559583
rect 675382 559519 675434 559525
rect 674134 555063 674186 555069
rect 674134 555005 674186 555011
rect 673846 533825 673898 533831
rect 673846 533767 673898 533773
rect 674146 485731 674174 555005
rect 674326 548921 674378 548927
rect 674326 548863 674378 548869
rect 674230 548255 674282 548261
rect 674230 548197 674282 548203
rect 674134 485725 674186 485731
rect 674134 485667 674186 485673
rect 674242 483733 674270 548197
rect 674338 486693 674366 548863
rect 674326 486687 674378 486693
rect 674326 486629 674378 486635
rect 674434 486619 674462 559519
rect 675490 558959 675518 559218
rect 675476 558950 675532 558959
rect 675476 558885 675532 558894
rect 674998 558837 675050 558843
rect 674998 558779 675050 558785
rect 674518 558097 674570 558103
rect 674518 558039 674570 558045
rect 674422 486613 674474 486619
rect 674422 486555 674474 486561
rect 674530 483807 674558 558039
rect 675010 553515 675038 558779
rect 675394 558103 675422 558626
rect 675382 558097 675434 558103
rect 675382 558039 675434 558045
rect 675298 557946 675408 557974
rect 675298 556105 675326 557946
rect 675286 556099 675338 556105
rect 675286 556041 675338 556047
rect 675286 555951 675338 555957
rect 675286 555893 675338 555899
rect 674998 553509 675050 553515
rect 674998 553451 675050 553457
rect 675298 551240 675326 555893
rect 675490 555069 675518 555444
rect 675478 555063 675530 555069
rect 675478 555005 675530 555011
rect 675394 554403 675422 554926
rect 675382 554397 675434 554403
rect 675382 554339 675434 554345
rect 675490 553959 675518 554260
rect 675478 553953 675530 553959
rect 675478 553895 675530 553901
rect 675382 553509 675434 553515
rect 675382 553451 675434 553457
rect 675394 553076 675422 553451
rect 675490 553367 675518 553631
rect 675478 553361 675530 553367
rect 675478 553303 675530 553309
rect 675490 551961 675518 552410
rect 675478 551955 675530 551961
rect 675478 551897 675530 551903
rect 675298 551212 675408 551240
rect 675298 550581 675408 550609
rect 675298 548927 675326 550581
rect 675286 548921 675338 548927
rect 675286 548863 675338 548869
rect 675298 548741 675408 548769
rect 675298 548261 675326 548741
rect 675286 548255 675338 548261
rect 675286 548197 675338 548203
rect 676148 534974 676204 534983
rect 676148 534909 676204 534918
rect 676052 534234 676108 534243
rect 676052 534169 676108 534178
rect 675958 533825 676010 533831
rect 675956 533790 675958 533799
rect 676010 533790 676012 533799
rect 675956 533725 676012 533734
rect 676066 533313 676094 534169
rect 676054 533307 676106 533313
rect 676054 533249 676106 533255
rect 676162 533165 676190 534909
rect 676244 534382 676300 534391
rect 676244 534317 676300 534326
rect 676150 533159 676202 533165
rect 676150 533101 676202 533107
rect 676258 533017 676286 534317
rect 676532 533050 676588 533059
rect 676246 533011 676298 533017
rect 676532 532985 676588 532994
rect 676246 532953 676298 532959
rect 676052 532754 676108 532763
rect 676052 532689 676054 532698
rect 676106 532689 676108 532698
rect 676054 532657 676106 532663
rect 676244 531570 676300 531579
rect 676244 531505 676246 531514
rect 676298 531505 676300 531514
rect 676246 531473 676298 531479
rect 676246 528053 676298 528059
rect 676244 528018 676246 528027
rect 676298 528018 676300 528027
rect 676244 527953 676300 527962
rect 676246 527461 676298 527467
rect 676244 527426 676246 527435
rect 676298 527426 676300 527435
rect 676244 527361 676300 527370
rect 676054 526721 676106 526727
rect 676052 526686 676054 526695
rect 676106 526686 676108 526695
rect 676052 526621 676108 526630
rect 676054 526351 676106 526357
rect 676052 526316 676054 526325
rect 676106 526316 676108 526325
rect 676052 526251 676108 526260
rect 676246 525981 676298 525987
rect 676244 525946 676246 525955
rect 676298 525946 676300 525955
rect 676244 525881 676300 525890
rect 676054 525241 676106 525247
rect 676052 525206 676054 525215
rect 676106 525206 676108 525215
rect 676052 525141 676108 525150
rect 676054 524871 676106 524877
rect 676052 524836 676054 524845
rect 676106 524836 676108 524845
rect 676052 524771 676108 524780
rect 676246 524501 676298 524507
rect 676244 524466 676246 524475
rect 676298 524466 676300 524475
rect 676244 524401 676300 524410
rect 676546 498311 676574 532985
rect 676628 532014 676684 532023
rect 676628 531949 676684 531958
rect 676534 498305 676586 498311
rect 676534 498247 676586 498253
rect 676244 490574 676300 490583
rect 676244 490509 676300 490518
rect 676148 490130 676204 490139
rect 676258 490097 676286 490509
rect 676148 490065 676204 490074
rect 676246 490091 676298 490097
rect 676162 489801 676190 490065
rect 676246 490033 676298 490039
rect 676244 489982 676300 489991
rect 676244 489917 676246 489926
rect 676298 489917 676300 489926
rect 676246 489885 676298 489891
rect 676150 489795 676202 489801
rect 676150 489737 676202 489743
rect 676246 489277 676298 489283
rect 676246 489219 676298 489225
rect 676052 488354 676108 488363
rect 676052 488289 676108 488298
rect 676066 488173 676094 488289
rect 676054 488167 676106 488173
rect 676054 488109 676106 488115
rect 676258 487179 676286 489219
rect 676642 488173 676670 531949
rect 676724 530978 676780 530987
rect 676724 530913 676780 530922
rect 676738 489283 676766 530913
rect 679796 523578 679852 523587
rect 679796 523513 679852 523522
rect 679810 522995 679838 523513
rect 679796 522986 679852 522995
rect 679796 522921 679852 522930
rect 685460 522986 685516 522995
rect 685460 522921 685516 522930
rect 679810 521325 679838 522921
rect 685474 522551 685502 522921
rect 685460 522542 685516 522551
rect 685460 522477 685516 522486
rect 679798 521319 679850 521325
rect 679798 521261 679850 521267
rect 679702 498305 679754 498311
rect 679702 498247 679754 498253
rect 676726 489277 676778 489283
rect 679714 489251 679742 498247
rect 676726 489219 676778 489225
rect 679700 489242 679756 489251
rect 679700 489177 679756 489186
rect 676724 488650 676780 488659
rect 676724 488585 676780 488594
rect 676630 488167 676682 488173
rect 676630 488109 676682 488115
rect 676244 487170 676300 487179
rect 676244 487105 676246 487114
rect 676298 487105 676300 487114
rect 676246 487073 676298 487079
rect 676054 486687 676106 486693
rect 676054 486629 676106 486635
rect 676066 485847 676094 486629
rect 676246 486613 676298 486619
rect 676246 486555 676298 486561
rect 676052 485838 676108 485847
rect 676052 485773 676108 485782
rect 676054 485725 676106 485731
rect 676054 485667 676106 485673
rect 676066 484367 676094 485667
rect 676258 485107 676286 486555
rect 676244 485098 676300 485107
rect 676244 485033 676300 485042
rect 676052 484358 676108 484367
rect 676052 484293 676108 484302
rect 674518 483801 674570 483807
rect 676054 483801 676106 483807
rect 674518 483743 674570 483749
rect 675956 483766 676012 483775
rect 674230 483727 674282 483733
rect 676054 483743 676106 483749
rect 675956 483701 675958 483710
rect 674230 483669 674282 483675
rect 676010 483701 676012 483710
rect 675958 483669 676010 483675
rect 676066 482295 676094 483743
rect 676052 482286 676108 482295
rect 676052 482221 676108 482230
rect 676054 481951 676106 481957
rect 676052 481916 676054 481925
rect 676106 481916 676108 481925
rect 676052 481851 676108 481860
rect 676246 481581 676298 481587
rect 676244 481546 676246 481555
rect 676298 481546 676300 481555
rect 676244 481481 676300 481490
rect 676054 480841 676106 480847
rect 676052 480806 676054 480815
rect 676106 480806 676108 480815
rect 676052 480741 676108 480750
rect 676054 480471 676106 480477
rect 676052 480436 676054 480445
rect 676106 480436 676108 480445
rect 676052 480371 676108 480380
rect 673750 480101 673802 480107
rect 676246 480101 676298 480107
rect 673750 480043 673802 480049
rect 676244 480066 676246 480075
rect 676298 480066 676300 480075
rect 676244 480001 676300 480010
rect 676630 440659 676682 440665
rect 676630 440601 676682 440607
rect 676534 434961 676586 434967
rect 676534 434903 676586 434909
rect 676148 402366 676204 402375
rect 676148 402301 676204 402310
rect 676052 401626 676108 401635
rect 676052 401561 676108 401570
rect 676066 400483 676094 401561
rect 676162 400631 676190 402301
rect 676244 401774 676300 401783
rect 676244 401709 676300 401718
rect 676150 400625 676202 400631
rect 676150 400567 676202 400573
rect 676258 400557 676286 401709
rect 676246 400551 676298 400557
rect 676246 400493 676298 400499
rect 676054 400477 676106 400483
rect 676054 400419 676106 400425
rect 676244 400442 676300 400451
rect 673846 400403 673898 400409
rect 676244 400377 676246 400386
rect 673846 400345 673898 400351
rect 676298 400377 676300 400386
rect 676246 400345 676298 400351
rect 673174 395593 673226 395599
rect 673174 395535 673226 395541
rect 673186 372141 673214 395535
rect 673366 385899 673418 385905
rect 673366 385841 673418 385847
rect 673270 385825 673322 385831
rect 673270 385767 673322 385773
rect 673174 372135 673226 372141
rect 673174 372077 673226 372083
rect 673282 354677 673310 385767
rect 673378 355713 673406 385841
rect 673858 356823 673886 400345
rect 676546 400303 676574 434903
rect 676532 400294 676588 400303
rect 676532 400229 676588 400238
rect 676052 399702 676108 399711
rect 676052 399637 676108 399646
rect 676066 398781 676094 399637
rect 674422 398775 674474 398781
rect 674422 398717 674474 398723
rect 676054 398775 676106 398781
rect 676054 398717 676106 398723
rect 674434 385905 674462 398717
rect 676052 398666 676108 398675
rect 676052 398601 676108 398610
rect 676066 397893 676094 398601
rect 676546 398485 676574 400229
rect 676642 399415 676670 440601
rect 676738 401043 676766 488585
rect 677876 487614 677932 487623
rect 677876 487549 677932 487558
rect 677782 475291 677834 475297
rect 677782 475233 677834 475239
rect 677794 440665 677822 475233
rect 677782 440659 677834 440665
rect 677782 440601 677834 440607
rect 677890 434967 677918 487549
rect 679796 486578 679852 486587
rect 679796 486513 679852 486522
rect 679700 478586 679756 478595
rect 679700 478521 679756 478530
rect 679714 478151 679742 478521
rect 679700 478142 679756 478151
rect 679700 478077 679756 478086
rect 679810 475297 679838 486513
rect 679892 479178 679948 479187
rect 679892 479113 679948 479122
rect 679906 478595 679934 479113
rect 679892 478586 679948 478595
rect 679892 478521 679948 478530
rect 679906 478183 679934 478521
rect 679894 478177 679946 478183
rect 679894 478119 679946 478125
rect 679798 475291 679850 475297
rect 679798 475233 679850 475239
rect 677878 434961 677930 434967
rect 677878 434903 677930 434909
rect 676724 401034 676780 401043
rect 676724 400969 676780 400978
rect 676628 399406 676684 399415
rect 676628 399341 676684 399350
rect 676642 398929 676670 399341
rect 676630 398923 676682 398929
rect 676630 398865 676682 398871
rect 676534 398479 676586 398485
rect 676534 398421 676586 398427
rect 674518 397887 674570 397893
rect 674518 397829 674570 397835
rect 676054 397887 676106 397893
rect 676054 397829 676106 397835
rect 674422 385899 674474 385905
rect 674422 385841 674474 385847
rect 674530 385831 674558 397829
rect 676052 395632 676108 395641
rect 676052 395567 676054 395576
rect 676106 395567 676108 395576
rect 676054 395535 676106 395541
rect 679796 390970 679852 390979
rect 679796 390905 679852 390914
rect 679810 390387 679838 390905
rect 679796 390378 679852 390387
rect 679796 390313 679852 390322
rect 685460 390378 685516 390387
rect 685460 390313 685516 390322
rect 679810 388865 679838 390313
rect 685474 389943 685502 390313
rect 685460 389934 685516 389943
rect 685460 389869 685516 389878
rect 679798 388859 679850 388865
rect 679798 388801 679850 388807
rect 675106 386266 675408 386294
rect 674518 385825 674570 385831
rect 674518 385767 674570 385773
rect 675106 381613 675134 386266
rect 675188 385938 675244 385947
rect 675188 385873 675244 385882
rect 675202 385737 675230 385873
rect 675202 385709 675408 385737
rect 675764 385642 675820 385651
rect 675764 385577 675820 385586
rect 675778 385096 675806 385577
rect 675188 384458 675244 384467
rect 675244 384416 675408 384444
rect 675188 384393 675244 384402
rect 675764 382978 675820 382987
rect 675764 382913 675820 382922
rect 675778 382580 675806 382913
rect 675476 382386 675532 382395
rect 675476 382321 675532 382330
rect 675490 382062 675518 382321
rect 675764 381794 675820 381803
rect 675764 381729 675820 381738
rect 675094 381607 675146 381613
rect 675094 381549 675146 381555
rect 675778 381396 675806 381729
rect 675764 381202 675820 381211
rect 675764 381137 675820 381146
rect 675778 380730 675806 381137
rect 675476 378834 675532 378843
rect 675476 378769 675532 378778
rect 675490 378288 675518 378769
rect 675572 378094 675628 378103
rect 675572 378029 675628 378038
rect 675586 377696 675614 378029
rect 675380 377206 675436 377215
rect 675380 377141 675436 377150
rect 675394 377075 675422 377141
rect 675764 376762 675820 376771
rect 675764 376697 675820 376706
rect 675778 376438 675806 376697
rect 675764 375726 675820 375735
rect 675764 375661 675820 375670
rect 675778 375254 675806 375661
rect 675476 373950 675532 373959
rect 675476 373885 675532 373894
rect 675490 373404 675518 373885
rect 675382 372135 675434 372141
rect 675382 372077 675434 372083
rect 675394 371554 675422 372077
rect 676340 358114 676396 358123
rect 676340 358049 676396 358058
rect 676148 357522 676204 357531
rect 676148 357457 676204 357466
rect 676162 357267 676190 357457
rect 676244 357374 676300 357383
rect 676244 357309 676246 357318
rect 676298 357309 676300 357318
rect 676246 357277 676298 357283
rect 676150 357261 676202 357267
rect 676150 357203 676202 357209
rect 676354 357193 676382 358049
rect 676342 357187 676394 357193
rect 676342 357129 676394 357135
rect 673846 356817 673898 356823
rect 676054 356817 676106 356823
rect 673846 356759 673898 356765
rect 676052 356782 676054 356791
rect 676106 356782 676108 356791
rect 676052 356717 676108 356726
rect 676052 355746 676108 355755
rect 673366 355707 673418 355713
rect 676052 355681 676054 355690
rect 673366 355649 673418 355655
rect 676106 355681 676108 355690
rect 676054 355649 676106 355655
rect 673270 354671 673322 354677
rect 673270 354613 673322 354619
rect 672502 354375 672554 354381
rect 672502 354317 672554 354323
rect 672404 278046 672460 278055
rect 672404 277981 672460 277990
rect 670484 277898 670540 277907
rect 670484 277833 670540 277842
rect 670292 277454 670348 277463
rect 670292 277389 670348 277398
rect 672514 276279 672542 354317
rect 673282 354307 673310 354613
rect 673378 354381 673406 355649
rect 676052 354710 676108 354719
rect 676052 354645 676054 354654
rect 676106 354645 676108 354654
rect 676054 354613 676106 354619
rect 673366 354375 673418 354381
rect 673366 354317 673418 354323
rect 672790 354301 672842 354307
rect 672790 354243 672842 354249
rect 673270 354301 673322 354307
rect 673270 354243 673322 354249
rect 672802 278351 672830 354243
rect 675572 352638 675628 352647
rect 675572 352573 675628 352582
rect 674998 351415 675050 351421
rect 674998 351357 675050 351363
rect 674230 348603 674282 348609
rect 674230 348545 674282 348551
rect 674242 336621 674270 348545
rect 674710 345791 674762 345797
rect 674710 345733 674762 345739
rect 674230 336615 674282 336621
rect 674230 336557 674282 336563
rect 674722 331589 674750 345733
rect 674806 345717 674858 345723
rect 674806 345659 674858 345665
rect 674818 332773 674846 345659
rect 674902 345643 674954 345649
rect 674902 345585 674954 345591
rect 674914 336103 674942 345585
rect 675010 337953 675038 351357
rect 675094 350379 675146 350385
rect 675094 350321 675146 350327
rect 675106 339877 675134 350321
rect 675190 348529 675242 348535
rect 675586 348494 675614 352573
rect 676052 352342 676108 352351
rect 676052 352277 676108 352286
rect 676066 351421 676094 352277
rect 676054 351415 676106 351421
rect 676054 351357 676106 351363
rect 676916 351010 676972 351019
rect 676916 350945 676972 350954
rect 676052 350862 676108 350871
rect 676052 350797 676108 350806
rect 676066 350385 676094 350797
rect 676054 350379 676106 350385
rect 676054 350321 676106 350327
rect 676052 350270 676108 350279
rect 676052 350205 676108 350214
rect 676066 348535 676094 350205
rect 676244 349530 676300 349539
rect 676244 349465 676300 349474
rect 676258 348609 676286 349465
rect 676820 349086 676876 349095
rect 676820 349021 676876 349030
rect 676246 348603 676298 348609
rect 676246 348545 676298 348551
rect 675190 348471 675242 348477
rect 675094 339871 675146 339877
rect 675094 339813 675146 339819
rect 674998 337947 675050 337953
rect 674998 337889 675050 337895
rect 675202 337287 675230 348471
rect 675490 348466 675614 348494
rect 676054 348529 676106 348535
rect 676054 348471 676106 348477
rect 675490 341431 675518 348466
rect 676244 348050 676300 348059
rect 676244 347985 676300 347994
rect 676052 347828 676108 347837
rect 676052 347763 676108 347772
rect 675956 347310 676012 347319
rect 675956 347245 676012 347254
rect 675970 345797 675998 347245
rect 675958 345791 676010 345797
rect 675958 345733 676010 345739
rect 676066 345723 676094 347763
rect 676054 345717 676106 345723
rect 676054 345659 676106 345665
rect 676258 345649 676286 347985
rect 676246 345643 676298 345649
rect 676246 345585 676298 345591
rect 676834 343027 676862 349021
rect 676820 343018 676876 343027
rect 676820 342953 676876 342962
rect 676930 342879 676958 350945
rect 679892 346570 679948 346579
rect 679892 346505 679948 346514
rect 679906 346135 679934 346505
rect 679892 346126 679948 346135
rect 679892 346061 679948 346070
rect 679700 345978 679756 345987
rect 679700 345913 679756 345922
rect 679714 345543 679742 345913
rect 679906 345871 679934 346061
rect 679894 345865 679946 345871
rect 679894 345807 679946 345813
rect 679700 345534 679756 345543
rect 679700 345469 679756 345478
rect 676916 342870 676972 342879
rect 676916 342805 676972 342814
rect 675478 341425 675530 341431
rect 675478 341367 675530 341373
rect 675298 341052 675408 341080
rect 675298 340025 675326 341052
rect 675382 340981 675434 340987
rect 675382 340923 675434 340929
rect 675394 340784 675422 340923
rect 675394 340756 675518 340784
rect 675490 340548 675518 340756
rect 675286 340019 675338 340025
rect 675286 339961 675338 339967
rect 675298 339877 675408 339896
rect 675286 339871 675408 339877
rect 675338 339868 675408 339871
rect 675286 339813 675338 339819
rect 675764 339614 675820 339623
rect 675764 339549 675820 339558
rect 675778 339216 675806 339549
rect 675478 337947 675530 337953
rect 675478 337889 675530 337895
rect 675490 337395 675518 337889
rect 675190 337281 675242 337287
rect 675190 337223 675242 337229
rect 675478 337281 675530 337287
rect 675478 337223 675530 337229
rect 675490 336848 675518 337223
rect 675382 336615 675434 336621
rect 675382 336557 675434 336563
rect 675394 336182 675422 336557
rect 674902 336097 674954 336103
rect 674902 336039 674954 336045
rect 675382 336097 675434 336103
rect 675382 336039 675434 336045
rect 675394 335555 675422 336039
rect 675380 333546 675436 333555
rect 675380 333481 675436 333490
rect 675394 333074 675422 333481
rect 674806 332767 674858 332773
rect 674806 332709 674858 332715
rect 675382 332767 675434 332773
rect 675382 332709 675434 332715
rect 675394 332519 675422 332709
rect 675476 332362 675532 332371
rect 675476 332297 675532 332306
rect 675490 331890 675518 332297
rect 674710 331583 674762 331589
rect 674710 331525 674762 331531
rect 675382 331583 675434 331589
rect 675382 331525 675434 331531
rect 675394 331224 675422 331525
rect 675764 330586 675820 330595
rect 675764 330521 675820 330530
rect 675778 330040 675806 330521
rect 675380 328366 675436 328375
rect 675380 328301 675436 328310
rect 675394 328190 675422 328301
rect 675764 326886 675820 326895
rect 675764 326821 675820 326830
rect 675778 326340 675806 326821
rect 676340 312234 676396 312243
rect 676340 312169 676396 312178
rect 676148 311642 676204 311651
rect 676148 311577 676204 311586
rect 676162 311165 676190 311577
rect 676246 311233 676298 311239
rect 676244 311198 676246 311207
rect 676298 311198 676300 311207
rect 676150 311159 676202 311165
rect 676244 311133 676300 311142
rect 676150 311101 676202 311107
rect 676354 311091 676382 312169
rect 676342 311085 676394 311091
rect 676342 311027 676394 311033
rect 676052 308016 676108 308025
rect 676052 307951 676108 307960
rect 676066 305393 676094 307951
rect 676820 307202 676876 307211
rect 676820 307137 676876 307146
rect 676244 306758 676300 306767
rect 676244 306693 676300 306702
rect 674518 305387 674570 305393
rect 674518 305329 674570 305335
rect 676054 305387 676106 305393
rect 676054 305329 676106 305335
rect 674326 302575 674378 302581
rect 674326 302517 674378 302523
rect 674338 291629 674366 302517
rect 674422 302501 674474 302507
rect 674422 302443 674474 302449
rect 674434 292073 674462 302443
rect 674530 294589 674558 305329
rect 676258 305319 676286 306693
rect 675094 305313 675146 305319
rect 675094 305255 675146 305261
rect 676246 305313 676298 305319
rect 676246 305255 676298 305261
rect 674710 302427 674762 302433
rect 674710 302369 674762 302375
rect 674722 295477 674750 302369
rect 674902 299689 674954 299695
rect 674902 299631 674954 299637
rect 674806 295693 674858 295699
rect 674806 295635 674858 295641
rect 674710 295471 674762 295477
rect 674710 295413 674762 295419
rect 674518 294583 674570 294589
rect 674518 294525 674570 294531
rect 674422 292067 674474 292073
rect 674422 292009 674474 292015
rect 674326 291623 674378 291629
rect 674326 291565 674378 291571
rect 674818 290889 674846 295635
rect 674806 290883 674858 290889
rect 674806 290825 674858 290831
rect 674914 286819 674942 299631
rect 674998 299615 675050 299621
rect 674998 299557 675050 299563
rect 675010 287781 675038 299557
rect 675106 295537 675134 305255
rect 676244 304834 676300 304843
rect 676244 304769 676300 304778
rect 676052 304464 676108 304473
rect 676052 304399 676108 304408
rect 675956 303946 676012 303955
rect 675956 303881 676012 303890
rect 675970 302581 675998 303881
rect 675958 302575 676010 302581
rect 675958 302517 676010 302523
rect 676066 302507 676094 304399
rect 676054 302501 676106 302507
rect 676054 302443 676106 302449
rect 676258 302433 676286 304769
rect 676246 302427 676298 302433
rect 676246 302369 676298 302375
rect 676052 302022 676108 302031
rect 676052 301957 676108 301966
rect 676066 299621 676094 301957
rect 676244 301282 676300 301291
rect 676244 301217 676300 301226
rect 676258 299695 676286 301217
rect 676246 299689 676298 299695
rect 676246 299631 676298 299637
rect 676054 299615 676106 299621
rect 676054 299557 676106 299563
rect 676834 299219 676862 307137
rect 679988 300690 680044 300699
rect 679988 300625 680044 300634
rect 680002 300255 680030 300625
rect 679796 300246 679852 300255
rect 679796 300181 679852 300190
rect 679988 300246 680044 300255
rect 679988 300181 680044 300190
rect 679810 299811 679838 300181
rect 679796 299802 679852 299811
rect 680002 299769 680030 300181
rect 679796 299737 679852 299746
rect 679990 299763 680042 299769
rect 679990 299705 680042 299711
rect 676820 299210 676876 299219
rect 676820 299145 676876 299154
rect 675202 296060 675408 296088
rect 675202 295699 675230 296060
rect 675190 295693 675242 295699
rect 675190 295635 675242 295641
rect 675106 295509 675408 295537
rect 675286 295471 675338 295477
rect 675286 295413 675338 295419
rect 675298 294904 675326 295413
rect 675298 294876 675408 294904
rect 675382 294583 675434 294589
rect 675382 294525 675434 294531
rect 675394 294224 675422 294525
rect 675668 292846 675724 292855
rect 675668 292781 675724 292790
rect 675682 292374 675710 292781
rect 675478 292067 675530 292073
rect 675478 292009 675530 292015
rect 675490 291856 675518 292009
rect 675382 291623 675434 291629
rect 675382 291565 675434 291571
rect 675394 291190 675422 291565
rect 675764 290774 675820 290783
rect 675764 290709 675820 290718
rect 675778 290555 675806 290709
rect 675476 288554 675532 288563
rect 675476 288489 675532 288498
rect 675490 288082 675518 288489
rect 674998 287775 675050 287781
rect 674998 287717 675050 287723
rect 675382 287775 675434 287781
rect 675382 287717 675434 287723
rect 675394 287519 675422 287717
rect 675476 287222 675532 287231
rect 675476 287157 675532 287166
rect 675490 286898 675518 287157
rect 674902 286813 674954 286819
rect 674902 286755 674954 286761
rect 675382 286813 675434 286819
rect 675382 286755 675434 286761
rect 675394 286232 675422 286755
rect 675476 285298 675532 285307
rect 675476 285233 675532 285242
rect 675490 285048 675518 285233
rect 675764 283670 675820 283679
rect 675764 283605 675820 283614
rect 675778 283198 675806 283605
rect 675380 281894 675436 281903
rect 675380 281829 675436 281838
rect 675394 281348 675422 281829
rect 672788 278342 672844 278351
rect 672788 278277 672844 278286
rect 676532 278194 676588 278203
rect 676532 278129 676588 278138
rect 676546 276681 676574 278129
rect 676534 276675 676586 276681
rect 676534 276617 676586 276623
rect 679798 276675 679850 276681
rect 679798 276617 679850 276623
rect 679700 276566 679756 276575
rect 679700 276501 679756 276510
rect 672500 276270 672556 276279
rect 672500 276205 672556 276214
rect 670196 270646 670252 270655
rect 670196 270581 670252 270590
rect 676244 266946 676300 266955
rect 676244 266881 676300 266890
rect 672788 266798 672844 266807
rect 672788 266733 672844 266742
rect 672404 266650 672460 266659
rect 672404 266585 672460 266594
rect 671638 266389 671690 266395
rect 671638 266331 671690 266337
rect 671650 265063 671678 266331
rect 671638 265057 671690 265063
rect 671638 264999 671690 265005
rect 669814 264983 669866 264989
rect 669814 264925 669866 264931
rect 669622 264909 669674 264915
rect 669622 264851 669674 264857
rect 666646 250701 666698 250707
rect 666646 250643 666698 250649
rect 666658 247673 666686 250643
rect 666646 247667 666698 247673
rect 666646 247609 666698 247615
rect 672418 174751 672446 266585
rect 672596 266354 672652 266363
rect 672596 266289 672652 266298
rect 672404 174742 672460 174751
rect 672404 174677 672460 174686
rect 672610 173567 672638 266289
rect 672802 217967 672830 266733
rect 672980 266502 673036 266511
rect 672980 266437 673036 266446
rect 676148 266502 676204 266511
rect 676148 266437 676204 266446
rect 672994 219151 673022 266437
rect 676052 266206 676108 266215
rect 676052 266141 676108 266150
rect 676066 265433 676094 266141
rect 676054 265427 676106 265433
rect 676054 265369 676106 265375
rect 676052 265244 676108 265253
rect 673270 265205 673322 265211
rect 676052 265179 676054 265188
rect 673270 265147 673322 265153
rect 676106 265179 676108 265188
rect 676054 265147 676106 265153
rect 673282 220663 673310 265147
rect 676162 265137 676190 266437
rect 676258 265285 676286 266881
rect 676246 265279 676298 265285
rect 676246 265221 676298 265227
rect 676150 265131 676202 265137
rect 676150 265073 676202 265079
rect 673366 265057 673418 265063
rect 673366 264999 673418 265005
rect 676054 265057 676106 265063
rect 676054 264999 676106 265005
rect 673270 220657 673322 220663
rect 673270 220599 673322 220605
rect 673378 219553 673406 264999
rect 676066 264291 676094 264999
rect 679714 264883 679742 276501
rect 679700 264874 679756 264883
rect 679700 264809 679756 264818
rect 676052 264282 676108 264291
rect 676052 264217 676108 264226
rect 679810 264143 679838 276617
rect 679796 264134 679852 264143
rect 679796 264069 679852 264078
rect 676916 262062 676972 262071
rect 676916 261997 676972 262006
rect 676052 261322 676108 261331
rect 676052 261257 676108 261266
rect 675284 259842 675340 259851
rect 675284 259777 675340 259786
rect 674710 259359 674762 259365
rect 674710 259301 674762 259307
rect 674614 256991 674666 256997
rect 674614 256933 674666 256939
rect 674626 246637 674654 256933
rect 674722 247303 674750 259301
rect 675190 259285 675242 259291
rect 675190 259227 675242 259233
rect 674806 256473 674858 256479
rect 674806 256415 674858 256421
rect 674710 247297 674762 247303
rect 674710 247239 674762 247245
rect 674614 246631 674666 246637
rect 674614 246573 674666 246579
rect 674818 242789 674846 256415
rect 674902 256399 674954 256405
rect 674902 256341 674954 256347
rect 674914 246119 674942 256341
rect 674998 253587 675050 253593
rect 674998 253529 675050 253535
rect 674902 246113 674954 246119
rect 674902 246055 674954 246061
rect 674806 242783 674858 242789
rect 674806 242725 674858 242731
rect 675010 241605 675038 253529
rect 675202 247969 675230 259227
rect 675298 250356 675326 259777
rect 675958 259359 676010 259365
rect 675958 259301 676010 259307
rect 675970 259259 675998 259301
rect 676066 259291 676094 261257
rect 676820 259990 676876 259999
rect 676820 259925 676876 259934
rect 676054 259285 676106 259291
rect 675956 259250 676012 259259
rect 676054 259227 676106 259233
rect 675956 259185 676012 259194
rect 676052 258732 676108 258741
rect 676052 258667 676108 258676
rect 676066 256997 676094 258667
rect 676244 257030 676300 257039
rect 676054 256991 676106 256997
rect 676244 256965 676300 256974
rect 676054 256933 676106 256939
rect 676052 256882 676108 256891
rect 676052 256817 676108 256826
rect 676066 256479 676094 256817
rect 676054 256473 676106 256479
rect 676054 256415 676106 256421
rect 676258 256405 676286 256965
rect 676246 256399 676298 256405
rect 676246 256341 676298 256347
rect 676052 256290 676108 256299
rect 676052 256225 676108 256234
rect 676066 253593 676094 256225
rect 676054 253587 676106 253593
rect 676054 253529 676106 253535
rect 676834 253339 676862 259925
rect 676820 253330 676876 253339
rect 676820 253265 676876 253274
rect 676930 253191 676958 261997
rect 679700 255550 679756 255559
rect 679700 255485 679756 255494
rect 679714 254967 679742 255485
rect 679700 254958 679756 254967
rect 679700 254893 679756 254902
rect 685460 254958 685516 254967
rect 685460 254893 685516 254902
rect 679714 253519 679742 254893
rect 685474 254523 685502 254893
rect 685460 254514 685516 254523
rect 685460 254449 685516 254458
rect 679702 253513 679754 253519
rect 679702 253455 679754 253461
rect 676916 253182 676972 253191
rect 676916 253117 676972 253126
rect 675394 250707 675422 251082
rect 675764 250814 675820 250823
rect 675764 250749 675820 250758
rect 675382 250701 675434 250707
rect 675382 250643 675434 250649
rect 675778 250523 675806 250749
rect 675298 250328 675518 250356
rect 675490 249898 675518 250328
rect 675572 249630 675628 249639
rect 675572 249565 675628 249574
rect 675586 249232 675614 249565
rect 675190 247963 675242 247969
rect 675190 247905 675242 247911
rect 675382 247963 675434 247969
rect 675382 247905 675434 247911
rect 675394 247382 675422 247905
rect 675478 247297 675530 247303
rect 675478 247239 675530 247245
rect 675490 246864 675518 247239
rect 675382 246631 675434 246637
rect 675382 246573 675434 246579
rect 675394 246198 675422 246573
rect 675382 246113 675434 246119
rect 675382 246055 675434 246061
rect 675394 245532 675422 246055
rect 675668 243562 675724 243571
rect 675668 243497 675724 243506
rect 675682 243090 675710 243497
rect 675382 242783 675434 242789
rect 675382 242725 675434 242731
rect 675394 242498 675422 242725
rect 675380 242082 675436 242091
rect 675380 242017 675436 242026
rect 675394 241875 675422 242017
rect 674998 241599 675050 241605
rect 674998 241541 675050 241547
rect 675478 241599 675530 241605
rect 675478 241541 675530 241547
rect 675490 241240 675518 241541
rect 675476 240602 675532 240611
rect 675476 240537 675532 240546
rect 675490 240056 675518 240537
rect 675764 238678 675820 238687
rect 675764 238613 675820 238622
rect 675778 238206 675806 238613
rect 675764 236902 675820 236911
rect 675764 236837 675820 236846
rect 675778 236356 675806 236837
rect 676246 221841 676298 221847
rect 676244 221806 676246 221815
rect 676298 221806 676300 221815
rect 676244 221741 676300 221750
rect 676148 221214 676204 221223
rect 676148 221149 676204 221158
rect 676054 220657 676106 220663
rect 676052 220622 676054 220631
rect 676106 220622 676108 220631
rect 676052 220557 676108 220566
rect 673366 219547 673418 219553
rect 676054 219547 676106 219553
rect 673366 219489 673418 219495
rect 676052 219512 676054 219521
rect 676106 219512 676108 219521
rect 676052 219447 676108 219456
rect 672980 219142 673036 219151
rect 676162 219109 676190 221149
rect 676244 220770 676300 220779
rect 676244 220705 676300 220714
rect 676258 219257 676286 220705
rect 676246 219251 676298 219257
rect 676246 219193 676298 219199
rect 672980 219077 673036 219086
rect 676150 219103 676202 219109
rect 676150 219045 676202 219051
rect 672788 217958 672844 217967
rect 672788 217893 672844 217902
rect 676916 216774 676972 216783
rect 676916 216709 676972 216718
rect 675764 216478 675820 216487
rect 675764 216413 675820 216422
rect 675094 213257 675146 213263
rect 675094 213199 675146 213205
rect 674710 212147 674762 212153
rect 674710 212089 674762 212095
rect 674722 197057 674750 212089
rect 674806 210445 674858 210451
rect 674806 210387 674858 210393
rect 674710 197051 674762 197057
rect 674710 196993 674762 196999
rect 674818 196613 674846 210387
rect 674902 210371 674954 210377
rect 674902 210313 674954 210319
rect 674914 197797 674942 210313
rect 674998 210297 675050 210303
rect 674998 210239 675050 210245
rect 675010 200905 675038 210239
rect 675106 205808 675134 213199
rect 675286 213183 675338 213189
rect 675286 213125 675338 213131
rect 675106 205780 675230 205808
rect 675094 205709 675146 205715
rect 675094 205651 675146 205657
rect 675106 201571 675134 205651
rect 675202 201941 675230 205780
rect 675298 204698 675326 213125
rect 675778 206159 675806 216413
rect 676820 214850 676876 214859
rect 676820 214785 676876 214794
rect 676052 214628 676108 214637
rect 676052 214563 676108 214572
rect 675956 214110 676012 214119
rect 675956 214045 676012 214054
rect 675970 213263 675998 214045
rect 675958 213257 676010 213263
rect 675958 213199 676010 213205
rect 676066 213189 676094 214563
rect 676054 213183 676106 213189
rect 676054 213125 676106 213131
rect 676052 212630 676108 212639
rect 676052 212565 676108 212574
rect 676066 212153 676094 212565
rect 676054 212147 676106 212153
rect 676054 212089 676106 212095
rect 676052 212038 676108 212047
rect 676052 211973 676108 211982
rect 675956 211076 676012 211085
rect 675956 211011 676012 211020
rect 675970 210451 675998 211011
rect 675958 210445 676010 210451
rect 675958 210387 676010 210393
rect 676066 210303 676094 211973
rect 676244 211446 676300 211455
rect 676244 211381 676300 211390
rect 676258 210377 676286 211381
rect 676246 210371 676298 210377
rect 676246 210313 676298 210319
rect 676054 210297 676106 210303
rect 676054 210239 676106 210245
rect 676834 207607 676862 214785
rect 676820 207598 676876 207607
rect 676820 207533 676876 207542
rect 676930 207459 676958 216709
rect 679796 210706 679852 210715
rect 679796 210641 679852 210650
rect 679810 209827 679838 210641
rect 679796 209818 679852 209827
rect 679796 209753 679852 209762
rect 685460 209818 685516 209827
rect 685460 209753 685516 209762
rect 676916 207450 676972 207459
rect 679810 207417 679838 209753
rect 685474 209383 685502 209753
rect 685460 209374 685516 209383
rect 685460 209309 685516 209318
rect 676916 207385 676972 207394
rect 679798 207411 679850 207417
rect 679798 207353 679850 207359
rect 675766 206153 675818 206159
rect 675766 206095 675818 206101
rect 675490 205715 675518 205868
rect 675478 205709 675530 205715
rect 675478 205651 675530 205657
rect 675766 205635 675818 205641
rect 675766 205577 675818 205583
rect 675778 205350 675806 205577
rect 675298 204670 675408 204698
rect 675764 204490 675820 204499
rect 675764 204425 675820 204434
rect 675778 204018 675806 204425
rect 675668 202714 675724 202723
rect 675668 202649 675724 202658
rect 675682 202168 675710 202649
rect 675190 201935 675242 201941
rect 675190 201877 675242 201883
rect 675478 201935 675530 201941
rect 675478 201877 675530 201883
rect 675490 201650 675518 201877
rect 675094 201565 675146 201571
rect 675094 201507 675146 201513
rect 675572 201382 675628 201391
rect 675572 201317 675628 201326
rect 675586 200984 675614 201317
rect 674998 200899 675050 200905
rect 674998 200841 675050 200847
rect 675382 200899 675434 200905
rect 675382 200841 675434 200847
rect 675394 200355 675422 200841
rect 675764 198422 675820 198431
rect 675764 198357 675820 198366
rect 675778 197876 675806 198357
rect 674902 197791 674954 197797
rect 674902 197733 674954 197739
rect 675382 197791 675434 197797
rect 675382 197733 675434 197739
rect 675394 197319 675422 197733
rect 675478 197051 675530 197057
rect 675478 196993 675530 196999
rect 675490 196692 675518 196993
rect 674806 196607 674858 196613
rect 674806 196549 674858 196555
rect 675382 196607 675434 196613
rect 675382 196549 675434 196555
rect 675394 196026 675422 196549
rect 675476 195314 675532 195323
rect 675476 195249 675532 195258
rect 675490 194842 675518 195249
rect 675764 193538 675820 193547
rect 675764 193473 675820 193482
rect 675778 192992 675806 193473
rect 675764 191614 675820 191623
rect 675764 191549 675820 191558
rect 675778 191142 675806 191549
rect 676340 177406 676396 177415
rect 676340 177341 676396 177350
rect 676148 176814 676204 176823
rect 676148 176749 676204 176758
rect 676162 175893 676190 176749
rect 676244 176370 676300 176379
rect 676244 176305 676300 176314
rect 676258 176189 676286 176305
rect 676246 176183 676298 176189
rect 676246 176125 676298 176131
rect 676354 176041 676382 177341
rect 676342 176035 676394 176041
rect 676342 175977 676394 175983
rect 676150 175887 676202 175893
rect 676150 175829 676202 175835
rect 672596 173558 672652 173567
rect 672596 173493 672652 173502
rect 676244 171930 676300 171939
rect 676244 171865 676300 171874
rect 676052 170228 676108 170237
rect 676052 170163 676108 170172
rect 675286 170041 675338 170047
rect 675286 169983 675338 169989
rect 675094 169967 675146 169973
rect 675094 169909 675146 169915
rect 674902 167155 674954 167161
rect 674902 167097 674954 167103
rect 674134 166267 674186 166273
rect 674134 166209 674186 166215
rect 674146 151473 674174 166209
rect 674914 156357 674942 167097
rect 674998 167081 675050 167087
rect 674998 167023 675050 167029
rect 675010 157097 675038 167023
rect 675106 160816 675134 169909
rect 675106 160788 675230 160816
rect 675094 160643 675146 160649
rect 675094 160585 675146 160591
rect 674998 157091 675050 157097
rect 674998 157033 675050 157039
rect 674902 156351 674954 156357
rect 674902 156293 674954 156299
rect 675106 155543 675134 160585
rect 675202 159706 675230 160788
rect 675298 160337 675326 169983
rect 676066 169973 676094 170163
rect 676258 170047 676286 171865
rect 676246 170041 676298 170047
rect 676246 169983 676298 169989
rect 676054 169967 676106 169973
rect 676054 169909 676106 169915
rect 676052 169710 676108 169719
rect 676052 169645 676108 169654
rect 676066 167087 676094 169645
rect 676244 168970 676300 168979
rect 676244 168905 676300 168914
rect 676258 167161 676286 168905
rect 676246 167155 676298 167161
rect 676246 167097 676298 167103
rect 676054 167081 676106 167087
rect 676054 167023 676106 167029
rect 676052 166676 676108 166685
rect 676052 166611 676108 166620
rect 676066 166273 676094 166611
rect 676054 166267 676106 166273
rect 676054 166209 676106 166215
rect 676052 166158 676108 166167
rect 676052 166093 676108 166102
rect 676066 164423 676094 166093
rect 676148 165566 676204 165575
rect 676148 165501 676204 165510
rect 676054 164417 676106 164423
rect 676054 164359 676106 164365
rect 676162 164275 676190 165501
rect 676244 164974 676300 164983
rect 676244 164909 676300 164918
rect 676258 164349 676286 164909
rect 676246 164343 676298 164349
rect 676246 164285 676298 164291
rect 676150 164269 676202 164275
rect 676150 164211 676202 164217
rect 675394 160649 675422 160876
rect 675382 160643 675434 160649
rect 675382 160585 675434 160591
rect 675298 160309 675408 160337
rect 675202 159678 675408 159706
rect 675764 159350 675820 159359
rect 675764 159285 675820 159294
rect 675778 159026 675806 159285
rect 675764 157722 675820 157731
rect 675764 157657 675820 157666
rect 675778 157176 675806 157657
rect 675478 157091 675530 157097
rect 675478 157033 675530 157039
rect 675490 156658 675518 157033
rect 675382 156351 675434 156357
rect 675382 156293 675434 156299
rect 675394 155992 675422 156293
rect 675094 155537 675146 155543
rect 675094 155479 675146 155485
rect 675764 155502 675820 155511
rect 675764 155437 675820 155446
rect 675778 155355 675806 155437
rect 675476 153430 675532 153439
rect 675476 153365 675532 153374
rect 675490 152884 675518 153365
rect 675380 152542 675436 152551
rect 675380 152477 675436 152486
rect 675394 152292 675422 152477
rect 675476 152246 675532 152255
rect 675476 152181 675532 152190
rect 675490 151700 675518 152181
rect 674134 151467 674186 151473
rect 674134 151409 674186 151415
rect 675382 151467 675434 151473
rect 675382 151409 675434 151415
rect 675394 151034 675422 151409
rect 675476 150322 675532 150331
rect 675476 150257 675532 150266
rect 675490 149850 675518 150257
rect 675476 148546 675532 148555
rect 675476 148481 675532 148490
rect 675490 148000 675518 148481
rect 675764 146622 675820 146631
rect 675764 146557 675820 146566
rect 675778 146150 675806 146557
rect 676148 131822 676204 131831
rect 676148 131757 676204 131766
rect 676162 130161 676190 131757
rect 676340 131230 676396 131239
rect 676340 131165 676396 131174
rect 676244 130786 676300 130795
rect 676244 130721 676300 130730
rect 676150 130155 676202 130161
rect 676150 130097 676202 130103
rect 676258 130013 676286 130721
rect 676246 130007 676298 130013
rect 676246 129949 676298 129955
rect 676354 129865 676382 131165
rect 676342 129859 676394 129865
rect 676342 129801 676394 129807
rect 676244 129750 676300 129759
rect 676244 129685 676300 129694
rect 676258 129643 676286 129685
rect 676246 129637 676298 129643
rect 676246 129579 676298 129585
rect 676148 128862 676204 128871
rect 676148 128797 676204 128806
rect 676052 127604 676108 127613
rect 676052 127539 676108 127548
rect 676066 126757 676094 127539
rect 676162 126831 676190 128797
rect 676244 127826 676300 127835
rect 676244 127761 676300 127770
rect 676258 126979 676286 127761
rect 676246 126973 676298 126979
rect 676246 126915 676298 126921
rect 676150 126825 676202 126831
rect 676150 126767 676202 126773
rect 676916 126790 676972 126799
rect 674326 126751 674378 126757
rect 674326 126693 674378 126699
rect 676054 126751 676106 126757
rect 676916 126725 676972 126734
rect 676054 126693 676106 126699
rect 665302 115281 665354 115287
rect 665302 115223 665354 115229
rect 670390 115281 670442 115287
rect 670390 115223 670442 115229
rect 663766 112987 663818 112993
rect 663766 112929 663818 112935
rect 665206 112987 665258 112993
rect 665206 112929 665258 112935
rect 665218 112327 665246 112929
rect 665206 112321 665258 112327
rect 665206 112263 665258 112269
rect 647060 111398 647116 111407
rect 647060 111333 647116 111342
rect 646676 109474 646732 109483
rect 646676 109409 646732 109418
rect 646582 77689 646634 77695
rect 646582 77631 646634 77637
rect 646690 77621 646718 109409
rect 646772 107994 646828 108003
rect 646772 107929 646828 107938
rect 646786 92717 646814 107929
rect 646774 92711 646826 92717
rect 646774 92653 646826 92659
rect 646870 92267 646922 92273
rect 646870 92209 646922 92215
rect 646774 83609 646826 83615
rect 646774 83551 646826 83557
rect 646678 77615 646730 77621
rect 646678 77557 646730 77563
rect 646786 57091 646814 83551
rect 646882 68635 646910 92209
rect 646966 92193 647018 92199
rect 646966 92135 647018 92141
rect 646978 71891 647006 92135
rect 647074 87093 647102 111333
rect 665204 105626 665260 105635
rect 665204 105561 665260 105570
rect 647924 104146 647980 104155
rect 647924 104081 647980 104090
rect 647938 103965 647966 104081
rect 647926 103959 647978 103965
rect 647926 103901 647978 103907
rect 661174 103959 661226 103965
rect 661174 103901 661226 103907
rect 657526 103737 657578 103743
rect 657526 103679 657578 103685
rect 652438 102109 652490 102115
rect 652438 102051 652490 102057
rect 647924 99706 647980 99715
rect 647924 99641 647980 99650
rect 647156 98078 647212 98087
rect 647156 98013 647212 98022
rect 647062 87087 647114 87093
rect 647062 87029 647114 87035
rect 647170 77769 647198 98013
rect 647938 97971 647966 99641
rect 647926 97965 647978 97971
rect 647926 97907 647978 97913
rect 647732 94082 647788 94091
rect 647732 94017 647788 94026
rect 647746 81617 647774 94017
rect 647828 92750 647884 92759
rect 647828 92685 647884 92694
rect 647842 81839 647870 92685
rect 650902 87531 650954 87537
rect 650902 87473 650954 87479
rect 647926 87309 647978 87315
rect 647926 87251 647978 87257
rect 647938 87135 647966 87251
rect 647924 87126 647980 87135
rect 647924 87061 647980 87070
rect 650914 86247 650942 87473
rect 650900 86238 650956 86247
rect 650900 86173 650956 86182
rect 652340 85350 652396 85359
rect 652340 85285 652396 85294
rect 651764 84314 651820 84323
rect 651764 84249 651820 84258
rect 651778 83615 651806 84249
rect 651766 83609 651818 83615
rect 651766 83551 651818 83557
rect 652244 83426 652300 83435
rect 652244 83361 652300 83370
rect 647924 82686 647980 82695
rect 647924 82621 647980 82630
rect 647938 81913 647966 82621
rect 647926 81907 647978 81913
rect 647926 81849 647978 81855
rect 647830 81833 647882 81839
rect 647830 81775 647882 81781
rect 647734 81611 647786 81617
rect 647734 81553 647786 81559
rect 647924 81058 647980 81067
rect 647924 80993 647980 81002
rect 647938 80803 647966 80993
rect 647926 80797 647978 80803
rect 647926 80739 647978 80745
rect 647158 77763 647210 77769
rect 647158 77705 647210 77711
rect 647926 77541 647978 77547
rect 647924 77506 647926 77515
rect 647978 77506 647980 77515
rect 647924 77441 647980 77450
rect 647062 74951 647114 74957
rect 647062 74893 647114 74899
rect 646964 71882 647020 71891
rect 646964 71817 647020 71826
rect 646868 68626 646924 68635
rect 646868 68561 646924 68570
rect 647074 60347 647102 74893
rect 647924 73658 647980 73667
rect 647924 73593 647980 73602
rect 647938 72219 647966 73593
rect 647926 72213 647978 72219
rect 647926 72155 647978 72161
rect 647924 69662 647980 69671
rect 647924 69597 647926 69606
rect 647978 69597 647980 69606
rect 647926 69565 647978 69571
rect 647924 64186 647980 64195
rect 647924 64121 647980 64130
rect 647938 63635 647966 64121
rect 647926 63629 647978 63635
rect 647926 63571 647978 63577
rect 647924 62262 647980 62271
rect 647924 62197 647980 62206
rect 647938 61045 647966 62197
rect 647926 61039 647978 61045
rect 647926 60981 647978 60987
rect 647060 60338 647116 60347
rect 647060 60273 647116 60282
rect 652258 59121 652286 83361
rect 652354 66225 652382 85285
rect 652450 82695 652478 102051
rect 653686 95967 653738 95973
rect 653686 95909 653738 95915
rect 653698 86987 653726 95909
rect 657538 88000 657566 103679
rect 660694 92415 660746 92421
rect 660694 92357 660746 92363
rect 659830 92267 659882 92273
rect 659830 92209 659882 92215
rect 658870 92193 658922 92199
rect 658870 92135 658922 92141
rect 657538 87972 657792 88000
rect 658882 87986 658910 92135
rect 659348 90826 659404 90835
rect 659348 90761 659404 90770
rect 659362 88000 659390 90761
rect 659842 88000 659870 92209
rect 659362 87972 659616 88000
rect 659842 87972 660144 88000
rect 660706 87986 660734 92357
rect 661186 88000 661214 103901
rect 662518 97965 662570 97971
rect 662518 97907 662570 97913
rect 661750 92341 661802 92347
rect 661750 92283 661802 92289
rect 661762 88000 661790 92283
rect 661186 87972 661440 88000
rect 661762 87972 662016 88000
rect 662530 87986 662558 97907
rect 665218 96491 665246 105561
rect 665314 105191 665342 115223
rect 670402 112327 670430 115223
rect 674338 114177 674366 126693
rect 675572 126494 675628 126503
rect 675572 126429 675628 126438
rect 674614 124235 674666 124241
rect 674614 124177 674666 124183
rect 674326 114171 674378 114177
rect 674326 114113 674378 114119
rect 674626 112549 674654 124177
rect 674806 124013 674858 124019
rect 674806 123955 674858 123961
rect 674710 121201 674762 121207
rect 674710 121143 674762 121149
rect 674614 112543 674666 112549
rect 674614 112485 674666 112491
rect 670390 112321 670442 112327
rect 670390 112263 670442 112269
rect 674722 106574 674750 121143
rect 674818 111883 674846 123955
rect 675286 123939 675338 123945
rect 675286 123881 675338 123887
rect 675094 122163 675146 122169
rect 675094 122105 675146 122111
rect 674902 121127 674954 121133
rect 674902 121069 674954 121075
rect 674806 111877 674858 111883
rect 674806 111819 674858 111825
rect 674914 107591 674942 121069
rect 674998 121053 675050 121059
rect 674998 120995 675050 121001
rect 675010 110699 675038 120995
rect 675106 115528 675134 122105
rect 675106 115500 675230 115528
rect 675202 111217 675230 115500
rect 675298 114492 675326 123881
rect 675586 116027 675614 126429
rect 676052 126124 676108 126133
rect 676052 126059 676108 126068
rect 676066 124241 676094 126059
rect 676820 124866 676876 124875
rect 676820 124801 676876 124810
rect 676244 124422 676300 124431
rect 676244 124357 676300 124366
rect 676054 124235 676106 124241
rect 676054 124177 676106 124183
rect 676052 124126 676108 124135
rect 676052 124061 676108 124070
rect 676066 124019 676094 124061
rect 676054 124013 676106 124019
rect 676054 123955 676106 123961
rect 676258 123945 676286 124357
rect 676246 123939 676298 123945
rect 676246 123881 676298 123887
rect 676052 123534 676108 123543
rect 676052 123469 676108 123478
rect 676066 122169 676094 123469
rect 676054 122163 676106 122169
rect 676054 122105 676106 122111
rect 676052 122054 676108 122063
rect 676052 121989 676108 121998
rect 675958 121201 676010 121207
rect 675958 121143 676010 121149
rect 675970 121101 675998 121143
rect 675956 121092 676012 121101
rect 676066 121059 676094 121989
rect 676244 121462 676300 121471
rect 676244 121397 676300 121406
rect 676258 121133 676286 121397
rect 676246 121127 676298 121133
rect 676246 121069 676298 121075
rect 675956 121027 676012 121036
rect 676054 121053 676106 121059
rect 676054 120995 676106 121001
rect 676052 120574 676108 120583
rect 676052 120509 676108 120518
rect 676066 118173 676094 120509
rect 676148 119834 676204 119843
rect 676148 119769 676204 119778
rect 676162 118247 676190 119769
rect 676244 119390 676300 119399
rect 676244 119325 676300 119334
rect 676258 118395 676286 119325
rect 676246 118389 676298 118395
rect 676246 118331 676298 118337
rect 676150 118241 676202 118247
rect 676150 118183 676202 118189
rect 676054 118167 676106 118173
rect 676054 118109 676106 118115
rect 676834 116143 676862 124801
rect 676930 116735 676958 126725
rect 676916 116726 676972 116735
rect 676916 116661 676972 116670
rect 676820 116134 676876 116143
rect 676820 116069 676876 116078
rect 675574 116021 675626 116027
rect 675574 115963 675626 115969
rect 675490 115287 675518 115662
rect 675574 115355 675626 115361
rect 675574 115297 675626 115303
rect 675478 115281 675530 115287
rect 675478 115223 675530 115229
rect 675586 115144 675614 115297
rect 675298 114464 675408 114492
rect 675382 114171 675434 114177
rect 675382 114113 675434 114119
rect 675394 113812 675422 114113
rect 675382 112543 675434 112549
rect 675382 112485 675434 112491
rect 675394 111995 675422 112485
rect 675382 111877 675434 111883
rect 675382 111819 675434 111825
rect 675394 111444 675422 111819
rect 675190 111211 675242 111217
rect 675190 111153 675242 111159
rect 675382 111211 675434 111217
rect 675382 111153 675434 111159
rect 675394 110778 675422 111153
rect 674998 110693 675050 110699
rect 674998 110635 675050 110641
rect 675382 110693 675434 110699
rect 675382 110635 675434 110641
rect 675394 110155 675422 110635
rect 675764 108142 675820 108151
rect 675764 108077 675820 108086
rect 675778 107670 675806 108077
rect 674902 107585 674954 107591
rect 674902 107527 674954 107533
rect 675382 107585 675434 107591
rect 675382 107527 675434 107533
rect 675394 107119 675422 107527
rect 675476 106662 675532 106671
rect 675476 106597 675532 106606
rect 674722 106546 674846 106574
rect 674818 106407 674846 106546
rect 675490 106486 675518 106597
rect 674806 106401 674858 106407
rect 674806 106343 674858 106349
rect 675382 106401 675434 106407
rect 675382 106343 675434 106349
rect 668276 106070 668332 106079
rect 668276 106005 668332 106014
rect 665300 105182 665356 105191
rect 665300 105117 665356 105126
rect 665206 96485 665258 96491
rect 665206 96427 665258 96433
rect 663094 92711 663146 92717
rect 663094 92653 663146 92659
rect 663106 87986 663134 92653
rect 658006 87309 658058 87315
rect 658058 87257 658320 87260
rect 658006 87251 658320 87257
rect 658018 87232 658320 87251
rect 663286 87087 663338 87093
rect 663286 87029 663338 87035
rect 653684 86978 653740 86987
rect 653684 86913 653740 86922
rect 663298 86395 663326 87029
rect 663284 86386 663340 86395
rect 663284 86321 663340 86330
rect 663284 84758 663340 84767
rect 663202 84716 663284 84744
rect 657046 84201 657098 84207
rect 657046 84143 657098 84149
rect 652436 82686 652492 82695
rect 652436 82621 652492 82630
rect 657058 81691 657086 84143
rect 657046 81685 657098 81691
rect 657046 81627 657098 81633
rect 658582 81685 658634 81691
rect 662420 81650 662476 81659
rect 658634 81633 658896 81636
rect 658582 81627 658896 81633
rect 658594 81608 658896 81627
rect 662420 81585 662422 81594
rect 662474 81585 662476 81594
rect 662422 81553 662474 81559
rect 656962 81016 657216 81044
rect 657538 81016 657792 81044
rect 656962 77547 656990 81016
rect 656950 77541 657002 77547
rect 656950 77483 657002 77489
rect 657538 76141 657566 81016
rect 658306 77769 658334 81030
rect 659602 80748 659630 81030
rect 659554 80729 659630 80748
rect 659446 80723 659498 80729
rect 659446 80665 659498 80671
rect 659542 80723 659630 80729
rect 659594 80720 659630 80723
rect 659542 80665 659594 80671
rect 658294 77763 658346 77769
rect 658294 77705 658346 77711
rect 659458 77695 659486 80665
rect 659446 77689 659498 77695
rect 659446 77631 659498 77637
rect 657526 76135 657578 76141
rect 657526 76077 657578 76083
rect 660130 74957 660158 81030
rect 660118 74951 660170 74957
rect 660118 74893 660170 74899
rect 660706 72219 660734 81030
rect 661440 81016 661502 81044
rect 660694 72213 660746 72219
rect 660694 72155 660746 72161
rect 661474 69629 661502 81016
rect 661762 81016 662016 81044
rect 661762 77621 661790 81016
rect 662530 80803 662558 81030
rect 662518 80797 662570 80803
rect 662518 80739 662570 80745
rect 661750 77615 661802 77621
rect 661750 77557 661802 77563
rect 661462 69623 661514 69629
rect 661462 69565 661514 69571
rect 652342 66219 652394 66225
rect 652342 66161 652394 66167
rect 663202 63635 663230 84716
rect 663284 84693 663340 84702
rect 663476 84018 663532 84027
rect 663476 83953 663532 83962
rect 663380 82834 663436 82843
rect 663380 82769 663436 82778
rect 663284 82094 663340 82103
rect 663284 82029 663340 82038
rect 663298 81913 663326 82029
rect 663286 81907 663338 81913
rect 663286 81849 663338 81855
rect 663394 81839 663422 82769
rect 663382 81833 663434 81839
rect 663382 81775 663434 81781
rect 663190 63629 663242 63635
rect 663190 63571 663242 63577
rect 663490 61045 663518 83953
rect 663478 61039 663530 61045
rect 663478 60981 663530 60987
rect 652246 59115 652298 59121
rect 652246 59057 652298 59063
rect 646772 57082 646828 57091
rect 646772 57017 646828 57026
rect 646484 54714 646540 54723
rect 646484 54649 646540 54658
rect 668290 53201 668318 106005
rect 675394 105820 675422 106343
rect 675380 105182 675436 105191
rect 675380 105117 675436 105126
rect 675394 104636 675422 105117
rect 675764 103258 675820 103267
rect 675764 103193 675820 103202
rect 675778 102786 675806 103193
rect 675764 101482 675820 101491
rect 675764 101417 675820 101426
rect 675778 100936 675806 101417
rect 668278 53195 668330 53201
rect 668278 53137 668330 53143
rect 633622 49051 633674 49057
rect 633622 48993 633674 48999
rect 640726 49051 640778 49057
rect 640726 48993 640778 48999
rect 562486 47941 562538 47947
rect 562486 47883 562538 47889
rect 539734 46239 539786 46245
rect 539734 46181 539786 46187
rect 545206 46239 545258 46245
rect 545206 46181 545258 46187
rect 512180 41838 512236 41847
rect 525908 41838 525964 41847
rect 514882 41805 515136 41824
rect 512180 41773 512236 41782
rect 514006 41799 514058 41805
rect 514006 41741 514058 41747
rect 514870 41799 515136 41805
rect 514922 41796 515136 41799
rect 525964 41796 526176 41824
rect 525908 41773 525964 41782
rect 514870 41741 514922 41747
rect 514018 37439 514046 41741
rect 539746 40515 539774 46181
rect 633634 43285 633662 48993
rect 629014 43279 629066 43285
rect 629014 43221 629066 43227
rect 633622 43279 633674 43285
rect 633622 43221 633674 43227
rect 629026 42027 629054 43221
rect 629014 42021 629066 42027
rect 629014 41963 629066 41969
rect 539732 40506 539788 40515
rect 539732 40441 539788 40450
rect 475510 37433 475562 37439
rect 475510 37375 475562 37381
rect 514006 37433 514058 37439
rect 514006 37375 514058 37381
rect 420790 34547 420842 34553
rect 420790 34489 420842 34495
rect 444886 34547 444938 34553
rect 444886 34489 444938 34495
rect 328342 31661 328394 31667
rect 311156 31626 311212 31635
rect 311156 31561 311212 31570
rect 328340 31626 328342 31635
rect 335446 31661 335498 31667
rect 328394 31626 328396 31635
rect 335446 31603 335498 31609
rect 328340 31561 328396 31570
<< via2 >>
rect 81140 1002302 81196 1002358
rect 184052 1002319 184108 1002358
rect 184052 1002302 184054 1002319
rect 184054 1002302 184106 1002319
rect 184106 1002302 184108 1002319
rect 482612 1002319 482668 1002358
rect 482612 1002302 482614 1002319
rect 482614 1002302 482666 1002319
rect 482666 1002302 482668 1002319
rect 132404 997122 132460 997178
rect 241172 997122 241228 997178
rect 80564 982914 80620 982970
rect 132404 982914 132460 982970
rect 184244 982914 184300 982970
rect 233204 982914 233260 982970
rect 240884 982953 240886 982970
rect 240886 982953 240938 982970
rect 240938 982953 240940 982970
rect 240884 982914 240940 982953
rect 241172 982914 241228 982970
rect 290804 997122 290860 997178
rect 290804 983210 290860 983266
rect 394580 997714 394636 997770
rect 397460 983210 397516 983266
rect 292148 983062 292204 983118
rect 535700 997714 535756 997770
rect 636500 997714 636556 997770
rect 636500 983062 636556 983118
rect 285044 982914 285100 982970
rect 391604 982931 391660 982970
rect 391604 982914 391606 982931
rect 391606 982914 391658 982931
rect 391658 982914 391660 982931
rect 394580 982914 394636 982970
rect 483860 982914 483916 982970
rect 538580 982914 538636 982970
rect 40148 959234 40204 959290
rect 60020 959103 60076 959142
rect 60020 959086 60022 959103
rect 60022 959086 60074 959103
rect 60074 959086 60076 959103
rect 653780 959086 653836 959142
rect 676820 950371 676876 950410
rect 676820 950354 676822 950371
rect 676822 950354 676874 950371
rect 676874 950354 676876 950371
rect 676148 894114 676204 894170
rect 676052 893374 676108 893430
rect 655220 868806 655276 868862
rect 655124 866438 655180 866494
rect 676244 893522 676300 893578
rect 676052 892429 676108 892468
rect 676052 892412 676054 892429
rect 676054 892412 676106 892429
rect 676106 892412 676108 892429
rect 655412 867622 655468 867678
rect 655316 865254 655372 865310
rect 654164 863922 654220 863978
rect 653780 862886 653836 862942
rect 41780 817933 41782 817950
rect 41782 817933 41834 817950
rect 41834 817933 41836 817950
rect 41780 817894 41836 817933
rect 41780 817319 41836 817358
rect 41780 817302 41782 817319
rect 41782 817302 41834 817319
rect 41834 817302 41836 817319
rect 41588 816579 41644 816618
rect 41588 816562 41590 816579
rect 41590 816562 41642 816579
rect 41642 816562 41644 816579
rect 41780 815839 41836 815878
rect 41780 815822 41782 815839
rect 41782 815822 41834 815839
rect 41834 815822 41836 815839
rect 41780 814877 41836 814916
rect 41780 814860 41782 814877
rect 41782 814860 41834 814877
rect 41834 814860 41836 814877
rect 41588 813619 41644 813658
rect 41588 813602 41590 813619
rect 41590 813602 41642 813619
rect 41642 813602 41644 813619
rect 41588 813158 41644 813214
rect 40244 812418 40300 812474
rect 42548 812862 42604 812918
rect 28820 805610 28876 805666
rect 28820 805166 28876 805222
rect 41588 811678 41644 811734
rect 41972 811308 42028 811364
rect 41876 810790 41932 810846
rect 41780 809845 41836 809884
rect 41780 809828 41782 809845
rect 41782 809828 41834 809845
rect 41834 809828 41836 809845
rect 41780 808866 41836 808922
rect 41684 808126 41740 808182
rect 41588 806663 41644 806702
rect 41588 806646 41590 806663
rect 41590 806646 41642 806663
rect 41642 806646 41644 806663
rect 41588 806054 41644 806110
rect 41588 805183 41644 805222
rect 41588 805166 41590 805183
rect 41590 805166 41642 805183
rect 41642 805166 41644 805183
rect 40244 802058 40300 802114
rect 41780 807403 41836 807442
rect 41780 807386 41782 807403
rect 41782 807386 41834 807403
rect 41834 807386 41836 807403
rect 41684 800430 41740 800486
rect 42068 809310 42124 809366
rect 42164 807830 42220 807886
rect 42068 800430 42124 800486
rect 41972 800282 42028 800338
rect 42740 800874 42796 800930
rect 41780 794214 41836 794270
rect 42740 793474 42796 793530
rect 41972 792882 42028 792938
rect 42164 790070 42220 790126
rect 42836 789330 42892 789386
rect 42740 789182 42796 789238
rect 41780 774695 41836 774734
rect 41780 774678 41782 774695
rect 41782 774678 41834 774695
rect 41834 774678 41836 774695
rect 41588 773955 41644 773994
rect 41588 773938 41590 773955
rect 41590 773938 41642 773955
rect 41642 773938 41644 773955
rect 41588 773363 41644 773402
rect 41588 773346 41590 773363
rect 41590 773346 41642 773363
rect 41642 773346 41644 773363
rect 41780 773237 41782 773254
rect 41782 773237 41834 773254
rect 41834 773237 41836 773254
rect 41780 773198 41836 773237
rect 41588 772902 41644 772958
rect 41780 772623 41836 772662
rect 41780 772606 41782 772623
rect 41782 772606 41834 772623
rect 41834 772606 41836 772623
rect 42740 771905 42742 771922
rect 42742 771905 42794 771922
rect 42794 771905 42796 771922
rect 42740 771866 42796 771905
rect 41588 770830 41644 770886
rect 41396 769942 41452 769998
rect 40244 768906 40300 768962
rect 28820 762394 28876 762450
rect 28820 761950 28876 762006
rect 40244 759878 40300 759934
rect 41972 769646 42028 769702
rect 41684 768462 41740 768518
rect 41492 766390 41548 766446
rect 41588 763447 41644 763486
rect 41588 763430 41590 763447
rect 41590 763430 41642 763447
rect 41642 763430 41644 763447
rect 41780 768183 41836 768222
rect 41780 768166 41782 768183
rect 41782 768166 41834 768183
rect 41834 768166 41836 768183
rect 41876 767574 41932 767630
rect 41780 765149 41836 765188
rect 41780 765132 41782 765149
rect 41782 765132 41834 765149
rect 41834 765132 41836 765149
rect 41780 764187 41836 764226
rect 41780 764170 41782 764187
rect 41782 764170 41834 764187
rect 41834 764170 41836 764187
rect 41780 762115 41836 762154
rect 41780 762098 41782 762115
rect 41782 762098 41834 762115
rect 41834 762098 41836 762115
rect 41684 757362 41740 757418
rect 42068 766094 42124 766150
rect 42164 765650 42220 765706
rect 42836 757806 42892 757862
rect 42068 757214 42124 757270
rect 41972 757066 42028 757122
rect 41972 754846 42028 754902
rect 42932 751294 42988 751350
rect 42452 747742 42508 747798
rect 41780 747446 41836 747502
rect 42164 746854 42220 746910
rect 42356 746558 42412 746614
rect 42932 747150 42988 747206
rect 41780 731479 41836 731518
rect 41780 731462 41782 731479
rect 41782 731462 41834 731479
rect 41834 731462 41836 731479
rect 41588 730739 41644 730778
rect 41588 730722 41590 730739
rect 41590 730722 41642 730739
rect 41642 730722 41644 730739
rect 41780 730369 41836 730408
rect 41780 730352 41782 730369
rect 41782 730352 41834 730369
rect 41834 730352 41836 730369
rect 41588 730169 41590 730186
rect 41590 730169 41642 730186
rect 41642 730169 41644 730186
rect 41588 730130 41644 730169
rect 41396 729242 41452 729298
rect 41588 729259 41644 729298
rect 41588 729242 41590 729259
rect 41590 729242 41642 729259
rect 41642 729242 41644 729259
rect 40436 728689 40438 728706
rect 40438 728689 40490 728706
rect 40490 728689 40492 728706
rect 40436 728650 40492 728689
rect 41780 728815 41836 728854
rect 41780 728798 41782 728815
rect 41782 728798 41834 728815
rect 41834 728798 41836 728815
rect 41780 727927 41836 727966
rect 41780 727910 41782 727927
rect 41782 727910 41834 727927
rect 41834 727910 41836 727927
rect 41492 726726 41548 726782
rect 34388 725690 34444 725746
rect 28820 719178 28876 719234
rect 28820 718734 28876 718790
rect 34484 723766 34540 723822
rect 34388 716662 34444 716718
rect 34484 716070 34540 716126
rect 42068 726430 42124 726486
rect 41972 725468 42028 725524
rect 41780 724358 41836 724414
rect 41684 722286 41740 722342
rect 41588 721694 41644 721750
rect 41588 720231 41644 720270
rect 41588 720214 41590 720231
rect 41590 720214 41642 720231
rect 41642 720214 41644 720231
rect 41588 718751 41644 718790
rect 41588 718734 41590 718751
rect 41590 718734 41642 718751
rect 41642 718734 41644 718751
rect 41492 714146 41548 714202
rect 41876 722917 41878 722934
rect 41878 722917 41930 722934
rect 41930 722917 41932 722934
rect 41876 722878 41932 722917
rect 41972 713998 42028 714054
rect 42164 724950 42220 725006
rect 42452 723470 42508 723526
rect 42068 713850 42124 713906
rect 42452 712222 42508 712278
rect 42068 711630 42124 711686
rect 43028 711630 43084 711686
rect 42932 711482 42988 711538
rect 42932 711186 42988 711242
rect 42452 708818 42508 708874
rect 41780 707338 41836 707394
rect 43028 711038 43084 711094
rect 42932 707930 42988 707986
rect 42932 705118 42988 705174
rect 42356 704822 42412 704878
rect 41780 699938 41836 699994
rect 43028 703490 43084 703546
rect 41780 688263 41836 688302
rect 41780 688246 41782 688263
rect 41782 688246 41834 688263
rect 41834 688246 41836 688263
rect 41588 687523 41644 687562
rect 41588 687506 41590 687523
rect 41590 687506 41642 687523
rect 41642 687506 41644 687523
rect 41780 687227 41836 687266
rect 41780 687210 41782 687227
rect 41782 687210 41834 687227
rect 41834 687210 41836 687227
rect 41588 686953 41590 686970
rect 41590 686953 41642 686970
rect 41642 686953 41644 686970
rect 41588 686914 41644 686953
rect 41588 686043 41644 686082
rect 41588 686026 41590 686043
rect 41590 686026 41642 686043
rect 41642 686026 41644 686043
rect 43316 711334 43372 711390
rect 41780 685325 41782 685342
rect 41782 685325 41834 685342
rect 41834 685325 41836 685342
rect 41780 685286 41836 685325
rect 43700 711334 43756 711390
rect 41780 684141 41782 684158
rect 41782 684141 41834 684158
rect 41834 684141 41836 684158
rect 41780 684102 41836 684141
rect 41972 683806 42028 683862
rect 41780 683214 41836 683270
rect 34388 682474 34444 682530
rect 28820 675962 28876 676018
rect 28820 675518 28876 675574
rect 37364 682030 37420 682086
rect 34484 679514 34540 679570
rect 34388 672410 34444 672466
rect 41876 681734 41932 681790
rect 41780 681142 41836 681198
rect 39764 680550 39820 680606
rect 39860 679958 39916 680014
rect 41588 679070 41644 679126
rect 41684 677590 41740 677646
rect 41588 677015 41644 677054
rect 41588 676998 41590 677015
rect 41590 676998 41642 677015
rect 41642 676998 41644 677015
rect 41588 675535 41644 675574
rect 41588 675518 41590 675535
rect 41590 675518 41642 675535
rect 41642 675518 41644 675535
rect 39764 671078 39820 671134
rect 42068 678774 42124 678830
rect 42260 678182 42316 678238
rect 41972 670634 42028 670690
rect 42740 665010 42796 665066
rect 42836 662346 42892 662402
rect 42932 660718 42988 660774
rect 43028 658794 43084 658850
rect 41588 644899 41644 644938
rect 41588 644882 41590 644899
rect 41590 644882 41642 644899
rect 41642 644882 41644 644899
rect 41492 644734 41548 644790
rect 41588 644307 41644 644346
rect 41588 644290 41590 644307
rect 41590 644290 41642 644307
rect 41642 644290 41644 644307
rect 41780 644011 41836 644050
rect 41780 643994 41782 644011
rect 41782 643994 41834 644011
rect 41834 643994 41836 644011
rect 41588 643737 41590 643754
rect 41590 643737 41642 643754
rect 41642 643737 41644 643754
rect 41588 643698 41644 643737
rect 41588 642827 41644 642866
rect 41588 642810 41590 642827
rect 41590 642810 41642 642827
rect 41642 642810 41644 642827
rect 41588 641347 41644 641386
rect 41588 641330 41590 641347
rect 41590 641330 41642 641347
rect 41642 641330 41644 641347
rect 41492 641182 41548 641238
rect 37364 640294 37420 640350
rect 34484 639258 34540 639314
rect 34388 636742 34444 636798
rect 28820 632746 28876 632802
rect 28820 632302 28876 632358
rect 34484 629194 34540 629250
rect 41972 639998 42028 640054
rect 40148 638814 40204 638870
rect 41684 638666 41740 638722
rect 40244 637334 40300 637390
rect 41588 635262 41644 635318
rect 41588 634374 41644 634430
rect 41876 637926 41932 637982
rect 41780 636076 41836 636132
rect 41780 634078 41836 634134
rect 41588 632319 41644 632358
rect 41588 632302 41590 632319
rect 41590 632302 41642 632319
rect 41642 632302 41644 632319
rect 40244 628306 40300 628362
rect 41780 627418 41836 627474
rect 42164 636446 42220 636502
rect 42068 627566 42124 627622
rect 42260 634966 42316 635022
rect 42164 627418 42220 627474
rect 42740 625198 42796 625254
rect 42836 622090 42892 622146
rect 42836 619130 42892 619186
rect 42740 616466 42796 616522
rect 42356 616318 42412 616374
rect 40340 601666 40396 601722
rect 41588 601683 41644 601722
rect 41588 601666 41590 601683
rect 41590 601666 41642 601683
rect 41642 601666 41644 601683
rect 41780 601387 41836 601426
rect 41780 601370 41782 601387
rect 41782 601370 41834 601387
rect 41834 601370 41836 601387
rect 41780 600795 41836 600834
rect 41780 600778 41782 600795
rect 41782 600778 41834 600795
rect 41834 600778 41836 600795
rect 41780 600373 41782 600390
rect 41782 600373 41834 600390
rect 41834 600373 41836 600390
rect 41780 600334 41836 600373
rect 41780 599833 41836 599872
rect 41780 599816 41782 599833
rect 41782 599816 41834 599833
rect 41834 599816 41836 599833
rect 40340 599446 40396 599502
rect 41780 599315 41836 599354
rect 41780 599298 41782 599315
rect 41782 599298 41834 599315
rect 41834 599298 41836 599315
rect 40340 598706 40396 598762
rect 41780 598353 41836 598392
rect 41780 598336 41782 598353
rect 41782 598336 41834 598353
rect 41834 598336 41836 598353
rect 41780 597857 41782 597874
rect 41782 597857 41834 597874
rect 41834 597857 41836 597874
rect 41780 597818 41836 597857
rect 37364 597078 37420 597134
rect 34292 596042 34348 596098
rect 28820 589530 28876 589586
rect 28820 589086 28876 589142
rect 34388 594118 34444 594174
rect 34484 593082 34540 593138
rect 34388 585682 34444 585738
rect 34292 585238 34348 585294
rect 41588 596651 41644 596690
rect 41588 596634 41590 596651
rect 41590 596634 41642 596651
rect 41642 596634 41644 596651
rect 40148 595598 40204 595654
rect 41972 595302 42028 595358
rect 41780 594784 41836 594840
rect 40244 593674 40300 593730
rect 41588 591027 41644 591066
rect 41588 591010 41590 591027
rect 41590 591010 41642 591027
rect 41642 591010 41644 591027
rect 41588 589086 41644 589142
rect 41876 592934 41932 592990
rect 41876 584202 41932 584258
rect 42068 592342 42124 592398
rect 42260 591750 42316 591806
rect 42164 591306 42220 591362
rect 42260 584794 42316 584850
rect 42260 584202 42316 584258
rect 42548 578282 42604 578338
rect 42356 575322 42412 575378
rect 41876 572658 41932 572714
rect 43028 578726 43084 578782
rect 43124 573990 43180 574046
rect 41780 539802 41836 539858
rect 41780 538026 41836 538082
rect 41780 536250 41836 536306
rect 41780 535066 41836 535122
rect 41780 534178 41836 534234
rect 41780 533882 41836 533938
rect 41780 533142 41836 533198
rect 41780 530774 41836 530830
rect 41876 530034 41932 530090
rect 42068 529294 42124 529350
rect 42164 528702 42220 528758
rect 42164 527074 42220 527130
rect 41780 476053 41782 476070
rect 41782 476053 41834 476070
rect 41834 476053 41836 476070
rect 41780 476014 41836 476053
rect 41780 475535 41782 475552
rect 41782 475535 41834 475552
rect 41834 475535 41836 475552
rect 41780 475496 41836 475535
rect 41780 474978 41836 475034
rect 40436 473794 40492 473850
rect 39668 473202 39724 473258
rect 37364 470686 37420 470742
rect 34484 464322 34540 464378
rect 23060 463730 23116 463786
rect 23060 463286 23116 463342
rect 39764 472314 39820 472370
rect 41876 474573 41878 474590
rect 41878 474573 41930 474590
rect 41930 474573 41932 474590
rect 41876 474534 41932 474573
rect 41588 472166 41644 472222
rect 43412 473054 43468 473110
rect 41588 468762 41644 468818
rect 41780 463599 41836 463638
rect 41780 463582 41782 463599
rect 41782 463582 41834 463599
rect 41834 463582 41836 463599
rect 41588 426895 41644 426934
rect 41588 426878 41590 426895
rect 41590 426878 41642 426895
rect 41642 426878 41644 426895
rect 41780 426525 41836 426564
rect 41780 426508 41782 426525
rect 41782 426508 41834 426525
rect 41834 426508 41836 426525
rect 41780 426007 41836 426046
rect 41780 425990 41782 426007
rect 41782 425990 41834 426007
rect 41834 425990 41836 426007
rect 40436 425250 40492 425306
rect 41588 424823 41644 424862
rect 41588 424806 41590 424823
rect 41590 424806 41642 424823
rect 41642 424806 41644 424823
rect 34484 424214 34540 424270
rect 39668 424214 39724 424270
rect 41780 423491 41836 423530
rect 41780 423474 41782 423491
rect 41782 423474 41834 423491
rect 41834 423474 41836 423491
rect 41588 422751 41644 422790
rect 41588 422734 41590 422751
rect 41590 422734 41642 422751
rect 41642 422734 41644 422751
rect 34484 421698 34540 421754
rect 39764 420810 39820 420866
rect 39668 419182 39724 419238
rect 39668 416370 39724 416426
rect 39956 420218 40012 420274
rect 39860 419774 39916 419830
rect 40244 418738 40300 418794
rect 40052 418294 40108 418350
rect 39956 416814 40012 416870
rect 40148 417850 40204 417906
rect 40244 417258 40300 417314
rect 41588 416370 41644 416426
rect 40052 416222 40108 416278
rect 39764 414890 39820 414946
rect 23060 414742 23116 414798
rect 23060 414298 23116 414354
rect 41588 414315 41644 414354
rect 41588 414298 41590 414315
rect 41590 414298 41642 414315
rect 41642 414298 41644 414315
rect 41876 416074 41932 416130
rect 41876 411190 41932 411246
rect 41780 407638 41836 407694
rect 42068 406010 42124 406066
rect 41780 403790 41836 403846
rect 42164 403050 42220 403106
rect 41876 402606 41932 402662
rect 41780 401866 41836 401922
rect 41780 400090 41836 400146
rect 41780 399350 41836 399406
rect 41780 398758 41836 398814
rect 41780 388694 41836 388750
rect 41780 386326 41836 386382
rect 41588 385921 41590 385938
rect 41590 385921 41642 385938
rect 41642 385921 41644 385938
rect 41588 385882 41644 385921
rect 41588 385307 41644 385346
rect 41588 385290 41590 385307
rect 41590 385290 41642 385307
rect 41642 385290 41644 385307
rect 41588 384737 41590 384754
rect 41590 384737 41642 384754
rect 41642 384737 41644 384754
rect 41588 384698 41644 384737
rect 41588 383827 41644 383866
rect 41588 383810 41590 383827
rect 41590 383810 41642 383827
rect 41642 383810 41644 383827
rect 34484 383218 34540 383274
rect 41876 385011 41932 385050
rect 41876 384994 41878 385011
rect 41878 384994 41930 385011
rect 41930 384994 41932 385011
rect 41780 383070 41836 383126
rect 41588 382347 41644 382386
rect 41588 382330 41590 382347
rect 41590 382330 41642 382347
rect 41642 382330 41644 382347
rect 41780 381999 41782 382016
rect 41782 381999 41834 382016
rect 41834 381999 41836 382016
rect 41780 381960 41836 381999
rect 39188 381294 39244 381350
rect 34484 378778 34540 378834
rect 28820 373746 28876 373802
rect 28820 373302 28876 373358
rect 39284 380850 39340 380906
rect 39476 379222 39532 379278
rect 40052 378334 40108 378390
rect 39764 377742 39820 377798
rect 39284 373746 39340 373802
rect 39956 377298 40012 377354
rect 42452 376854 42508 376910
rect 41492 376262 41548 376318
rect 41684 375226 41740 375282
rect 41588 374782 41644 374838
rect 40052 373894 40108 373950
rect 39956 373302 40012 373358
rect 39764 373154 39820 373210
rect 39188 372266 39244 372322
rect 41780 374486 41836 374542
rect 41780 373541 41836 373580
rect 41780 373524 41782 373541
rect 41782 373524 41834 373541
rect 41834 373524 41836 373541
rect 41780 368122 41836 368178
rect 41780 362794 41836 362850
rect 41780 360574 41836 360630
rect 41972 359834 42028 359890
rect 42068 359242 42124 359298
rect 41780 358798 41836 358854
rect 41876 356874 41932 356930
rect 41780 356134 41836 356190
rect 42164 355542 42220 355598
rect 41684 343110 41740 343166
rect 41588 340611 41644 340650
rect 41588 340594 41590 340611
rect 41590 340594 41642 340611
rect 41642 340594 41644 340611
rect 41780 342831 41836 342870
rect 41780 342814 41782 342831
rect 41782 342814 41834 342831
rect 41834 342814 41836 342831
rect 41780 342313 41836 342352
rect 41780 342296 41782 342313
rect 41782 342296 41834 342313
rect 41834 342296 41836 342313
rect 41780 341795 41836 341834
rect 41780 341778 41782 341795
rect 41782 341778 41834 341795
rect 41834 341778 41836 341795
rect 41780 341373 41782 341390
rect 41782 341373 41834 341390
rect 41834 341373 41836 341390
rect 41780 341334 41836 341373
rect 41780 340315 41836 340354
rect 41780 340298 41782 340315
rect 41782 340298 41834 340315
rect 41834 340298 41836 340315
rect 41684 340002 41740 340058
rect 41588 339131 41644 339170
rect 41588 339114 41590 339131
rect 41590 339114 41642 339131
rect 41642 339114 41644 339131
rect 41780 338818 41836 338874
rect 28724 338078 28780 338134
rect 39764 337634 39820 337690
rect 39284 337042 39340 337098
rect 41780 335710 41836 335766
rect 41492 333638 41548 333694
rect 41396 333046 41452 333102
rect 39764 331122 39820 331178
rect 41588 331566 41644 331622
rect 39284 330678 39340 330734
rect 28820 330530 28876 330586
rect 28820 330086 28876 330142
rect 28724 329050 28780 329106
rect 41876 331270 41932 331326
rect 41876 330399 41932 330438
rect 41876 330382 41878 330399
rect 41878 330382 41930 330399
rect 41930 330382 41932 330399
rect 41780 324906 41836 324962
rect 41780 320466 41836 320522
rect 41780 319726 41836 319782
rect 41876 317358 41932 317414
rect 41780 316618 41836 316674
rect 41780 316174 41836 316230
rect 41780 315434 41836 315490
rect 42068 313658 42124 313714
rect 41780 313066 41836 313122
rect 42164 312474 42220 312530
rect 39668 298710 39724 298766
rect 28724 294862 28780 294918
rect 41780 299615 41836 299654
rect 41780 299598 41782 299615
rect 41782 299598 41834 299615
rect 41834 299598 41836 299615
rect 41780 299171 41836 299210
rect 41780 299154 41782 299171
rect 41782 299154 41834 299171
rect 41834 299154 41836 299171
rect 41780 298157 41782 298174
rect 41782 298157 41834 298174
rect 41834 298157 41836 298174
rect 41780 298118 41836 298157
rect 41780 297617 41836 297656
rect 41780 297600 41782 297617
rect 41782 297600 41834 297617
rect 41834 297600 41836 297617
rect 41780 297099 41836 297138
rect 41780 297082 41782 297099
rect 41782 297082 41834 297099
rect 41834 297082 41836 297099
rect 39764 296490 39820 296546
rect 39956 295898 40012 295954
rect 41588 295915 41644 295954
rect 41588 295898 41590 295915
rect 41590 295898 41642 295915
rect 41642 295898 41644 295915
rect 41780 292568 41836 292624
rect 41492 290422 41548 290478
rect 28820 287314 28876 287370
rect 28820 286870 28876 286926
rect 41684 288794 41740 288850
rect 41588 288350 41644 288406
rect 28724 285094 28780 285150
rect 42452 290126 42508 290182
rect 41876 287183 41932 287222
rect 41876 287166 41878 287183
rect 41878 287166 41930 287183
rect 41930 287166 41932 287183
rect 41876 281690 41932 281746
rect 42452 281542 42508 281598
rect 42164 277990 42220 278046
rect 41780 276510 41836 276566
rect 41780 274142 41836 274198
rect 41780 273550 41836 273606
rect 41780 272810 41836 272866
rect 41780 272366 41836 272422
rect 42068 270590 42124 270646
rect 41780 269998 41836 270054
rect 41876 269258 41932 269314
rect 23156 254162 23212 254218
rect 23060 253274 23116 253330
rect 43316 263486 43372 263542
rect 40244 256234 40300 256290
rect 41588 255642 41644 255698
rect 41780 255385 41782 255402
rect 41782 255385 41834 255402
rect 41834 255385 41836 255402
rect 41780 255346 41836 255385
rect 41780 254941 41782 254958
rect 41782 254941 41834 254958
rect 41834 254941 41836 254958
rect 41780 254902 41836 254941
rect 41780 254475 41836 254514
rect 41780 254458 41782 254475
rect 41782 254458 41834 254475
rect 41834 254458 41836 254475
rect 23348 253274 23404 253330
rect 23252 252682 23308 252738
rect 41876 249426 41932 249482
rect 41684 247206 41740 247262
rect 41300 246762 41356 246818
rect 41396 245578 41452 245634
rect 41492 245134 41548 245190
rect 41588 244690 41644 244746
rect 41588 243654 41644 243710
rect 41780 244855 41836 244894
rect 41780 244838 41782 244855
rect 41782 244838 41834 244855
rect 41834 244838 41836 244855
rect 41780 237882 41836 237938
rect 41780 233294 41836 233350
rect 41780 231074 41836 231130
rect 41780 230334 41836 230390
rect 41780 229742 41836 229798
rect 41780 229002 41836 229058
rect 41780 227374 41836 227430
rect 41780 226634 41836 226690
rect 42068 226190 42124 226246
rect 41780 213279 41782 213296
rect 41782 213279 41834 213296
rect 41834 213279 41836 213296
rect 41780 213240 41836 213279
rect 41588 212909 41590 212926
rect 41590 212909 41642 212926
rect 41642 212909 41644 212926
rect 41588 212870 41644 212909
rect 41780 212169 41782 212186
rect 41782 212169 41834 212186
rect 41834 212169 41836 212186
rect 41780 212130 41836 212169
rect 41780 211725 41782 211742
rect 41782 211725 41834 211742
rect 41834 211725 41836 211742
rect 41780 211686 41836 211725
rect 41588 211429 41590 211446
rect 41590 211429 41642 211446
rect 41642 211429 41644 211446
rect 41588 211390 41644 211429
rect 41780 210689 41782 210706
rect 41782 210689 41834 210706
rect 41834 210689 41836 210706
rect 41780 210650 41836 210689
rect 41780 210223 41836 210262
rect 43508 266890 43564 266946
rect 41780 210206 41782 210223
rect 41782 210206 41834 210223
rect 41834 210206 41836 210223
rect 41588 209949 41590 209966
rect 41590 209949 41642 209966
rect 41642 209949 41644 209966
rect 41588 209910 41644 209949
rect 57716 790810 57772 790866
rect 57620 789626 57676 789682
rect 58196 788442 58252 788498
rect 58388 787258 58444 787314
rect 59636 785482 59692 785538
rect 59156 784890 59212 784946
rect 45236 702010 45292 702066
rect 44756 275326 44812 275382
rect 44660 267038 44716 267094
rect 45236 473054 45292 473110
rect 45140 278286 45196 278342
rect 45236 276214 45292 276270
rect 45044 274142 45100 274198
rect 45332 273550 45388 273606
rect 44852 263042 44908 263098
rect 41588 209357 41590 209374
rect 41590 209357 41642 209374
rect 41642 209357 41644 209374
rect 41588 209318 41644 209357
rect 25556 208430 25612 208486
rect 25748 207986 25804 208042
rect 25652 206358 25708 206414
rect 25556 199994 25612 200050
rect 25844 207838 25900 207894
rect 41972 206210 42028 206266
rect 41684 203990 41740 204046
rect 41492 202510 41548 202566
rect 41588 202066 41644 202122
rect 25844 200882 25900 200938
rect 41492 200921 41494 200938
rect 41494 200921 41546 200938
rect 41546 200921 41548 200938
rect 41492 200882 41548 200921
rect 25748 200438 25804 200494
rect 25652 199550 25708 199606
rect 41780 203694 41836 203750
rect 41876 201661 41878 201678
rect 41878 201661 41930 201678
rect 41930 201661 41932 201678
rect 41876 201622 41932 201661
rect 41876 201365 41878 201382
rect 41878 201365 41930 201382
rect 41930 201365 41932 201382
rect 41876 201326 41932 201365
rect 41780 195258 41836 195314
rect 58676 747594 58732 747650
rect 54740 745983 54796 746022
rect 54740 745966 54742 745983
rect 54742 745966 54794 745983
rect 54794 745966 54796 745983
rect 54644 745818 54700 745874
rect 59636 745374 59692 745430
rect 57620 745226 57676 745282
rect 58196 744042 58252 744098
rect 59636 742858 59692 742914
rect 59732 741674 59788 741730
rect 59636 704378 59692 704434
rect 58772 702641 58774 702658
rect 58774 702641 58826 702658
rect 58826 702641 58828 702658
rect 58772 702602 58828 702641
rect 58676 700826 58732 700882
rect 59252 699642 59308 699698
rect 58868 698458 58924 698514
rect 59636 661162 59692 661218
rect 58772 659425 58774 659442
rect 58774 659425 58826 659442
rect 58826 659425 58828 659442
rect 58772 659386 58828 659425
rect 58676 657610 58732 657666
rect 58196 656426 58252 656482
rect 58388 655242 58444 655298
rect 58964 617946 59020 618002
rect 58196 615578 58252 615634
rect 59636 616209 59638 616226
rect 59638 616209 59690 616226
rect 59690 616209 59692 616226
rect 59636 616170 59692 616209
rect 58964 614394 59020 614450
rect 59636 613210 59692 613266
rect 59540 612026 59596 612082
rect 41780 190078 41836 190134
rect 41876 187858 41932 187914
rect 42164 187118 42220 187174
rect 41780 186378 41836 186434
rect 41780 185786 41836 185842
rect 41780 184158 41836 184214
rect 41780 183418 41836 183474
rect 42068 182974 42124 183030
rect 50420 275178 50476 275234
rect 50612 275030 50668 275086
rect 58964 574730 59020 574786
rect 58196 572362 58252 572418
rect 59636 572993 59638 573010
rect 59638 572993 59690 573010
rect 59690 572993 59692 573010
rect 59636 572954 59692 572993
rect 58964 571178 59020 571234
rect 59348 569994 59404 570050
rect 59540 568810 59596 568866
rect 57716 531662 57772 531718
rect 57620 530478 57676 530534
rect 58196 529294 58252 529350
rect 58964 527074 59020 527130
rect 58580 525890 58636 525946
rect 59348 524706 59404 524762
rect 58484 404086 58540 404142
rect 59348 402310 59404 402366
rect 57716 400534 57772 400590
rect 59636 399942 59692 399998
rect 59732 399350 59788 399406
rect 59540 398166 59596 398222
rect 59252 360870 59308 360926
rect 59156 359686 59212 359742
rect 57620 357466 57676 357522
rect 58196 356134 58252 356190
rect 59636 356726 59692 356782
rect 58580 354950 58636 355006
rect 58484 317654 58540 317710
rect 59156 316470 59212 316526
rect 59348 314102 59404 314158
rect 58196 312918 58252 312974
rect 59636 313510 59692 313566
rect 59732 311734 59788 311790
rect 59636 295158 59692 295214
rect 58388 292790 58444 292846
rect 58772 292642 58828 292698
rect 60308 293974 60364 294030
rect 60212 291458 60268 291514
rect 58004 289551 58060 289590
rect 58004 289534 58006 289551
rect 58006 289534 58058 289551
rect 58058 289534 58060 289551
rect 59636 288071 59692 288110
rect 59636 288054 59638 288071
rect 59638 288054 59690 288071
rect 59690 288054 59692 288071
rect 58964 286870 59020 286926
rect 59060 285686 59116 285742
rect 57620 284502 57676 284558
rect 58964 282430 59020 282486
rect 59636 283318 59692 283374
rect 59540 280950 59596 281006
rect 59348 279766 59404 279822
rect 61940 278138 61996 278194
rect 62132 536990 62188 537046
rect 62132 276066 62188 276122
rect 62036 266594 62092 266650
rect 62324 277842 62380 277898
rect 64724 386326 64780 386382
rect 62612 343110 62668 343166
rect 62612 277990 62668 278046
rect 62804 277694 62860 277750
rect 62996 277546 63052 277602
rect 64724 277398 64780 277454
rect 62516 270590 62572 270646
rect 65876 269258 65932 269314
rect 70580 272070 70636 272126
rect 69428 269554 69484 269610
rect 72980 272218 73036 272274
rect 71732 269406 71788 269462
rect 78836 272366 78892 272422
rect 77588 269702 77644 269758
rect 62420 266742 62476 266798
rect 62228 266446 62284 266502
rect 61844 266298 61900 266354
rect 88340 272514 88396 272570
rect 91892 272662 91948 272718
rect 139124 269850 139180 269906
rect 148340 244542 148396 244598
rect 148244 239658 148300 239714
rect 147860 232258 147916 232314
rect 146900 229890 146956 229946
rect 147092 226338 147148 226394
rect 147284 221454 147340 221510
rect 147284 214071 147340 214110
rect 147284 214054 147286 214071
rect 147286 214054 147338 214071
rect 147338 214054 147340 214071
rect 146900 212887 146956 212926
rect 146900 212870 146902 212887
rect 146902 212870 146954 212887
rect 146954 212870 146956 212887
rect 147092 211686 147148 211742
rect 147476 210371 147532 210410
rect 147476 210354 147478 210371
rect 147478 210354 147530 210371
rect 147530 210354 147532 210371
rect 146900 209170 146956 209226
rect 147188 207986 147244 208042
rect 147092 206358 147148 206414
rect 147476 199550 147532 199606
rect 147380 190966 147436 191022
rect 147764 176462 147820 176518
rect 148724 243358 148780 243414
rect 148532 242026 148588 242082
rect 148436 238474 148492 238530
rect 148628 233590 148684 233646
rect 148532 169062 148588 169118
rect 148340 168026 148396 168082
rect 148244 164326 148300 164382
rect 147476 159442 147532 159498
rect 146900 156926 146956 156982
rect 147668 146122 147724 146178
rect 147476 144494 147532 144550
rect 147476 143606 147532 143662
rect 147668 142439 147724 142478
rect 147668 142422 147670 142439
rect 147670 142422 147722 142439
rect 147722 142422 147724 142439
rect 147476 139906 147532 139962
rect 147476 138722 147532 138778
rect 147476 130286 147532 130342
rect 147476 127918 147532 127974
rect 148436 166250 148492 166306
rect 148340 122442 148396 122498
rect 147860 120535 147916 120574
rect 147860 120518 147862 120535
rect 147862 120518 147914 120535
rect 147914 120518 147916 120535
rect 148244 111934 148300 111990
rect 147188 108382 147244 108438
rect 149012 240842 149068 240898
rect 148916 236698 148972 236754
rect 148820 234774 148876 234830
rect 149108 235958 149164 236014
rect 149396 231074 149452 231130
rect 149396 228114 149452 228170
rect 149396 227374 149452 227430
rect 149492 225154 149548 225210
rect 149492 223822 149548 223878
rect 149396 222638 149452 222694
rect 149492 219678 149548 219734
rect 149396 218955 149452 218994
rect 149396 218938 149398 218955
rect 149398 218938 149450 218955
rect 149450 218938 149452 218955
rect 149396 217754 149452 217810
rect 149492 216570 149548 216626
rect 149396 214942 149452 214998
rect 149396 205618 149452 205674
rect 149300 204434 149356 204490
rect 149492 203250 149548 203306
rect 149396 201918 149452 201974
rect 149396 200734 149452 200790
rect 149492 198366 149548 198422
rect 149396 197034 149452 197090
rect 149396 195867 149452 195906
rect 149396 195850 149398 195867
rect 149398 195850 149450 195867
rect 149450 195850 149452 195867
rect 149492 194666 149548 194722
rect 149396 193334 149452 193390
rect 149396 192150 149452 192206
rect 149396 189782 149452 189838
rect 149300 187414 149356 187470
rect 149204 186230 149260 186286
rect 149492 188006 149548 188062
rect 149396 183714 149452 183770
rect 149588 184454 149644 184510
rect 149492 182530 149548 182586
rect 149300 181346 149356 181402
rect 149492 179570 149548 179626
rect 149396 178830 149452 178886
rect 149396 177646 149452 177702
rect 149396 175130 149452 175186
rect 149108 173946 149164 174002
rect 149012 170246 149068 170302
rect 148724 165510 148780 165566
rect 148628 161810 148684 161866
rect 148916 163142 148972 163198
rect 148820 160626 148876 160682
rect 149588 172762 149644 172818
rect 149492 170986 149548 171042
rect 149300 157666 149356 157722
rect 149396 155742 149452 155798
rect 148532 121702 148588 121758
rect 148436 107198 148492 107254
rect 148820 133838 148876 133894
rect 149012 132654 149068 132710
rect 148820 115190 148876 115246
rect 148628 109583 148684 109622
rect 148628 109566 148630 109583
rect 148630 109566 148682 109583
rect 148682 109566 148684 109583
rect 148820 106014 148876 106070
rect 148628 104682 148684 104738
rect 148724 103498 148780 103554
rect 149300 154558 149356 154614
rect 149396 153078 149452 153134
rect 149204 152042 149260 152098
rect 149396 150858 149452 150914
rect 149300 149822 149356 149878
rect 149300 148490 149356 148546
rect 149396 147306 149452 147362
rect 149684 141255 149740 141294
rect 149684 141238 149686 141255
rect 149686 141238 149738 141255
rect 149738 141238 149740 141255
rect 149588 137538 149644 137594
rect 149684 135910 149740 135966
rect 149684 135022 149740 135078
rect 149684 130878 149740 130934
rect 149108 129102 149164 129158
rect 149300 126586 149356 126642
rect 148916 102314 148972 102370
rect 148820 86495 148876 86534
rect 148820 86478 148822 86495
rect 148822 86478 148874 86495
rect 148874 86478 148876 86495
rect 149588 125402 149644 125458
rect 149396 124235 149452 124274
rect 149396 124218 149398 124235
rect 149398 124218 149450 124235
rect 149450 124218 149452 124235
rect 149492 119334 149548 119390
rect 149396 118189 149398 118206
rect 149398 118189 149450 118206
rect 149450 118189 149452 118206
rect 149396 118150 149452 118189
rect 149492 116818 149548 116874
rect 149396 115634 149452 115690
rect 149396 115190 149452 115246
rect 149396 114450 149452 114506
rect 149396 113118 149452 113174
rect 149396 110898 149452 110954
rect 149396 100851 149452 100890
rect 149396 100834 149398 100851
rect 149398 100834 149450 100851
rect 149450 100834 149452 100851
rect 149492 99798 149548 99854
rect 149396 98614 149452 98670
rect 149492 97430 149548 97486
rect 149396 95654 149452 95710
rect 149588 94914 149644 94970
rect 149492 93730 149548 93786
rect 149396 92546 149452 92602
rect 149300 91362 149356 91418
rect 148820 85294 148876 85350
rect 147092 84110 147148 84166
rect 148436 81594 148492 81650
rect 149108 82334 149164 82390
rect 148916 77894 148972 77950
rect 149396 90178 149452 90234
rect 149396 88994 149452 89050
rect 149492 87218 149548 87274
rect 149588 80410 149644 80466
rect 149396 76710 149452 76766
rect 149204 75526 149260 75582
rect 149012 73010 149068 73066
rect 149108 71974 149164 72030
rect 149300 73750 149356 73806
rect 149684 79226 149740 79282
rect 184340 219530 184396 219586
rect 184340 218829 184342 218846
rect 184342 218829 184394 218846
rect 184394 218829 184396 218846
rect 184340 218790 184396 218829
rect 184340 199698 184396 199754
rect 184244 197626 184300 197682
rect 194420 272218 194476 272274
rect 193748 272070 193804 272126
rect 193076 269554 193132 269610
rect 192404 269258 192460 269314
rect 185588 220270 185644 220326
rect 185492 198218 185548 198274
rect 184436 196738 184492 196794
rect 184340 195998 184396 196054
rect 184340 195258 184396 195314
rect 184436 194370 184492 194426
rect 184532 193778 184588 193834
rect 184436 192890 184492 192946
rect 184340 192298 184396 192354
rect 184532 191410 184588 191466
rect 184628 190670 184684 190726
rect 184340 189969 184342 189986
rect 184342 189969 184394 189986
rect 184394 189969 184396 189986
rect 184340 189930 184396 189969
rect 184340 188450 184396 188506
rect 184532 189190 184588 189246
rect 184436 187562 184492 187618
rect 184340 186822 184396 186878
rect 184436 186082 184492 186138
rect 184628 185342 184684 185398
rect 184532 184602 184588 184658
rect 184340 183862 184396 183918
rect 184436 181494 184492 181550
rect 184340 180754 184396 180810
rect 184436 180014 184492 180070
rect 184628 179274 184684 179330
rect 184532 178534 184588 178590
rect 184436 177646 184492 177702
rect 184340 177054 184396 177110
rect 184532 176166 184588 176222
rect 184340 175613 184342 175630
rect 184342 175613 184394 175630
rect 184394 175613 184396 175630
rect 184340 175574 184396 175613
rect 184436 173946 184492 174002
rect 184340 171726 184396 171782
rect 184532 172466 184588 172522
rect 184436 170838 184492 170894
rect 184628 170246 184684 170302
rect 184340 169358 184396 169414
rect 184532 168618 184588 168674
rect 184436 167878 184492 167934
rect 184628 167138 184684 167194
rect 184340 166398 184396 166454
rect 184436 165658 184492 165714
rect 184532 164770 184588 164826
rect 184340 164047 184396 164086
rect 184340 164030 184342 164047
rect 184342 164030 184394 164047
rect 184394 164030 184396 164047
rect 184340 162550 184396 162606
rect 184532 163290 184588 163346
rect 184436 161810 184492 161866
rect 184436 160922 184492 160978
rect 184532 160330 184588 160386
rect 184340 159442 184396 159498
rect 184628 158850 184684 158906
rect 184340 157962 184396 158018
rect 184436 157370 184492 157426
rect 184532 156482 184588 156538
rect 184628 155594 184684 155650
rect 186068 211982 186124 212038
rect 185972 204286 186028 204342
rect 186356 210502 186412 210558
rect 186260 207246 186316 207302
rect 186548 213462 186604 213518
rect 186932 221010 186988 221066
rect 187124 243358 187180 243414
rect 187028 218050 187084 218106
rect 186836 216422 186892 216478
rect 186740 214942 186796 214998
rect 186644 209022 186700 209078
rect 186452 205914 186508 205970
rect 186164 202806 186220 202862
rect 194228 269406 194284 269462
rect 196628 272366 196684 272422
rect 196148 269702 196204 269758
rect 199220 272514 199276 272570
rect 200468 272662 200524 272718
rect 209684 270442 209740 270498
rect 213332 269850 213388 269906
rect 214292 270442 214348 270498
rect 341684 274290 341740 274346
rect 347636 274438 347692 274494
rect 350228 274586 350284 274642
rect 353396 274734 353452 274790
rect 370100 271922 370156 271978
rect 369620 271774 369676 271830
rect 367892 269110 367948 269166
rect 368372 268962 368428 269018
rect 374324 270442 374380 270498
rect 375572 273402 375628 273458
rect 377012 270294 377068 270350
rect 379124 274882 379180 274938
rect 378644 273254 378700 273310
rect 383444 275918 383500 275974
rect 382964 273106 383020 273162
rect 385556 270146 385612 270202
rect 388436 269998 388492 270054
rect 390356 275770 390412 275826
rect 390164 272958 390220 273014
rect 391508 269850 391564 269906
rect 392756 272810 392812 272866
rect 395156 276510 395212 276566
rect 397076 268814 397132 268870
rect 398900 275622 398956 275678
rect 398708 272662 398764 272718
rect 402548 276658 402604 276714
rect 403028 269702 403084 269758
rect 404180 272514 404236 272570
rect 405428 276806 405484 276862
rect 405620 269554 405676 269610
rect 407828 275474 407884 275530
rect 407252 272366 407308 272422
rect 410900 272218 410956 272274
rect 410420 269406 410476 269462
rect 411764 272070 411820 272126
rect 411572 269258 411628 269314
rect 474836 274290 474892 274346
rect 489044 274438 489100 274494
rect 496052 274586 496108 274642
rect 503156 274734 503212 274790
rect 522548 276806 522604 276862
rect 523796 268814 523852 268870
rect 529844 276658 529900 276714
rect 539828 269110 539884 269166
rect 540980 268962 541036 269018
rect 544532 271922 544588 271978
rect 543380 271774 543436 271830
rect 558740 273402 558796 273458
rect 555188 270442 555244 270498
rect 566996 274882 567052 274938
rect 565844 273254 565900 273310
rect 562292 270294 562348 270350
rect 577652 275918 577708 275974
rect 576500 273106 576556 273162
rect 583604 270146 583660 270202
rect 595412 275770 595468 275826
rect 594164 272958 594220 273014
rect 590612 269998 590668 270054
rect 601268 272810 601324 272866
rect 597716 269850 597772 269906
rect 607220 276510 607276 276566
rect 616628 275622 616684 275678
rect 615476 272662 615532 272718
rect 626132 269702 626188 269758
rect 629684 272514 629740 272570
rect 633236 269554 633292 269610
rect 637940 275474 637996 275530
rect 636788 272366 636844 272422
rect 646484 275326 646540 275382
rect 646196 272218 646252 272274
rect 645044 269406 645100 269462
rect 420404 262171 420460 262210
rect 420404 262154 420406 262171
rect 420406 262154 420458 262171
rect 420458 262154 420460 262171
rect 420404 259786 420460 259842
rect 191540 259342 191596 259398
rect 190196 251646 190252 251702
rect 420404 256974 420460 257030
rect 420404 255198 420460 255254
rect 420404 252830 420460 252886
rect 420308 250462 420364 250518
rect 420404 248094 420460 248150
rect 420404 245282 420460 245338
rect 420308 243506 420364 243562
rect 420308 241138 420364 241194
rect 412244 240250 412300 240306
rect 412148 240102 412204 240158
rect 412052 239971 412108 240010
rect 412052 239954 412054 239971
rect 412054 239954 412106 239971
rect 412106 239954 412108 239971
rect 292148 228854 292204 228910
rect 298964 231814 299020 231870
rect 299444 234922 299500 234978
rect 299348 234626 299404 234682
rect 301652 234774 301708 234830
rect 307604 231074 307660 231130
rect 313460 228114 313516 228170
rect 316724 231222 316780 231278
rect 318932 225154 318988 225210
rect 322484 231370 322540 231426
rect 327092 231518 327148 231574
rect 325940 225302 325996 225358
rect 327956 225598 328012 225654
rect 330260 231666 330316 231722
rect 331028 225746 331084 225802
rect 333044 228262 333100 228318
rect 333812 225894 333868 225950
rect 334868 233146 334924 233202
rect 336884 227374 336940 227430
rect 338612 234182 338668 234238
rect 339380 228410 339436 228466
rect 339860 230334 339916 230390
rect 341588 234330 341644 234386
rect 342164 228706 342220 228762
rect 343124 227226 343180 227282
rect 344372 235070 344428 235126
rect 345332 234774 345388 234830
rect 345428 228558 345484 228614
rect 344756 227078 344812 227134
rect 347636 234774 347692 234830
rect 352724 230817 352726 230834
rect 352726 230817 352778 230834
rect 352778 230817 352780 230834
rect 352724 230778 352780 230817
rect 354356 234922 354412 234978
rect 354260 230334 354316 230390
rect 354260 225450 354316 225506
rect 354164 224414 354220 224470
rect 356756 235218 356812 235274
rect 356852 234922 356908 234978
rect 359060 232998 359116 233054
rect 359060 230778 359116 230834
rect 358964 229890 359020 229946
rect 357428 222934 357484 222990
rect 359444 224562 359500 224618
rect 359828 228854 359884 228910
rect 359732 224118 359788 224174
rect 361748 236994 361804 237050
rect 360884 230334 360940 230390
rect 360980 224266 361036 224322
rect 363572 230038 363628 230094
rect 363476 223970 363532 224026
rect 364052 234478 364108 234534
rect 365684 233294 365740 233350
rect 367220 235958 367276 236014
rect 366164 223822 366220 223878
rect 368948 236994 369004 237050
rect 367604 223674 367660 223730
rect 370388 236846 370444 236902
rect 370772 232850 370828 232906
rect 372212 236254 372268 236310
rect 373460 236550 373516 236606
rect 373076 229742 373132 229798
rect 374900 236698 374956 236754
rect 375380 232702 375436 232758
rect 376532 236254 376588 236310
rect 376724 236254 376780 236310
rect 376340 233590 376396 233646
rect 376820 229594 376876 229650
rect 377204 233294 377260 233350
rect 377780 236994 377836 237050
rect 377972 236994 378028 237050
rect 379124 233886 379180 233942
rect 378740 232554 378796 232610
rect 377588 223526 377644 223582
rect 379796 223378 379852 223434
rect 382100 233738 382156 233794
rect 381716 232406 381772 232462
rect 381332 229446 381388 229502
rect 381236 223230 381292 223286
rect 382964 231962 383020 232018
rect 383540 229298 383596 229354
rect 384980 232258 385036 232314
rect 385364 232110 385420 232166
rect 384404 229150 384460 229206
rect 384308 223082 384364 223138
rect 385844 231814 385900 231870
rect 385748 222786 385804 222842
rect 388436 236994 388492 237050
rect 388724 236994 388780 237050
rect 391220 226930 391276 226986
rect 391604 226782 391660 226838
rect 393044 235810 393100 235866
rect 394484 226634 394540 226690
rect 394100 226486 394156 226542
rect 397076 236402 397132 236458
rect 396788 235662 396844 235718
rect 396980 235070 397036 235126
rect 397460 236994 397516 237050
rect 397556 236846 397612 236902
rect 397364 236441 397366 236458
rect 397366 236441 397418 236458
rect 397418 236441 397420 236458
rect 397364 236402 397420 236441
rect 397748 236994 397804 237050
rect 397748 236885 397750 236902
rect 397750 236885 397802 236902
rect 397802 236885 397804 236902
rect 397748 236846 397804 236885
rect 398132 229002 398188 229058
rect 399860 235514 399916 235570
rect 399476 228854 399532 228910
rect 400436 235958 400492 236014
rect 401396 235366 401452 235422
rect 400052 222638 400108 222694
rect 402548 235218 402604 235274
rect 402740 235218 402796 235274
rect 403412 234922 403468 234978
rect 402644 226338 402700 226394
rect 403988 236106 404044 236162
rect 403412 222490 403468 222546
rect 405428 235958 405484 236014
rect 405332 234626 405388 234682
rect 405236 231814 405292 231870
rect 405524 234626 405580 234682
rect 405908 234478 405964 234534
rect 405812 226042 405868 226098
rect 407444 234774 407500 234830
rect 407252 234034 407308 234090
rect 407636 230186 407692 230242
rect 408116 235070 408172 235126
rect 408500 234922 408556 234978
rect 409940 234774 409996 234830
rect 408788 233590 408844 233646
rect 407540 226190 407596 226246
rect 411380 237033 411382 237050
rect 411382 237033 411434 237050
rect 411434 237033 411436 237050
rect 411380 236994 411436 237033
rect 411572 236994 411628 237050
rect 411572 236254 411628 236310
rect 411284 234626 411340 234682
rect 411476 233886 411532 233942
rect 411764 236254 411820 236310
rect 411764 233738 411820 233794
rect 581780 240250 581836 240306
rect 567380 239954 567436 240010
rect 413396 238918 413452 238974
rect 414644 238770 414700 238826
rect 413684 238622 413740 238678
rect 413972 238326 414028 238382
rect 414260 238178 414316 238234
rect 414452 238030 414508 238086
rect 419156 237142 419212 237198
rect 419156 236846 419212 236902
rect 424724 231074 424780 231130
rect 436916 228114 436972 228170
rect 442868 231222 442924 231278
rect 445172 225154 445228 225210
rect 455156 231370 455212 231426
rect 457268 225302 457324 225358
rect 464084 231518 464140 231574
rect 463316 225598 463372 225654
rect 466484 234182 466540 234238
rect 470132 231666 470188 231722
rect 469364 225746 469420 225802
rect 476180 228262 476236 228318
rect 475316 225894 475372 225950
rect 479060 233146 479116 233202
rect 481460 227374 481516 227430
rect 488276 228410 488332 228466
rect 487508 225450 487564 225506
rect 490484 234330 490540 234386
rect 494228 228706 494284 228762
rect 493460 227226 493516 227282
rect 497972 228558 498028 228614
rect 498836 227078 498892 227134
rect 506804 234034 506860 234090
rect 514004 221732 514060 221788
rect 513908 221602 513964 221658
rect 518420 224414 518476 224470
rect 525236 232998 525292 233054
rect 524468 222934 524524 222990
rect 523796 222638 523852 222694
rect 522932 222490 522988 222546
rect 528308 230334 528364 230390
rect 527540 229890 527596 229946
rect 526676 224562 526732 224618
rect 528980 224118 529036 224174
rect 530516 224266 530572 224322
rect 532052 222786 532108 222842
rect 533492 238326 533548 238382
rect 538004 238030 538060 238086
rect 534260 230038 534316 230094
rect 544340 238622 544396 238678
rect 536564 223970 536620 224026
rect 541076 223822 541132 223878
rect 544052 223674 544108 223730
rect 550196 238918 550252 238974
rect 559892 238178 559948 238234
rect 559220 236698 559276 236754
rect 557012 236550 557068 236606
rect 553940 236402 553996 236458
rect 551636 232850 551692 232906
rect 553940 229742 553996 229798
rect 565268 236994 565324 237050
rect 562196 236846 562252 236902
rect 560756 232702 560812 232758
rect 564500 232554 564556 232610
rect 563636 229594 563692 229650
rect 562964 223526 563020 223582
rect 573140 238770 573196 238826
rect 570452 232406 570508 232462
rect 568244 223378 568300 223434
rect 571316 223230 571372 223286
rect 572756 229446 572812 229502
rect 573524 229298 573580 229354
rect 576596 232258 576652 232314
rect 575828 231962 575884 232018
rect 575060 230186 575116 230242
rect 578036 232110 578092 232166
rect 577268 223082 577324 223138
rect 578900 229150 578956 229206
rect 587348 236106 587404 236162
rect 588980 235958 589036 236014
rect 587828 235810 587884 235866
rect 587444 234478 587500 234534
rect 590900 226930 590956 226986
rect 591668 226782 591724 226838
rect 596948 226634 597004 226690
rect 596180 226486 596236 226542
rect 599924 229002 599980 229058
rect 602228 235662 602284 235718
rect 604532 231814 604588 231870
rect 627188 240102 627244 240158
rect 621140 236254 621196 236310
rect 608276 235514 608332 235570
rect 607508 228854 607564 228910
rect 611252 235366 611308 235422
rect 614324 235218 614380 235274
rect 613556 226338 613612 226394
rect 620372 226042 620428 226098
rect 624884 235070 624940 235126
rect 623348 226190 623404 226246
rect 625556 234922 625612 234978
rect 627860 234774 627916 234830
rect 630932 234626 630988 234682
rect 640148 212278 640204 212334
rect 640148 211538 640204 211594
rect 190292 201326 190348 201382
rect 640148 200882 640204 200938
rect 190292 200512 190348 200568
rect 640148 200142 640204 200198
rect 187220 199106 187276 199162
rect 185780 182382 185836 182438
rect 185684 174686 185740 174742
rect 184340 155002 184396 155058
rect 184436 154114 184492 154170
rect 184532 153522 184588 153578
rect 184628 152634 184684 152690
rect 184340 151894 184396 151950
rect 184436 151154 184492 151210
rect 184532 150414 184588 150470
rect 184340 149674 184396 149730
rect 184436 148934 184492 148990
rect 184724 148046 184780 148102
rect 184532 147306 184588 147362
rect 184340 145826 184396 145882
rect 184436 145086 184492 145142
rect 184628 146605 184630 146622
rect 184630 146605 184682 146622
rect 184682 146605 184684 146622
rect 184628 146566 184684 146605
rect 184532 144346 184588 144402
rect 184340 143606 184396 143662
rect 184436 142718 184492 142774
rect 184628 142126 184684 142182
rect 184532 141238 184588 141294
rect 184340 140498 184396 140554
rect 184436 139758 184492 139814
rect 184532 138870 184588 138926
rect 184340 134430 184396 134486
rect 185972 138278 186028 138334
rect 186068 137390 186124 137446
rect 185780 135170 185836 135226
rect 640244 185638 640300 185694
rect 640244 184898 640300 184954
rect 186740 183122 186796 183178
rect 645140 182974 645196 183030
rect 186356 173206 186412 173262
rect 186260 136798 186316 136854
rect 645140 179274 645196 179330
rect 645140 174873 645142 174890
rect 645142 174873 645194 174890
rect 645194 174873 645196 174890
rect 645140 174834 645196 174873
rect 645140 171025 645142 171042
rect 645142 171025 645194 171042
rect 645194 171025 645196 171042
rect 645140 170986 645196 171025
rect 645140 167730 645196 167786
rect 645140 163329 645142 163346
rect 645142 163329 645194 163346
rect 645194 163329 645196 163346
rect 645140 163290 645196 163329
rect 645140 159442 645196 159498
rect 645140 155446 645196 155502
rect 645140 152525 645142 152542
rect 645142 152525 645194 152542
rect 645194 152525 645196 152542
rect 645140 152486 645196 152525
rect 645140 148046 645196 148102
rect 186452 135910 186508 135966
rect 186164 133690 186220 133746
rect 184436 132950 184492 133006
rect 184340 132227 184396 132266
rect 184340 132210 184342 132227
rect 184342 132210 184394 132227
rect 184394 132210 184396 132227
rect 184436 131470 184492 131526
rect 184532 130582 184588 130638
rect 184628 129842 184684 129898
rect 184340 128362 184396 128418
rect 184436 127622 184492 127678
rect 184532 126882 184588 126938
rect 184340 125994 184396 126050
rect 184436 125402 184492 125458
rect 184532 124514 184588 124570
rect 184436 123774 184492 123830
rect 184340 123034 184396 123090
rect 184628 122146 184684 122202
rect 184532 121554 184588 121610
rect 184340 120666 184396 120722
rect 184532 120074 184588 120130
rect 184436 119186 184492 119242
rect 184724 118594 184780 118650
rect 184340 117706 184396 117762
rect 184436 116966 184492 117022
rect 184532 116226 184588 116282
rect 184628 115338 184684 115394
rect 184340 114746 184396 114802
rect 184436 113858 184492 113914
rect 184532 113118 184588 113174
rect 184628 112378 184684 112434
rect 184340 111638 184396 111694
rect 184436 110898 184492 110954
rect 184532 110158 184588 110214
rect 184340 109309 184342 109326
rect 184342 109309 184394 109326
rect 184394 109309 184396 109326
rect 184340 109270 184396 109309
rect 186740 129102 186796 129158
rect 645716 128954 645772 129010
rect 648596 272070 648652 272126
rect 647348 269258 647404 269314
rect 646580 267038 646636 267094
rect 185588 108678 185644 108734
rect 646676 144198 646732 144254
rect 655220 778230 655276 778286
rect 655124 775862 655180 775918
rect 654356 773494 654412 773550
rect 654068 730130 654124 730186
rect 655124 734422 655180 734478
rect 654164 728502 654220 728558
rect 653780 686914 653836 686970
rect 654164 685286 654220 685342
rect 654068 684546 654124 684602
rect 655412 777638 655468 777694
rect 655316 731610 655372 731666
rect 655220 689430 655276 689486
rect 649748 263486 649804 263542
rect 646772 140942 646828 140998
rect 655124 642366 655180 642422
rect 654164 640590 654220 640646
rect 653972 594118 654028 594174
rect 655604 776010 655660 776066
rect 655508 732646 655564 732702
rect 655412 688394 655468 688450
rect 655316 642958 655372 643014
rect 655220 597818 655276 597874
rect 655124 553270 655180 553326
rect 654164 548534 654220 548590
rect 656564 774678 656620 774734
rect 655700 731314 655756 731370
rect 655604 687062 655660 687118
rect 655508 640738 655564 640794
rect 655412 596634 655468 596690
rect 655316 550902 655372 550958
rect 655796 639110 655852 639166
rect 655988 638222 656044 638278
rect 655604 595450 655660 595506
rect 655508 552086 655564 552142
rect 655796 595302 655852 595358
rect 656564 592934 656620 592990
rect 655700 550754 655756 550810
rect 656564 549718 656620 549774
rect 655124 373302 655180 373358
rect 655508 374338 655564 374394
rect 655316 372118 655372 372174
rect 656564 370934 656620 370990
rect 655220 329790 655276 329846
rect 655124 328014 655180 328070
rect 655316 327422 655372 327478
rect 654164 326238 654220 326294
rect 654164 303298 654220 303354
rect 654068 302114 654124 302170
rect 654260 300930 654316 300986
rect 656564 298710 656620 298766
rect 656084 297526 656140 297582
rect 655892 293974 655948 294030
rect 655796 292790 655852 292846
rect 655604 289238 655660 289294
rect 655412 288054 655468 288110
rect 653780 284502 653836 284558
rect 655124 283318 655180 283374
rect 654164 279766 654220 279822
rect 652244 266890 652300 266946
rect 647060 134726 647116 134782
rect 647828 130878 647884 130934
rect 646964 127622 647020 127678
rect 646868 125698 646924 125754
rect 646580 123774 646636 123830
rect 646484 121998 646540 122054
rect 655316 282282 655372 282338
rect 655220 280950 655276 281006
rect 655508 286870 655564 286926
rect 655700 285686 655756 285742
rect 655988 290866 656044 290922
rect 656276 296786 656332 296842
rect 656180 291606 656236 291662
rect 656372 295158 656428 295214
rect 647924 119482 647980 119538
rect 645236 117558 645292 117614
rect 647924 115634 647980 115690
rect 646580 113118 646636 113174
rect 186164 107790 186220 107846
rect 184436 107050 184492 107106
rect 184340 105570 184396 105626
rect 185300 106349 185302 106366
rect 185302 106349 185354 106366
rect 185354 106349 185356 106366
rect 185300 106310 185356 106349
rect 645908 106014 645964 106070
rect 184532 104830 184588 104886
rect 184436 103942 184492 103998
rect 184436 103350 184492 103406
rect 184340 102462 184396 102518
rect 184532 101870 184588 101926
rect 184628 100982 184684 101038
rect 184340 100242 184396 100298
rect 184436 99502 184492 99558
rect 184628 98614 184684 98670
rect 184532 98022 184588 98078
rect 184340 97134 184396 97190
rect 184436 96394 184492 96450
rect 645140 102166 645196 102222
rect 184724 95654 184780 95710
rect 184340 94783 184396 94822
rect 184340 94766 184342 94783
rect 184342 94766 184394 94783
rect 184394 94766 184396 94783
rect 184436 94174 184492 94230
rect 184532 93434 184588 93490
rect 184628 92694 184684 92750
rect 184340 91971 184396 92010
rect 184340 91954 184342 91971
rect 184342 91954 184394 91971
rect 184394 91954 184396 91971
rect 184436 90326 184492 90382
rect 184628 91066 184684 91122
rect 184532 89586 184588 89642
rect 184340 88846 184396 88902
rect 184436 88106 184492 88162
rect 184532 87218 184588 87274
rect 184628 86626 184684 86682
rect 184340 85738 184396 85794
rect 184436 85146 184492 85202
rect 184532 84258 184588 84314
rect 184340 83409 184342 83426
rect 184342 83409 184394 83426
rect 184394 83409 184396 83426
rect 184340 83370 184396 83409
rect 184244 81890 184300 81946
rect 645428 95967 645484 96006
rect 645428 95950 645430 95967
rect 645430 95950 645482 95967
rect 645482 95950 645484 95967
rect 186164 82778 186220 82834
rect 184436 81298 184492 81354
rect 184436 79818 184492 79874
rect 184340 78930 184396 78986
rect 184628 80427 184684 80466
rect 184628 80410 184630 80427
rect 184630 80410 184682 80427
rect 184682 80410 184684 80427
rect 184532 78190 184588 78246
rect 184436 77450 184492 77506
rect 184340 76710 184396 76766
rect 184532 75970 184588 76026
rect 184628 75082 184684 75138
rect 184340 74342 184396 74398
rect 184532 73602 184588 73658
rect 184436 72862 184492 72918
rect 184628 72122 184684 72178
rect 149492 70790 149548 70846
rect 149396 69458 149452 69514
rect 149204 68274 149260 68330
rect 184436 71382 184492 71438
rect 184340 70494 184396 70550
rect 184532 69902 184588 69958
rect 184340 69031 184396 69070
rect 184340 69014 184342 69031
rect 184342 69014 184394 69031
rect 184394 69014 184396 69031
rect 149588 67090 149644 67146
rect 149492 65314 149548 65370
rect 149396 64574 149452 64630
rect 149300 63390 149356 63446
rect 184532 68422 184588 68478
rect 184436 67534 184492 67590
rect 184340 66794 184396 66850
rect 184340 66054 184396 66110
rect 184532 65166 184588 65222
rect 184436 64574 184492 64630
rect 184628 63686 184684 63742
rect 184436 63094 184492 63150
rect 149396 62206 149452 62262
rect 184340 62206 184396 62262
rect 184532 61466 184588 61522
rect 184628 60726 184684 60782
rect 149492 60578 149548 60634
rect 149396 59690 149452 59746
rect 184436 59986 184492 60042
rect 184340 59246 184396 59302
rect 149396 58506 149452 58562
rect 184532 58358 184588 58414
rect 184340 57618 184396 57674
rect 149492 57322 149548 57378
rect 149396 56177 149398 56194
rect 149398 56177 149450 56194
rect 149450 56177 149452 56194
rect 149396 56138 149452 56177
rect 184340 56878 184396 56934
rect 184340 56155 184396 56194
rect 184340 56138 184342 56155
rect 184342 56138 184394 56155
rect 184394 56138 184396 56155
rect 184436 55398 184492 55454
rect 149684 54806 149740 54862
rect 184340 54675 184396 54714
rect 184340 54658 184342 54675
rect 184342 54658 184394 54675
rect 184394 54658 184396 54675
rect 184340 53918 184396 53974
rect 149396 53770 149452 53826
rect 142100 40154 142156 40210
rect 311060 37194 311116 37250
rect 331220 37194 331276 37250
rect 417524 44890 417580 44946
rect 415220 41930 415276 41986
rect 416852 41782 416908 41838
rect 420788 40450 420844 40506
rect 472244 44890 472300 44946
rect 464852 41782 464908 41838
rect 470324 41782 470380 41838
rect 645908 88846 645964 88902
rect 645908 84406 645964 84462
rect 645524 79374 645580 79430
rect 646004 75526 646060 75582
rect 646004 66219 646060 66258
rect 646004 66202 646006 66219
rect 646006 66202 646058 66219
rect 646058 66202 646060 66219
rect 646004 58950 646060 59006
rect 669524 275178 669580 275234
rect 669716 275030 669772 275086
rect 669908 277546 669964 277602
rect 670100 277694 670156 277750
rect 670004 273550 670060 273606
rect 672308 278582 672364 278638
rect 676052 891467 676108 891506
rect 676052 891450 676054 891467
rect 676054 891450 676106 891467
rect 676106 891450 676108 891467
rect 676052 890431 676108 890470
rect 676052 890414 676054 890431
rect 676054 890414 676106 890431
rect 676106 890414 676108 890431
rect 680180 890118 680236 890174
rect 676244 889230 676300 889286
rect 679988 888638 680044 888694
rect 676244 887750 676300 887806
rect 676052 887380 676108 887436
rect 679700 886714 679756 886770
rect 676052 885456 676108 885512
rect 676052 884938 676108 884994
rect 675764 884346 675820 884402
rect 676052 883976 676108 884032
rect 676052 883458 676108 883514
rect 679796 886122 679852 886178
rect 679700 882718 679756 882774
rect 679700 882126 679756 882182
rect 679892 885678 679948 885734
rect 680084 888194 680140 888250
rect 685460 882126 685516 882182
rect 685460 881682 685516 881738
rect 675380 787998 675436 788054
rect 675764 787406 675820 787462
rect 675476 786666 675532 786722
rect 675380 784742 675436 784798
rect 675476 784150 675532 784206
rect 675284 783410 675340 783466
rect 675764 782966 675820 783022
rect 675668 780598 675724 780654
rect 675764 779858 675820 779914
rect 675764 779118 675820 779174
rect 675476 777638 675532 777694
rect 675764 775418 675820 775474
rect 674420 730574 674476 730630
rect 674996 772014 675052 772070
rect 674900 771866 674956 771922
rect 675476 742414 675532 742470
rect 675188 741082 675244 741138
rect 675476 740342 675532 740398
rect 675476 739158 675532 739214
rect 675764 735458 675820 735514
rect 676340 715478 676396 715534
rect 676148 714886 676204 714942
rect 676244 714755 676300 714794
rect 676244 714738 676246 714755
rect 676246 714738 676298 714755
rect 676298 714738 676300 714755
rect 676052 714185 676054 714202
rect 676054 714185 676106 714202
rect 676106 714185 676108 714202
rect 676052 714146 676108 714185
rect 676244 713423 676300 713462
rect 676244 713406 676246 713423
rect 676246 713406 676298 713423
rect 676298 713406 676300 713423
rect 676052 713127 676108 713166
rect 676052 713110 676054 713127
rect 676054 713110 676106 713127
rect 676106 713110 676108 713127
rect 676052 712683 676108 712722
rect 676052 712666 676054 712683
rect 676054 712666 676106 712683
rect 676106 712666 676108 712683
rect 676244 711943 676300 711982
rect 676244 711926 676246 711943
rect 676246 711926 676298 711943
rect 676298 711926 676300 711943
rect 676052 711573 676108 711612
rect 676052 711556 676054 711573
rect 676054 711556 676106 711573
rect 676106 711556 676108 711573
rect 676052 711186 676108 711242
rect 676052 708522 676108 708578
rect 676052 708152 676108 708208
rect 676244 704861 676246 704878
rect 676246 704861 676298 704878
rect 676298 704861 676300 704878
rect 676244 704822 676300 704861
rect 679988 704378 680044 704434
rect 679796 703342 679852 703398
rect 679988 703342 680044 703398
rect 679796 702898 679852 702954
rect 675380 697866 675436 697922
rect 675188 697126 675244 697182
rect 675188 696978 675244 697034
rect 675668 694906 675724 694962
rect 675284 694610 675340 694666
rect 676148 670338 676204 670394
rect 676052 669193 676054 669210
rect 676054 669193 676106 669210
rect 676106 669193 676108 669210
rect 676052 669154 676108 669193
rect 676052 668562 676108 668618
rect 676340 669746 676396 669802
rect 676244 669302 676300 669358
rect 675956 668061 676012 668100
rect 675956 668044 675958 668061
rect 675958 668044 676010 668061
rect 676010 668044 676012 668061
rect 675956 667691 676012 667730
rect 675956 667674 675958 667691
rect 675958 667674 676010 667691
rect 676010 667674 676012 667691
rect 676244 666934 676300 666990
rect 676244 666359 676300 666398
rect 676244 666342 676246 666359
rect 676246 666342 676298 666359
rect 676298 666342 676300 666359
rect 676052 665602 676108 665658
rect 676052 663530 676108 663586
rect 676052 662089 676054 662106
rect 676054 662089 676106 662106
rect 676106 662089 676108 662106
rect 676052 662050 676108 662089
rect 676052 661645 676054 661662
rect 676054 661645 676106 661662
rect 676106 661645 676108 661662
rect 676052 661606 676108 661645
rect 676244 661349 676246 661366
rect 676246 661349 676298 661366
rect 676298 661349 676300 661366
rect 676244 661310 676300 661349
rect 676052 660609 676054 660626
rect 676054 660609 676106 660626
rect 676106 660609 676108 660626
rect 676052 660570 676108 660609
rect 676052 660165 676054 660182
rect 676054 660165 676106 660182
rect 676106 660165 676108 660182
rect 676052 660126 676108 660165
rect 676244 659869 676246 659886
rect 676246 659869 676298 659886
rect 676298 659869 676300 659886
rect 676244 659830 676300 659869
rect 679796 659238 679852 659294
rect 679796 658350 679852 658406
rect 685460 658350 685516 658406
rect 685460 657906 685516 657962
rect 675380 652726 675436 652782
rect 675476 652134 675532 652190
rect 675380 651394 675436 651450
rect 675380 649618 675436 649674
rect 675476 645326 675532 645382
rect 675764 640294 675820 640350
rect 675764 638518 675820 638574
rect 676244 625050 676300 625106
rect 676148 624606 676204 624662
rect 676052 623979 676054 623996
rect 676054 623979 676106 623996
rect 676106 623979 676108 623996
rect 676052 623940 676108 623979
rect 676052 623439 676108 623478
rect 676052 623422 676054 623439
rect 676054 623422 676106 623439
rect 676106 623422 676108 623439
rect 676052 622830 676108 622886
rect 676052 622477 676108 622516
rect 676052 622460 676054 622477
rect 676054 622460 676106 622477
rect 676106 622460 676108 622477
rect 676244 624162 676300 624218
rect 676052 621959 676108 621998
rect 676052 621942 676054 621959
rect 676054 621942 676106 621959
rect 676106 621942 676108 621959
rect 676052 621367 676108 621406
rect 676052 621350 676054 621367
rect 676054 621350 676106 621367
rect 676106 621350 676108 621367
rect 676244 620610 676300 620666
rect 676052 618908 676108 618964
rect 676244 618538 676300 618594
rect 676244 617097 676246 617114
rect 676246 617097 676298 617114
rect 676298 617097 676300 617114
rect 676244 617058 676300 617097
rect 676052 616505 676054 616522
rect 676054 616505 676106 616522
rect 676106 616505 676108 616522
rect 676052 616466 676108 616505
rect 676052 615913 676054 615930
rect 676054 615913 676106 615930
rect 676106 615913 676108 615930
rect 676052 615874 676108 615913
rect 676244 615617 676246 615634
rect 676246 615617 676298 615634
rect 676298 615617 676300 615634
rect 676244 615578 676300 615617
rect 676244 615173 676246 615190
rect 676246 615173 676298 615190
rect 676298 615173 676300 615190
rect 676244 615134 676300 615173
rect 676052 614433 676054 614450
rect 676054 614433 676106 614450
rect 676106 614433 676108 614450
rect 676052 614394 676108 614433
rect 679988 613654 680044 613710
rect 679796 613210 679852 613266
rect 679988 613210 680044 613266
rect 679796 612766 679852 612822
rect 675188 607734 675244 607790
rect 675188 605958 675244 606014
rect 675284 604774 675340 604830
rect 675476 600186 675532 600242
rect 675764 595302 675820 595358
rect 675668 593378 675724 593434
rect 676340 578282 676396 578338
rect 676148 577542 676204 577598
rect 676052 576989 676054 577006
rect 676054 576989 676106 577006
rect 676106 576989 676108 577006
rect 676052 576950 676108 576989
rect 676244 577098 676300 577154
rect 676244 576210 676300 576266
rect 676052 575931 676108 575970
rect 676052 575914 676054 575931
rect 676054 575914 676106 575931
rect 676106 575914 676108 575931
rect 676052 575487 676108 575526
rect 676052 575470 676054 575487
rect 676054 575470 676106 575487
rect 676106 575470 676108 575487
rect 676052 574917 676054 574934
rect 676054 574917 676106 574934
rect 676106 574917 676108 574934
rect 676052 574878 676108 574917
rect 676052 574377 676108 574416
rect 676052 574360 676054 574377
rect 676054 574360 676106 574377
rect 676106 574360 676108 574377
rect 676244 570625 676246 570642
rect 676246 570625 676298 570642
rect 676298 570625 676300 570642
rect 676244 570586 676300 570625
rect 676052 569885 676054 569902
rect 676054 569885 676106 569902
rect 676106 569885 676108 569902
rect 676052 569846 676108 569885
rect 676052 569515 676054 569532
rect 676054 569515 676106 569532
rect 676106 569515 676108 569532
rect 676052 569476 676108 569515
rect 676244 569145 676246 569162
rect 676246 569145 676298 569162
rect 676298 569145 676300 569162
rect 676244 569106 676300 569145
rect 676052 568405 676054 568422
rect 676054 568405 676106 568422
rect 676106 568405 676108 568422
rect 676052 568366 676108 568405
rect 676052 567961 676054 567978
rect 676054 567961 676106 567978
rect 676106 567961 676108 567978
rect 676052 567922 676108 567961
rect 676244 567665 676246 567682
rect 676246 567665 676298 567682
rect 676298 567665 676300 567682
rect 676244 567626 676300 567665
rect 679796 567034 679852 567090
rect 679796 566146 679852 566202
rect 685460 566146 685516 566202
rect 685460 565702 685516 565758
rect 675476 562446 675532 562502
rect 675188 561706 675244 561762
rect 675380 561410 675436 561466
rect 675476 558894 675532 558950
rect 676148 534918 676204 534974
rect 676052 534178 676108 534234
rect 675956 533773 675958 533790
rect 675958 533773 676010 533790
rect 676010 533773 676012 533790
rect 675956 533734 676012 533773
rect 676244 534326 676300 534382
rect 676532 532994 676588 533050
rect 676052 532715 676108 532754
rect 676052 532698 676054 532715
rect 676054 532698 676106 532715
rect 676106 532698 676108 532715
rect 676244 531531 676300 531570
rect 676244 531514 676246 531531
rect 676246 531514 676298 531531
rect 676298 531514 676300 531531
rect 676244 528001 676246 528018
rect 676246 528001 676298 528018
rect 676298 528001 676300 528018
rect 676244 527962 676300 528001
rect 676244 527409 676246 527426
rect 676246 527409 676298 527426
rect 676298 527409 676300 527426
rect 676244 527370 676300 527409
rect 676052 526669 676054 526686
rect 676054 526669 676106 526686
rect 676106 526669 676108 526686
rect 676052 526630 676108 526669
rect 676052 526299 676054 526316
rect 676054 526299 676106 526316
rect 676106 526299 676108 526316
rect 676052 526260 676108 526299
rect 676244 525929 676246 525946
rect 676246 525929 676298 525946
rect 676298 525929 676300 525946
rect 676244 525890 676300 525929
rect 676052 525189 676054 525206
rect 676054 525189 676106 525206
rect 676106 525189 676108 525206
rect 676052 525150 676108 525189
rect 676052 524819 676054 524836
rect 676054 524819 676106 524836
rect 676106 524819 676108 524836
rect 676052 524780 676108 524819
rect 676244 524449 676246 524466
rect 676246 524449 676298 524466
rect 676298 524449 676300 524466
rect 676244 524410 676300 524449
rect 676628 531958 676684 532014
rect 676244 490518 676300 490574
rect 676148 490074 676204 490130
rect 676244 489943 676300 489982
rect 676244 489926 676246 489943
rect 676246 489926 676298 489943
rect 676298 489926 676300 489943
rect 676052 488298 676108 488354
rect 676724 530922 676780 530978
rect 679796 523522 679852 523578
rect 679796 522930 679852 522986
rect 685460 522930 685516 522986
rect 685460 522486 685516 522542
rect 679700 489186 679756 489242
rect 676724 488594 676780 488650
rect 676244 487131 676300 487170
rect 676244 487114 676246 487131
rect 676246 487114 676298 487131
rect 676298 487114 676300 487131
rect 676052 485782 676108 485838
rect 676244 485042 676300 485098
rect 676052 484302 676108 484358
rect 675956 483727 676012 483766
rect 675956 483710 675958 483727
rect 675958 483710 676010 483727
rect 676010 483710 676012 483727
rect 676052 482230 676108 482286
rect 676052 481899 676054 481916
rect 676054 481899 676106 481916
rect 676106 481899 676108 481916
rect 676052 481860 676108 481899
rect 676244 481529 676246 481546
rect 676246 481529 676298 481546
rect 676298 481529 676300 481546
rect 676244 481490 676300 481529
rect 676052 480789 676054 480806
rect 676054 480789 676106 480806
rect 676106 480789 676108 480806
rect 676052 480750 676108 480789
rect 676052 480419 676054 480436
rect 676054 480419 676106 480436
rect 676106 480419 676108 480436
rect 676052 480380 676108 480419
rect 676244 480049 676246 480066
rect 676246 480049 676298 480066
rect 676298 480049 676300 480066
rect 676244 480010 676300 480049
rect 676148 402310 676204 402366
rect 676052 401570 676108 401626
rect 676244 401718 676300 401774
rect 676244 400403 676300 400442
rect 676244 400386 676246 400403
rect 676246 400386 676298 400403
rect 676298 400386 676300 400403
rect 676532 400238 676588 400294
rect 676052 399646 676108 399702
rect 676052 398610 676108 398666
rect 677876 487558 677932 487614
rect 679796 486522 679852 486578
rect 679700 478530 679756 478586
rect 679700 478086 679756 478142
rect 679892 479122 679948 479178
rect 679892 478530 679948 478586
rect 676724 400978 676780 401034
rect 676628 399350 676684 399406
rect 676052 395593 676108 395632
rect 676052 395576 676054 395593
rect 676054 395576 676106 395593
rect 676106 395576 676108 395593
rect 679796 390914 679852 390970
rect 679796 390322 679852 390378
rect 685460 390322 685516 390378
rect 685460 389878 685516 389934
rect 675188 385882 675244 385938
rect 675764 385586 675820 385642
rect 675188 384402 675244 384458
rect 675764 382922 675820 382978
rect 675476 382330 675532 382386
rect 675764 381738 675820 381794
rect 675764 381146 675820 381202
rect 675476 378778 675532 378834
rect 675572 378038 675628 378094
rect 675380 377150 675436 377206
rect 675764 376706 675820 376762
rect 675764 375670 675820 375726
rect 675476 373894 675532 373950
rect 676340 358058 676396 358114
rect 676148 357466 676204 357522
rect 676244 357335 676300 357374
rect 676244 357318 676246 357335
rect 676246 357318 676298 357335
rect 676298 357318 676300 357335
rect 676052 356765 676054 356782
rect 676054 356765 676106 356782
rect 676106 356765 676108 356782
rect 676052 356726 676108 356765
rect 676052 355707 676108 355746
rect 676052 355690 676054 355707
rect 676054 355690 676106 355707
rect 676106 355690 676108 355707
rect 672404 277990 672460 278046
rect 670484 277842 670540 277898
rect 670292 277398 670348 277454
rect 676052 354671 676108 354710
rect 676052 354654 676054 354671
rect 676054 354654 676106 354671
rect 676106 354654 676108 354671
rect 675572 352582 675628 352638
rect 676052 352286 676108 352342
rect 676916 350954 676972 351010
rect 676052 350806 676108 350862
rect 676052 350214 676108 350270
rect 676244 349474 676300 349530
rect 676820 349030 676876 349086
rect 676244 347994 676300 348050
rect 676052 347772 676108 347828
rect 675956 347254 676012 347310
rect 676820 342962 676876 343018
rect 679892 346514 679948 346570
rect 679892 346070 679948 346126
rect 679700 345922 679756 345978
rect 679700 345478 679756 345534
rect 676916 342814 676972 342870
rect 675764 339558 675820 339614
rect 675380 333490 675436 333546
rect 675476 332306 675532 332362
rect 675764 330530 675820 330586
rect 675380 328310 675436 328366
rect 675764 326830 675820 326886
rect 676340 312178 676396 312234
rect 676148 311586 676204 311642
rect 676244 311181 676246 311198
rect 676246 311181 676298 311198
rect 676298 311181 676300 311198
rect 676244 311142 676300 311181
rect 676052 307960 676108 308016
rect 676820 307146 676876 307202
rect 676244 306702 676300 306758
rect 676244 304778 676300 304834
rect 676052 304408 676108 304464
rect 675956 303890 676012 303946
rect 676052 301966 676108 302022
rect 676244 301226 676300 301282
rect 679988 300634 680044 300690
rect 679796 300190 679852 300246
rect 679988 300190 680044 300246
rect 679796 299746 679852 299802
rect 676820 299154 676876 299210
rect 675668 292790 675724 292846
rect 675764 290718 675820 290774
rect 675476 288498 675532 288554
rect 675476 287166 675532 287222
rect 675476 285242 675532 285298
rect 675764 283614 675820 283670
rect 675380 281838 675436 281894
rect 672788 278286 672844 278342
rect 676532 278138 676588 278194
rect 679700 276510 679756 276566
rect 672500 276214 672556 276270
rect 670196 270590 670252 270646
rect 676244 266890 676300 266946
rect 672788 266742 672844 266798
rect 672404 266594 672460 266650
rect 672596 266298 672652 266354
rect 672404 174686 672460 174742
rect 672980 266446 673036 266502
rect 676148 266446 676204 266502
rect 676052 266150 676108 266206
rect 676052 265205 676108 265244
rect 676052 265188 676054 265205
rect 676054 265188 676106 265205
rect 676106 265188 676108 265205
rect 679700 264818 679756 264874
rect 676052 264226 676108 264282
rect 679796 264078 679852 264134
rect 676916 262006 676972 262062
rect 676052 261266 676108 261322
rect 675284 259786 675340 259842
rect 676820 259934 676876 259990
rect 675956 259194 676012 259250
rect 676052 258676 676108 258732
rect 676244 256974 676300 257030
rect 676052 256826 676108 256882
rect 676052 256234 676108 256290
rect 676820 253274 676876 253330
rect 679700 255494 679756 255550
rect 679700 254902 679756 254958
rect 685460 254902 685516 254958
rect 685460 254458 685516 254514
rect 676916 253126 676972 253182
rect 675764 250758 675820 250814
rect 675572 249574 675628 249630
rect 675668 243506 675724 243562
rect 675380 242026 675436 242082
rect 675476 240546 675532 240602
rect 675764 238622 675820 238678
rect 675764 236846 675820 236902
rect 676244 221789 676246 221806
rect 676246 221789 676298 221806
rect 676298 221789 676300 221806
rect 676244 221750 676300 221789
rect 676148 221158 676204 221214
rect 676052 220605 676054 220622
rect 676054 220605 676106 220622
rect 676106 220605 676108 220622
rect 676052 220566 676108 220605
rect 676052 219495 676054 219512
rect 676054 219495 676106 219512
rect 676106 219495 676108 219512
rect 676052 219456 676108 219495
rect 672980 219086 673036 219142
rect 676244 220714 676300 220770
rect 672788 217902 672844 217958
rect 676916 216718 676972 216774
rect 675764 216422 675820 216478
rect 676820 214794 676876 214850
rect 676052 214572 676108 214628
rect 675956 214054 676012 214110
rect 676052 212574 676108 212630
rect 676052 211982 676108 212038
rect 675956 211020 676012 211076
rect 676244 211390 676300 211446
rect 676820 207542 676876 207598
rect 679796 210650 679852 210706
rect 679796 209762 679852 209818
rect 685460 209762 685516 209818
rect 676916 207394 676972 207450
rect 685460 209318 685516 209374
rect 675764 204434 675820 204490
rect 675668 202658 675724 202714
rect 675572 201326 675628 201382
rect 675764 198366 675820 198422
rect 675476 195258 675532 195314
rect 675764 193482 675820 193538
rect 675764 191558 675820 191614
rect 676340 177350 676396 177406
rect 676148 176758 676204 176814
rect 676244 176314 676300 176370
rect 672596 173502 672652 173558
rect 676244 171874 676300 171930
rect 676052 170172 676108 170228
rect 676052 169654 676108 169710
rect 676244 168914 676300 168970
rect 676052 166620 676108 166676
rect 676052 166102 676108 166158
rect 676148 165510 676204 165566
rect 676244 164918 676300 164974
rect 675764 159294 675820 159350
rect 675764 157666 675820 157722
rect 675764 155446 675820 155502
rect 675476 153374 675532 153430
rect 675380 152486 675436 152542
rect 675476 152190 675532 152246
rect 675476 150266 675532 150322
rect 675476 148490 675532 148546
rect 675764 146566 675820 146622
rect 676148 131766 676204 131822
rect 676340 131174 676396 131230
rect 676244 130730 676300 130786
rect 676244 129694 676300 129750
rect 676148 128806 676204 128862
rect 676052 127548 676108 127604
rect 676244 127770 676300 127826
rect 676916 126734 676972 126790
rect 647060 111342 647116 111398
rect 646676 109418 646732 109474
rect 646772 107938 646828 107994
rect 665204 105570 665260 105626
rect 647924 104090 647980 104146
rect 647924 99650 647980 99706
rect 647156 98022 647212 98078
rect 647732 94026 647788 94082
rect 647828 92694 647884 92750
rect 647924 87070 647980 87126
rect 650900 86182 650956 86238
rect 652340 85294 652396 85350
rect 651764 84258 651820 84314
rect 652244 83370 652300 83426
rect 647924 82630 647980 82686
rect 647924 81002 647980 81058
rect 647924 77489 647926 77506
rect 647926 77489 647978 77506
rect 647978 77489 647980 77506
rect 647924 77450 647980 77489
rect 646964 71826 647020 71882
rect 646868 68570 646924 68626
rect 647924 73602 647980 73658
rect 647924 69623 647980 69662
rect 647924 69606 647926 69623
rect 647926 69606 647978 69623
rect 647978 69606 647980 69623
rect 647924 64130 647980 64186
rect 647924 62206 647980 62262
rect 647060 60282 647116 60338
rect 659348 90770 659404 90826
rect 675572 126438 675628 126494
rect 676052 126068 676108 126124
rect 676820 124810 676876 124866
rect 676244 124366 676300 124422
rect 676052 124070 676108 124126
rect 676052 123478 676108 123534
rect 676052 121998 676108 122054
rect 675956 121036 676012 121092
rect 676244 121406 676300 121462
rect 676052 120518 676108 120574
rect 676148 119778 676204 119834
rect 676244 119334 676300 119390
rect 676916 116670 676972 116726
rect 676820 116078 676876 116134
rect 675764 108086 675820 108142
rect 675476 106606 675532 106662
rect 668276 106014 668332 106070
rect 665300 105126 665356 105182
rect 653684 86922 653740 86978
rect 663284 86330 663340 86386
rect 652436 82630 652492 82686
rect 662420 81611 662476 81650
rect 662420 81594 662422 81611
rect 662422 81594 662474 81611
rect 662474 81594 662476 81611
rect 663284 84702 663340 84758
rect 663476 83962 663532 84018
rect 663380 82778 663436 82834
rect 663284 82038 663340 82094
rect 646772 57026 646828 57082
rect 646484 54658 646540 54714
rect 675380 105126 675436 105182
rect 675764 103202 675820 103258
rect 675764 101426 675820 101482
rect 512180 41782 512236 41838
rect 525908 41782 525964 41838
rect 539732 40450 539788 40506
rect 311156 31570 311212 31626
rect 328340 31609 328342 31626
rect 328342 31609 328394 31626
rect 328394 31609 328396 31626
rect 328340 31570 328396 31609
<< metal3 >>
rect 81135 1002360 81201 1002363
rect 184047 1002360 184113 1002363
rect 482607 1002360 482673 1002363
rect 81135 1002358 81312 1002360
rect 81135 1002302 81140 1002358
rect 81196 1002302 81312 1002358
rect 81135 1002300 81312 1002302
rect 184032 1002358 184113 1002360
rect 184032 1002302 184052 1002358
rect 184108 1002302 184113 1002358
rect 184032 1002300 184113 1002302
rect 482592 1002358 482673 1002360
rect 482592 1002302 482612 1002358
rect 482668 1002302 482673 1002358
rect 482592 1002300 482673 1002302
rect 81135 1002297 81201 1002300
rect 184047 1002297 184113 1002300
rect 482607 1002297 482673 1002300
rect 394575 997772 394641 997775
rect 535695 997772 535761 997775
rect 636495 997772 636561 997775
rect 393696 997770 394641 997772
rect 132399 997180 132465 997183
rect 132546 997180 132606 997742
rect 241218 997183 241278 997742
rect 132399 997178 132606 997180
rect 132399 997122 132404 997178
rect 132460 997122 132606 997178
rect 132399 997120 132606 997122
rect 241167 997178 241278 997183
rect 241167 997122 241172 997178
rect 241228 997122 241278 997178
rect 241167 997120 241278 997122
rect 290799 997180 290865 997183
rect 292098 997180 292158 997742
rect 393696 997714 394580 997770
rect 394636 997714 394641 997770
rect 393696 997712 394641 997714
rect 534048 997770 535761 997772
rect 534048 997714 535700 997770
rect 535756 997714 535761 997770
rect 534048 997712 535761 997714
rect 635808 997770 636561 997772
rect 635808 997714 636500 997770
rect 636556 997714 636561 997770
rect 635808 997712 636561 997714
rect 394575 997709 394641 997712
rect 535695 997709 535761 997712
rect 636495 997709 636561 997712
rect 290799 997178 292158 997180
rect 290799 997122 290804 997178
rect 290860 997122 292158 997178
rect 290799 997120 292158 997122
rect 132399 997117 132465 997120
rect 241167 997117 241233 997120
rect 290799 997117 290865 997120
rect 290799 983268 290865 983271
rect 397455 983268 397521 983271
rect 290799 983266 293118 983268
rect 290799 983210 290804 983266
rect 290860 983210 293118 983266
rect 290799 983208 293118 983210
rect 290799 983205 290865 983208
rect 292143 983120 292209 983123
rect 292098 983118 292209 983120
rect 292098 983062 292148 983118
rect 292204 983062 292209 983118
rect 292098 983057 292209 983062
rect 80559 982972 80625 982975
rect 132399 982972 132465 982975
rect 184239 982972 184305 982975
rect 233199 982972 233265 982975
rect 240879 982972 240945 982975
rect 80559 982970 81726 982972
rect 80559 982914 80564 982970
rect 80620 982914 81726 982970
rect 80559 982912 81726 982914
rect 80559 982909 80625 982912
rect 81666 982646 81726 982912
rect 132399 982970 133566 982972
rect 132399 982914 132404 982970
rect 132460 982914 133566 982970
rect 132399 982912 133566 982914
rect 132399 982909 132465 982912
rect 133506 982646 133566 982912
rect 184239 982970 185598 982972
rect 184239 982914 184244 982970
rect 184300 982914 185598 982970
rect 184239 982912 185598 982914
rect 184239 982909 184305 982912
rect 185538 982646 185598 982912
rect 233199 982970 236286 982972
rect 233199 982914 233204 982970
rect 233260 982914 236286 982970
rect 233199 982912 236286 982914
rect 233199 982909 233265 982912
rect 236226 982646 236286 982912
rect 240834 982970 240945 982972
rect 240834 982914 240884 982970
rect 240940 982914 240945 982970
rect 240834 982909 240945 982914
rect 241167 982972 241233 982975
rect 285039 982972 285105 982975
rect 241167 982970 241278 982972
rect 241167 982914 241172 982970
rect 241228 982914 241278 982970
rect 241167 982909 241278 982914
rect 285039 982970 288126 982972
rect 285039 982914 285044 982970
rect 285100 982914 288126 982970
rect 285039 982912 288126 982914
rect 285039 982909 285105 982912
rect 240834 982646 240894 982909
rect 241218 982646 241278 982909
rect 288066 982646 288126 982912
rect 292098 982646 292158 983057
rect 293058 982646 293118 983208
rect 397455 983266 397566 983268
rect 397455 983210 397460 983266
rect 397516 983210 397566 983266
rect 397455 983205 397566 983210
rect 391599 982972 391665 982975
rect 394575 982972 394641 982975
rect 391554 982970 391665 982972
rect 391554 982914 391604 982970
rect 391660 982914 391665 982970
rect 391554 982909 391665 982914
rect 394242 982970 394641 982972
rect 394242 982914 394580 982970
rect 394636 982914 394641 982970
rect 394242 982912 394641 982914
rect 391554 982646 391614 982909
rect 394242 982646 394302 982912
rect 394575 982909 394641 982912
rect 397506 982646 397566 983205
rect 636495 983120 636561 983123
rect 636495 983118 636606 983120
rect 636495 983062 636500 983118
rect 636556 983062 636606 983118
rect 636495 983057 636606 983062
rect 483855 982972 483921 982975
rect 538575 982972 538641 982975
rect 483522 982970 483921 982972
rect 483522 982914 483860 982970
rect 483916 982914 483921 982970
rect 483522 982912 483921 982914
rect 483522 982646 483582 982912
rect 483855 982909 483921 982912
rect 535554 982970 538641 982972
rect 535554 982914 538580 982970
rect 538636 982914 538641 982970
rect 535554 982912 538641 982914
rect 535554 982646 535614 982912
rect 538575 982909 538641 982912
rect 636546 982646 636606 983057
rect 40143 959292 40209 959295
rect 39840 959290 40209 959292
rect 39840 959234 40148 959290
rect 40204 959234 40209 959290
rect 39840 959232 40209 959234
rect 40143 959229 40209 959232
rect 60015 959144 60081 959147
rect 653775 959144 653841 959147
rect 60015 959142 65376 959144
rect 60015 959086 60020 959142
rect 60076 959086 65376 959142
rect 60015 959084 65376 959086
rect 649248 959142 653841 959144
rect 649248 959086 653780 959142
rect 653836 959086 653841 959142
rect 649248 959084 653841 959086
rect 60015 959081 60081 959084
rect 653775 959081 653841 959084
rect 676815 950412 676881 950415
rect 676815 950410 677664 950412
rect 676815 950354 676820 950410
rect 676876 950354 677664 950410
rect 676815 950352 677664 950354
rect 676815 950349 676881 950352
rect 676143 894172 676209 894175
rect 676290 894172 676350 894438
rect 676143 894170 676350 894172
rect 676143 894114 676148 894170
rect 676204 894114 676350 894170
rect 676143 894112 676350 894114
rect 676143 894109 676209 894112
rect 676290 893583 676350 893920
rect 676239 893578 676350 893583
rect 676239 893522 676244 893578
rect 676300 893522 676350 893578
rect 676239 893520 676350 893522
rect 676239 893517 676305 893520
rect 676047 893432 676113 893435
rect 676047 893430 676320 893432
rect 676047 893374 676052 893430
rect 676108 893374 676320 893430
rect 676047 893372 676320 893374
rect 676047 893369 676113 893372
rect 676047 892470 676113 892473
rect 676047 892468 676320 892470
rect 676047 892412 676052 892468
rect 676108 892412 676320 892468
rect 676047 892410 676320 892412
rect 676047 892407 676113 892410
rect 676047 891508 676113 891511
rect 676047 891506 676320 891508
rect 676047 891450 676052 891506
rect 676108 891450 676320 891506
rect 676047 891448 676320 891450
rect 676047 891445 676113 891448
rect 676047 890472 676113 890475
rect 676047 890470 676320 890472
rect 676047 890414 676052 890470
rect 676108 890414 676320 890470
rect 676047 890412 676320 890414
rect 676047 890409 676113 890412
rect 680175 890176 680241 890179
rect 680130 890174 680241 890176
rect 680130 890118 680180 890174
rect 680236 890118 680241 890174
rect 680130 890113 680241 890118
rect 680130 889998 680190 890113
rect 676290 889291 676350 889406
rect 676239 889286 676350 889291
rect 676239 889230 676244 889286
rect 676300 889230 676350 889286
rect 676239 889228 676350 889230
rect 676239 889225 676305 889228
rect 679938 888699 679998 888888
rect 679938 888694 680049 888699
rect 679938 888638 679988 888694
rect 680044 888638 680049 888694
rect 679938 888636 680049 888638
rect 679983 888633 680049 888636
rect 680130 888255 680190 888518
rect 680079 888250 680190 888255
rect 680079 888194 680084 888250
rect 680140 888194 680190 888250
rect 680079 888192 680190 888194
rect 680079 888189 680145 888192
rect 676290 887811 676350 887926
rect 676239 887806 676350 887811
rect 676239 887750 676244 887806
rect 676300 887750 676350 887806
rect 676239 887748 676350 887750
rect 676239 887745 676305 887748
rect 676047 887438 676113 887441
rect 676047 887436 676320 887438
rect 676047 887380 676052 887436
rect 676108 887380 676320 887436
rect 676047 887378 676320 887380
rect 676047 887375 676113 887378
rect 679746 886775 679806 887038
rect 679695 886770 679806 886775
rect 679695 886714 679700 886770
rect 679756 886714 679806 886770
rect 679695 886712 679806 886714
rect 679695 886709 679761 886712
rect 679746 886183 679806 886446
rect 679746 886178 679857 886183
rect 679746 886122 679796 886178
rect 679852 886122 679857 886178
rect 679746 886120 679857 886122
rect 679791 886117 679857 886120
rect 679938 885739 679998 885854
rect 679887 885734 679998 885739
rect 679887 885678 679892 885734
rect 679948 885678 679998 885734
rect 679887 885676 679998 885678
rect 679887 885673 679953 885676
rect 676047 885514 676113 885517
rect 676047 885512 676320 885514
rect 676047 885456 676052 885512
rect 676108 885456 676320 885512
rect 676047 885454 676320 885456
rect 676047 885451 676113 885454
rect 676047 884996 676113 884999
rect 676047 884994 676320 884996
rect 676047 884938 676052 884994
rect 676108 884938 676320 884994
rect 676047 884936 676320 884938
rect 676047 884933 676113 884936
rect 675759 884404 675825 884407
rect 675759 884402 676320 884404
rect 675759 884346 675764 884402
rect 675820 884346 676320 884402
rect 675759 884344 676320 884346
rect 675759 884341 675825 884344
rect 676047 884034 676113 884037
rect 676047 884032 676320 884034
rect 676047 883976 676052 884032
rect 676108 883976 676320 884032
rect 676047 883974 676320 883976
rect 676047 883971 676113 883974
rect 676047 883516 676113 883519
rect 676047 883514 676320 883516
rect 676047 883458 676052 883514
rect 676108 883458 676320 883514
rect 676047 883456 676320 883458
rect 676047 883453 676113 883456
rect 679746 882779 679806 882894
rect 679695 882774 679806 882779
rect 679695 882718 679700 882774
rect 679756 882718 679806 882774
rect 679695 882716 679806 882718
rect 679695 882713 679761 882716
rect 685506 882187 685566 882450
rect 679695 882184 679761 882187
rect 679695 882182 679806 882184
rect 679695 882126 679700 882182
rect 679756 882126 679806 882182
rect 679695 882121 679806 882126
rect 685455 882182 685566 882187
rect 685455 882126 685460 882182
rect 685516 882126 685566 882182
rect 685455 882124 685566 882126
rect 685455 882121 685521 882124
rect 679746 882006 679806 882121
rect 685455 881740 685521 881743
rect 685455 881738 685566 881740
rect 685455 881682 685460 881738
rect 685516 881682 685566 881738
rect 685455 881677 685566 881682
rect 685506 881414 685566 881677
rect 655215 868864 655281 868867
rect 649986 868862 655281 868864
rect 649986 868806 655220 868862
rect 655276 868806 655281 868862
rect 649986 868804 655281 868806
rect 649986 868246 650046 868804
rect 655215 868801 655281 868804
rect 655407 867680 655473 867683
rect 649986 867678 655473 867680
rect 649986 867622 655412 867678
rect 655468 867622 655473 867678
rect 649986 867620 655473 867622
rect 649986 867064 650046 867620
rect 655407 867617 655473 867620
rect 655119 866496 655185 866499
rect 649986 866494 655185 866496
rect 649986 866438 655124 866494
rect 655180 866438 655185 866494
rect 649986 866436 655185 866438
rect 649986 865882 650046 866436
rect 655119 866433 655185 866436
rect 655311 865312 655377 865315
rect 649986 865310 655377 865312
rect 649986 865254 655316 865310
rect 655372 865254 655377 865310
rect 649986 865252 655377 865254
rect 649986 864700 650046 865252
rect 655311 865249 655377 865252
rect 654159 863980 654225 863983
rect 649986 863978 654225 863980
rect 649986 863922 654164 863978
rect 654220 863922 654225 863978
rect 649986 863920 654225 863922
rect 649986 863518 650046 863920
rect 654159 863917 654225 863920
rect 653775 862944 653841 862947
rect 649986 862942 653841 862944
rect 649986 862886 653780 862942
rect 653836 862886 653841 862942
rect 649986 862884 653841 862886
rect 649986 862336 650046 862884
rect 653775 862881 653841 862884
rect 41775 817952 41841 817955
rect 41568 817950 41841 817952
rect 41568 817894 41780 817950
rect 41836 817894 41841 817950
rect 41568 817892 41841 817894
rect 41775 817889 41841 817892
rect 41775 817360 41841 817363
rect 41568 817358 41841 817360
rect 41568 817302 41780 817358
rect 41836 817302 41841 817358
rect 41568 817300 41841 817302
rect 41775 817297 41841 817300
rect 41538 816623 41598 816738
rect 41538 816618 41649 816623
rect 41538 816562 41588 816618
rect 41644 816562 41649 816618
rect 41538 816560 41649 816562
rect 41583 816557 41649 816560
rect 41775 815880 41841 815883
rect 41568 815878 41841 815880
rect 41568 815822 41780 815878
rect 41836 815822 41841 815878
rect 41568 815820 41841 815822
rect 41775 815817 41841 815820
rect 40386 815142 40446 815258
rect 40378 815078 40384 815142
rect 40448 815078 40454 815142
rect 41775 814918 41841 814921
rect 41568 814916 41841 814918
rect 41568 814860 41780 814916
rect 41836 814860 41841 814916
rect 41568 814858 41841 814860
rect 41775 814855 41841 814858
rect 40578 814106 40638 814370
rect 40570 814042 40576 814106
rect 40640 814042 40646 814106
rect 41538 813663 41598 813778
rect 41538 813658 41649 813663
rect 41538 813602 41588 813658
rect 41644 813602 41649 813658
rect 41538 813600 41649 813602
rect 41583 813597 41649 813600
rect 41538 813219 41598 813334
rect 41538 813214 41649 813219
rect 41538 813158 41588 813214
rect 41644 813158 41649 813214
rect 41538 813156 41649 813158
rect 41583 813153 41649 813156
rect 42543 812920 42609 812923
rect 41568 812918 42609 812920
rect 41568 812862 42548 812918
rect 42604 812862 42609 812918
rect 41568 812860 42609 812862
rect 42543 812857 42609 812860
rect 40239 812476 40305 812479
rect 40194 812474 40305 812476
rect 40194 812418 40244 812474
rect 40300 812418 40305 812474
rect 40194 812413 40305 812418
rect 40194 812298 40254 812413
rect 41538 811739 41598 811854
rect 41538 811734 41649 811739
rect 41538 811678 41588 811734
rect 41644 811678 41649 811734
rect 41538 811676 41649 811678
rect 41583 811673 41649 811676
rect 41967 811366 42033 811369
rect 41568 811364 42033 811366
rect 41568 811308 41972 811364
rect 42028 811308 42033 811364
rect 41568 811306 42033 811308
rect 41967 811303 42033 811306
rect 41871 810848 41937 810851
rect 41568 810846 41937 810848
rect 41568 810790 41876 810846
rect 41932 810790 41937 810846
rect 41568 810788 41937 810790
rect 41871 810785 41937 810788
rect 41538 810258 41598 810374
rect 41530 810194 41536 810258
rect 41600 810194 41606 810258
rect 41775 809886 41841 809889
rect 41568 809884 41841 809886
rect 41568 809828 41780 809884
rect 41836 809828 41841 809884
rect 41568 809826 41841 809828
rect 41775 809823 41841 809826
rect 42063 809368 42129 809371
rect 41568 809366 42129 809368
rect 41568 809310 42068 809366
rect 42124 809310 42129 809366
rect 41568 809308 42129 809310
rect 42063 809305 42129 809308
rect 41775 808924 41841 808927
rect 41568 808922 41841 808924
rect 41568 808866 41780 808922
rect 41836 808866 41841 808922
rect 41568 808864 41841 808866
rect 41775 808861 41841 808864
rect 41538 808184 41598 808302
rect 41679 808184 41745 808187
rect 41538 808182 41745 808184
rect 41538 808126 41684 808182
rect 41740 808126 41745 808182
rect 41538 808124 41745 808126
rect 41679 808121 41745 808124
rect 42159 807888 42225 807891
rect 41568 807886 42225 807888
rect 41568 807830 42164 807886
rect 42220 807830 42225 807886
rect 41568 807828 42225 807830
rect 42159 807825 42225 807828
rect 41775 807444 41841 807447
rect 41568 807442 41841 807444
rect 41568 807386 41780 807442
rect 41836 807386 41841 807442
rect 41568 807384 41841 807386
rect 41775 807381 41841 807384
rect 41538 806707 41598 806822
rect 41538 806702 41649 806707
rect 41538 806646 41588 806702
rect 41644 806646 41649 806702
rect 41538 806644 41649 806646
rect 41583 806641 41649 806644
rect 41538 806115 41598 806304
rect 41538 806110 41649 806115
rect 41538 806054 41588 806110
rect 41644 806054 41649 806110
rect 41538 806052 41649 806054
rect 41583 806049 41649 806052
rect 28866 805671 28926 805934
rect 28815 805666 28926 805671
rect 28815 805610 28820 805666
rect 28876 805610 28926 805666
rect 28815 805608 28926 805610
rect 28815 805605 28881 805608
rect 41538 805227 41598 805342
rect 28815 805224 28881 805227
rect 28815 805222 28926 805224
rect 28815 805166 28820 805222
rect 28876 805166 28926 805222
rect 28815 805161 28926 805166
rect 41538 805222 41649 805227
rect 41538 805166 41588 805222
rect 41644 805166 41649 805222
rect 41538 805164 41649 805166
rect 41583 805161 41649 805164
rect 28866 804824 28926 805161
rect 40239 802116 40305 802119
rect 41338 802116 41344 802118
rect 40239 802114 41344 802116
rect 40239 802058 40244 802114
rect 40300 802058 41344 802114
rect 40239 802056 41344 802058
rect 40239 802053 40305 802056
rect 41338 802054 41344 802056
rect 41408 802054 41414 802118
rect 42735 800934 42801 800935
rect 42682 800870 42688 800934
rect 42752 800932 42801 800934
rect 42752 800930 42844 800932
rect 42796 800874 42844 800930
rect 42752 800872 42844 800874
rect 42752 800870 42801 800872
rect 42735 800869 42801 800870
rect 41679 800490 41745 800491
rect 42063 800490 42129 800491
rect 41679 800488 41728 800490
rect 41636 800486 41728 800488
rect 41636 800430 41684 800486
rect 41636 800428 41728 800430
rect 41679 800426 41728 800428
rect 41792 800426 41798 800490
rect 42063 800488 42112 800490
rect 42020 800486 42112 800488
rect 42020 800430 42068 800486
rect 42020 800428 42112 800430
rect 42063 800426 42112 800428
rect 42176 800426 42182 800490
rect 41679 800425 41745 800426
rect 42063 800425 42129 800426
rect 41967 800342 42033 800343
rect 41914 800278 41920 800342
rect 41984 800340 42033 800342
rect 41984 800338 42076 800340
rect 42028 800282 42076 800338
rect 41984 800280 42076 800282
rect 41984 800278 42033 800280
rect 41967 800277 42033 800278
rect 41775 794274 41841 794275
rect 41722 794272 41728 794274
rect 41684 794212 41728 794272
rect 41792 794270 41841 794274
rect 41836 794214 41841 794270
rect 41722 794210 41728 794212
rect 41792 794210 41841 794214
rect 41775 794209 41841 794210
rect 42735 793534 42801 793535
rect 42682 793532 42688 793534
rect 42644 793472 42688 793532
rect 42752 793530 42801 793534
rect 42796 793474 42801 793530
rect 42682 793470 42688 793472
rect 42752 793470 42801 793474
rect 42735 793469 42801 793470
rect 41967 792942 42033 792943
rect 41914 792940 41920 792942
rect 41876 792880 41920 792940
rect 41984 792938 42033 792942
rect 42028 792882 42033 792938
rect 41914 792878 41920 792880
rect 41984 792878 42033 792882
rect 41967 792877 42033 792878
rect 57711 790868 57777 790871
rect 57711 790866 64638 790868
rect 57711 790810 57716 790866
rect 57772 790810 64638 790866
rect 57711 790808 64638 790810
rect 57711 790805 57777 790808
rect 64578 790304 64638 790808
rect 42159 790130 42225 790131
rect 42106 790128 42112 790130
rect 42068 790068 42112 790128
rect 42176 790126 42225 790130
rect 42220 790070 42225 790126
rect 42106 790066 42112 790068
rect 42176 790066 42225 790070
rect 42159 790065 42225 790066
rect 57615 789684 57681 789687
rect 57615 789682 64638 789684
rect 57615 789626 57620 789682
rect 57676 789626 64638 789682
rect 57615 789624 64638 789626
rect 57615 789621 57681 789624
rect 41338 789326 41344 789390
rect 41408 789388 41414 789390
rect 42831 789388 42897 789391
rect 41408 789386 42897 789388
rect 41408 789330 42836 789386
rect 42892 789330 42897 789386
rect 41408 789328 42897 789330
rect 41408 789326 41414 789328
rect 42831 789325 42897 789328
rect 41530 789178 41536 789242
rect 41600 789240 41606 789242
rect 42735 789240 42801 789243
rect 41600 789238 42801 789240
rect 41600 789182 42740 789238
rect 42796 789182 42801 789238
rect 41600 789180 42801 789182
rect 41600 789178 41606 789180
rect 42735 789177 42801 789180
rect 64578 789122 64638 789624
rect 58191 788500 58257 788503
rect 58191 788498 64638 788500
rect 58191 788442 58196 788498
rect 58252 788442 64638 788498
rect 58191 788440 64638 788442
rect 58191 788437 58257 788440
rect 64578 787940 64638 788440
rect 674746 787994 674752 788058
rect 674816 788056 674822 788058
rect 675375 788056 675441 788059
rect 674816 788054 675441 788056
rect 674816 787998 675380 788054
rect 675436 787998 675441 788054
rect 674816 787996 675441 787998
rect 674816 787994 674822 787996
rect 675375 787993 675441 787996
rect 675759 787464 675825 787467
rect 676090 787464 676096 787466
rect 675759 787462 676096 787464
rect 675759 787406 675764 787462
rect 675820 787406 676096 787462
rect 675759 787404 676096 787406
rect 675759 787401 675825 787404
rect 676090 787402 676096 787404
rect 676160 787402 676166 787466
rect 58383 787316 58449 787319
rect 58383 787314 64638 787316
rect 58383 787258 58388 787314
rect 58444 787258 64638 787314
rect 58383 787256 64638 787258
rect 58383 787253 58449 787256
rect 64578 786758 64638 787256
rect 675471 786726 675537 786727
rect 675471 786722 675520 786726
rect 675584 786724 675590 786726
rect 675471 786666 675476 786722
rect 675471 786662 675520 786666
rect 675584 786664 675628 786724
rect 675584 786662 675590 786664
rect 675471 786661 675537 786662
rect 59631 785540 59697 785543
rect 64578 785540 64638 785576
rect 59631 785538 64638 785540
rect 59631 785482 59636 785538
rect 59692 785482 64638 785538
rect 59631 785480 64638 785482
rect 59631 785477 59697 785480
rect 59151 784948 59217 784951
rect 59151 784946 64638 784948
rect 59151 784890 59156 784946
rect 59212 784890 64638 784946
rect 59151 784888 64638 784890
rect 59151 784885 59217 784888
rect 64578 784394 64638 784888
rect 675130 784738 675136 784802
rect 675200 784800 675206 784802
rect 675375 784800 675441 784803
rect 675200 784798 675441 784800
rect 675200 784742 675380 784798
rect 675436 784742 675441 784798
rect 675200 784740 675441 784742
rect 675200 784738 675206 784740
rect 675375 784737 675441 784740
rect 674362 784146 674368 784210
rect 674432 784208 674438 784210
rect 675471 784208 675537 784211
rect 674432 784206 675537 784208
rect 674432 784150 675476 784206
rect 675532 784150 675537 784206
rect 674432 784148 675537 784150
rect 674432 784146 674438 784148
rect 675471 784145 675537 784148
rect 673978 783406 673984 783470
rect 674048 783468 674054 783470
rect 675279 783468 675345 783471
rect 674048 783466 675345 783468
rect 674048 783410 675284 783466
rect 675340 783410 675345 783466
rect 674048 783408 675345 783410
rect 674048 783406 674054 783408
rect 675279 783405 675345 783408
rect 675759 783024 675825 783027
rect 676474 783024 676480 783026
rect 675759 783022 676480 783024
rect 675759 782966 675764 783022
rect 675820 782966 676480 783022
rect 675759 782964 676480 782966
rect 675759 782961 675825 782964
rect 676474 782962 676480 782964
rect 676544 782962 676550 783026
rect 675663 780658 675729 780659
rect 675663 780654 675712 780658
rect 675776 780656 675782 780658
rect 675663 780598 675668 780654
rect 675663 780594 675712 780598
rect 675776 780596 675820 780656
rect 675776 780594 675782 780596
rect 675663 780593 675729 780594
rect 675759 779916 675825 779919
rect 676282 779916 676288 779918
rect 675759 779914 676288 779916
rect 675759 779858 675764 779914
rect 675820 779858 676288 779914
rect 675759 779856 676288 779858
rect 675759 779853 675825 779856
rect 676282 779854 676288 779856
rect 676352 779854 676358 779918
rect 675759 779176 675825 779179
rect 676666 779176 676672 779178
rect 675759 779174 676672 779176
rect 675759 779118 675764 779174
rect 675820 779118 676672 779174
rect 675759 779116 676672 779118
rect 675759 779113 675825 779116
rect 676666 779114 676672 779116
rect 676736 779114 676742 779178
rect 649986 778288 650046 778824
rect 655215 778288 655281 778291
rect 649986 778286 655281 778288
rect 649986 778230 655220 778286
rect 655276 778230 655281 778286
rect 649986 778228 655281 778230
rect 655215 778225 655281 778228
rect 655407 777696 655473 777699
rect 649986 777694 655473 777696
rect 649986 777638 655412 777694
rect 655468 777638 655473 777694
rect 649986 777636 655473 777638
rect 655407 777633 655473 777636
rect 675322 777634 675328 777698
rect 675392 777696 675398 777698
rect 675471 777696 675537 777699
rect 675392 777694 675537 777696
rect 675392 777638 675476 777694
rect 675532 777638 675537 777694
rect 675392 777636 675537 777638
rect 675392 777634 675398 777636
rect 675471 777633 675537 777636
rect 649986 776068 650046 776460
rect 655599 776068 655665 776071
rect 649986 776066 655665 776068
rect 649986 776010 655604 776066
rect 655660 776010 655665 776066
rect 649986 776008 655665 776010
rect 655599 776005 655665 776008
rect 655119 775920 655185 775923
rect 649986 775918 655185 775920
rect 649986 775862 655124 775918
rect 655180 775862 655185 775918
rect 649986 775860 655185 775862
rect 649986 775278 650046 775860
rect 655119 775857 655185 775860
rect 675759 775476 675825 775479
rect 675898 775476 675904 775478
rect 675759 775474 675904 775476
rect 675759 775418 675764 775474
rect 675820 775418 675904 775474
rect 675759 775416 675904 775418
rect 675759 775413 675825 775416
rect 675898 775414 675904 775416
rect 675968 775414 675974 775478
rect 41775 774736 41841 774739
rect 656559 774736 656625 774739
rect 41568 774734 41841 774736
rect 41568 774678 41780 774734
rect 41836 774678 41841 774734
rect 41568 774676 41841 774678
rect 41775 774673 41841 774676
rect 649986 774734 656625 774736
rect 649986 774678 656564 774734
rect 656620 774678 656625 774734
rect 649986 774676 656625 774678
rect 41538 773999 41598 774114
rect 649986 774096 650046 774676
rect 656559 774673 656625 774676
rect 41538 773994 41649 773999
rect 41538 773938 41588 773994
rect 41644 773938 41649 773994
rect 41538 773936 41649 773938
rect 41583 773933 41649 773936
rect 654351 773552 654417 773555
rect 649986 773550 654417 773552
rect 41538 773407 41598 773522
rect 649986 773494 654356 773550
rect 654412 773494 654417 773550
rect 649986 773492 654417 773494
rect 41538 773402 41649 773407
rect 41538 773346 41588 773402
rect 41644 773346 41649 773402
rect 41538 773344 41649 773346
rect 41583 773341 41649 773344
rect 41775 773256 41841 773259
rect 41568 773254 41841 773256
rect 41568 773198 41780 773254
rect 41836 773198 41841 773254
rect 41568 773196 41841 773198
rect 41775 773193 41841 773196
rect 40570 772898 40576 772962
rect 40640 772960 40646 772962
rect 41583 772960 41649 772963
rect 40640 772958 41649 772960
rect 40640 772902 41588 772958
rect 41644 772902 41649 772958
rect 649986 772914 650046 773492
rect 654351 773489 654417 773492
rect 40640 772900 41649 772902
rect 40640 772898 40646 772900
rect 41583 772897 41649 772900
rect 41775 772664 41841 772667
rect 41568 772662 41841 772664
rect 41568 772606 41780 772662
rect 41836 772606 41841 772662
rect 41568 772604 41841 772606
rect 41775 772601 41841 772604
rect 674991 772072 675057 772075
rect 676090 772072 676096 772074
rect 674991 772070 676096 772072
rect 40386 771872 40446 772042
rect 674991 772014 674996 772070
rect 675052 772014 676096 772070
rect 674991 772012 676096 772014
rect 674991 772009 675057 772012
rect 676090 772010 676096 772012
rect 676160 772010 676166 772074
rect 40378 771808 40384 771872
rect 40448 771808 40454 771872
rect 40570 771862 40576 771926
rect 40640 771924 40646 771926
rect 42735 771924 42801 771927
rect 40640 771922 42801 771924
rect 40640 771866 42740 771922
rect 42796 771866 42801 771922
rect 40640 771864 42801 771866
rect 40640 771862 40646 771864
rect 41538 771672 41598 771864
rect 42735 771861 42801 771864
rect 674895 771924 674961 771927
rect 675514 771924 675520 771926
rect 674895 771922 675520 771924
rect 674895 771866 674900 771922
rect 674956 771866 675520 771922
rect 674895 771864 675520 771866
rect 674895 771861 674961 771864
rect 675514 771862 675520 771864
rect 675584 771862 675590 771926
rect 40578 770890 40638 771154
rect 40570 770826 40576 770890
rect 40640 770826 40646 770890
rect 41583 770888 41649 770891
rect 41538 770886 41649 770888
rect 41538 770830 41588 770886
rect 41644 770830 41649 770886
rect 41538 770825 41649 770830
rect 41538 770562 41598 770825
rect 41346 770003 41406 770192
rect 41346 769998 41457 770003
rect 41346 769942 41396 769998
rect 41452 769942 41457 769998
rect 41346 769940 41457 769942
rect 41391 769937 41457 769940
rect 41967 769704 42033 769707
rect 41568 769702 42033 769704
rect 41568 769646 41972 769702
rect 42028 769646 42033 769702
rect 41568 769644 42033 769646
rect 41967 769641 42033 769644
rect 40194 768967 40254 769082
rect 40194 768962 40305 768967
rect 40194 768906 40244 768962
rect 40300 768906 40305 768962
rect 40194 768904 40305 768906
rect 40239 768901 40305 768904
rect 41538 768520 41598 768638
rect 41679 768520 41745 768523
rect 41538 768518 41745 768520
rect 41538 768462 41684 768518
rect 41740 768462 41745 768518
rect 41538 768460 41745 768462
rect 41679 768457 41745 768460
rect 41775 768224 41841 768227
rect 41568 768222 41841 768224
rect 41568 768166 41780 768222
rect 41836 768166 41841 768222
rect 41568 768164 41841 768166
rect 41775 768161 41841 768164
rect 41871 767632 41937 767635
rect 41568 767630 41937 767632
rect 41568 767574 41876 767630
rect 41932 767574 41937 767630
rect 41568 767572 41937 767574
rect 41871 767569 41937 767572
rect 40770 767042 40830 767158
rect 40762 766978 40768 767042
rect 40832 766978 40838 767042
rect 41538 766451 41598 766640
rect 41487 766446 41598 766451
rect 41487 766390 41492 766446
rect 41548 766390 41598 766446
rect 41487 766388 41598 766390
rect 41487 766385 41553 766388
rect 42063 766152 42129 766155
rect 41568 766150 42129 766152
rect 41568 766094 42068 766150
rect 42124 766094 42129 766150
rect 41568 766092 42129 766094
rect 42063 766089 42129 766092
rect 42159 765708 42225 765711
rect 41568 765706 42225 765708
rect 41568 765650 42164 765706
rect 42220 765650 42225 765706
rect 41568 765648 42225 765650
rect 42159 765645 42225 765648
rect 41775 765190 41841 765193
rect 41568 765188 41841 765190
rect 41568 765132 41780 765188
rect 41836 765132 41841 765188
rect 41568 765130 41841 765132
rect 41775 765127 41841 765130
rect 41722 764672 41728 764674
rect 41568 764612 41728 764672
rect 41722 764610 41728 764612
rect 41792 764610 41798 764674
rect 41775 764228 41841 764231
rect 41568 764226 41841 764228
rect 41568 764170 41780 764226
rect 41836 764170 41841 764226
rect 41568 764168 41841 764170
rect 41775 764165 41841 764168
rect 41538 763491 41598 763606
rect 41538 763486 41649 763491
rect 41538 763430 41588 763486
rect 41644 763430 41649 763486
rect 41538 763428 41649 763430
rect 41583 763425 41649 763428
rect 41538 762896 41598 763162
rect 41538 762836 41790 762896
rect 28866 762455 28926 762718
rect 28815 762450 28926 762455
rect 41730 762452 41790 762836
rect 28815 762394 28820 762450
rect 28876 762394 28926 762450
rect 28815 762392 28926 762394
rect 41538 762392 41790 762452
rect 28815 762389 28881 762392
rect 41538 762156 41598 762392
rect 41775 762156 41841 762159
rect 41538 762154 41841 762156
rect 41538 762126 41780 762154
rect 41568 762098 41780 762126
rect 41836 762098 41841 762154
rect 41568 762096 41841 762098
rect 41775 762093 41841 762096
rect 28815 762008 28881 762011
rect 28815 762006 28926 762008
rect 28815 761950 28820 762006
rect 28876 761950 28926 762006
rect 28815 761945 28926 761950
rect 28866 761608 28926 761945
rect 40239 759936 40305 759939
rect 40954 759936 40960 759938
rect 40239 759934 40960 759936
rect 40239 759878 40244 759934
rect 40300 759878 40960 759934
rect 40239 759876 40960 759878
rect 40239 759873 40305 759876
rect 40954 759874 40960 759876
rect 41024 759874 41030 759938
rect 42831 757866 42897 757867
rect 42831 757864 42880 757866
rect 42788 757862 42880 757864
rect 42788 757806 42836 757862
rect 42788 757804 42880 757806
rect 42831 757802 42880 757804
rect 42944 757802 42950 757866
rect 42831 757801 42897 757802
rect 41679 757420 41745 757423
rect 42106 757420 42112 757422
rect 41679 757418 42112 757420
rect 41679 757362 41684 757418
rect 41740 757362 42112 757418
rect 41679 757360 42112 757362
rect 41679 757357 41745 757360
rect 42106 757358 42112 757360
rect 42176 757358 42182 757422
rect 42063 757272 42129 757275
rect 42298 757272 42304 757274
rect 42063 757270 42304 757272
rect 42063 757214 42068 757270
rect 42124 757214 42304 757270
rect 42063 757212 42304 757214
rect 42063 757209 42129 757212
rect 42298 757210 42304 757212
rect 42368 757210 42374 757274
rect 41967 757126 42033 757127
rect 41914 757062 41920 757126
rect 41984 757124 42033 757126
rect 41984 757122 42076 757124
rect 42028 757066 42076 757122
rect 41984 757064 42076 757066
rect 41984 757062 42033 757064
rect 41967 757061 42033 757062
rect 41967 754906 42033 754907
rect 41914 754904 41920 754906
rect 41876 754844 41920 754904
rect 41984 754902 42033 754906
rect 42028 754846 42033 754902
rect 41914 754842 41920 754844
rect 41984 754842 42033 754846
rect 41967 754841 42033 754842
rect 42927 751354 42993 751355
rect 42874 751290 42880 751354
rect 42944 751352 42993 751354
rect 42944 751350 43036 751352
rect 42988 751294 43036 751350
rect 42944 751292 43036 751294
rect 42944 751290 42993 751292
rect 42927 751289 42993 751290
rect 42106 747738 42112 747802
rect 42176 747800 42182 747802
rect 42447 747800 42513 747803
rect 42176 747798 42513 747800
rect 42176 747742 42452 747798
rect 42508 747742 42513 747798
rect 42176 747740 42513 747742
rect 42176 747738 42182 747740
rect 42447 747737 42513 747740
rect 58671 747652 58737 747655
rect 58671 747650 64638 747652
rect 58671 747594 58676 747650
rect 58732 747594 64638 747650
rect 58671 747592 64638 747594
rect 58671 747589 58737 747592
rect 41775 747506 41841 747507
rect 41722 747504 41728 747506
rect 41684 747444 41728 747504
rect 41792 747502 41841 747506
rect 41836 747446 41841 747502
rect 41722 747442 41728 747444
rect 41792 747442 41841 747446
rect 41775 747441 41841 747442
rect 40762 747146 40768 747210
rect 40832 747208 40838 747210
rect 42927 747208 42993 747211
rect 40832 747206 42993 747208
rect 40832 747150 42932 747206
rect 42988 747150 42993 747206
rect 40832 747148 42993 747150
rect 40832 747146 40838 747148
rect 42927 747145 42993 747148
rect 64578 747082 64638 747592
rect 42159 746912 42225 746915
rect 42298 746912 42304 746914
rect 42159 746910 42304 746912
rect 42159 746854 42164 746910
rect 42220 746854 42304 746910
rect 42159 746852 42304 746854
rect 42159 746849 42225 746852
rect 42298 746850 42304 746852
rect 42368 746850 42374 746914
rect 40954 746554 40960 746618
rect 41024 746616 41030 746618
rect 42351 746616 42417 746619
rect 41024 746614 42417 746616
rect 41024 746558 42356 746614
rect 42412 746558 42417 746614
rect 41024 746556 42417 746558
rect 41024 746554 41030 746556
rect 42351 746553 42417 746556
rect 54735 746024 54801 746027
rect 54690 746022 54801 746024
rect 54690 745966 54740 746022
rect 54796 745966 54801 746022
rect 54690 745961 54801 745966
rect 54690 745879 54750 745961
rect 54639 745874 54750 745879
rect 54639 745818 54644 745874
rect 54700 745818 54750 745874
rect 54639 745816 54750 745818
rect 54639 745813 54705 745816
rect 59631 745432 59697 745435
rect 64578 745432 64638 745900
rect 676282 745814 676288 745878
rect 676352 745876 676358 745878
rect 677242 745876 677248 745878
rect 676352 745816 677248 745876
rect 676352 745814 676358 745816
rect 677242 745814 677248 745816
rect 677312 745814 677318 745878
rect 59631 745430 64638 745432
rect 59631 745374 59636 745430
rect 59692 745374 64638 745430
rect 59631 745372 64638 745374
rect 59631 745369 59697 745372
rect 57615 745284 57681 745287
rect 57615 745282 64638 745284
rect 57615 745226 57620 745282
rect 57676 745226 64638 745282
rect 57615 745224 64638 745226
rect 57615 745221 57681 745224
rect 64578 744718 64638 745224
rect 58191 744100 58257 744103
rect 58191 744098 64638 744100
rect 58191 744042 58196 744098
rect 58252 744042 64638 744098
rect 58191 744040 64638 744042
rect 58191 744037 58257 744040
rect 64578 743536 64638 744040
rect 676474 743002 676480 743066
rect 676544 743064 676550 743066
rect 676858 743064 676864 743066
rect 676544 743004 676864 743064
rect 676544 743002 676550 743004
rect 676858 743002 676864 743004
rect 676928 743002 676934 743066
rect 59631 742916 59697 742919
rect 59631 742914 64638 742916
rect 59631 742858 59636 742914
rect 59692 742858 64638 742914
rect 59631 742856 64638 742858
rect 59631 742853 59697 742856
rect 64578 742354 64638 742856
rect 674170 742410 674176 742474
rect 674240 742472 674246 742474
rect 675471 742472 675537 742475
rect 674240 742470 675537 742472
rect 674240 742414 675476 742470
rect 675532 742414 675537 742470
rect 674240 742412 675537 742414
rect 674240 742410 674246 742412
rect 675471 742409 675537 742412
rect 59727 741732 59793 741735
rect 59727 741730 64638 741732
rect 59727 741674 59732 741730
rect 59788 741674 64638 741730
rect 59727 741672 64638 741674
rect 59727 741669 59793 741672
rect 64578 741172 64638 741672
rect 674938 741078 674944 741142
rect 675008 741140 675014 741142
rect 675183 741140 675249 741143
rect 675008 741138 675249 741140
rect 675008 741082 675188 741138
rect 675244 741082 675249 741138
rect 675008 741080 675249 741082
rect 675008 741078 675014 741080
rect 675183 741077 675249 741080
rect 674554 740338 674560 740402
rect 674624 740400 674630 740402
rect 675471 740400 675537 740403
rect 674624 740398 675537 740400
rect 674624 740342 675476 740398
rect 675532 740342 675537 740398
rect 674624 740340 675537 740342
rect 674624 740338 674630 740340
rect 675471 740337 675537 740340
rect 675471 739218 675537 739219
rect 675471 739214 675520 739218
rect 675584 739216 675590 739218
rect 675471 739158 675476 739214
rect 675471 739154 675520 739158
rect 675584 739156 675628 739216
rect 675584 739154 675590 739156
rect 675471 739153 675537 739154
rect 675759 735516 675825 735519
rect 676282 735516 676288 735518
rect 675759 735514 676288 735516
rect 675759 735458 675764 735514
rect 675820 735458 676288 735514
rect 675759 735456 676288 735458
rect 675759 735453 675825 735456
rect 676282 735454 676288 735456
rect 676352 735454 676358 735518
rect 655119 734480 655185 734483
rect 649986 734478 655185 734480
rect 649986 734422 655124 734478
rect 655180 734422 655185 734478
rect 649986 734420 655185 734422
rect 649986 734402 650046 734420
rect 655119 734417 655185 734420
rect 649986 732704 650046 733220
rect 655503 732704 655569 732707
rect 649986 732702 655569 732704
rect 649986 732646 655508 732702
rect 655564 732646 655569 732702
rect 649986 732644 655569 732646
rect 655503 732641 655569 732644
rect 649986 731668 650046 732038
rect 655311 731668 655377 731671
rect 649986 731666 655377 731668
rect 649986 731610 655316 731666
rect 655372 731610 655377 731666
rect 649986 731608 655377 731610
rect 655311 731605 655377 731608
rect 41775 731520 41841 731523
rect 41568 731518 41841 731520
rect 41568 731462 41780 731518
rect 41836 731462 41841 731518
rect 41568 731460 41841 731462
rect 41775 731457 41841 731460
rect 655695 731372 655761 731375
rect 649986 731370 655761 731372
rect 649986 731314 655700 731370
rect 655756 731314 655761 731370
rect 649986 731312 655761 731314
rect 41538 730783 41598 730898
rect 649986 730856 650046 731312
rect 655695 731309 655761 731312
rect 41538 730778 41649 730783
rect 41538 730722 41588 730778
rect 41644 730722 41649 730778
rect 41538 730720 41649 730722
rect 41583 730717 41649 730720
rect 674415 730632 674481 730635
rect 676090 730632 676096 730634
rect 674415 730630 676096 730632
rect 674415 730574 674420 730630
rect 674476 730574 676096 730630
rect 674415 730572 676096 730574
rect 674415 730569 674481 730572
rect 676090 730570 676096 730572
rect 676160 730570 676166 730634
rect 41775 730410 41841 730413
rect 41568 730408 41841 730410
rect 41568 730352 41780 730408
rect 41836 730352 41841 730408
rect 41568 730350 41841 730352
rect 41775 730347 41841 730350
rect 41583 730188 41649 730191
rect 654063 730188 654129 730191
rect 41538 730186 41649 730188
rect 41538 730130 41588 730186
rect 41644 730130 41649 730186
rect 41538 730125 41649 730130
rect 649986 730186 654129 730188
rect 649986 730130 654068 730186
rect 654124 730130 654129 730186
rect 649986 730128 654129 730130
rect 41538 730010 41598 730125
rect 649986 729674 650046 730128
rect 654063 730125 654129 730128
rect 676858 729830 676864 729894
rect 676928 729830 676934 729894
rect 676866 729448 676926 729830
rect 677050 729448 677056 729450
rect 41538 729303 41598 729418
rect 676866 729388 677056 729448
rect 677050 729386 677056 729388
rect 677120 729386 677126 729450
rect 40570 729238 40576 729302
rect 40640 729300 40646 729302
rect 41391 729300 41457 729303
rect 40640 729298 41457 729300
rect 40640 729242 41396 729298
rect 41452 729242 41457 729298
rect 40640 729240 41457 729242
rect 41538 729298 41649 729303
rect 41538 729242 41588 729298
rect 41644 729242 41649 729298
rect 41538 729240 41649 729242
rect 40640 729238 40646 729240
rect 41391 729237 41457 729240
rect 41583 729237 41649 729240
rect 41775 728856 41841 728859
rect 41568 728854 41841 728856
rect 41568 728798 41780 728854
rect 41836 728798 41841 728854
rect 41568 728796 41841 728798
rect 41775 728793 41841 728796
rect 40431 728710 40497 728711
rect 40378 728646 40384 728710
rect 40448 728708 40497 728710
rect 40448 728706 40576 728708
rect 40492 728650 40576 728706
rect 40448 728648 40576 728650
rect 40448 728646 40497 728648
rect 40386 728645 40497 728646
rect 40386 728530 40446 728645
rect 654159 728560 654225 728563
rect 649986 728558 654225 728560
rect 649986 728502 654164 728558
rect 654220 728502 654225 728558
rect 649986 728500 654225 728502
rect 649986 728492 650046 728500
rect 654159 728497 654225 728500
rect 676666 728054 676672 728118
rect 676736 728116 676742 728118
rect 677242 728116 677248 728118
rect 676736 728056 677248 728116
rect 676736 728054 676742 728056
rect 677242 728054 677248 728056
rect 677312 728054 677318 728118
rect 41775 727968 41841 727971
rect 41568 727966 41841 727968
rect 41568 727910 41780 727966
rect 41836 727910 41841 727966
rect 41568 727908 41841 727910
rect 41775 727905 41841 727908
rect 40570 727610 40576 727674
rect 40640 727610 40646 727674
rect 40578 727346 40638 727610
rect 41538 726787 41598 726976
rect 41487 726782 41598 726787
rect 41487 726726 41492 726782
rect 41548 726726 41598 726782
rect 41487 726724 41598 726726
rect 41487 726721 41553 726724
rect 42063 726488 42129 726491
rect 41568 726486 42129 726488
rect 41568 726430 42068 726486
rect 42124 726430 42129 726486
rect 41568 726428 42129 726430
rect 42063 726425 42129 726428
rect 34434 725751 34494 725866
rect 34383 725746 34494 725751
rect 34383 725690 34388 725746
rect 34444 725690 34494 725746
rect 34383 725688 34494 725690
rect 34383 725685 34449 725688
rect 41967 725526 42033 725529
rect 41568 725524 42033 725526
rect 41568 725468 41972 725524
rect 42028 725468 42033 725524
rect 41568 725466 42033 725468
rect 41967 725463 42033 725466
rect 42159 725008 42225 725011
rect 41568 725006 42225 725008
rect 41568 724950 42164 725006
rect 42220 724950 42225 725006
rect 41568 724948 42225 724950
rect 42159 724945 42225 724948
rect 41775 724416 41841 724419
rect 41568 724414 41841 724416
rect 41568 724358 41780 724414
rect 41836 724358 41841 724414
rect 41568 724356 41841 724358
rect 41775 724353 41841 724356
rect 34434 723827 34494 723942
rect 34434 723822 34545 723827
rect 34434 723766 34484 723822
rect 34540 723766 34545 723822
rect 34434 723764 34545 723766
rect 34479 723761 34545 723764
rect 42447 723528 42513 723531
rect 41568 723526 42513 723528
rect 41568 723470 42452 723526
rect 42508 723470 42513 723526
rect 41568 723468 42513 723470
rect 42447 723465 42513 723468
rect 41871 722936 41937 722939
rect 41568 722934 41937 722936
rect 41568 722878 41876 722934
rect 41932 722878 41937 722934
rect 41568 722876 41937 722878
rect 41871 722873 41937 722876
rect 41538 722344 41598 722462
rect 41679 722344 41745 722347
rect 41538 722342 41745 722344
rect 41538 722286 41684 722342
rect 41740 722286 41745 722342
rect 41538 722284 41745 722286
rect 41679 722281 41745 722284
rect 41538 721755 41598 721944
rect 41538 721750 41649 721755
rect 41538 721694 41588 721750
rect 41644 721694 41649 721750
rect 41538 721692 41649 721694
rect 41583 721689 41649 721692
rect 41914 721456 41920 721458
rect 41568 721396 41920 721456
rect 41914 721394 41920 721396
rect 41984 721394 41990 721458
rect 41722 721012 41728 721014
rect 41568 720952 41728 721012
rect 41722 720950 41728 720952
rect 41792 720950 41798 721014
rect 41538 720275 41598 720464
rect 41538 720270 41649 720275
rect 41538 720214 41588 720270
rect 41644 720214 41649 720270
rect 41538 720212 41649 720214
rect 41583 720209 41649 720212
rect 41538 719680 41598 719946
rect 41538 719620 41790 719680
rect 28866 719239 28926 719502
rect 28815 719234 28926 719239
rect 41730 719236 41790 719620
rect 28815 719178 28820 719234
rect 28876 719178 28926 719234
rect 28815 719176 28926 719178
rect 41538 719176 41790 719236
rect 28815 719173 28881 719176
rect 41538 718795 41598 719176
rect 28815 718792 28881 718795
rect 28815 718790 28926 718792
rect 28815 718734 28820 718790
rect 28876 718734 28926 718790
rect 28815 718729 28926 718734
rect 41538 718790 41649 718795
rect 41538 718734 41588 718790
rect 41644 718734 41649 718790
rect 41538 718732 41649 718734
rect 41583 718729 41649 718732
rect 28866 718466 28926 718729
rect 34383 716720 34449 716723
rect 40570 716720 40576 716722
rect 34383 716718 40576 716720
rect 34383 716662 34388 716718
rect 34444 716662 40576 716718
rect 34383 716660 40576 716662
rect 34383 716657 34449 716660
rect 40570 716658 40576 716660
rect 40640 716658 40646 716722
rect 34479 716128 34545 716131
rect 40378 716128 40384 716130
rect 34479 716126 40384 716128
rect 34479 716070 34484 716126
rect 34540 716070 40384 716126
rect 34479 716068 40384 716070
rect 34479 716065 34545 716068
rect 40378 716066 40384 716068
rect 40448 716066 40454 716130
rect 676290 715539 676350 715654
rect 676290 715534 676401 715539
rect 676290 715478 676340 715534
rect 676396 715478 676401 715534
rect 676290 715476 676401 715478
rect 676335 715473 676401 715476
rect 676143 714944 676209 714947
rect 676290 714944 676350 715136
rect 676143 714942 676350 714944
rect 676143 714886 676148 714942
rect 676204 714886 676350 714942
rect 676143 714884 676350 714886
rect 676143 714881 676209 714884
rect 676239 714796 676305 714799
rect 676239 714794 676350 714796
rect 676239 714738 676244 714794
rect 676300 714738 676350 714794
rect 676239 714733 676350 714738
rect 676290 714618 676350 714733
rect 41487 714204 41553 714207
rect 43066 714204 43072 714206
rect 41487 714202 43072 714204
rect 41487 714146 41492 714202
rect 41548 714146 43072 714202
rect 41487 714144 43072 714146
rect 41487 714141 41553 714144
rect 43066 714142 43072 714144
rect 43136 714142 43142 714206
rect 676047 714204 676113 714207
rect 676047 714202 676320 714204
rect 676047 714146 676052 714202
rect 676108 714146 676320 714202
rect 676047 714144 676320 714146
rect 676047 714141 676113 714144
rect 41967 714056 42033 714059
rect 42874 714056 42880 714058
rect 41967 714054 42880 714056
rect 41967 713998 41972 714054
rect 42028 713998 42880 714054
rect 41967 713996 42880 713998
rect 41967 713993 42033 713996
rect 42874 713994 42880 713996
rect 42944 713994 42950 714058
rect 42063 713910 42129 713911
rect 42063 713908 42112 713910
rect 42020 713906 42112 713908
rect 42020 713850 42068 713906
rect 42020 713848 42112 713850
rect 42063 713846 42112 713848
rect 42176 713846 42182 713910
rect 42063 713845 42129 713846
rect 676290 713467 676350 713582
rect 676239 713462 676350 713467
rect 676239 713406 676244 713462
rect 676300 713406 676350 713462
rect 676239 713404 676350 713406
rect 676239 713401 676305 713404
rect 676047 713168 676113 713171
rect 676047 713166 676320 713168
rect 676047 713110 676052 713166
rect 676108 713110 676320 713166
rect 676047 713108 676320 713110
rect 676047 713105 676113 713108
rect 676047 712724 676113 712727
rect 676047 712722 676320 712724
rect 676047 712666 676052 712722
rect 676108 712666 676320 712722
rect 676047 712664 676320 712666
rect 676047 712661 676113 712664
rect 42447 712282 42513 712283
rect 42447 712278 42496 712282
rect 42560 712280 42566 712282
rect 42447 712222 42452 712278
rect 42447 712218 42496 712222
rect 42560 712220 42604 712280
rect 42560 712218 42566 712220
rect 42447 712217 42513 712218
rect 676290 711987 676350 712102
rect 676239 711982 676350 711987
rect 676239 711926 676244 711982
rect 676300 711926 676350 711982
rect 676239 711924 676350 711926
rect 676239 711921 676305 711924
rect 42063 711690 42129 711691
rect 42063 711686 42112 711690
rect 42176 711688 42182 711690
rect 42063 711630 42068 711686
rect 42063 711626 42112 711630
rect 42176 711628 42220 711688
rect 42176 711626 42182 711628
rect 42682 711626 42688 711690
rect 42752 711688 42758 711690
rect 43023 711688 43089 711691
rect 42752 711686 43089 711688
rect 42752 711630 43028 711686
rect 43084 711630 43089 711686
rect 42752 711628 43089 711630
rect 42752 711626 42758 711628
rect 42063 711625 42129 711626
rect 43023 711625 43089 711628
rect 676047 711614 676113 711617
rect 676047 711612 676320 711614
rect 676047 711556 676052 711612
rect 676108 711556 676320 711612
rect 676047 711554 676320 711556
rect 676047 711551 676113 711554
rect 42298 711478 42304 711542
rect 42368 711540 42374 711542
rect 42927 711540 42993 711543
rect 42368 711538 42993 711540
rect 42368 711482 42932 711538
rect 42988 711482 42993 711538
rect 42368 711480 42993 711482
rect 42368 711478 42374 711480
rect 42927 711477 42993 711480
rect 43311 711392 43377 711395
rect 43695 711392 43761 711395
rect 43311 711390 43761 711392
rect 43311 711334 43316 711390
rect 43372 711334 43700 711390
rect 43756 711334 43761 711390
rect 43311 711332 43761 711334
rect 43311 711329 43377 711332
rect 43695 711329 43761 711332
rect 42682 711182 42688 711246
rect 42752 711244 42758 711246
rect 42927 711244 42993 711247
rect 42752 711242 42993 711244
rect 42752 711186 42932 711242
rect 42988 711186 42993 711242
rect 42752 711184 42993 711186
rect 42752 711182 42758 711184
rect 42927 711181 42993 711184
rect 676047 711244 676113 711247
rect 676047 711242 676320 711244
rect 676047 711186 676052 711242
rect 676108 711186 676320 711242
rect 676047 711184 676320 711186
rect 676047 711181 676113 711184
rect 42298 711034 42304 711098
rect 42368 711096 42374 711098
rect 43023 711096 43089 711099
rect 42368 711094 43089 711096
rect 42368 711038 43028 711094
rect 43084 711038 43089 711094
rect 42368 711036 43089 711038
rect 42368 711034 42374 711036
rect 43023 711033 43089 711036
rect 675898 710590 675904 710654
rect 675968 710652 675974 710654
rect 675968 710592 676320 710652
rect 675968 710590 675974 710592
rect 674746 710442 674752 710506
rect 674816 710504 674822 710506
rect 674816 710444 676350 710504
rect 674816 710442 674822 710444
rect 676290 710104 676350 710444
rect 675130 709702 675136 709766
rect 675200 709764 675206 709766
rect 675200 709704 676320 709764
rect 675200 709702 675206 709704
rect 675706 709110 675712 709174
rect 675776 709172 675782 709174
rect 675776 709112 676320 709172
rect 675776 709110 675782 709112
rect 41914 708814 41920 708878
rect 41984 708876 41990 708878
rect 42447 708876 42513 708879
rect 41984 708874 42513 708876
rect 41984 708818 42452 708874
rect 42508 708818 42513 708874
rect 41984 708816 42513 708818
rect 41984 708814 41990 708816
rect 42447 708813 42513 708816
rect 676047 708580 676113 708583
rect 676047 708578 676320 708580
rect 676047 708522 676052 708578
rect 676108 708522 676320 708578
rect 676047 708520 676320 708522
rect 676047 708517 676113 708520
rect 676047 708210 676113 708213
rect 676047 708208 676320 708210
rect 676047 708152 676052 708208
rect 676108 708152 676320 708208
rect 676047 708150 676320 708152
rect 676047 708147 676113 708150
rect 42927 707990 42993 707991
rect 42874 707926 42880 707990
rect 42944 707988 42993 707990
rect 42944 707986 43036 707988
rect 42988 707930 43036 707986
rect 42944 707928 43036 707930
rect 42944 707926 42993 707928
rect 42927 707925 42993 707926
rect 674362 707630 674368 707694
rect 674432 707692 674438 707694
rect 674432 707632 676320 707692
rect 674432 707630 674438 707632
rect 41775 707398 41841 707399
rect 41722 707396 41728 707398
rect 41684 707336 41728 707396
rect 41792 707394 41841 707398
rect 41836 707338 41841 707394
rect 41722 707334 41728 707336
rect 41792 707334 41841 707338
rect 41775 707333 41841 707334
rect 673978 707038 673984 707102
rect 674048 707100 674054 707102
rect 674048 707040 676320 707100
rect 674048 707038 674054 707040
rect 675322 706890 675328 706954
rect 675392 706952 675398 706954
rect 675392 706892 676350 706952
rect 675392 706890 675398 706892
rect 676290 706700 676350 706892
rect 677242 706446 677248 706510
rect 677312 706446 677318 706510
rect 677250 706182 677310 706446
rect 677050 705854 677056 705918
rect 677120 705854 677126 705918
rect 677058 705590 677118 705854
rect 676858 705410 676864 705474
rect 676928 705410 676934 705474
rect 40570 705114 40576 705178
rect 40640 705176 40646 705178
rect 42927 705176 42993 705179
rect 40640 705174 42993 705176
rect 40640 705118 42932 705174
rect 42988 705118 42993 705174
rect 676866 705146 676926 705410
rect 40640 705116 42993 705118
rect 40640 705114 40646 705116
rect 42927 705113 42993 705116
rect 42351 704880 42417 704883
rect 42490 704880 42496 704882
rect 42351 704878 42496 704880
rect 42351 704822 42356 704878
rect 42412 704822 42496 704878
rect 42351 704820 42496 704822
rect 42351 704817 42417 704820
rect 42490 704818 42496 704820
rect 42560 704818 42566 704882
rect 676239 704880 676305 704883
rect 676239 704878 676350 704880
rect 676239 704822 676244 704878
rect 676300 704822 676350 704878
rect 676239 704817 676350 704822
rect 676290 704702 676350 704817
rect 59631 704436 59697 704439
rect 679983 704436 680049 704439
rect 59631 704434 64638 704436
rect 59631 704378 59636 704434
rect 59692 704378 64638 704434
rect 59631 704376 64638 704378
rect 59631 704373 59697 704376
rect 64578 703860 64638 704376
rect 679938 704434 680049 704436
rect 679938 704378 679988 704434
rect 680044 704378 680049 704434
rect 679938 704373 680049 704378
rect 679938 704110 679998 704373
rect 43023 703550 43089 703551
rect 43023 703548 43072 703550
rect 42980 703546 43072 703548
rect 42980 703490 43028 703546
rect 42980 703488 43072 703490
rect 43023 703486 43072 703488
rect 43136 703486 43142 703550
rect 43023 703485 43089 703486
rect 679746 703403 679806 703666
rect 679746 703398 679857 703403
rect 679983 703400 680049 703403
rect 679746 703342 679796 703398
rect 679852 703342 679857 703398
rect 679746 703340 679857 703342
rect 679791 703337 679857 703340
rect 679938 703398 680049 703400
rect 679938 703342 679988 703398
rect 680044 703342 680049 703398
rect 679938 703337 680049 703342
rect 679938 703148 679998 703337
rect 679791 702956 679857 702959
rect 679746 702954 679857 702956
rect 679746 702898 679796 702954
rect 679852 702898 679857 702954
rect 679746 702893 679857 702898
rect 58767 702660 58833 702663
rect 64578 702660 64638 702678
rect 58767 702658 64638 702660
rect 58767 702602 58772 702658
rect 58828 702602 64638 702658
rect 679746 702630 679806 702893
rect 58767 702600 64638 702602
rect 58767 702597 58833 702600
rect 45231 702068 45297 702071
rect 45231 702066 64638 702068
rect 45231 702010 45236 702066
rect 45292 702010 64638 702066
rect 45231 702008 64638 702010
rect 45231 702005 45297 702008
rect 64578 701496 64638 702008
rect 58671 700884 58737 700887
rect 58671 700882 64638 700884
rect 58671 700826 58676 700882
rect 58732 700826 64638 700882
rect 58671 700824 64638 700826
rect 58671 700821 58737 700824
rect 64578 700314 64638 700824
rect 40378 699934 40384 699998
rect 40448 699996 40454 699998
rect 41775 699996 41841 699999
rect 40448 699994 41841 699996
rect 40448 699938 41780 699994
rect 41836 699938 41841 699994
rect 40448 699936 41841 699938
rect 40448 699934 40454 699936
rect 41775 699933 41841 699936
rect 59247 699700 59313 699703
rect 59247 699698 64638 699700
rect 59247 699642 59252 699698
rect 59308 699642 64638 699698
rect 59247 699640 64638 699642
rect 59247 699637 59313 699640
rect 64578 699132 64638 699640
rect 58863 698516 58929 698519
rect 58863 698514 64638 698516
rect 58863 698458 58868 698514
rect 58924 698458 64638 698514
rect 58863 698456 64638 698458
rect 58863 698453 58929 698456
rect 64578 697950 64638 698456
rect 675130 697862 675136 697926
rect 675200 697924 675206 697926
rect 675375 697924 675441 697927
rect 675200 697922 675441 697924
rect 675200 697866 675380 697922
rect 675436 697866 675441 697922
rect 675200 697864 675441 697866
rect 675200 697862 675206 697864
rect 675375 697861 675441 697864
rect 674362 697122 674368 697186
rect 674432 697184 674438 697186
rect 675183 697184 675249 697187
rect 674432 697182 675249 697184
rect 674432 697126 675188 697182
rect 675244 697126 675249 697182
rect 674432 697124 675249 697126
rect 674432 697122 674438 697124
rect 675183 697121 675249 697124
rect 674746 696974 674752 697038
rect 674816 697036 674822 697038
rect 675183 697036 675249 697039
rect 674816 697034 675249 697036
rect 674816 696978 675188 697034
rect 675244 696978 675249 697034
rect 674816 696976 675249 696978
rect 674816 696974 674822 696976
rect 675183 696973 675249 696976
rect 675663 694966 675729 694967
rect 675663 694962 675712 694966
rect 675776 694964 675782 694966
rect 675663 694906 675668 694962
rect 675663 694902 675712 694906
rect 675776 694904 675820 694964
rect 675776 694902 675782 694904
rect 675663 694901 675729 694902
rect 675279 694670 675345 694671
rect 675279 694666 675328 694670
rect 675392 694668 675398 694670
rect 675279 694610 675284 694666
rect 675279 694606 675328 694610
rect 675392 694608 675436 694668
rect 675392 694606 675398 694608
rect 675279 694605 675345 694606
rect 649986 689488 650046 689980
rect 655215 689488 655281 689491
rect 649986 689486 655281 689488
rect 649986 689430 655220 689486
rect 655276 689430 655281 689486
rect 649986 689428 655281 689430
rect 655215 689425 655281 689428
rect 649986 688452 650046 688798
rect 655407 688452 655473 688455
rect 649986 688450 655473 688452
rect 649986 688394 655412 688450
rect 655468 688394 655473 688450
rect 649986 688392 655473 688394
rect 655407 688389 655473 688392
rect 41775 688304 41841 688307
rect 41568 688302 41841 688304
rect 41568 688246 41780 688302
rect 41836 688246 41841 688302
rect 41568 688244 41841 688246
rect 41775 688241 41841 688244
rect 41538 687567 41598 687682
rect 41538 687562 41649 687567
rect 41538 687506 41588 687562
rect 41644 687506 41649 687562
rect 41538 687504 41649 687506
rect 41583 687501 41649 687504
rect 41775 687268 41841 687271
rect 41568 687266 41841 687268
rect 41568 687210 41780 687266
rect 41836 687210 41841 687266
rect 41568 687208 41841 687210
rect 41775 687205 41841 687208
rect 649986 687120 650046 687616
rect 655599 687120 655665 687123
rect 649986 687118 655665 687120
rect 649986 687062 655604 687118
rect 655660 687062 655665 687118
rect 649986 687060 655665 687062
rect 655599 687057 655665 687060
rect 41583 686972 41649 686975
rect 653775 686972 653841 686975
rect 41538 686970 41649 686972
rect 41538 686914 41588 686970
rect 41644 686914 41649 686970
rect 41538 686909 41649 686914
rect 649986 686970 653841 686972
rect 649986 686914 653780 686970
rect 653836 686914 653841 686970
rect 649986 686912 653841 686914
rect 41538 686794 41598 686909
rect 649986 686434 650046 686912
rect 653775 686909 653841 686912
rect 41538 686087 41598 686202
rect 41538 686082 41649 686087
rect 41538 686026 41588 686082
rect 41644 686026 41649 686082
rect 41538 686024 41649 686026
rect 41583 686021 41649 686024
rect 40386 685494 40446 685684
rect 40378 685430 40384 685494
rect 40448 685430 40454 685494
rect 41775 685344 41841 685347
rect 654159 685344 654225 685347
rect 41568 685342 41841 685344
rect 41568 685286 41780 685342
rect 41836 685286 41841 685342
rect 41568 685284 41841 685286
rect 41775 685281 41841 685284
rect 649986 685342 654225 685344
rect 649986 685286 654164 685342
rect 654220 685286 654225 685342
rect 649986 685284 654225 685286
rect 649986 685252 650046 685284
rect 654159 685281 654225 685284
rect 40578 684458 40638 684722
rect 654063 684604 654129 684607
rect 649986 684602 654129 684604
rect 649986 684546 654068 684602
rect 654124 684546 654129 684602
rect 649986 684544 654129 684546
rect 40570 684394 40576 684458
rect 40640 684394 40646 684458
rect 41775 684160 41841 684163
rect 41568 684158 41841 684160
rect 41568 684102 41780 684158
rect 41836 684102 41841 684158
rect 41568 684100 41841 684102
rect 41775 684097 41841 684100
rect 649986 684070 650046 684544
rect 654063 684541 654129 684544
rect 41967 683864 42033 683867
rect 41568 683862 42033 683864
rect 41568 683806 41972 683862
rect 42028 683806 42033 683862
rect 41568 683804 42033 683806
rect 41967 683801 42033 683804
rect 41775 683272 41841 683275
rect 41568 683270 41841 683272
rect 41568 683214 41780 683270
rect 41836 683214 41841 683270
rect 41568 683212 41841 683214
rect 41775 683209 41841 683212
rect 34434 682535 34494 682650
rect 34383 682530 34494 682535
rect 34383 682474 34388 682530
rect 34444 682474 34494 682530
rect 34383 682472 34494 682474
rect 34383 682469 34449 682472
rect 37314 682091 37374 682280
rect 37314 682086 37425 682091
rect 37314 682030 37364 682086
rect 37420 682030 37425 682086
rect 37314 682028 37425 682030
rect 37359 682025 37425 682028
rect 41871 681792 41937 681795
rect 41568 681790 41937 681792
rect 41568 681734 41876 681790
rect 41932 681734 41937 681790
rect 41568 681732 41937 681734
rect 41871 681729 41937 681732
rect 41775 681200 41841 681203
rect 41568 681198 41841 681200
rect 41568 681142 41780 681198
rect 41836 681142 41841 681198
rect 41568 681140 41841 681142
rect 41775 681137 41841 681140
rect 39810 680611 39870 680800
rect 39759 680606 39870 680611
rect 39759 680550 39764 680606
rect 39820 680550 39870 680606
rect 39759 680548 39870 680550
rect 39759 680545 39825 680548
rect 39810 680019 39870 680282
rect 39810 680014 39921 680019
rect 39810 679958 39860 680014
rect 39916 679958 39921 680014
rect 39810 679956 39921 679958
rect 39855 679953 39921 679956
rect 34434 679575 34494 679710
rect 34434 679570 34545 679575
rect 34434 679514 34484 679570
rect 34540 679514 34545 679570
rect 34434 679512 34545 679514
rect 34479 679509 34545 679512
rect 41538 679131 41598 679246
rect 41538 679126 41649 679131
rect 41538 679070 41588 679126
rect 41644 679070 41649 679126
rect 41538 679068 41649 679070
rect 41583 679065 41649 679068
rect 42063 678832 42129 678835
rect 41568 678830 42129 678832
rect 41568 678774 42068 678830
rect 42124 678774 42129 678830
rect 41568 678772 42129 678774
rect 42063 678769 42129 678772
rect 42255 678240 42321 678243
rect 41568 678238 42321 678240
rect 41568 678182 42260 678238
rect 42316 678182 42321 678238
rect 41568 678180 42321 678182
rect 42255 678177 42321 678180
rect 41538 677648 41598 677766
rect 41679 677648 41745 677651
rect 41538 677646 41745 677648
rect 41538 677590 41684 677646
rect 41740 677590 41745 677646
rect 41538 677588 41745 677590
rect 41679 677585 41745 677588
rect 41538 677059 41598 677248
rect 41538 677054 41649 677059
rect 41538 676998 41588 677054
rect 41644 676998 41649 677054
rect 41538 676996 41649 676998
rect 41583 676993 41649 676996
rect 41568 676700 41790 676760
rect 28866 676023 28926 676286
rect 41730 676168 41790 676700
rect 28815 676018 28926 676023
rect 28815 675962 28820 676018
rect 28876 675962 28926 676018
rect 28815 675960 28926 675962
rect 41538 676108 41790 676168
rect 28815 675957 28881 675960
rect 41538 675579 41598 676108
rect 28815 675576 28881 675579
rect 28815 675574 28926 675576
rect 28815 675518 28820 675574
rect 28876 675518 28926 675574
rect 28815 675513 28926 675518
rect 41538 675574 41649 675579
rect 41538 675518 41588 675574
rect 41644 675518 41649 675574
rect 41538 675516 41649 675518
rect 41583 675513 41649 675516
rect 28866 675250 28926 675513
rect 34383 672468 34449 672471
rect 40570 672468 40576 672470
rect 34383 672466 40576 672468
rect 34383 672410 34388 672466
rect 34444 672410 40576 672466
rect 34383 672408 40576 672410
rect 34383 672405 34449 672408
rect 40570 672406 40576 672408
rect 40640 672406 40646 672470
rect 39759 671136 39825 671139
rect 41146 671136 41152 671138
rect 39759 671134 41152 671136
rect 39759 671078 39764 671134
rect 39820 671078 41152 671134
rect 39759 671076 41152 671078
rect 39759 671073 39825 671076
rect 41146 671074 41152 671076
rect 41216 671074 41222 671138
rect 41967 670692 42033 670695
rect 42298 670692 42304 670694
rect 41967 670690 42304 670692
rect 41967 670634 41972 670690
rect 42028 670634 42304 670690
rect 41967 670632 42304 670634
rect 41967 670629 42033 670632
rect 42298 670630 42304 670632
rect 42368 670630 42374 670694
rect 676143 670396 676209 670399
rect 676290 670396 676350 670662
rect 676143 670394 676350 670396
rect 676143 670338 676148 670394
rect 676204 670338 676350 670394
rect 676143 670336 676350 670338
rect 676143 670333 676209 670336
rect 676290 669807 676350 670070
rect 676290 669802 676401 669807
rect 676290 669746 676340 669802
rect 676396 669746 676401 669802
rect 676290 669744 676401 669746
rect 676335 669741 676401 669744
rect 676290 669363 676350 669626
rect 676239 669358 676350 669363
rect 676239 669302 676244 669358
rect 676300 669302 676350 669358
rect 676239 669300 676350 669302
rect 676239 669297 676305 669300
rect 676047 669212 676113 669215
rect 676047 669210 676320 669212
rect 676047 669154 676052 669210
rect 676108 669154 676320 669210
rect 676047 669152 676320 669154
rect 676047 669149 676113 669152
rect 676047 668620 676113 668623
rect 676047 668618 676320 668620
rect 676047 668562 676052 668618
rect 676108 668562 676320 668618
rect 676047 668560 676320 668562
rect 676047 668557 676113 668560
rect 675951 668102 676017 668105
rect 675951 668100 676320 668102
rect 675951 668044 675956 668100
rect 676012 668044 676320 668100
rect 675951 668042 676320 668044
rect 675951 668039 676017 668042
rect 675951 667732 676017 667735
rect 675951 667730 676320 667732
rect 675951 667674 675956 667730
rect 676012 667674 676320 667730
rect 675951 667672 676320 667674
rect 675951 667669 676017 667672
rect 676290 666995 676350 667110
rect 676239 666990 676350 666995
rect 676239 666934 676244 666990
rect 676300 666934 676350 666990
rect 676239 666932 676350 666934
rect 676239 666929 676305 666932
rect 676290 666403 676350 666592
rect 676239 666398 676350 666403
rect 676239 666342 676244 666398
rect 676300 666342 676350 666398
rect 676239 666340 676350 666342
rect 676239 666337 676305 666340
rect 674938 666190 674944 666254
rect 675008 666252 675014 666254
rect 675008 666192 676320 666252
rect 675008 666190 675014 666192
rect 676047 665660 676113 665663
rect 676047 665658 676320 665660
rect 676047 665602 676052 665658
rect 676108 665602 676320 665658
rect 676047 665600 676320 665602
rect 676047 665597 676113 665600
rect 42298 665006 42304 665070
rect 42368 665068 42374 665070
rect 42735 665068 42801 665071
rect 42368 665066 42801 665068
rect 42368 665010 42740 665066
rect 42796 665010 42801 665066
rect 42368 665008 42801 665010
rect 42368 665006 42374 665008
rect 42735 665005 42801 665008
rect 676090 664858 676096 664922
rect 676160 664920 676166 664922
rect 676290 664920 676350 665038
rect 676160 664860 676350 664920
rect 676160 664858 676166 664860
rect 674554 664710 674560 664774
rect 674624 664772 674630 664774
rect 674624 664712 676320 664772
rect 674624 664710 674630 664712
rect 676282 664414 676288 664478
rect 676352 664414 676358 664478
rect 676290 664150 676350 664414
rect 676047 663588 676113 663591
rect 676047 663586 676320 663588
rect 676047 663530 676052 663586
rect 676108 663530 676320 663586
rect 676047 663528 676320 663530
rect 676047 663525 676113 663528
rect 674170 663378 674176 663442
rect 674240 663440 674246 663442
rect 674240 663380 676350 663440
rect 674240 663378 674246 663380
rect 676290 663188 676350 663380
rect 675514 662638 675520 662702
rect 675584 662700 675590 662702
rect 675584 662640 676320 662700
rect 675584 662638 675590 662640
rect 41146 662342 41152 662406
rect 41216 662404 41222 662406
rect 42831 662404 42897 662407
rect 41216 662402 42897 662404
rect 41216 662346 42836 662402
rect 42892 662346 42897 662402
rect 41216 662344 42897 662346
rect 41216 662342 41222 662344
rect 42831 662341 42897 662344
rect 676047 662108 676113 662111
rect 676047 662106 676320 662108
rect 676047 662050 676052 662106
rect 676108 662050 676320 662106
rect 676047 662048 676320 662050
rect 676047 662045 676113 662048
rect 676047 661664 676113 661667
rect 676047 661662 676320 661664
rect 676047 661606 676052 661662
rect 676108 661606 676320 661662
rect 676047 661604 676320 661606
rect 676047 661601 676113 661604
rect 676239 661368 676305 661371
rect 676239 661366 676350 661368
rect 676239 661310 676244 661366
rect 676300 661310 676350 661366
rect 676239 661305 676350 661310
rect 59631 661220 59697 661223
rect 59631 661218 64638 661220
rect 59631 661162 59636 661218
rect 59692 661162 64638 661218
rect 676290 661190 676350 661305
rect 59631 661160 64638 661162
rect 59631 661157 59697 661160
rect 40570 660714 40576 660778
rect 40640 660776 40646 660778
rect 42927 660776 42993 660779
rect 40640 660774 42993 660776
rect 40640 660718 42932 660774
rect 42988 660718 42993 660774
rect 40640 660716 42993 660718
rect 40640 660714 40646 660716
rect 42927 660713 42993 660716
rect 64578 660638 64638 661160
rect 676047 660628 676113 660631
rect 676047 660626 676320 660628
rect 676047 660570 676052 660626
rect 676108 660570 676320 660626
rect 676047 660568 676320 660570
rect 676047 660565 676113 660568
rect 676047 660184 676113 660187
rect 676047 660182 676320 660184
rect 676047 660126 676052 660182
rect 676108 660126 676320 660182
rect 676047 660124 676320 660126
rect 676047 660121 676113 660124
rect 676239 659888 676305 659891
rect 676239 659886 676350 659888
rect 676239 659830 676244 659886
rect 676300 659830 676350 659886
rect 676239 659825 676350 659830
rect 676290 659710 676350 659825
rect 58767 659444 58833 659447
rect 64578 659444 64638 659456
rect 58767 659442 64638 659444
rect 58767 659386 58772 659442
rect 58828 659386 64638 659442
rect 58767 659384 64638 659386
rect 58767 659381 58833 659384
rect 679791 659296 679857 659299
rect 679746 659294 679857 659296
rect 679746 659238 679796 659294
rect 679852 659238 679857 659294
rect 679746 659233 679857 659238
rect 679746 659118 679806 659233
rect 43023 658852 43089 658855
rect 43023 658850 64638 658852
rect 43023 658794 43028 658850
rect 43084 658794 64638 658850
rect 43023 658792 64638 658794
rect 43023 658789 43089 658792
rect 64578 658274 64638 658792
rect 685506 658411 685566 658674
rect 679791 658408 679857 658411
rect 679746 658406 679857 658408
rect 679746 658350 679796 658406
rect 679852 658350 679857 658406
rect 679746 658345 679857 658350
rect 685455 658406 685566 658411
rect 685455 658350 685460 658406
rect 685516 658350 685566 658406
rect 685455 658348 685566 658350
rect 685455 658345 685521 658348
rect 679746 658156 679806 658345
rect 685455 657964 685521 657967
rect 685455 657962 685566 657964
rect 685455 657906 685460 657962
rect 685516 657906 685566 657962
rect 685455 657901 685566 657906
rect 58671 657668 58737 657671
rect 58671 657666 64638 657668
rect 58671 657610 58676 657666
rect 58732 657610 64638 657666
rect 685506 657638 685566 657901
rect 58671 657608 64638 657610
rect 58671 657605 58737 657608
rect 64578 657092 64638 657608
rect 58191 656484 58257 656487
rect 58191 656482 64638 656484
rect 58191 656426 58196 656482
rect 58252 656426 64638 656482
rect 58191 656424 64638 656426
rect 58191 656421 58257 656424
rect 64578 655910 64638 656424
rect 58383 655300 58449 655303
rect 58383 655298 64638 655300
rect 58383 655242 58388 655298
rect 58444 655242 64638 655298
rect 58383 655240 64638 655242
rect 58383 655237 58449 655240
rect 64578 654728 64638 655240
rect 673978 652722 673984 652786
rect 674048 652784 674054 652786
rect 675375 652784 675441 652787
rect 674048 652782 675441 652784
rect 674048 652726 675380 652782
rect 675436 652726 675441 652782
rect 674048 652724 675441 652726
rect 674048 652722 674054 652724
rect 675375 652721 675441 652724
rect 674170 652130 674176 652194
rect 674240 652192 674246 652194
rect 675471 652192 675537 652195
rect 674240 652190 675537 652192
rect 674240 652134 675476 652190
rect 675532 652134 675537 652190
rect 674240 652132 675537 652134
rect 674240 652130 674246 652132
rect 675471 652129 675537 652132
rect 674938 651390 674944 651454
rect 675008 651452 675014 651454
rect 675375 651452 675441 651455
rect 675008 651450 675441 651452
rect 675008 651394 675380 651450
rect 675436 651394 675441 651450
rect 675008 651392 675441 651394
rect 675008 651390 675014 651392
rect 675375 651389 675441 651392
rect 674554 649614 674560 649678
rect 674624 649676 674630 649678
rect 675375 649676 675441 649679
rect 674624 649674 675441 649676
rect 674624 649618 675380 649674
rect 675436 649618 675441 649674
rect 674624 649616 675441 649618
rect 674624 649614 674630 649616
rect 675375 649613 675441 649616
rect 675471 645386 675537 645387
rect 675471 645382 675520 645386
rect 675584 645384 675590 645386
rect 675471 645326 675476 645382
rect 675471 645322 675520 645326
rect 675584 645324 675628 645384
rect 675584 645322 675590 645324
rect 675471 645321 675537 645322
rect 41538 644943 41598 645058
rect 41538 644938 41649 644943
rect 41538 644882 41588 644938
rect 41644 644882 41649 644938
rect 41538 644880 41649 644882
rect 41583 644877 41649 644880
rect 40762 644730 40768 644794
rect 40832 644792 40838 644794
rect 41487 644792 41553 644795
rect 40832 644790 41553 644792
rect 40832 644734 41492 644790
rect 41548 644734 41553 644790
rect 40832 644732 41553 644734
rect 40832 644730 40838 644732
rect 41487 644729 41553 644732
rect 41538 644351 41598 644466
rect 41538 644346 41649 644351
rect 41538 644290 41588 644346
rect 41644 644290 41649 644346
rect 41538 644288 41649 644290
rect 41583 644285 41649 644288
rect 41775 644052 41841 644055
rect 41568 644050 41841 644052
rect 41568 643994 41780 644050
rect 41836 643994 41841 644050
rect 41568 643992 41841 643994
rect 41775 643989 41841 643992
rect 41583 643756 41649 643759
rect 41538 643754 41649 643756
rect 41538 643698 41588 643754
rect 41644 643698 41649 643754
rect 41538 643693 41649 643698
rect 41538 643578 41598 643693
rect 649986 643016 650046 643558
rect 655311 643016 655377 643019
rect 649986 643014 655377 643016
rect 41538 642871 41598 642986
rect 649986 642958 655316 643014
rect 655372 642958 655377 643014
rect 649986 642956 655377 642958
rect 655311 642953 655377 642956
rect 41538 642866 41649 642871
rect 41538 642810 41588 642866
rect 41644 642810 41649 642866
rect 41538 642808 41649 642810
rect 41583 642805 41649 642808
rect 40386 642278 40446 642542
rect 655119 642424 655185 642427
rect 649986 642422 655185 642424
rect 649986 642366 655124 642422
rect 655180 642366 655185 642422
rect 649986 642364 655185 642366
rect 655119 642361 655185 642364
rect 40378 642214 40384 642278
rect 40448 642214 40454 642278
rect 40570 642214 40576 642278
rect 40640 642276 40646 642278
rect 42874 642276 42880 642278
rect 40640 642216 42880 642276
rect 40640 642214 40646 642216
rect 42874 642214 42880 642216
rect 42944 642214 42950 642278
rect 40578 642098 40638 642214
rect 41538 641391 41598 641506
rect 41538 641386 41649 641391
rect 41538 641330 41588 641386
rect 41644 641330 41649 641386
rect 41538 641328 41649 641330
rect 41583 641325 41649 641328
rect 41487 641240 41553 641243
rect 41487 641238 41598 641240
rect 41487 641182 41492 641238
rect 41548 641182 41598 641238
rect 41487 641177 41598 641182
rect 41538 640988 41598 641177
rect 649986 640796 650046 641194
rect 655503 640796 655569 640799
rect 649986 640794 655569 640796
rect 649986 640738 655508 640794
rect 655564 640738 655569 640794
rect 649986 640736 655569 640738
rect 655503 640733 655569 640736
rect 654159 640648 654225 640651
rect 649986 640646 654225 640648
rect 37314 640355 37374 640618
rect 649986 640590 654164 640646
rect 654220 640590 654225 640646
rect 649986 640588 654225 640590
rect 37314 640350 37425 640355
rect 37314 640294 37364 640350
rect 37420 640294 37425 640350
rect 37314 640292 37425 640294
rect 37359 640289 37425 640292
rect 41967 640056 42033 640059
rect 41568 640054 42033 640056
rect 41568 639998 41972 640054
rect 42028 639998 42033 640054
rect 649986 640012 650046 640588
rect 654159 640585 654225 640588
rect 675759 640352 675825 640355
rect 676090 640352 676096 640354
rect 675759 640350 676096 640352
rect 675759 640294 675764 640350
rect 675820 640294 676096 640350
rect 675759 640292 676096 640294
rect 675759 640289 675825 640292
rect 676090 640290 676096 640292
rect 676160 640290 676166 640354
rect 41568 639996 42033 639998
rect 41967 639993 42033 639996
rect 34434 639319 34494 639434
rect 34434 639314 34545 639319
rect 34434 639258 34484 639314
rect 34540 639258 34545 639314
rect 34434 639256 34545 639258
rect 34479 639253 34545 639256
rect 655791 639168 655857 639171
rect 649986 639166 655857 639168
rect 40194 638875 40254 639138
rect 40143 638870 40254 638875
rect 40143 638814 40148 638870
rect 40204 638814 40254 638870
rect 649986 639110 655796 639166
rect 655852 639110 655857 639166
rect 649986 639108 655857 639110
rect 649986 638830 650046 639108
rect 655791 639105 655857 639108
rect 40143 638812 40254 638814
rect 40143 638809 40209 638812
rect 41679 638724 41745 638727
rect 41538 638722 41745 638724
rect 41538 638666 41684 638722
rect 41740 638666 41745 638722
rect 41538 638664 41745 638666
rect 41538 638546 41598 638664
rect 41679 638661 41745 638664
rect 675759 638576 675825 638579
rect 675898 638576 675904 638578
rect 675759 638574 675904 638576
rect 675759 638518 675764 638574
rect 675820 638518 675904 638574
rect 675759 638516 675904 638518
rect 675759 638513 675825 638516
rect 675898 638514 675904 638516
rect 675968 638514 675974 638578
rect 655983 638280 656049 638283
rect 649986 638278 656049 638280
rect 649986 638222 655988 638278
rect 656044 638222 656049 638278
rect 649986 638220 656049 638222
rect 41871 637984 41937 637987
rect 41568 637982 41937 637984
rect 41568 637926 41876 637982
rect 41932 637926 41937 637982
rect 41568 637924 41937 637926
rect 41871 637921 41937 637924
rect 649986 637648 650046 638220
rect 655983 638217 656049 638220
rect 40194 637395 40254 637584
rect 40194 637390 40305 637395
rect 40194 637334 40244 637390
rect 40300 637334 40305 637390
rect 40194 637332 40305 637334
rect 40239 637329 40305 637332
rect 34434 636803 34494 637066
rect 34383 636798 34494 636803
rect 34383 636742 34388 636798
rect 34444 636742 34494 636798
rect 34383 636740 34494 636742
rect 34383 636737 34449 636740
rect 42159 636504 42225 636507
rect 41568 636502 42225 636504
rect 41568 636446 42164 636502
rect 42220 636446 42225 636502
rect 41568 636444 42225 636446
rect 42159 636441 42225 636444
rect 41775 636134 41841 636137
rect 41568 636132 41841 636134
rect 41568 636076 41780 636132
rect 41836 636076 41841 636132
rect 41568 636074 41841 636076
rect 41775 636071 41841 636074
rect 41538 635323 41598 635586
rect 41538 635318 41649 635323
rect 41538 635262 41588 635318
rect 41644 635262 41649 635318
rect 41538 635260 41649 635262
rect 41583 635257 41649 635260
rect 42255 635024 42321 635027
rect 41568 635022 42321 635024
rect 41568 634966 42260 635022
rect 42316 634966 42321 635022
rect 41568 634964 42321 634966
rect 42255 634961 42321 634964
rect 41538 634435 41598 634550
rect 41538 634430 41649 634435
rect 41538 634374 41588 634430
rect 41644 634374 41649 634430
rect 41538 634372 41649 634374
rect 41583 634369 41649 634372
rect 41775 634136 41841 634139
rect 41568 634134 41841 634136
rect 41568 634078 41780 634134
rect 41836 634078 41841 634134
rect 41568 634076 41841 634078
rect 41775 634073 41841 634076
rect 41568 633484 41790 633544
rect 28866 632807 28926 633070
rect 41730 632952 41790 633484
rect 28815 632802 28926 632807
rect 28815 632746 28820 632802
rect 28876 632746 28926 632802
rect 28815 632744 28926 632746
rect 41538 632892 41790 632952
rect 28815 632741 28881 632744
rect 41538 632363 41598 632892
rect 28815 632360 28881 632363
rect 28815 632358 28926 632360
rect 28815 632302 28820 632358
rect 28876 632302 28926 632358
rect 28815 632297 28926 632302
rect 41538 632358 41649 632363
rect 41538 632302 41588 632358
rect 41644 632302 41649 632358
rect 41538 632300 41649 632302
rect 41583 632297 41649 632300
rect 28866 632034 28926 632297
rect 34479 629252 34545 629255
rect 40762 629252 40768 629254
rect 34479 629250 40768 629252
rect 34479 629194 34484 629250
rect 34540 629194 40768 629250
rect 34479 629192 40768 629194
rect 34479 629189 34545 629192
rect 40762 629190 40768 629192
rect 40832 629190 40838 629254
rect 40239 628364 40305 628367
rect 40570 628364 40576 628366
rect 40239 628362 40576 628364
rect 40239 628306 40244 628362
rect 40300 628306 40576 628362
rect 40239 628304 40576 628306
rect 40239 628301 40305 628304
rect 40570 628302 40576 628304
rect 40640 628302 40646 628366
rect 42063 627624 42129 627627
rect 43066 627624 43072 627626
rect 42063 627622 43072 627624
rect 42063 627566 42068 627622
rect 42124 627566 43072 627622
rect 42063 627564 43072 627566
rect 42063 627561 42129 627564
rect 43066 627562 43072 627564
rect 43136 627562 43142 627626
rect 41775 627476 41841 627479
rect 41914 627476 41920 627478
rect 41775 627474 41920 627476
rect 41775 627418 41780 627474
rect 41836 627418 41920 627474
rect 41775 627416 41920 627418
rect 41775 627413 41841 627416
rect 41914 627414 41920 627416
rect 41984 627414 41990 627478
rect 42159 627476 42225 627479
rect 42298 627476 42304 627478
rect 42159 627474 42304 627476
rect 42159 627418 42164 627474
rect 42220 627418 42304 627474
rect 42159 627416 42304 627418
rect 42159 627413 42225 627416
rect 42298 627414 42304 627416
rect 42368 627414 42374 627478
rect 41914 625194 41920 625258
rect 41984 625256 41990 625258
rect 42735 625256 42801 625259
rect 41984 625254 42801 625256
rect 41984 625198 42740 625254
rect 42796 625198 42801 625254
rect 41984 625196 42801 625198
rect 41984 625194 41990 625196
rect 42735 625193 42801 625196
rect 676290 625111 676350 625522
rect 676239 625106 676350 625111
rect 676239 625050 676244 625106
rect 676300 625050 676350 625106
rect 676239 625048 676350 625050
rect 676239 625045 676305 625048
rect 676143 624664 676209 624667
rect 676290 624664 676350 624930
rect 676143 624662 676350 624664
rect 676143 624606 676148 624662
rect 676204 624606 676350 624662
rect 676143 624604 676350 624606
rect 676143 624601 676209 624604
rect 676290 624223 676350 624338
rect 676239 624218 676350 624223
rect 676239 624162 676244 624218
rect 676300 624162 676350 624218
rect 676239 624160 676350 624162
rect 676239 624157 676305 624160
rect 676047 623998 676113 624001
rect 676047 623996 676320 623998
rect 676047 623940 676052 623996
rect 676108 623940 676320 623996
rect 676047 623938 676320 623940
rect 676047 623935 676113 623938
rect 676047 623480 676113 623483
rect 676047 623478 676320 623480
rect 676047 623422 676052 623478
rect 676108 623422 676320 623478
rect 676047 623420 676320 623422
rect 676047 623417 676113 623420
rect 676047 622888 676113 622891
rect 676047 622886 676320 622888
rect 676047 622830 676052 622886
rect 676108 622830 676320 622886
rect 676047 622828 676320 622830
rect 676047 622825 676113 622828
rect 676047 622518 676113 622521
rect 676047 622516 676320 622518
rect 676047 622460 676052 622516
rect 676108 622460 676320 622516
rect 676047 622458 676320 622460
rect 676047 622455 676113 622458
rect 42298 622086 42304 622150
rect 42368 622148 42374 622150
rect 42831 622148 42897 622151
rect 42368 622146 42897 622148
rect 42368 622090 42836 622146
rect 42892 622090 42897 622146
rect 42368 622088 42897 622090
rect 42368 622086 42374 622088
rect 42831 622085 42897 622088
rect 676047 622000 676113 622003
rect 676047 621998 676320 622000
rect 676047 621942 676052 621998
rect 676108 621942 676320 621998
rect 676047 621940 676320 621942
rect 676047 621937 676113 621940
rect 676047 621408 676113 621411
rect 676047 621406 676320 621408
rect 676047 621350 676052 621406
rect 676108 621350 676320 621406
rect 676047 621348 676320 621350
rect 676047 621345 676113 621348
rect 674746 620902 674752 620966
rect 674816 620964 674822 620966
rect 674816 620904 676320 620964
rect 674816 620902 674822 620904
rect 676239 620668 676305 620671
rect 676239 620666 676350 620668
rect 676239 620610 676244 620666
rect 676300 620610 676350 620666
rect 676239 620605 676350 620610
rect 676290 620490 676350 620605
rect 675130 619866 675136 619930
rect 675200 619928 675206 619930
rect 675200 619868 676320 619928
rect 675200 619866 675206 619868
rect 675706 619422 675712 619486
rect 675776 619484 675782 619486
rect 675776 619424 676320 619484
rect 675776 619422 675782 619424
rect 42831 619188 42897 619191
rect 43066 619188 43072 619190
rect 42831 619186 43072 619188
rect 42831 619130 42836 619186
rect 42892 619130 43072 619186
rect 42831 619128 43072 619130
rect 42831 619125 42897 619128
rect 43066 619126 43072 619128
rect 43136 619126 43142 619190
rect 676047 618966 676113 618969
rect 676047 618964 676320 618966
rect 676047 618908 676052 618964
rect 676108 618908 676320 618964
rect 676047 618906 676320 618908
rect 676047 618903 676113 618906
rect 676239 618596 676305 618599
rect 676239 618594 676350 618596
rect 676239 618538 676244 618594
rect 676300 618538 676350 618594
rect 676239 618533 676350 618538
rect 676290 618418 676350 618533
rect 58959 618004 59025 618007
rect 58959 618002 64638 618004
rect 58959 617946 58964 618002
rect 59020 617946 64638 618002
rect 58959 617944 64638 617946
rect 58959 617941 59025 617944
rect 64578 617416 64638 617944
rect 674362 617942 674368 618006
rect 674432 618004 674438 618006
rect 674432 617944 676320 618004
rect 674432 617942 674438 617944
rect 675322 617794 675328 617858
rect 675392 617856 675398 617858
rect 675392 617796 676350 617856
rect 675392 617794 675398 617796
rect 676290 617456 676350 617796
rect 676239 617116 676305 617119
rect 676239 617114 676350 617116
rect 676239 617058 676244 617114
rect 676300 617058 676350 617114
rect 676239 617053 676350 617058
rect 676290 616938 676350 617053
rect 40570 616462 40576 616526
rect 40640 616524 40646 616526
rect 42735 616524 42801 616527
rect 40640 616522 42801 616524
rect 40640 616466 42740 616522
rect 42796 616466 42801 616522
rect 40640 616464 42801 616466
rect 40640 616462 40646 616464
rect 42735 616461 42801 616464
rect 676047 616524 676113 616527
rect 676047 616522 676320 616524
rect 676047 616466 676052 616522
rect 676108 616466 676320 616522
rect 676047 616464 676320 616466
rect 676047 616461 676113 616464
rect 40762 616314 40768 616378
rect 40832 616376 40838 616378
rect 42351 616376 42417 616379
rect 40832 616374 42417 616376
rect 40832 616318 42356 616374
rect 42412 616318 42417 616374
rect 40832 616316 42417 616318
rect 40832 616314 40838 616316
rect 42351 616313 42417 616316
rect 59631 616228 59697 616231
rect 64578 616228 64638 616234
rect 59631 616226 64638 616228
rect 59631 616170 59636 616226
rect 59692 616170 64638 616226
rect 59631 616168 64638 616170
rect 59631 616165 59697 616168
rect 676047 615932 676113 615935
rect 676047 615930 676320 615932
rect 676047 615874 676052 615930
rect 676108 615874 676320 615930
rect 676047 615872 676320 615874
rect 676047 615869 676113 615872
rect 58191 615636 58257 615639
rect 676239 615636 676305 615639
rect 58191 615634 64638 615636
rect 58191 615578 58196 615634
rect 58252 615578 64638 615634
rect 58191 615576 64638 615578
rect 58191 615573 58257 615576
rect 64578 615052 64638 615576
rect 676239 615634 676350 615636
rect 676239 615578 676244 615634
rect 676300 615578 676350 615634
rect 676239 615573 676350 615578
rect 676290 615458 676350 615573
rect 676239 615192 676305 615195
rect 676239 615190 676350 615192
rect 676239 615134 676244 615190
rect 676300 615134 676350 615190
rect 676239 615129 676350 615134
rect 676290 615014 676350 615129
rect 58959 614452 59025 614455
rect 676047 614452 676113 614455
rect 58959 614450 64638 614452
rect 58959 614394 58964 614450
rect 59020 614394 64638 614450
rect 58959 614392 64638 614394
rect 58959 614389 59025 614392
rect 64578 613870 64638 614392
rect 676047 614450 676320 614452
rect 676047 614394 676052 614450
rect 676108 614394 676320 614450
rect 676047 614392 676320 614394
rect 676047 614389 676113 614392
rect 679938 613715 679998 613904
rect 679938 613710 680049 613715
rect 679938 613654 679988 613710
rect 680044 613654 680049 613710
rect 679938 613652 680049 613654
rect 679983 613649 680049 613652
rect 679746 613271 679806 613534
rect 59631 613268 59697 613271
rect 59631 613266 64638 613268
rect 59631 613210 59636 613266
rect 59692 613210 64638 613266
rect 59631 613208 64638 613210
rect 679746 613266 679857 613271
rect 679983 613268 680049 613271
rect 679746 613210 679796 613266
rect 679852 613210 679857 613266
rect 679746 613208 679857 613210
rect 59631 613205 59697 613208
rect 64578 612688 64638 613208
rect 679791 613205 679857 613208
rect 679938 613266 680049 613268
rect 679938 613210 679988 613266
rect 680044 613210 680049 613266
rect 679938 613205 680049 613210
rect 679938 612942 679998 613205
rect 679791 612824 679857 612827
rect 679746 612822 679857 612824
rect 679746 612766 679796 612822
rect 679852 612766 679857 612822
rect 679746 612761 679857 612766
rect 679746 612424 679806 612761
rect 59535 612084 59601 612087
rect 59535 612082 64638 612084
rect 59535 612026 59540 612082
rect 59596 612026 64638 612082
rect 59535 612024 64638 612026
rect 59535 612021 59601 612024
rect 64578 611506 64638 612024
rect 674362 607730 674368 607794
rect 674432 607792 674438 607794
rect 675183 607792 675249 607795
rect 674432 607790 675249 607792
rect 674432 607734 675188 607790
rect 675244 607734 675249 607790
rect 674432 607732 675249 607734
rect 674432 607730 674438 607732
rect 675183 607729 675249 607732
rect 675183 606018 675249 606019
rect 675130 606016 675136 606018
rect 675092 605956 675136 606016
rect 675200 606014 675249 606018
rect 675244 605958 675249 606014
rect 675130 605954 675136 605956
rect 675200 605954 675249 605958
rect 675183 605953 675249 605954
rect 674746 604770 674752 604834
rect 674816 604832 674822 604834
rect 675279 604832 675345 604835
rect 674816 604830 675345 604832
rect 674816 604774 675284 604830
rect 675340 604774 675345 604830
rect 674816 604772 675345 604774
rect 674816 604770 674822 604772
rect 675279 604769 675345 604772
rect 41538 601727 41598 601842
rect 40335 601726 40401 601727
rect 40335 601724 40384 601726
rect 40292 601722 40384 601724
rect 40292 601666 40340 601722
rect 40292 601664 40384 601666
rect 40335 601662 40384 601664
rect 40448 601662 40454 601726
rect 41538 601722 41649 601727
rect 41538 601666 41588 601722
rect 41644 601666 41649 601722
rect 41538 601664 41649 601666
rect 40335 601661 40401 601662
rect 41583 601661 41649 601664
rect 41775 601428 41841 601431
rect 41568 601426 41841 601428
rect 41568 601370 41780 601426
rect 41836 601370 41841 601426
rect 41568 601368 41841 601370
rect 41775 601365 41841 601368
rect 41775 600836 41841 600839
rect 41568 600834 41841 600836
rect 41568 600778 41780 600834
rect 41836 600778 41841 600834
rect 41568 600776 41841 600778
rect 41775 600773 41841 600776
rect 41775 600392 41841 600395
rect 41568 600390 41841 600392
rect 41568 600334 41780 600390
rect 41836 600334 41841 600390
rect 41568 600332 41841 600334
rect 41775 600329 41841 600332
rect 675322 600182 675328 600246
rect 675392 600244 675398 600246
rect 675471 600244 675537 600247
rect 675392 600242 675537 600244
rect 675392 600186 675476 600242
rect 675532 600186 675537 600242
rect 675392 600184 675537 600186
rect 675392 600182 675398 600184
rect 675471 600181 675537 600184
rect 41775 599874 41841 599877
rect 41568 599872 41841 599874
rect 41568 599816 41780 599872
rect 41836 599816 41841 599872
rect 41568 599814 41841 599816
rect 41775 599811 41841 599814
rect 40335 599504 40401 599507
rect 43066 599504 43072 599506
rect 40335 599502 43072 599504
rect 40335 599446 40340 599502
rect 40396 599446 43072 599502
rect 40335 599444 43072 599446
rect 40335 599441 40401 599444
rect 43066 599442 43072 599444
rect 43136 599442 43142 599506
rect 41775 599356 41841 599359
rect 41568 599354 41841 599356
rect 41568 599298 41780 599354
rect 41836 599298 41841 599354
rect 41568 599296 41841 599298
rect 41775 599293 41841 599296
rect 40386 598767 40446 598882
rect 40335 598762 40446 598767
rect 40335 598706 40340 598762
rect 40396 598706 40446 598762
rect 40335 598704 40446 598706
rect 40335 598701 40401 598704
rect 41775 598394 41841 598397
rect 41568 598392 41841 598394
rect 41568 598336 41780 598392
rect 41836 598336 41841 598392
rect 41568 598334 41841 598336
rect 41775 598331 41841 598334
rect 41775 597876 41841 597879
rect 41568 597874 41841 597876
rect 41568 597818 41780 597874
rect 41836 597818 41841 597874
rect 41568 597816 41841 597818
rect 649986 597876 650046 598336
rect 655215 597876 655281 597879
rect 649986 597874 655281 597876
rect 649986 597818 655220 597874
rect 655276 597818 655281 597874
rect 649986 597816 655281 597818
rect 41775 597813 41841 597816
rect 655215 597813 655281 597816
rect 37314 597139 37374 597402
rect 37314 597134 37425 597139
rect 37314 597078 37364 597134
rect 37420 597078 37425 597134
rect 37314 597076 37425 597078
rect 37359 597073 37425 597076
rect 41538 596695 41598 596810
rect 41538 596690 41649 596695
rect 41538 596634 41588 596690
rect 41644 596634 41649 596690
rect 41538 596632 41649 596634
rect 649986 596692 650046 597154
rect 655407 596692 655473 596695
rect 649986 596690 655473 596692
rect 649986 596634 655412 596690
rect 655468 596634 655473 596690
rect 649986 596632 655473 596634
rect 41583 596629 41649 596632
rect 655407 596629 655473 596632
rect 34242 596103 34302 596366
rect 34242 596098 34353 596103
rect 34242 596042 34292 596098
rect 34348 596042 34353 596098
rect 34242 596040 34353 596042
rect 34287 596037 34353 596040
rect 40194 595659 40254 595922
rect 40143 595654 40254 595659
rect 40143 595598 40148 595654
rect 40204 595598 40254 595654
rect 40143 595596 40254 595598
rect 40143 595593 40209 595596
rect 649986 595508 650046 595972
rect 655599 595508 655665 595511
rect 649986 595506 655665 595508
rect 649986 595450 655604 595506
rect 655660 595450 655665 595506
rect 649986 595448 655665 595450
rect 655599 595445 655665 595448
rect 41967 595360 42033 595363
rect 655791 595360 655857 595363
rect 41568 595358 42033 595360
rect 41568 595302 41972 595358
rect 42028 595302 42033 595358
rect 41568 595300 42033 595302
rect 41967 595297 42033 595300
rect 649986 595358 655857 595360
rect 649986 595302 655796 595358
rect 655852 595302 655857 595358
rect 649986 595300 655857 595302
rect 41775 594842 41841 594845
rect 41568 594840 41841 594842
rect 41568 594784 41780 594840
rect 41836 594784 41841 594840
rect 649986 594790 650046 595300
rect 655791 595297 655857 595300
rect 675759 595360 675825 595363
rect 676282 595360 676288 595362
rect 675759 595358 676288 595360
rect 675759 595302 675764 595358
rect 675820 595302 676288 595358
rect 675759 595300 676288 595302
rect 675759 595297 675825 595300
rect 676282 595298 676288 595300
rect 676352 595298 676358 595362
rect 41568 594782 41841 594784
rect 41775 594779 41841 594782
rect 34434 594179 34494 594442
rect 34383 594174 34494 594179
rect 653967 594176 654033 594179
rect 34383 594118 34388 594174
rect 34444 594118 34494 594174
rect 34383 594116 34494 594118
rect 649986 594174 654033 594176
rect 649986 594118 653972 594174
rect 654028 594118 654033 594174
rect 649986 594116 654033 594118
rect 34383 594113 34449 594116
rect 40194 593735 40254 593850
rect 40194 593730 40305 593735
rect 40194 593674 40244 593730
rect 40300 593674 40305 593730
rect 40194 593672 40305 593674
rect 40239 593669 40305 593672
rect 649986 593608 650046 594116
rect 653967 594113 654033 594116
rect 675663 593438 675729 593439
rect 675663 593434 675712 593438
rect 675776 593436 675782 593438
rect 675663 593378 675668 593434
rect 675663 593374 675712 593378
rect 675776 593376 675820 593436
rect 675776 593374 675782 593376
rect 675663 593373 675729 593374
rect 34434 593143 34494 593332
rect 34434 593138 34545 593143
rect 34434 593082 34484 593138
rect 34540 593082 34545 593138
rect 34434 593080 34545 593082
rect 34479 593077 34545 593080
rect 41871 592992 41937 592995
rect 656559 592992 656625 592995
rect 41568 592990 41937 592992
rect 41568 592934 41876 592990
rect 41932 592934 41937 592990
rect 41568 592932 41937 592934
rect 41871 592929 41937 592932
rect 649986 592990 656625 592992
rect 649986 592934 656564 592990
rect 656620 592934 656625 592990
rect 649986 592932 656625 592934
rect 649986 592426 650046 592932
rect 656559 592929 656625 592932
rect 42063 592400 42129 592403
rect 41568 592398 42129 592400
rect 41568 592342 42068 592398
rect 42124 592342 42129 592398
rect 41568 592340 42129 592342
rect 42063 592337 42129 592340
rect 42255 591808 42321 591811
rect 41568 591806 42321 591808
rect 41568 591750 42260 591806
rect 42316 591750 42321 591806
rect 41568 591748 42321 591750
rect 42255 591745 42321 591748
rect 41538 591364 41598 591408
rect 42159 591364 42225 591367
rect 41538 591362 42225 591364
rect 41538 591306 42164 591362
rect 42220 591306 42225 591362
rect 41538 591304 42225 591306
rect 42159 591301 42225 591304
rect 41583 591068 41649 591071
rect 41538 591066 41649 591068
rect 41538 591010 41588 591066
rect 41644 591010 41649 591066
rect 41538 591005 41649 591010
rect 41538 590890 41598 591005
rect 41538 590180 41598 590298
rect 41538 590120 41790 590180
rect 28866 589591 28926 589928
rect 41730 589736 41790 590120
rect 28815 589586 28926 589591
rect 28815 589530 28820 589586
rect 28876 589530 28926 589586
rect 28815 589528 28926 589530
rect 41538 589676 41790 589736
rect 28815 589525 28881 589528
rect 41538 589147 41598 589676
rect 28815 589144 28881 589147
rect 28815 589142 28926 589144
rect 28815 589086 28820 589142
rect 28876 589086 28926 589142
rect 28815 589081 28926 589086
rect 41538 589142 41649 589147
rect 41538 589086 41588 589142
rect 41644 589086 41649 589142
rect 41538 589084 41649 589086
rect 41583 589081 41649 589084
rect 28866 588818 28926 589081
rect 34383 585740 34449 585743
rect 40378 585740 40384 585742
rect 34383 585738 40384 585740
rect 34383 585682 34388 585738
rect 34444 585682 40384 585738
rect 34383 585680 40384 585682
rect 34383 585677 34449 585680
rect 40378 585678 40384 585680
rect 40448 585678 40454 585742
rect 34287 585296 34353 585299
rect 40570 585296 40576 585298
rect 34287 585294 40576 585296
rect 34287 585238 34292 585294
rect 34348 585238 40576 585294
rect 34287 585236 40576 585238
rect 34287 585233 34353 585236
rect 40570 585234 40576 585236
rect 40640 585234 40646 585298
rect 42255 584852 42321 584855
rect 42682 584852 42688 584854
rect 42255 584850 42688 584852
rect 42255 584794 42260 584850
rect 42316 584794 42688 584850
rect 42255 584792 42688 584794
rect 42255 584789 42321 584792
rect 42682 584790 42688 584792
rect 42752 584790 42758 584854
rect 41871 584262 41937 584263
rect 42255 584262 42321 584263
rect 41871 584260 41920 584262
rect 41828 584258 41920 584260
rect 41828 584202 41876 584258
rect 41828 584200 41920 584202
rect 41871 584198 41920 584200
rect 41984 584198 41990 584262
rect 42255 584260 42304 584262
rect 42212 584258 42304 584260
rect 42212 584202 42260 584258
rect 42212 584200 42304 584202
rect 42255 584198 42304 584200
rect 42368 584198 42374 584262
rect 41871 584197 41937 584198
rect 42255 584197 42321 584198
rect 42682 578722 42688 578786
rect 42752 578784 42758 578786
rect 43023 578784 43089 578787
rect 42752 578782 43089 578784
rect 42752 578726 43028 578782
rect 43084 578726 43089 578782
rect 42752 578724 43089 578726
rect 42752 578722 42758 578724
rect 43023 578721 43089 578724
rect 676290 578343 676350 578458
rect 42298 578278 42304 578342
rect 42368 578340 42374 578342
rect 42543 578340 42609 578343
rect 42368 578338 42609 578340
rect 42368 578282 42548 578338
rect 42604 578282 42609 578338
rect 42368 578280 42609 578282
rect 676290 578338 676401 578343
rect 676290 578282 676340 578338
rect 676396 578282 676401 578338
rect 676290 578280 676401 578282
rect 42368 578278 42374 578280
rect 42543 578277 42609 578280
rect 676335 578277 676401 578280
rect 676143 577600 676209 577603
rect 676290 577600 676350 577866
rect 676143 577598 676350 577600
rect 676143 577542 676148 577598
rect 676204 577542 676350 577598
rect 676143 577540 676350 577542
rect 676143 577537 676209 577540
rect 676290 577159 676350 577422
rect 676239 577154 676350 577159
rect 676239 577098 676244 577154
rect 676300 577098 676350 577154
rect 676239 577096 676350 577098
rect 676239 577093 676305 577096
rect 676047 577008 676113 577011
rect 676047 577006 676320 577008
rect 676047 576950 676052 577006
rect 676108 576950 676320 577006
rect 676047 576948 676320 576950
rect 676047 576945 676113 576948
rect 676290 576271 676350 576386
rect 676239 576266 676350 576271
rect 676239 576210 676244 576266
rect 676300 576210 676350 576266
rect 676239 576208 676350 576210
rect 676239 576205 676305 576208
rect 676047 575972 676113 575975
rect 676047 575970 676320 575972
rect 676047 575914 676052 575970
rect 676108 575914 676320 575970
rect 676047 575912 676320 575914
rect 676047 575909 676113 575912
rect 676047 575528 676113 575531
rect 676047 575526 676320 575528
rect 676047 575470 676052 575526
rect 676108 575470 676320 575526
rect 676047 575468 676320 575470
rect 676047 575465 676113 575468
rect 40570 575318 40576 575382
rect 40640 575380 40646 575382
rect 42351 575380 42417 575383
rect 40640 575378 42417 575380
rect 40640 575322 42356 575378
rect 42412 575322 42417 575378
rect 40640 575320 42417 575322
rect 40640 575318 40646 575320
rect 42351 575317 42417 575320
rect 676047 574936 676113 574939
rect 676047 574934 676320 574936
rect 676047 574878 676052 574934
rect 676108 574878 676320 574934
rect 676047 574876 676320 574878
rect 676047 574873 676113 574876
rect 58959 574788 59025 574791
rect 58959 574786 64638 574788
rect 58959 574730 58964 574786
rect 59020 574730 64638 574786
rect 58959 574728 64638 574730
rect 58959 574725 59025 574728
rect 64578 574194 64638 574728
rect 676047 574418 676113 574421
rect 676047 574416 676320 574418
rect 676047 574360 676052 574416
rect 676108 574360 676320 574416
rect 676047 574358 676320 574360
rect 676047 574355 676113 574358
rect 40378 573986 40384 574050
rect 40448 574048 40454 574050
rect 43119 574048 43185 574051
rect 40448 574046 43185 574048
rect 40448 573990 43124 574046
rect 43180 573990 43185 574046
rect 40448 573988 43185 573990
rect 40448 573986 40454 573988
rect 43119 573985 43185 573988
rect 674938 573986 674944 574050
rect 675008 574048 675014 574050
rect 675008 573988 676320 574048
rect 675008 573986 675014 573988
rect 676090 573690 676096 573754
rect 676160 573752 676166 573754
rect 676160 573692 676350 573752
rect 676160 573690 676166 573692
rect 676290 573426 676350 573692
rect 59631 573012 59697 573015
rect 59631 573010 64638 573012
rect 59631 572954 59636 573010
rect 59692 572954 64638 573010
rect 59631 572952 64638 572954
rect 59631 572949 59697 572952
rect 673978 572802 673984 572866
rect 674048 572864 674054 572866
rect 674048 572804 676320 572864
rect 674048 572802 674054 572804
rect 41871 572718 41937 572719
rect 41871 572714 41920 572718
rect 41984 572716 41990 572718
rect 41871 572658 41876 572714
rect 41871 572654 41920 572658
rect 41984 572656 42028 572716
rect 41984 572654 41990 572656
rect 41871 572653 41937 572654
rect 674554 572506 674560 572570
rect 674624 572568 674630 572570
rect 674624 572508 676320 572568
rect 674624 572506 674630 572508
rect 58191 572420 58257 572423
rect 58191 572418 64638 572420
rect 58191 572362 58196 572418
rect 58252 572362 64638 572418
rect 58191 572360 64638 572362
rect 58191 572357 58257 572360
rect 64578 571830 64638 572360
rect 675514 571914 675520 571978
rect 675584 571976 675590 571978
rect 675584 571916 676320 571976
rect 675584 571914 675590 571916
rect 675898 571322 675904 571386
rect 675968 571384 675974 571386
rect 675968 571324 676320 571384
rect 675968 571322 675974 571324
rect 58959 571236 59025 571239
rect 58959 571234 64638 571236
rect 58959 571178 58964 571234
rect 59020 571178 64638 571234
rect 58959 571176 64638 571178
rect 58959 571173 59025 571176
rect 64578 570648 64638 571176
rect 674170 571174 674176 571238
rect 674240 571236 674246 571238
rect 674240 571176 676350 571236
rect 674240 571174 674246 571176
rect 676290 570984 676350 571176
rect 676239 570644 676305 570647
rect 676239 570642 676350 570644
rect 676239 570586 676244 570642
rect 676300 570586 676350 570642
rect 676239 570581 676350 570586
rect 676290 570466 676350 570581
rect 59343 570052 59409 570055
rect 59343 570050 64638 570052
rect 59343 569994 59348 570050
rect 59404 569994 64638 570050
rect 59343 569992 64638 569994
rect 59343 569989 59409 569992
rect 64578 569466 64638 569992
rect 676047 569904 676113 569907
rect 676047 569902 676320 569904
rect 676047 569846 676052 569902
rect 676108 569846 676320 569902
rect 676047 569844 676320 569846
rect 676047 569841 676113 569844
rect 676047 569534 676113 569537
rect 676047 569532 676320 569534
rect 676047 569476 676052 569532
rect 676108 569476 676320 569532
rect 676047 569474 676320 569476
rect 676047 569471 676113 569474
rect 676239 569164 676305 569167
rect 676239 569162 676350 569164
rect 676239 569106 676244 569162
rect 676300 569106 676350 569162
rect 676239 569101 676350 569106
rect 676290 568986 676350 569101
rect 59535 568868 59601 568871
rect 59535 568866 64638 568868
rect 59535 568810 59540 568866
rect 59596 568810 64638 568866
rect 59535 568808 64638 568810
rect 59535 568805 59601 568808
rect 64578 568284 64638 568808
rect 676047 568424 676113 568427
rect 676047 568422 676320 568424
rect 676047 568366 676052 568422
rect 676108 568366 676320 568422
rect 676047 568364 676320 568366
rect 676047 568361 676113 568364
rect 676047 567980 676113 567983
rect 676047 567978 676320 567980
rect 676047 567922 676052 567978
rect 676108 567922 676320 567978
rect 676047 567920 676320 567922
rect 676047 567917 676113 567920
rect 676239 567684 676305 567687
rect 676239 567682 676350 567684
rect 676239 567626 676244 567682
rect 676300 567626 676350 567682
rect 676239 567621 676350 567626
rect 676290 567506 676350 567621
rect 679791 567092 679857 567095
rect 679746 567090 679857 567092
rect 679746 567034 679796 567090
rect 679852 567034 679857 567090
rect 679746 567029 679857 567034
rect 679746 566914 679806 567029
rect 685506 566207 685566 566470
rect 679791 566204 679857 566207
rect 679746 566202 679857 566204
rect 679746 566146 679796 566202
rect 679852 566146 679857 566202
rect 679746 566141 679857 566146
rect 685455 566202 685566 566207
rect 685455 566146 685460 566202
rect 685516 566146 685566 566202
rect 685455 566144 685566 566146
rect 685455 566141 685521 566144
rect 679746 565952 679806 566141
rect 685455 565760 685521 565763
rect 685455 565758 685566 565760
rect 685455 565702 685460 565758
rect 685516 565702 685566 565758
rect 685455 565697 685566 565702
rect 685506 565434 685566 565697
rect 675471 562506 675537 562507
rect 675471 562502 675520 562506
rect 675584 562504 675590 562506
rect 675471 562446 675476 562502
rect 675471 562442 675520 562446
rect 675584 562444 675628 562504
rect 675584 562442 675590 562444
rect 675471 562441 675537 562442
rect 674170 561702 674176 561766
rect 674240 561764 674246 561766
rect 675183 561764 675249 561767
rect 674240 561762 675249 561764
rect 674240 561706 675188 561762
rect 675244 561706 675249 561762
rect 674240 561704 675249 561706
rect 674240 561702 674246 561704
rect 675183 561701 675249 561704
rect 674938 561406 674944 561470
rect 675008 561468 675014 561470
rect 675375 561468 675441 561471
rect 675008 561466 675441 561468
rect 675008 561410 675380 561466
rect 675436 561410 675441 561466
rect 675008 561408 675441 561410
rect 675008 561406 675014 561408
rect 675375 561405 675441 561408
rect 674554 558890 674560 558954
rect 674624 558952 674630 558954
rect 675471 558952 675537 558955
rect 674624 558950 675537 558952
rect 674624 558894 675476 558950
rect 675532 558894 675537 558950
rect 674624 558892 675537 558894
rect 674624 558890 674630 558892
rect 675471 558889 675537 558892
rect 649986 553328 650046 553914
rect 655119 553328 655185 553331
rect 649986 553326 655185 553328
rect 649986 553270 655124 553326
rect 655180 553270 655185 553326
rect 649986 553268 655185 553270
rect 655119 553265 655185 553268
rect 649986 552144 650046 552732
rect 655503 552144 655569 552147
rect 649986 552142 655569 552144
rect 649986 552086 655508 552142
rect 655564 552086 655569 552142
rect 649986 552084 655569 552086
rect 655503 552081 655569 552084
rect 649986 550960 650046 551550
rect 655311 550960 655377 550963
rect 649986 550958 655377 550960
rect 649986 550902 655316 550958
rect 655372 550902 655377 550958
rect 649986 550900 655377 550902
rect 655311 550897 655377 550900
rect 655695 550812 655761 550815
rect 649986 550810 655761 550812
rect 649986 550754 655700 550810
rect 655756 550754 655761 550810
rect 649986 550752 655761 550754
rect 649986 550368 650046 550752
rect 655695 550749 655761 550752
rect 656559 549776 656625 549779
rect 649986 549774 656625 549776
rect 649986 549718 656564 549774
rect 656620 549718 656625 549774
rect 649986 549716 656625 549718
rect 649986 549186 650046 549716
rect 656559 549713 656625 549716
rect 654159 548592 654225 548595
rect 649986 548590 654225 548592
rect 649986 548534 654164 548590
rect 654220 548534 654225 548590
rect 649986 548532 654225 548534
rect 649986 548004 650046 548532
rect 654159 548529 654225 548532
rect 40378 539798 40384 539862
rect 40448 539860 40454 539862
rect 41775 539860 41841 539863
rect 40448 539858 41841 539860
rect 40448 539802 41780 539858
rect 41836 539802 41841 539858
rect 40448 539800 41841 539802
rect 40448 539798 40454 539800
rect 41775 539797 41841 539800
rect 41146 538022 41152 538086
rect 41216 538084 41222 538086
rect 41775 538084 41841 538087
rect 41216 538082 41841 538084
rect 41216 538026 41780 538082
rect 41836 538026 41841 538082
rect 41216 538024 41841 538026
rect 41216 538022 41222 538024
rect 41775 538021 41841 538024
rect 42874 536986 42880 537050
rect 42944 537048 42950 537050
rect 62127 537048 62193 537051
rect 42944 537046 62193 537048
rect 42944 536990 62132 537046
rect 62188 536990 62193 537046
rect 42944 536988 62193 536990
rect 42944 536986 42950 536988
rect 62127 536985 62193 536988
rect 40954 536246 40960 536310
rect 41024 536308 41030 536310
rect 41775 536308 41841 536311
rect 41024 536306 41841 536308
rect 41024 536250 41780 536306
rect 41836 536250 41841 536306
rect 41024 536248 41841 536250
rect 41024 536246 41030 536248
rect 41775 536245 41841 536248
rect 40762 535062 40768 535126
rect 40832 535124 40838 535126
rect 41775 535124 41841 535127
rect 40832 535122 41841 535124
rect 40832 535066 41780 535122
rect 41836 535066 41841 535122
rect 40832 535064 41841 535066
rect 40832 535062 40838 535064
rect 41775 535061 41841 535064
rect 676143 534976 676209 534979
rect 676290 534976 676350 535242
rect 676143 534974 676350 534976
rect 676143 534918 676148 534974
rect 676204 534918 676350 534974
rect 676143 534916 676350 534918
rect 676143 534913 676209 534916
rect 676290 534387 676350 534724
rect 676239 534382 676350 534387
rect 676239 534326 676244 534382
rect 676300 534326 676350 534382
rect 676239 534324 676350 534326
rect 676239 534321 676305 534324
rect 41530 534174 41536 534238
rect 41600 534236 41606 534238
rect 41775 534236 41841 534239
rect 41600 534234 41841 534236
rect 41600 534178 41780 534234
rect 41836 534178 41841 534234
rect 41600 534176 41841 534178
rect 41600 534174 41606 534176
rect 41775 534173 41841 534176
rect 676047 534236 676113 534239
rect 676047 534234 676320 534236
rect 676047 534178 676052 534234
rect 676108 534178 676320 534234
rect 676047 534176 676320 534178
rect 676047 534173 676113 534176
rect 40570 533878 40576 533942
rect 40640 533940 40646 533942
rect 41775 533940 41841 533943
rect 40640 533938 41841 533940
rect 40640 533882 41780 533938
rect 41836 533882 41841 533938
rect 40640 533880 41841 533882
rect 40640 533878 40646 533880
rect 41775 533877 41841 533880
rect 675951 533792 676017 533795
rect 675951 533790 676320 533792
rect 675951 533734 675956 533790
rect 676012 533734 676320 533790
rect 675951 533732 676320 533734
rect 675951 533729 676017 533732
rect 41775 533202 41841 533203
rect 41722 533200 41728 533202
rect 41684 533140 41728 533200
rect 41792 533198 41841 533202
rect 41836 533142 41841 533198
rect 41722 533138 41728 533140
rect 41792 533138 41841 533142
rect 41775 533137 41841 533138
rect 676482 533055 676542 533170
rect 676482 533050 676593 533055
rect 676482 532994 676532 533050
rect 676588 532994 676593 533050
rect 676482 532992 676593 532994
rect 676527 532989 676593 532992
rect 676047 532756 676113 532759
rect 676047 532754 676320 532756
rect 676047 532698 676052 532754
rect 676108 532698 676320 532754
rect 676047 532696 676320 532698
rect 676047 532693 676113 532696
rect 676674 532019 676734 532282
rect 676623 532014 676734 532019
rect 676623 531958 676628 532014
rect 676684 531958 676734 532014
rect 676623 531956 676734 531958
rect 676623 531953 676689 531956
rect 57711 531720 57777 531723
rect 57711 531718 64638 531720
rect 57711 531662 57716 531718
rect 57772 531662 64638 531718
rect 57711 531660 64638 531662
rect 57711 531657 57777 531660
rect 64578 531172 64638 531660
rect 676290 531575 676350 531690
rect 676239 531570 676350 531575
rect 676239 531514 676244 531570
rect 676300 531514 676350 531570
rect 676239 531512 676350 531514
rect 676239 531509 676305 531512
rect 676674 530983 676734 531246
rect 676674 530978 676785 530983
rect 676674 530922 676724 530978
rect 676780 530922 676785 530978
rect 676674 530920 676785 530922
rect 676719 530917 676785 530920
rect 41338 530770 41344 530834
rect 41408 530832 41414 530834
rect 41775 530832 41841 530835
rect 41408 530830 41841 530832
rect 41408 530774 41780 530830
rect 41836 530774 41841 530830
rect 41408 530772 41841 530774
rect 41408 530770 41414 530772
rect 41775 530769 41841 530772
rect 675130 530770 675136 530834
rect 675200 530832 675206 530834
rect 675200 530772 676320 530832
rect 675200 530770 675206 530772
rect 57615 530536 57681 530539
rect 57615 530534 64638 530536
rect 57615 530478 57620 530534
rect 57676 530478 64638 530534
rect 57615 530476 64638 530478
rect 57615 530473 57681 530476
rect 41871 530094 41937 530095
rect 41871 530090 41920 530094
rect 41984 530092 41990 530094
rect 41871 530034 41876 530090
rect 41871 530030 41920 530034
rect 41984 530032 42028 530092
rect 41984 530030 41990 530032
rect 41871 530029 41937 530030
rect 64578 529990 64638 530476
rect 676282 530474 676288 530538
rect 676352 530474 676358 530538
rect 676290 530210 676350 530474
rect 674362 529882 674368 529946
rect 674432 529944 674438 529946
rect 674432 529884 676350 529944
rect 674432 529882 674438 529884
rect 676290 529692 676350 529884
rect 42063 529354 42129 529355
rect 42063 529350 42112 529354
rect 42176 529352 42182 529354
rect 58191 529352 58257 529355
rect 42063 529294 42068 529350
rect 42063 529290 42112 529294
rect 42176 529292 42220 529352
rect 58191 529350 64638 529352
rect 58191 529294 58196 529350
rect 58252 529294 64638 529350
rect 58191 529292 64638 529294
rect 42176 529290 42182 529292
rect 42063 529289 42129 529290
rect 58191 529289 58257 529292
rect 64578 528808 64638 529292
rect 674746 529290 674752 529354
rect 674816 529352 674822 529354
rect 674816 529292 676320 529352
rect 674816 529290 674822 529292
rect 42159 528760 42225 528763
rect 42298 528760 42304 528762
rect 42159 528758 42304 528760
rect 42159 528702 42164 528758
rect 42220 528702 42304 528758
rect 42159 528700 42304 528702
rect 42159 528697 42225 528700
rect 42298 528698 42304 528700
rect 42368 528698 42374 528762
rect 675322 528698 675328 528762
rect 675392 528760 675398 528762
rect 675392 528700 676320 528760
rect 675392 528698 675398 528700
rect 675706 528106 675712 528170
rect 675776 528168 675782 528170
rect 675776 528108 676320 528168
rect 675776 528106 675782 528108
rect 676239 528020 676305 528023
rect 676239 528018 676350 528020
rect 676239 527962 676244 528018
rect 676300 527962 676350 528018
rect 676239 527957 676350 527962
rect 676290 527842 676350 527957
rect 42159 527132 42225 527135
rect 42490 527132 42496 527134
rect 42159 527130 42496 527132
rect 42159 527074 42164 527130
rect 42220 527074 42496 527130
rect 42159 527072 42496 527074
rect 42159 527069 42225 527072
rect 42490 527070 42496 527072
rect 42560 527070 42566 527134
rect 58959 527132 59025 527135
rect 64578 527132 64638 527626
rect 676239 527428 676305 527431
rect 676239 527426 676350 527428
rect 676239 527370 676244 527426
rect 676300 527370 676350 527426
rect 676239 527365 676350 527370
rect 676290 527250 676350 527365
rect 58959 527130 64638 527132
rect 58959 527074 58964 527130
rect 59020 527074 64638 527130
rect 58959 527072 64638 527074
rect 58959 527069 59025 527072
rect 676047 526688 676113 526691
rect 676047 526686 676320 526688
rect 676047 526630 676052 526686
rect 676108 526630 676320 526686
rect 676047 526628 676320 526630
rect 676047 526625 676113 526628
rect 58575 525948 58641 525951
rect 64578 525948 64638 526444
rect 676047 526318 676113 526321
rect 676047 526316 676320 526318
rect 676047 526260 676052 526316
rect 676108 526260 676320 526316
rect 676047 526258 676320 526260
rect 676047 526255 676113 526258
rect 58575 525946 64638 525948
rect 58575 525890 58580 525946
rect 58636 525890 64638 525946
rect 58575 525888 64638 525890
rect 676239 525948 676305 525951
rect 676239 525946 676350 525948
rect 676239 525890 676244 525946
rect 676300 525890 676350 525946
rect 58575 525885 58641 525888
rect 676239 525885 676350 525890
rect 676290 525770 676350 525885
rect 59343 524764 59409 524767
rect 64578 524764 64638 525262
rect 676047 525208 676113 525211
rect 676047 525206 676320 525208
rect 676047 525150 676052 525206
rect 676108 525150 676320 525206
rect 676047 525148 676320 525150
rect 676047 525145 676113 525148
rect 676047 524838 676113 524841
rect 676047 524836 676320 524838
rect 676047 524780 676052 524836
rect 676108 524780 676320 524836
rect 676047 524778 676320 524780
rect 676047 524775 676113 524778
rect 59343 524762 64638 524764
rect 59343 524706 59348 524762
rect 59404 524706 64638 524762
rect 59343 524704 64638 524706
rect 59343 524701 59409 524704
rect 676239 524468 676305 524471
rect 676239 524466 676350 524468
rect 676239 524410 676244 524466
rect 676300 524410 676350 524466
rect 676239 524405 676350 524410
rect 676290 524290 676350 524405
rect 679746 523583 679806 523698
rect 679746 523578 679857 523583
rect 679746 523522 679796 523578
rect 679852 523522 679857 523578
rect 679746 523520 679857 523522
rect 679791 523517 679857 523520
rect 685506 522991 685566 523254
rect 679791 522988 679857 522991
rect 679746 522986 679857 522988
rect 679746 522930 679796 522986
rect 679852 522930 679857 522986
rect 679746 522925 679857 522930
rect 685455 522986 685566 522991
rect 685455 522930 685460 522986
rect 685516 522930 685566 522986
rect 685455 522928 685566 522930
rect 685455 522925 685521 522928
rect 679746 522810 679806 522925
rect 685455 522544 685521 522547
rect 685455 522542 685566 522544
rect 685455 522486 685460 522542
rect 685516 522486 685566 522542
rect 685455 522481 685566 522486
rect 685506 522218 685566 522481
rect 676290 490579 676350 490842
rect 676239 490574 676350 490579
rect 676239 490518 676244 490574
rect 676300 490518 676350 490574
rect 676239 490516 676350 490518
rect 676239 490513 676305 490516
rect 676143 490132 676209 490135
rect 676290 490132 676350 490324
rect 676143 490130 676350 490132
rect 676143 490074 676148 490130
rect 676204 490074 676350 490130
rect 676143 490072 676350 490074
rect 676143 490069 676209 490072
rect 676239 489984 676305 489987
rect 676239 489982 676350 489984
rect 676239 489926 676244 489982
rect 676300 489926 676350 489982
rect 676239 489921 676350 489926
rect 676290 489806 676350 489921
rect 679746 489247 679806 489362
rect 679695 489242 679806 489247
rect 679695 489186 679700 489242
rect 679756 489186 679806 489242
rect 679695 489184 679806 489186
rect 679695 489181 679761 489184
rect 676674 488655 676734 488770
rect 676674 488650 676785 488655
rect 676674 488594 676724 488650
rect 676780 488594 676785 488650
rect 676674 488592 676785 488594
rect 676719 488589 676785 488592
rect 676047 488356 676113 488359
rect 676047 488354 676320 488356
rect 676047 488298 676052 488354
rect 676108 488298 676320 488354
rect 676047 488296 676320 488298
rect 676047 488293 676113 488296
rect 677826 487619 677886 487882
rect 677826 487614 677937 487619
rect 677826 487558 677876 487614
rect 677932 487558 677937 487614
rect 677826 487556 677937 487558
rect 677871 487553 677937 487556
rect 676290 487175 676350 487290
rect 676239 487170 676350 487175
rect 676239 487114 676244 487170
rect 676300 487114 676350 487170
rect 676239 487112 676350 487114
rect 676239 487109 676305 487112
rect 679746 486583 679806 486846
rect 679746 486578 679857 486583
rect 679746 486522 679796 486578
rect 679852 486522 679857 486578
rect 679746 486520 679857 486522
rect 679791 486517 679857 486520
rect 674938 486370 674944 486434
rect 675008 486432 675014 486434
rect 675008 486372 676320 486432
rect 675008 486370 675014 486372
rect 676047 485840 676113 485843
rect 676047 485838 676320 485840
rect 676047 485782 676052 485838
rect 676108 485782 676320 485838
rect 676047 485780 676320 485782
rect 676047 485777 676113 485780
rect 675514 485630 675520 485694
rect 675584 485692 675590 485694
rect 675584 485632 676350 485692
rect 675584 485630 675590 485632
rect 676290 485292 676350 485632
rect 676239 485100 676305 485103
rect 676239 485098 676350 485100
rect 676239 485042 676244 485098
rect 676300 485042 676350 485098
rect 676239 485037 676350 485042
rect 676290 484922 676350 485037
rect 676047 484360 676113 484363
rect 676047 484358 676320 484360
rect 676047 484302 676052 484358
rect 676108 484302 676320 484358
rect 676047 484300 676320 484302
rect 676047 484297 676113 484300
rect 675951 483768 676017 483771
rect 675951 483766 676320 483768
rect 675951 483710 675956 483766
rect 676012 483710 676320 483766
rect 675951 483708 676320 483710
rect 675951 483705 676017 483708
rect 674170 483410 674176 483474
rect 674240 483472 674246 483474
rect 674240 483412 676320 483472
rect 674240 483410 674246 483412
rect 674554 482818 674560 482882
rect 674624 482880 674630 482882
rect 674624 482820 676320 482880
rect 674624 482818 674630 482820
rect 676047 482288 676113 482291
rect 676047 482286 676320 482288
rect 676047 482230 676052 482286
rect 676108 482230 676320 482286
rect 676047 482228 676320 482230
rect 676047 482225 676113 482228
rect 676047 481918 676113 481921
rect 676047 481916 676320 481918
rect 676047 481860 676052 481916
rect 676108 481860 676320 481916
rect 676047 481858 676320 481860
rect 676047 481855 676113 481858
rect 676239 481548 676305 481551
rect 676239 481546 676350 481548
rect 676239 481490 676244 481546
rect 676300 481490 676350 481546
rect 676239 481485 676350 481490
rect 676290 481370 676350 481485
rect 676047 480808 676113 480811
rect 676047 480806 676320 480808
rect 676047 480750 676052 480806
rect 676108 480750 676320 480806
rect 676047 480748 676320 480750
rect 676047 480745 676113 480748
rect 676047 480438 676113 480441
rect 676047 480436 676320 480438
rect 676047 480380 676052 480436
rect 676108 480380 676320 480436
rect 676047 480378 676320 480380
rect 676047 480375 676113 480378
rect 676239 480068 676305 480071
rect 676239 480066 676350 480068
rect 676239 480010 676244 480066
rect 676300 480010 676350 480066
rect 676239 480005 676350 480010
rect 676290 479890 676350 480005
rect 679938 479183 679998 479298
rect 679887 479178 679998 479183
rect 679887 479122 679892 479178
rect 679948 479122 679998 479178
rect 679887 479120 679998 479122
rect 679887 479117 679953 479120
rect 679746 478591 679806 478854
rect 679695 478586 679806 478591
rect 679695 478530 679700 478586
rect 679756 478530 679806 478586
rect 679695 478528 679806 478530
rect 679887 478588 679953 478591
rect 679887 478586 679998 478588
rect 679887 478530 679892 478586
rect 679948 478530 679998 478586
rect 679695 478525 679761 478528
rect 679887 478525 679998 478530
rect 679938 478410 679998 478525
rect 679695 478144 679761 478147
rect 679695 478142 679806 478144
rect 679695 478086 679700 478142
rect 679756 478086 679806 478142
rect 679695 478081 679806 478086
rect 679746 477818 679806 478081
rect 41775 476072 41841 476075
rect 41568 476070 41841 476072
rect 41568 476014 41780 476070
rect 41836 476014 41841 476070
rect 41568 476012 41841 476014
rect 41775 476009 41841 476012
rect 41775 475554 41841 475557
rect 41568 475552 41841 475554
rect 41568 475496 41780 475552
rect 41836 475496 41841 475552
rect 41568 475494 41841 475496
rect 41775 475491 41841 475494
rect 41775 475036 41841 475039
rect 41568 475034 41841 475036
rect 41568 474978 41780 475034
rect 41836 474978 41841 475034
rect 41568 474976 41841 474978
rect 41775 474973 41841 474976
rect 41871 474592 41937 474595
rect 41568 474590 41937 474592
rect 41568 474534 41876 474590
rect 41932 474534 41937 474590
rect 41568 474532 41937 474534
rect 41871 474529 41937 474532
rect 40386 473855 40446 473970
rect 40386 473850 40497 473855
rect 40386 473794 40436 473850
rect 40492 473794 40497 473850
rect 40386 473792 40497 473794
rect 40431 473789 40497 473792
rect 39618 473263 39678 473526
rect 39618 473258 39729 473263
rect 39618 473202 39668 473258
rect 39724 473202 39729 473258
rect 39618 473200 39729 473202
rect 39663 473197 39729 473200
rect 43407 473112 43473 473115
rect 45231 473112 45297 473115
rect 41568 473110 45297 473112
rect 41568 473054 43412 473110
rect 43468 473054 45236 473110
rect 45292 473054 45297 473110
rect 41568 473052 45297 473054
rect 43407 473049 43473 473052
rect 45231 473049 45297 473052
rect 39810 472375 39870 472490
rect 39759 472370 39870 472375
rect 39759 472314 39764 472370
rect 39820 472314 39870 472370
rect 39759 472312 39870 472314
rect 39759 472309 39825 472312
rect 41583 472224 41649 472227
rect 41538 472222 41649 472224
rect 41538 472166 41588 472222
rect 41644 472166 41649 472222
rect 41538 472161 41649 472166
rect 41538 472046 41598 472161
rect 42490 471632 42496 471634
rect 41568 471572 42496 471632
rect 42490 471570 42496 471572
rect 42560 471570 42566 471634
rect 41146 471274 41152 471338
rect 41216 471274 41222 471338
rect 41154 471010 41214 471274
rect 37359 470744 37425 470747
rect 37314 470742 37425 470744
rect 37314 470686 37364 470742
rect 37420 470686 37425 470742
rect 37314 470681 37425 470686
rect 37314 470492 37374 470681
rect 42298 470152 42304 470154
rect 41568 470092 42304 470152
rect 42298 470090 42304 470092
rect 42368 470090 42374 470154
rect 41722 469560 41728 469562
rect 41568 469500 41728 469560
rect 41722 469498 41728 469500
rect 41792 469498 41798 469562
rect 40378 469350 40384 469414
rect 40448 469350 40454 469414
rect 40386 468938 40446 469350
rect 41583 468820 41649 468823
rect 41538 468818 41649 468820
rect 41538 468762 41588 468818
rect 41644 468762 41649 468818
rect 41538 468757 41649 468762
rect 41538 468642 41598 468757
rect 42106 468080 42112 468082
rect 41568 468020 42112 468080
rect 42106 468018 42112 468020
rect 42176 468018 42182 468082
rect 41914 467488 41920 467490
rect 41568 467428 41920 467488
rect 41914 467426 41920 467428
rect 41984 467426 41990 467490
rect 40954 467278 40960 467342
rect 41024 467278 41030 467342
rect 40962 467088 41022 467278
rect 41530 466834 41536 466898
rect 41600 466834 41606 466898
rect 41538 466570 41598 466834
rect 41338 466242 41344 466306
rect 41408 466242 41414 466306
rect 41346 465978 41406 466242
rect 40570 465798 40576 465862
rect 40640 465798 40646 465862
rect 40578 465608 40638 465798
rect 40762 465354 40768 465418
rect 40832 465354 40838 465418
rect 40770 465090 40830 465354
rect 34434 464383 34494 464498
rect 34434 464378 34545 464383
rect 34434 464322 34484 464378
rect 34540 464322 34545 464378
rect 34434 464320 34545 464322
rect 34479 464317 34545 464320
rect 23106 463791 23166 464054
rect 23055 463786 23166 463791
rect 23055 463730 23060 463786
rect 23116 463730 23166 463786
rect 23055 463728 23166 463730
rect 23055 463725 23121 463728
rect 41775 463640 41841 463643
rect 41568 463638 41841 463640
rect 41568 463582 41780 463638
rect 41836 463582 41841 463638
rect 41568 463580 41841 463582
rect 41775 463577 41841 463580
rect 23055 463344 23121 463347
rect 23055 463342 23166 463344
rect 23055 463286 23060 463342
rect 23116 463286 23166 463342
rect 23055 463281 23166 463286
rect 23106 463018 23166 463281
rect 41538 426939 41598 427054
rect 41538 426934 41649 426939
rect 41538 426878 41588 426934
rect 41644 426878 41649 426934
rect 41538 426876 41649 426878
rect 41583 426873 41649 426876
rect 41775 426566 41841 426569
rect 41568 426564 41841 426566
rect 41568 426508 41780 426564
rect 41836 426508 41841 426564
rect 41568 426506 41841 426508
rect 41775 426503 41841 426506
rect 41775 426048 41841 426051
rect 41568 426046 41841 426048
rect 41568 425990 41780 426046
rect 41836 425990 41841 426046
rect 41568 425988 41841 425990
rect 41775 425985 41841 425988
rect 40386 425311 40446 425574
rect 40386 425306 40497 425311
rect 40386 425250 40436 425306
rect 40492 425250 40497 425306
rect 40386 425248 40497 425250
rect 40431 425245 40497 425248
rect 41538 424867 41598 424982
rect 41538 424862 41649 424867
rect 41538 424806 41588 424862
rect 41644 424806 41649 424862
rect 41538 424804 41649 424806
rect 41583 424801 41649 424804
rect 34434 424275 34494 424538
rect 34434 424270 34545 424275
rect 39663 424272 39729 424275
rect 34434 424214 34484 424270
rect 34540 424214 34545 424270
rect 34434 424212 34545 424214
rect 34479 424209 34545 424212
rect 39618 424270 39729 424272
rect 39618 424214 39668 424270
rect 39724 424214 39729 424270
rect 39618 424209 39729 424214
rect 39618 424094 39678 424209
rect 41775 423532 41841 423535
rect 41568 423530 41841 423532
rect 41568 423474 41780 423530
rect 41836 423474 41841 423530
rect 41568 423472 41841 423474
rect 41775 423469 41841 423472
rect 41538 422795 41598 422984
rect 41538 422790 41649 422795
rect 41538 422734 41588 422790
rect 41644 422734 41649 422790
rect 41538 422732 41649 422734
rect 41583 422729 41649 422732
rect 41538 422350 41598 422614
rect 41530 422286 41536 422350
rect 41600 422286 41606 422350
rect 40386 421906 40446 422022
rect 40378 421842 40384 421906
rect 40448 421842 40454 421906
rect 34479 421756 34545 421759
rect 42490 421756 42496 421758
rect 34479 421754 42496 421756
rect 34479 421698 34484 421754
rect 34540 421698 42496 421754
rect 34479 421696 42496 421698
rect 34479 421693 34545 421696
rect 42490 421694 42496 421696
rect 42560 421694 42566 421758
rect 40578 421314 40638 421504
rect 40570 421250 40576 421314
rect 40640 421250 40646 421314
rect 39810 420871 39870 421134
rect 39759 420866 39870 420871
rect 39759 420810 39764 420866
rect 39820 420810 39870 420866
rect 39759 420808 39870 420810
rect 39759 420805 39825 420808
rect 40002 420279 40062 420542
rect 39951 420274 40062 420279
rect 39951 420218 39956 420274
rect 40012 420218 40062 420274
rect 39951 420216 40062 420218
rect 39951 420213 40017 420216
rect 39810 419835 39870 419950
rect 39810 419830 39921 419835
rect 39810 419774 39860 419830
rect 39916 419774 39921 419830
rect 39810 419772 39921 419774
rect 39855 419769 39921 419772
rect 39618 419243 39678 419580
rect 39618 419238 39729 419243
rect 39618 419182 39668 419238
rect 39724 419182 39729 419238
rect 39618 419180 39729 419182
rect 39663 419177 39729 419180
rect 40194 418799 40254 419062
rect 40194 418794 40305 418799
rect 40194 418738 40244 418794
rect 40300 418738 40305 418794
rect 40194 418736 40305 418738
rect 40239 418733 40305 418736
rect 40002 418355 40062 418470
rect 40002 418350 40113 418355
rect 40002 418294 40052 418350
rect 40108 418294 40113 418350
rect 40002 418292 40113 418294
rect 40047 418289 40113 418292
rect 40194 417911 40254 418100
rect 40143 417906 40254 417911
rect 40143 417850 40148 417906
rect 40204 417850 40254 417906
rect 40143 417848 40254 417850
rect 40143 417845 40209 417848
rect 40954 417698 40960 417762
rect 41024 417698 41030 417762
rect 40962 417582 41022 417698
rect 40239 417316 40305 417319
rect 41914 417316 41920 417318
rect 40239 417314 41920 417316
rect 40239 417258 40244 417314
rect 40300 417258 41920 417314
rect 40239 417256 41920 417258
rect 40239 417253 40305 417256
rect 41914 417254 41920 417256
rect 41984 417254 41990 417318
rect 41722 417020 41728 417022
rect 41568 416960 41728 417020
rect 41722 416958 41728 416960
rect 41792 416958 41798 417022
rect 39951 416872 40017 416875
rect 42106 416872 42112 416874
rect 39951 416870 42112 416872
rect 39951 416814 39956 416870
rect 40012 416814 42112 416870
rect 39951 416812 42112 416814
rect 39951 416809 40017 416812
rect 42106 416810 42112 416812
rect 42176 416810 42182 416874
rect 41538 416431 41598 416546
rect 39663 416428 39729 416431
rect 41146 416428 41152 416430
rect 39663 416426 41152 416428
rect 39663 416370 39668 416426
rect 39724 416370 41152 416426
rect 39663 416368 41152 416370
rect 39663 416365 39729 416368
rect 41146 416366 41152 416368
rect 41216 416366 41222 416430
rect 41538 416426 41649 416431
rect 41538 416370 41588 416426
rect 41644 416370 41649 416426
rect 41538 416368 41649 416370
rect 41583 416365 41649 416368
rect 40047 416280 40113 416283
rect 42298 416280 42304 416282
rect 40047 416278 42304 416280
rect 40047 416222 40052 416278
rect 40108 416222 42304 416278
rect 40047 416220 42304 416222
rect 40047 416217 40113 416220
rect 42298 416218 42304 416220
rect 42368 416218 42374 416282
rect 41871 416132 41937 416135
rect 41568 416130 41937 416132
rect 41568 416074 41876 416130
rect 41932 416074 41937 416130
rect 41568 416072 41937 416074
rect 41871 416069 41937 416072
rect 41568 415480 41790 415540
rect 23106 414803 23166 415066
rect 39759 414948 39825 414951
rect 41338 414948 41344 414950
rect 39759 414946 41344 414948
rect 39759 414890 39764 414946
rect 39820 414890 41344 414946
rect 39759 414888 41344 414890
rect 39759 414885 39825 414888
rect 41338 414886 41344 414888
rect 41408 414886 41414 414950
rect 41730 414948 41790 415480
rect 41538 414888 41790 414948
rect 23055 414798 23166 414803
rect 23055 414742 23060 414798
rect 23116 414742 23166 414798
rect 23055 414740 23166 414742
rect 23055 414737 23121 414740
rect 41538 414359 41598 414888
rect 23055 414356 23121 414359
rect 23055 414354 23166 414356
rect 23055 414298 23060 414354
rect 23116 414298 23166 414354
rect 23055 414293 23166 414298
rect 41538 414354 41649 414359
rect 41538 414298 41588 414354
rect 41644 414298 41649 414354
rect 41538 414296 41649 414298
rect 41583 414293 41649 414296
rect 23106 414030 23166 414293
rect 40378 411186 40384 411250
rect 40448 411248 40454 411250
rect 41871 411248 41937 411251
rect 40448 411246 41937 411248
rect 40448 411190 41876 411246
rect 41932 411190 41937 411246
rect 40448 411188 41937 411190
rect 40448 411186 40454 411188
rect 41871 411185 41937 411188
rect 40954 407634 40960 407698
rect 41024 407696 41030 407698
rect 41775 407696 41841 407699
rect 41024 407694 41841 407696
rect 41024 407638 41780 407694
rect 41836 407638 41841 407694
rect 41024 407636 41841 407638
rect 41024 407634 41030 407636
rect 41775 407633 41841 407636
rect 42063 406070 42129 406071
rect 42063 406066 42112 406070
rect 42176 406068 42182 406070
rect 42063 406010 42068 406066
rect 42063 406006 42112 406010
rect 42176 406008 42220 406068
rect 42176 406006 42182 406008
rect 42063 406005 42129 406006
rect 58479 404144 58545 404147
rect 58479 404142 64638 404144
rect 58479 404086 58484 404142
rect 58540 404086 64638 404142
rect 58479 404084 64638 404086
rect 58479 404081 58545 404084
rect 41775 403850 41841 403851
rect 41722 403848 41728 403850
rect 41684 403788 41728 403848
rect 41792 403846 41841 403850
rect 41836 403790 41841 403846
rect 41722 403786 41728 403788
rect 41792 403786 41841 403790
rect 41775 403785 41841 403786
rect 64578 403550 64638 404084
rect 42159 403108 42225 403111
rect 42298 403108 42304 403110
rect 42159 403106 42304 403108
rect 42159 403050 42164 403106
rect 42220 403050 42304 403106
rect 42159 403048 42304 403050
rect 42159 403045 42225 403048
rect 42298 403046 42304 403048
rect 42368 403046 42374 403110
rect 41871 402666 41937 402667
rect 41871 402662 41920 402666
rect 41984 402664 41990 402666
rect 41871 402606 41876 402662
rect 41871 402602 41920 402606
rect 41984 402604 42028 402664
rect 41984 402602 41990 402604
rect 41871 402601 41937 402602
rect 59343 402368 59409 402371
rect 676143 402368 676209 402371
rect 676290 402368 676350 402634
rect 59343 402366 64638 402368
rect 59343 402310 59348 402366
rect 59404 402310 64638 402366
rect 59343 402308 64638 402310
rect 676143 402366 676350 402368
rect 676143 402310 676148 402366
rect 676204 402310 676350 402366
rect 676143 402308 676350 402310
rect 59343 402305 59409 402308
rect 676143 402305 676209 402308
rect 41338 401862 41344 401926
rect 41408 401924 41414 401926
rect 41775 401924 41841 401927
rect 41408 401922 41841 401924
rect 41408 401866 41780 401922
rect 41836 401866 41841 401922
rect 41408 401864 41841 401866
rect 41408 401862 41414 401864
rect 41775 401861 41841 401864
rect 676290 401779 676350 402116
rect 676239 401774 676350 401779
rect 676239 401718 676244 401774
rect 676300 401718 676350 401774
rect 676239 401716 676350 401718
rect 676239 401713 676305 401716
rect 676047 401628 676113 401631
rect 676047 401626 676320 401628
rect 676047 401570 676052 401626
rect 676108 401570 676320 401626
rect 676047 401568 676320 401570
rect 676047 401565 676113 401568
rect 57711 400592 57777 400595
rect 64578 400592 64638 401186
rect 676674 401039 676734 401154
rect 676674 401034 676785 401039
rect 676674 400978 676724 401034
rect 676780 400978 676785 401034
rect 676674 400976 676785 400978
rect 676719 400973 676785 400976
rect 57711 400590 64638 400592
rect 57711 400534 57716 400590
rect 57772 400534 64638 400590
rect 57711 400532 64638 400534
rect 57711 400529 57777 400532
rect 676290 400447 676350 400636
rect 676239 400442 676350 400447
rect 676239 400386 676244 400442
rect 676300 400386 676350 400442
rect 676239 400384 676350 400386
rect 676239 400381 676305 400384
rect 676527 400296 676593 400299
rect 676482 400294 676593 400296
rect 676482 400238 676532 400294
rect 676588 400238 676593 400294
rect 676482 400233 676593 400238
rect 41530 400086 41536 400150
rect 41600 400148 41606 400150
rect 41775 400148 41841 400151
rect 41600 400146 41841 400148
rect 41600 400090 41780 400146
rect 41836 400090 41841 400146
rect 676482 400118 676542 400233
rect 41600 400088 41841 400090
rect 41600 400086 41606 400088
rect 41775 400085 41841 400088
rect 59631 400000 59697 400003
rect 64578 400000 64638 400004
rect 59631 399998 64638 400000
rect 59631 399942 59636 399998
rect 59692 399942 64638 399998
rect 59631 399940 64638 399942
rect 59631 399937 59697 399940
rect 676047 399704 676113 399707
rect 676047 399702 676320 399704
rect 676047 399646 676052 399702
rect 676108 399646 676320 399702
rect 676047 399644 676320 399646
rect 676047 399641 676113 399644
rect 41146 399346 41152 399410
rect 41216 399408 41222 399410
rect 41775 399408 41841 399411
rect 41216 399406 41841 399408
rect 41216 399350 41780 399406
rect 41836 399350 41841 399406
rect 41216 399348 41841 399350
rect 41216 399346 41222 399348
rect 41775 399345 41841 399348
rect 59727 399408 59793 399411
rect 676623 399408 676689 399411
rect 59727 399406 64638 399408
rect 59727 399350 59732 399406
rect 59788 399350 64638 399406
rect 59727 399348 64638 399350
rect 59727 399345 59793 399348
rect 64578 398822 64638 399348
rect 676623 399406 676734 399408
rect 676623 399350 676628 399406
rect 676684 399350 676734 399406
rect 676623 399345 676734 399350
rect 676674 399082 676734 399345
rect 40570 398754 40576 398818
rect 40640 398816 40646 398818
rect 41775 398816 41841 398819
rect 40640 398814 41841 398816
rect 40640 398758 41780 398814
rect 41836 398758 41841 398814
rect 40640 398756 41841 398758
rect 40640 398754 40646 398756
rect 41775 398753 41841 398756
rect 676047 398668 676113 398671
rect 676047 398666 676320 398668
rect 676047 398610 676052 398666
rect 676108 398610 676320 398666
rect 676047 398608 676320 398610
rect 676047 398605 676113 398608
rect 59535 398224 59601 398227
rect 59535 398222 64638 398224
rect 59535 398166 59540 398222
rect 59596 398166 64638 398222
rect 59535 398164 64638 398166
rect 59535 398161 59601 398164
rect 64578 397640 64638 398164
rect 676674 397930 676734 398194
rect 676666 397866 676672 397930
rect 676736 397866 676742 397930
rect 673978 397570 673984 397634
rect 674048 397632 674054 397634
rect 674048 397572 676320 397632
rect 674048 397570 674054 397572
rect 675130 396830 675136 396894
rect 675200 396892 675206 396894
rect 676290 396892 676350 397084
rect 675200 396832 676350 396892
rect 675200 396830 675206 396832
rect 676674 396450 676734 396714
rect 676666 396386 676672 396450
rect 676736 396386 676742 396450
rect 674746 396090 674752 396154
rect 674816 396152 674822 396154
rect 674816 396092 676320 396152
rect 674816 396090 674822 396092
rect 676047 395634 676113 395637
rect 676047 395632 676320 395634
rect 676047 395576 676052 395632
rect 676108 395576 676320 395632
rect 676047 395574 676320 395576
rect 676047 395571 676113 395574
rect 675898 395202 675904 395266
rect 675968 395264 675974 395266
rect 675968 395204 676320 395264
rect 675968 395202 675974 395204
rect 675322 394610 675328 394674
rect 675392 394672 675398 394674
rect 675392 394612 676320 394672
rect 675392 394610 675398 394612
rect 676482 393934 676542 394050
rect 676474 393870 676480 393934
rect 676544 393870 676550 393934
rect 676090 393278 676096 393342
rect 676160 393340 676166 393342
rect 676290 393340 676350 393680
rect 676160 393280 676350 393340
rect 676160 393278 676166 393280
rect 674362 393130 674368 393194
rect 674432 393192 674438 393194
rect 674432 393132 676320 393192
rect 674432 393130 674438 393132
rect 675706 392538 675712 392602
rect 675776 392600 675782 392602
rect 675776 392540 676320 392600
rect 675776 392538 675782 392540
rect 675514 391798 675520 391862
rect 675584 391860 675590 391862
rect 676290 391860 676350 392200
rect 675584 391800 676350 391860
rect 675584 391798 675590 391800
rect 676290 391418 676350 391682
rect 676282 391354 676288 391418
rect 676352 391354 676358 391418
rect 679746 390975 679806 391090
rect 679746 390970 679857 390975
rect 679746 390914 679796 390970
rect 679852 390914 679857 390970
rect 679746 390912 679857 390914
rect 679791 390909 679857 390912
rect 685506 390383 685566 390646
rect 679791 390380 679857 390383
rect 679746 390378 679857 390380
rect 679746 390322 679796 390378
rect 679852 390322 679857 390378
rect 679746 390317 679857 390322
rect 685455 390378 685566 390383
rect 685455 390322 685460 390378
rect 685516 390322 685566 390378
rect 685455 390320 685566 390322
rect 685455 390317 685521 390320
rect 679746 390202 679806 390317
rect 685455 389936 685521 389939
rect 685455 389934 685566 389936
rect 685455 389878 685460 389934
rect 685516 389878 685566 389934
rect 685455 389873 685566 389878
rect 685506 389610 685566 389873
rect 41775 388752 41841 388755
rect 42490 388752 42496 388754
rect 41775 388750 42496 388752
rect 41775 388694 41780 388750
rect 41836 388694 42496 388750
rect 41775 388692 42496 388694
rect 41775 388689 41841 388692
rect 42490 388690 42496 388692
rect 42560 388690 42566 388754
rect 41775 386384 41841 386387
rect 64719 386384 64785 386387
rect 41775 386382 64785 386384
rect 41775 386326 41780 386382
rect 41836 386326 64724 386382
rect 64780 386326 64785 386382
rect 41775 386324 64785 386326
rect 41775 386321 41841 386324
rect 64719 386321 64785 386324
rect 41538 385943 41598 386058
rect 41538 385938 41649 385943
rect 675183 385942 675249 385943
rect 41538 385882 41588 385938
rect 41644 385882 41649 385938
rect 41538 385880 41649 385882
rect 41583 385877 41649 385880
rect 675130 385878 675136 385942
rect 675200 385940 675249 385942
rect 675200 385938 675292 385940
rect 675244 385882 675292 385938
rect 675200 385880 675292 385882
rect 675200 385878 675249 385880
rect 675183 385877 675249 385878
rect 675759 385644 675825 385647
rect 675898 385644 675904 385646
rect 675759 385642 675904 385644
rect 675759 385586 675764 385642
rect 675820 385586 675904 385642
rect 675759 385584 675904 385586
rect 675759 385581 675825 385584
rect 675898 385582 675904 385584
rect 675968 385582 675974 385646
rect 41538 385351 41598 385466
rect 41538 385346 41649 385351
rect 41538 385290 41588 385346
rect 41644 385290 41649 385346
rect 41538 385288 41649 385290
rect 41583 385285 41649 385288
rect 41871 385052 41937 385055
rect 41568 385050 41937 385052
rect 41568 384994 41876 385050
rect 41932 384994 41937 385050
rect 41568 384992 41937 384994
rect 41871 384989 41937 384992
rect 41583 384756 41649 384759
rect 41538 384754 41649 384756
rect 41538 384698 41588 384754
rect 41644 384698 41649 384754
rect 41538 384693 41649 384698
rect 41538 384578 41598 384693
rect 674938 384398 674944 384462
rect 675008 384460 675014 384462
rect 675183 384460 675249 384463
rect 675008 384458 675249 384460
rect 675008 384402 675188 384458
rect 675244 384402 675249 384458
rect 675008 384400 675249 384402
rect 675008 384398 675014 384400
rect 675183 384397 675249 384400
rect 41538 383871 41598 383986
rect 41538 383866 41649 383871
rect 41538 383810 41588 383866
rect 41644 383810 41649 383866
rect 41538 383808 41649 383810
rect 41583 383805 41649 383808
rect 34434 383279 34494 383542
rect 34434 383274 34545 383279
rect 34434 383218 34484 383274
rect 34540 383218 34545 383274
rect 34434 383216 34545 383218
rect 34479 383213 34545 383216
rect 41775 383128 41841 383131
rect 41568 383126 41841 383128
rect 41568 383070 41780 383126
rect 41836 383070 41841 383126
rect 41568 383068 41841 383070
rect 41775 383065 41841 383068
rect 675759 382980 675825 382983
rect 676666 382980 676672 382982
rect 675759 382978 676672 382980
rect 675759 382922 675764 382978
rect 675820 382922 676672 382978
rect 675759 382920 676672 382922
rect 675759 382917 675825 382920
rect 676666 382918 676672 382920
rect 676736 382918 676742 382982
rect 41538 382391 41598 382506
rect 41538 382386 41649 382391
rect 41538 382330 41588 382386
rect 41644 382330 41649 382386
rect 41538 382328 41649 382330
rect 41583 382325 41649 382328
rect 675322 382326 675328 382390
rect 675392 382388 675398 382390
rect 675471 382388 675537 382391
rect 675392 382386 675537 382388
rect 675392 382330 675476 382386
rect 675532 382330 675537 382386
rect 675392 382328 675537 382330
rect 675392 382326 675398 382328
rect 675471 382325 675537 382328
rect 41775 382018 41841 382021
rect 41568 382016 41841 382018
rect 41568 381960 41780 382016
rect 41836 381960 41841 382016
rect 41568 381958 41841 381960
rect 41775 381955 41841 381958
rect 675759 381796 675825 381799
rect 676474 381796 676480 381798
rect 675759 381794 676480 381796
rect 675759 381738 675764 381794
rect 675820 381738 676480 381794
rect 675759 381736 676480 381738
rect 675759 381733 675825 381736
rect 676474 381734 676480 381736
rect 676544 381734 676550 381798
rect 39234 381355 39294 381618
rect 39183 381350 39294 381355
rect 39183 381294 39188 381350
rect 39244 381294 39294 381350
rect 39183 381292 39294 381294
rect 39183 381289 39249 381292
rect 675759 381206 675825 381207
rect 675706 381142 675712 381206
rect 675776 381204 675825 381206
rect 675776 381202 675868 381204
rect 675820 381146 675868 381202
rect 675776 381144 675868 381146
rect 675776 381142 675825 381144
rect 675759 381141 675825 381142
rect 39234 380911 39294 381026
rect 39234 380906 39345 380911
rect 39234 380850 39284 380906
rect 39340 380850 39345 380906
rect 39234 380848 39345 380850
rect 39279 380845 39345 380848
rect 39810 380318 39870 380434
rect 39802 380254 39808 380318
rect 39872 380254 39878 380318
rect 40578 379874 40638 380138
rect 40570 379810 40576 379874
rect 40640 379810 40646 379874
rect 39471 379280 39537 379283
rect 40002 379282 40062 379546
rect 39426 379278 39537 379280
rect 39426 379222 39476 379278
rect 39532 379222 39537 379278
rect 39426 379217 39537 379222
rect 39994 379218 40000 379282
rect 40064 379218 40070 379282
rect 39426 378954 39486 379217
rect 34479 378836 34545 378839
rect 42298 378836 42304 378838
rect 34479 378834 42304 378836
rect 34479 378778 34484 378834
rect 34540 378778 42304 378834
rect 34479 378776 42304 378778
rect 34479 378773 34545 378776
rect 42298 378774 42304 378776
rect 42368 378774 42374 378838
rect 674746 378774 674752 378838
rect 674816 378836 674822 378838
rect 675471 378836 675537 378839
rect 674816 378834 675537 378836
rect 674816 378778 675476 378834
rect 675532 378778 675537 378834
rect 674816 378776 675537 378778
rect 674816 378774 674822 378776
rect 675471 378773 675537 378776
rect 40002 378395 40062 378584
rect 40002 378390 40113 378395
rect 40002 378334 40052 378390
rect 40108 378334 40113 378390
rect 40002 378332 40113 378334
rect 40047 378329 40113 378332
rect 675567 378098 675633 378099
rect 39810 377803 39870 378066
rect 675514 378034 675520 378098
rect 675584 378096 675633 378098
rect 675584 378094 675676 378096
rect 675628 378038 675676 378094
rect 675584 378036 675676 378038
rect 675584 378034 675633 378036
rect 675567 378033 675633 378034
rect 39759 377798 39870 377803
rect 39759 377742 39764 377798
rect 39820 377742 39870 377798
rect 39759 377740 39870 377742
rect 39759 377737 39825 377740
rect 40002 377359 40062 377474
rect 39951 377354 40062 377359
rect 39951 377298 39956 377354
rect 40012 377298 40062 377354
rect 39951 377296 40062 377298
rect 39951 377293 40017 377296
rect 674362 377146 674368 377210
rect 674432 377208 674438 377210
rect 675375 377208 675441 377211
rect 674432 377206 675441 377208
rect 674432 377150 675380 377206
rect 675436 377150 675441 377206
rect 674432 377148 675441 377150
rect 674432 377146 674438 377148
rect 675375 377145 675441 377148
rect 41538 376912 41598 377104
rect 42447 376912 42513 376915
rect 41538 376910 42513 376912
rect 41538 376854 42452 376910
rect 42508 376854 42513 376910
rect 41538 376852 42513 376854
rect 42447 376849 42513 376852
rect 675759 376764 675825 376767
rect 676282 376764 676288 376766
rect 675759 376762 676288 376764
rect 675759 376706 675764 376762
rect 675820 376706 676288 376762
rect 675759 376704 676288 376706
rect 675759 376701 675825 376704
rect 676282 376702 676288 376704
rect 676352 376702 676358 376766
rect 41538 376323 41598 376586
rect 41487 376318 41598 376323
rect 41487 376262 41492 376318
rect 41548 376262 41598 376318
rect 41487 376260 41598 376262
rect 41487 376257 41553 376260
rect 41346 375878 41406 375994
rect 41338 375814 41344 375878
rect 41408 375814 41414 375878
rect 675759 375728 675825 375731
rect 676090 375728 676096 375730
rect 675759 375726 676096 375728
rect 675759 375670 675764 375726
rect 675820 375670 676096 375726
rect 675759 375668 676096 375670
rect 675759 375665 675825 375668
rect 676090 375666 676096 375668
rect 676160 375666 676166 375730
rect 41538 375284 41598 375550
rect 41679 375284 41745 375287
rect 41538 375282 41745 375284
rect 41538 375226 41684 375282
rect 41740 375226 41745 375282
rect 41538 375224 41745 375226
rect 41679 375221 41745 375224
rect 41538 374843 41598 375106
rect 41538 374838 41649 374843
rect 41538 374782 41588 374838
rect 41644 374782 41649 374838
rect 41538 374780 41649 374782
rect 41583 374777 41649 374780
rect 41775 374544 41841 374547
rect 41568 374542 41841 374544
rect 41568 374486 41780 374542
rect 41836 374486 41841 374542
rect 41568 374484 41841 374486
rect 41775 374481 41841 374484
rect 655503 374396 655569 374399
rect 649986 374394 655569 374396
rect 649986 374338 655508 374394
rect 655564 374338 655569 374394
rect 649986 374336 655569 374338
rect 28866 373807 28926 374070
rect 40047 373952 40113 373955
rect 40954 373952 40960 373954
rect 40047 373950 40960 373952
rect 40047 373894 40052 373950
rect 40108 373894 40960 373950
rect 40047 373892 40960 373894
rect 40047 373889 40113 373892
rect 40954 373890 40960 373892
rect 41024 373890 41030 373954
rect 649986 373892 650046 374336
rect 655503 374333 655569 374336
rect 673978 373890 673984 373954
rect 674048 373952 674054 373954
rect 675471 373952 675537 373955
rect 674048 373950 675537 373952
rect 674048 373894 675476 373950
rect 675532 373894 675537 373950
rect 674048 373892 675537 373894
rect 674048 373890 674054 373892
rect 675471 373889 675537 373892
rect 28815 373802 28926 373807
rect 28815 373746 28820 373802
rect 28876 373746 28926 373802
rect 28815 373744 28926 373746
rect 39279 373804 39345 373807
rect 41722 373804 41728 373806
rect 39279 373802 41728 373804
rect 39279 373746 39284 373802
rect 39340 373746 41728 373802
rect 39279 373744 41728 373746
rect 28815 373741 28881 373744
rect 39279 373741 39345 373744
rect 41722 373742 41728 373744
rect 41792 373742 41798 373806
rect 41775 373582 41841 373585
rect 41568 373580 41841 373582
rect 41568 373524 41780 373580
rect 41836 373524 41841 373580
rect 41568 373522 41841 373524
rect 41775 373519 41841 373522
rect 28815 373360 28881 373363
rect 39951 373360 40017 373363
rect 41914 373360 41920 373362
rect 28815 373358 28926 373360
rect 28815 373302 28820 373358
rect 28876 373302 28926 373358
rect 28815 373297 28926 373302
rect 39951 373358 41920 373360
rect 39951 373302 39956 373358
rect 40012 373302 41920 373358
rect 39951 373300 41920 373302
rect 39951 373297 40017 373300
rect 41914 373298 41920 373300
rect 41984 373298 41990 373362
rect 655119 373360 655185 373363
rect 649986 373358 655185 373360
rect 649986 373302 655124 373358
rect 655180 373302 655185 373358
rect 649986 373300 655185 373302
rect 28866 373034 28926 373297
rect 39759 373212 39825 373215
rect 42106 373212 42112 373214
rect 39759 373210 42112 373212
rect 39759 373154 39764 373210
rect 39820 373154 42112 373210
rect 39759 373152 42112 373154
rect 39759 373149 39825 373152
rect 42106 373150 42112 373152
rect 42176 373150 42182 373214
rect 649986 372710 650046 373300
rect 655119 373297 655185 373300
rect 39802 372410 39808 372474
rect 39872 372472 39878 372474
rect 42490 372472 42496 372474
rect 39872 372412 42496 372472
rect 39872 372410 39878 372412
rect 42490 372410 42496 372412
rect 42560 372410 42566 372474
rect 39183 372324 39249 372327
rect 40762 372324 40768 372326
rect 39183 372322 40768 372324
rect 39183 372266 39188 372322
rect 39244 372266 40768 372322
rect 39183 372264 40768 372266
rect 39183 372261 39249 372264
rect 40762 372262 40768 372264
rect 40832 372262 40838 372326
rect 655311 372176 655377 372179
rect 649986 372174 655377 372176
rect 649986 372118 655316 372174
rect 655372 372118 655377 372174
rect 649986 372116 655377 372118
rect 649986 371528 650046 372116
rect 655311 372113 655377 372116
rect 656559 370992 656625 370995
rect 649986 370990 656625 370992
rect 649986 370934 656564 370990
rect 656620 370934 656625 370990
rect 649986 370932 656625 370934
rect 649986 370346 650046 370932
rect 656559 370929 656625 370932
rect 41775 368182 41841 368183
rect 41722 368180 41728 368182
rect 41684 368120 41728 368180
rect 41792 368178 41841 368182
rect 41836 368122 41841 368178
rect 41722 368118 41728 368120
rect 41792 368118 41841 368122
rect 41775 368117 41841 368118
rect 40378 362790 40384 362854
rect 40448 362852 40454 362854
rect 41775 362852 41841 362855
rect 40448 362850 41841 362852
rect 40448 362794 41780 362850
rect 41836 362794 41841 362850
rect 40448 362792 41841 362794
rect 40448 362790 40454 362792
rect 41775 362789 41841 362792
rect 59247 360928 59313 360931
rect 59247 360926 64638 360928
rect 59247 360870 59252 360926
rect 59308 360870 64638 360926
rect 59247 360868 64638 360870
rect 59247 360865 59313 360868
rect 41338 360570 41344 360634
rect 41408 360632 41414 360634
rect 41775 360632 41841 360635
rect 41408 360630 41841 360632
rect 41408 360574 41780 360630
rect 41836 360574 41841 360630
rect 41408 360572 41841 360574
rect 41408 360570 41414 360572
rect 41775 360569 41841 360572
rect 64578 360328 64638 360868
rect 41967 359894 42033 359895
rect 41914 359892 41920 359894
rect 41876 359832 41920 359892
rect 41984 359890 42033 359894
rect 42028 359834 42033 359890
rect 41914 359830 41920 359832
rect 41984 359830 42033 359834
rect 41967 359829 42033 359830
rect 59151 359744 59217 359747
rect 59151 359742 64638 359744
rect 59151 359686 59156 359742
rect 59212 359686 64638 359742
rect 59151 359684 64638 359686
rect 59151 359681 59217 359684
rect 42063 359302 42129 359303
rect 42063 359298 42112 359302
rect 42176 359300 42182 359302
rect 42063 359242 42068 359298
rect 42063 359238 42112 359242
rect 42176 359240 42220 359300
rect 42176 359238 42182 359240
rect 42063 359237 42129 359238
rect 64578 359146 64638 359684
rect 40570 358794 40576 358858
rect 40640 358856 40646 358858
rect 41775 358856 41841 358859
rect 40640 358854 41841 358856
rect 40640 358798 41780 358854
rect 41836 358798 41841 358854
rect 40640 358796 41841 358798
rect 40640 358794 40646 358796
rect 41775 358793 41841 358796
rect 676290 358119 676350 358234
rect 676290 358114 676401 358119
rect 676290 358058 676340 358114
rect 676396 358058 676401 358114
rect 676290 358056 676401 358058
rect 676335 358053 676401 358056
rect 57615 357524 57681 357527
rect 64578 357524 64638 357964
rect 57615 357522 64638 357524
rect 57615 357466 57620 357522
rect 57676 357466 64638 357522
rect 57615 357464 64638 357466
rect 676143 357524 676209 357527
rect 676290 357524 676350 357716
rect 676143 357522 676350 357524
rect 676143 357466 676148 357522
rect 676204 357466 676350 357522
rect 676143 357464 676350 357466
rect 57615 357461 57681 357464
rect 676143 357461 676209 357464
rect 676239 357376 676305 357379
rect 676239 357374 676350 357376
rect 676239 357318 676244 357374
rect 676300 357318 676350 357374
rect 676239 357313 676350 357318
rect 40762 357166 40768 357230
rect 40832 357228 40838 357230
rect 41914 357228 41920 357230
rect 40832 357168 41920 357228
rect 40832 357166 40838 357168
rect 41914 357166 41920 357168
rect 41984 357166 41990 357230
rect 676290 357198 676350 357313
rect 41871 356934 41937 356935
rect 41871 356930 41920 356934
rect 41984 356932 41990 356934
rect 41871 356874 41876 356930
rect 41871 356870 41920 356874
rect 41984 356872 42028 356932
rect 41984 356870 41990 356872
rect 41871 356869 41937 356870
rect 59631 356784 59697 356787
rect 676047 356784 676113 356787
rect 59631 356782 64638 356784
rect 59631 356726 59636 356782
rect 59692 356726 64638 356782
rect 59631 356724 64638 356726
rect 676047 356782 676320 356784
rect 676047 356726 676052 356782
rect 676108 356726 676320 356782
rect 676047 356724 676320 356726
rect 59631 356721 59697 356724
rect 676047 356721 676113 356724
rect 40954 356130 40960 356194
rect 41024 356192 41030 356194
rect 41775 356192 41841 356195
rect 41024 356190 41841 356192
rect 41024 356134 41780 356190
rect 41836 356134 41841 356190
rect 41024 356132 41841 356134
rect 41024 356130 41030 356132
rect 41775 356129 41841 356132
rect 58191 356192 58257 356195
rect 58191 356190 64638 356192
rect 58191 356134 58196 356190
rect 58252 356134 64638 356190
rect 58191 356132 64638 356134
rect 58191 356129 58257 356132
rect 42159 355600 42225 355603
rect 42490 355600 42496 355602
rect 42159 355598 42496 355600
rect 42159 355542 42164 355598
rect 42220 355542 42496 355598
rect 42159 355540 42496 355542
rect 42159 355537 42225 355540
rect 42490 355538 42496 355540
rect 42560 355538 42566 355602
rect 64578 355600 64638 356132
rect 674170 355834 674176 355898
rect 674240 355896 674246 355898
rect 676290 355896 676350 356236
rect 674240 355836 676350 355896
rect 674240 355834 674246 355836
rect 676047 355748 676113 355751
rect 676047 355746 676320 355748
rect 676047 355690 676052 355746
rect 676108 355690 676320 355746
rect 676047 355688 676320 355690
rect 676047 355685 676113 355688
rect 673978 355242 673984 355306
rect 674048 355304 674054 355306
rect 674048 355244 676320 355304
rect 674048 355242 674054 355244
rect 58575 355008 58641 355011
rect 58575 355006 64638 355008
rect 58575 354950 58580 355006
rect 58636 354950 64638 355006
rect 58575 354948 64638 354950
rect 58575 354945 58641 354948
rect 64578 354418 64638 354948
rect 676047 354712 676113 354715
rect 676047 354710 676320 354712
rect 676047 354654 676052 354710
rect 676108 354654 676320 354710
rect 676047 354652 676320 354654
rect 676047 354649 676113 354652
rect 674362 354206 674368 354270
rect 674432 354268 674438 354270
rect 674432 354208 676320 354268
rect 674432 354206 674438 354208
rect 675898 353762 675904 353826
rect 675968 353824 675974 353826
rect 675968 353764 676320 353824
rect 675968 353762 675974 353764
rect 674554 353170 674560 353234
rect 674624 353232 674630 353234
rect 674624 353172 676320 353232
rect 674624 353170 674630 353172
rect 675567 352640 675633 352643
rect 676290 352640 676350 352684
rect 675567 352638 676350 352640
rect 675567 352582 675572 352638
rect 675628 352582 676350 352638
rect 675567 352580 676350 352582
rect 675567 352577 675633 352580
rect 676047 352344 676113 352347
rect 676047 352342 676320 352344
rect 676047 352286 676052 352342
rect 676108 352286 676320 352342
rect 676047 352284 676320 352286
rect 676047 352281 676113 352284
rect 674746 351690 674752 351754
rect 674816 351752 674822 351754
rect 674816 351692 676320 351752
rect 674816 351690 674822 351692
rect 676866 351015 676926 351204
rect 676866 351010 676977 351015
rect 676866 350954 676916 351010
rect 676972 350954 676977 351010
rect 676866 350952 676977 350954
rect 676911 350949 676977 350952
rect 676047 350864 676113 350867
rect 676047 350862 676320 350864
rect 676047 350806 676052 350862
rect 676108 350806 676320 350862
rect 676047 350804 676320 350806
rect 676047 350801 676113 350804
rect 676047 350272 676113 350275
rect 676047 350270 676320 350272
rect 676047 350214 676052 350270
rect 676108 350214 676320 350270
rect 676047 350212 676320 350214
rect 676047 350209 676113 350212
rect 676290 349535 676350 349650
rect 676239 349530 676350 349535
rect 676239 349474 676244 349530
rect 676300 349474 676350 349530
rect 676239 349472 676350 349474
rect 676239 349469 676305 349472
rect 676866 349091 676926 349280
rect 676815 349086 676926 349091
rect 676815 349030 676820 349086
rect 676876 349030 676926 349086
rect 676815 349028 676926 349030
rect 676815 349025 676881 349028
rect 674938 348730 674944 348794
rect 675008 348792 675014 348794
rect 675008 348732 676320 348792
rect 675008 348730 675014 348732
rect 676290 348055 676350 348170
rect 676239 348050 676350 348055
rect 676239 347994 676244 348050
rect 676300 347994 676350 348050
rect 676239 347992 676350 347994
rect 676239 347989 676305 347992
rect 676047 347830 676113 347833
rect 676047 347828 676320 347830
rect 676047 347772 676052 347828
rect 676108 347772 676320 347828
rect 676047 347770 676320 347772
rect 676047 347767 676113 347770
rect 675951 347312 676017 347315
rect 675951 347310 676320 347312
rect 675951 347254 675956 347310
rect 676012 347254 676320 347310
rect 675951 347252 676320 347254
rect 675951 347249 676017 347252
rect 679938 346575 679998 346690
rect 679887 346570 679998 346575
rect 679887 346514 679892 346570
rect 679948 346514 679998 346570
rect 679887 346512 679998 346514
rect 679887 346509 679953 346512
rect 679746 345983 679806 346246
rect 679887 346128 679953 346131
rect 679887 346126 679998 346128
rect 679887 346070 679892 346126
rect 679948 346070 679998 346126
rect 679887 346065 679998 346070
rect 679695 345978 679806 345983
rect 679695 345922 679700 345978
rect 679756 345922 679806 345978
rect 679695 345920 679806 345922
rect 679695 345917 679761 345920
rect 679938 345802 679998 346065
rect 679695 345536 679761 345539
rect 679695 345534 679806 345536
rect 679695 345478 679700 345534
rect 679756 345478 679806 345534
rect 679695 345473 679806 345478
rect 679746 345210 679806 345473
rect 41679 343170 41745 343171
rect 41679 343168 41728 343170
rect 41600 343166 41728 343168
rect 41792 343168 41798 343170
rect 62607 343168 62673 343171
rect 41792 343166 62673 343168
rect 41600 343110 41684 343166
rect 41792 343110 62612 343166
rect 62668 343110 62673 343166
rect 41600 343108 41728 343110
rect 41679 343106 41728 343108
rect 41792 343108 62673 343110
rect 41792 343106 41798 343108
rect 41679 343105 41745 343106
rect 62607 343105 62673 343108
rect 675706 342958 675712 343022
rect 675776 343020 675782 343022
rect 676815 343020 676881 343023
rect 675776 343018 676881 343020
rect 675776 342962 676820 343018
rect 676876 342962 676881 343018
rect 675776 342960 676881 342962
rect 675776 342958 675782 342960
rect 676815 342957 676881 342960
rect 41775 342872 41841 342875
rect 41568 342870 41841 342872
rect 41568 342814 41780 342870
rect 41836 342814 41841 342870
rect 41568 342812 41841 342814
rect 41775 342809 41841 342812
rect 676666 342810 676672 342874
rect 676736 342872 676742 342874
rect 676911 342872 676977 342875
rect 676736 342870 676977 342872
rect 676736 342814 676916 342870
rect 676972 342814 676977 342870
rect 676736 342812 676977 342814
rect 676736 342810 676742 342812
rect 676911 342809 676977 342812
rect 41775 342354 41841 342357
rect 41568 342352 41841 342354
rect 41568 342296 41780 342352
rect 41836 342296 41841 342352
rect 41568 342294 41841 342296
rect 41775 342291 41841 342294
rect 41775 341836 41841 341839
rect 41568 341834 41841 341836
rect 41568 341778 41780 341834
rect 41836 341778 41841 341834
rect 41568 341776 41841 341778
rect 41775 341773 41841 341776
rect 41775 341392 41841 341395
rect 41568 341390 41841 341392
rect 41568 341334 41780 341390
rect 41836 341334 41841 341390
rect 41568 341332 41841 341334
rect 41775 341329 41841 341332
rect 41538 340655 41598 340770
rect 41538 340650 41649 340655
rect 41538 340594 41588 340650
rect 41644 340594 41649 340650
rect 41538 340592 41649 340594
rect 41583 340589 41649 340592
rect 41775 340356 41841 340359
rect 41568 340354 41841 340356
rect 41568 340298 41780 340354
rect 41836 340298 41841 340354
rect 41568 340296 41841 340298
rect 41775 340293 41841 340296
rect 41679 340060 41745 340063
rect 41538 340058 41745 340060
rect 41538 340002 41684 340058
rect 41740 340002 41745 340058
rect 41538 340000 41745 340002
rect 41538 339882 41598 340000
rect 41679 339997 41745 340000
rect 675759 339616 675825 339619
rect 675898 339616 675904 339618
rect 675759 339614 675904 339616
rect 675759 339558 675764 339614
rect 675820 339558 675904 339614
rect 675759 339556 675904 339558
rect 675759 339553 675825 339556
rect 675898 339554 675904 339556
rect 675968 339554 675974 339618
rect 41538 339175 41598 339290
rect 41538 339170 41649 339175
rect 41538 339114 41588 339170
rect 41644 339114 41649 339170
rect 41538 339112 41649 339114
rect 41583 339109 41649 339112
rect 41775 338876 41841 338879
rect 41914 338876 41920 338878
rect 41568 338874 41920 338876
rect 41568 338818 41780 338874
rect 41836 338818 41920 338874
rect 41568 338816 41920 338818
rect 41775 338813 41841 338816
rect 41914 338814 41920 338816
rect 41984 338814 41990 338878
rect 28674 338139 28734 338402
rect 28674 338134 28785 338139
rect 28674 338078 28724 338134
rect 28780 338078 28785 338134
rect 28674 338076 28785 338078
rect 28719 338073 28785 338076
rect 39810 337695 39870 337810
rect 39759 337690 39870 337695
rect 39759 337634 39764 337690
rect 39820 337634 39870 337690
rect 39759 337632 39870 337634
rect 39759 337629 39825 337632
rect 39234 337103 39294 337292
rect 39234 337098 39345 337103
rect 39234 337042 39284 337098
rect 39340 337042 39345 337098
rect 39234 337040 39345 337042
rect 39279 337037 39345 337040
rect 40386 336658 40446 336922
rect 40378 336594 40384 336658
rect 40448 336594 40454 336658
rect 40770 336066 40830 336330
rect 40762 336002 40768 336066
rect 40832 336002 40838 336066
rect 41775 335768 41841 335771
rect 41568 335766 41841 335768
rect 41568 335710 41780 335766
rect 41836 335710 41841 335766
rect 41568 335708 41841 335710
rect 41775 335705 41841 335708
rect 40962 335178 41022 335442
rect 40954 335114 40960 335178
rect 41024 335114 41030 335178
rect 41346 334586 41406 334850
rect 41338 334522 41344 334586
rect 41408 334522 41414 334586
rect 41154 334142 41214 334258
rect 41146 334078 41152 334142
rect 41216 334078 41222 334142
rect 41538 333699 41598 333888
rect 41487 333694 41598 333699
rect 41487 333638 41492 333694
rect 41548 333638 41598 333694
rect 41487 333636 41598 333638
rect 41487 333633 41553 333636
rect 674746 333486 674752 333550
rect 674816 333548 674822 333550
rect 675375 333548 675441 333551
rect 674816 333546 675441 333548
rect 674816 333490 675380 333546
rect 675436 333490 675441 333546
rect 674816 333488 675441 333490
rect 674816 333486 674822 333488
rect 675375 333485 675441 333488
rect 41346 333107 41406 333370
rect 41346 333102 41457 333107
rect 41346 333046 41396 333102
rect 41452 333046 41457 333102
rect 41346 333044 41457 333046
rect 41391 333041 41457 333044
rect 41538 332662 41598 332778
rect 41530 332598 41536 332662
rect 41600 332598 41606 332662
rect 40578 332070 40638 332408
rect 674938 332302 674944 332366
rect 675008 332364 675014 332366
rect 675471 332364 675537 332367
rect 675008 332362 675537 332364
rect 675008 332306 675476 332362
rect 675532 332306 675537 332362
rect 675008 332304 675537 332306
rect 675008 332302 675014 332304
rect 675471 332301 675537 332304
rect 40570 332006 40576 332070
rect 40640 332006 40646 332070
rect 41538 331627 41598 331890
rect 41538 331622 41649 331627
rect 41538 331566 41588 331622
rect 41644 331566 41649 331622
rect 41538 331564 41649 331566
rect 41583 331561 41649 331564
rect 41871 331328 41937 331331
rect 41568 331326 41937 331328
rect 41568 331270 41876 331326
rect 41932 331270 41937 331326
rect 41568 331268 41937 331270
rect 41871 331265 41937 331268
rect 39759 331180 39825 331183
rect 41722 331180 41728 331182
rect 39759 331178 41728 331180
rect 39759 331122 39764 331178
rect 39820 331122 41728 331178
rect 39759 331120 41728 331122
rect 39759 331117 39825 331120
rect 41722 331118 41728 331120
rect 41792 331118 41798 331182
rect 28866 330591 28926 330854
rect 39279 330736 39345 330739
rect 42298 330736 42304 330738
rect 39279 330734 42304 330736
rect 39279 330678 39284 330734
rect 39340 330678 42304 330734
rect 39279 330676 42304 330678
rect 39279 330673 39345 330676
rect 42298 330674 42304 330676
rect 42368 330674 42374 330738
rect 28815 330586 28926 330591
rect 675759 330590 675825 330591
rect 28815 330530 28820 330586
rect 28876 330530 28926 330586
rect 28815 330528 28926 330530
rect 28815 330525 28881 330528
rect 675706 330526 675712 330590
rect 675776 330588 675825 330590
rect 675776 330586 675868 330588
rect 675820 330530 675868 330586
rect 675776 330528 675868 330530
rect 675776 330526 675825 330528
rect 675759 330525 675825 330526
rect 41871 330440 41937 330443
rect 41568 330438 41937 330440
rect 41568 330382 41876 330438
rect 41932 330382 41937 330438
rect 41568 330380 41937 330382
rect 41871 330377 41937 330380
rect 28815 330144 28881 330147
rect 28815 330142 28926 330144
rect 28815 330086 28820 330142
rect 28876 330086 28926 330142
rect 28815 330081 28926 330086
rect 28866 329818 28926 330081
rect 655215 329848 655281 329851
rect 649986 329846 655281 329848
rect 649986 329790 655220 329846
rect 655276 329790 655281 329846
rect 649986 329788 655281 329790
rect 649986 329234 650046 329788
rect 655215 329785 655281 329788
rect 28719 329108 28785 329111
rect 42106 329108 42112 329110
rect 28719 329106 42112 329108
rect 28719 329050 28724 329106
rect 28780 329050 42112 329106
rect 28719 329048 42112 329050
rect 28719 329045 28785 329048
rect 42106 329046 42112 329048
rect 42176 329046 42182 329110
rect 674554 328306 674560 328370
rect 674624 328368 674630 328370
rect 675375 328368 675441 328371
rect 674624 328366 675441 328368
rect 674624 328310 675380 328366
rect 675436 328310 675441 328366
rect 674624 328308 675441 328310
rect 674624 328306 674630 328308
rect 675375 328305 675441 328308
rect 655119 328072 655185 328075
rect 649986 328070 655185 328072
rect 649986 328014 655124 328070
rect 655180 328014 655185 328070
rect 649986 328012 655185 328014
rect 655119 328009 655185 328012
rect 655311 327480 655377 327483
rect 649986 327478 655377 327480
rect 649986 327422 655316 327478
rect 655372 327422 655377 327478
rect 649986 327420 655377 327422
rect 649986 326870 650046 327420
rect 655311 327417 655377 327420
rect 675759 326888 675825 326891
rect 676666 326888 676672 326890
rect 675759 326886 676672 326888
rect 675759 326830 675764 326886
rect 675820 326830 676672 326886
rect 675759 326828 676672 326830
rect 675759 326825 675825 326828
rect 676666 326826 676672 326828
rect 676736 326826 676742 326890
rect 654159 326296 654225 326299
rect 649986 326294 654225 326296
rect 649986 326238 654164 326294
rect 654220 326238 654225 326294
rect 649986 326236 654225 326238
rect 649986 325688 650046 326236
rect 654159 326233 654225 326236
rect 41775 324966 41841 324967
rect 41722 324964 41728 324966
rect 41684 324904 41728 324964
rect 41792 324962 41841 324966
rect 41836 324906 41841 324962
rect 41722 324902 41728 324904
rect 41792 324902 41841 324906
rect 41775 324901 41841 324902
rect 40570 320462 40576 320526
rect 40640 320524 40646 320526
rect 41775 320524 41841 320527
rect 40640 320522 41841 320524
rect 40640 320466 41780 320522
rect 41836 320466 41841 320522
rect 40640 320464 41841 320466
rect 40640 320462 40646 320464
rect 41775 320461 41841 320464
rect 40762 319722 40768 319786
rect 40832 319784 40838 319786
rect 41775 319784 41841 319787
rect 40832 319782 41841 319784
rect 40832 319726 41780 319782
rect 41836 319726 41841 319782
rect 40832 319724 41841 319726
rect 40832 319722 40838 319724
rect 41775 319721 41841 319724
rect 58479 317712 58545 317715
rect 58479 317710 64638 317712
rect 58479 317654 58484 317710
rect 58540 317654 64638 317710
rect 58479 317652 64638 317654
rect 58479 317649 58545 317652
rect 41530 317354 41536 317418
rect 41600 317416 41606 317418
rect 41871 317416 41937 317419
rect 41600 317414 41937 317416
rect 41600 317358 41876 317414
rect 41932 317358 41937 317414
rect 41600 317356 41937 317358
rect 41600 317354 41606 317356
rect 41871 317353 41937 317356
rect 64578 317106 64638 317652
rect 41146 316614 41152 316678
rect 41216 316676 41222 316678
rect 41775 316676 41841 316679
rect 41216 316674 41841 316676
rect 41216 316618 41780 316674
rect 41836 316618 41841 316674
rect 41216 316616 41841 316618
rect 41216 316614 41222 316616
rect 41775 316613 41841 316616
rect 59151 316528 59217 316531
rect 59151 316526 64638 316528
rect 59151 316470 59156 316526
rect 59212 316470 64638 316526
rect 59151 316468 64638 316470
rect 59151 316465 59217 316468
rect 41338 316170 41344 316234
rect 41408 316232 41414 316234
rect 41775 316232 41841 316235
rect 41408 316230 41841 316232
rect 41408 316174 41780 316230
rect 41836 316174 41841 316230
rect 41408 316172 41841 316174
rect 41408 316170 41414 316172
rect 41775 316169 41841 316172
rect 64578 315924 64638 316468
rect 40378 315430 40384 315494
rect 40448 315492 40454 315494
rect 41775 315492 41841 315495
rect 40448 315490 41841 315492
rect 40448 315434 41780 315490
rect 41836 315434 41841 315490
rect 40448 315432 41841 315434
rect 40448 315430 40454 315432
rect 41775 315429 41841 315432
rect 59343 314160 59409 314163
rect 64578 314160 64638 314742
rect 59343 314158 64638 314160
rect 59343 314102 59348 314158
rect 59404 314102 64638 314158
rect 59343 314100 64638 314102
rect 59343 314097 59409 314100
rect 42063 313718 42129 313719
rect 42063 313714 42112 313718
rect 42176 313716 42182 313718
rect 42063 313658 42068 313714
rect 42063 313654 42112 313658
rect 42176 313656 42220 313716
rect 42176 313654 42182 313656
rect 42063 313653 42129 313654
rect 59631 313568 59697 313571
rect 59631 313566 64638 313568
rect 59631 313510 59636 313566
rect 59692 313510 64638 313566
rect 59631 313508 64638 313510
rect 59631 313505 59697 313508
rect 40954 313062 40960 313126
rect 41024 313124 41030 313126
rect 41775 313124 41841 313127
rect 41024 313122 41841 313124
rect 41024 313066 41780 313122
rect 41836 313066 41841 313122
rect 41024 313064 41841 313066
rect 41024 313062 41030 313064
rect 41775 313061 41841 313064
rect 58191 312976 58257 312979
rect 58191 312974 64638 312976
rect 58191 312918 58196 312974
rect 58252 312918 64638 312974
rect 58191 312916 64638 312918
rect 58191 312913 58257 312916
rect 42159 312532 42225 312535
rect 42298 312532 42304 312534
rect 42159 312530 42304 312532
rect 42159 312474 42164 312530
rect 42220 312474 42304 312530
rect 42159 312472 42304 312474
rect 42159 312469 42225 312472
rect 42298 312470 42304 312472
rect 42368 312470 42374 312534
rect 64578 312378 64638 312916
rect 676290 312239 676350 312502
rect 676290 312234 676401 312239
rect 676290 312178 676340 312234
rect 676396 312178 676401 312234
rect 676290 312176 676401 312178
rect 676335 312173 676401 312176
rect 59727 311792 59793 311795
rect 59727 311790 64638 311792
rect 59727 311734 59732 311790
rect 59788 311734 64638 311790
rect 59727 311732 64638 311734
rect 59727 311729 59793 311732
rect 64578 311196 64638 311732
rect 676143 311644 676209 311647
rect 676290 311644 676350 311910
rect 676143 311642 676350 311644
rect 676143 311586 676148 311642
rect 676204 311586 676350 311642
rect 676143 311584 676350 311586
rect 676143 311581 676209 311584
rect 676290 311203 676350 311392
rect 676239 311198 676350 311203
rect 676239 311142 676244 311198
rect 676300 311142 676350 311198
rect 676239 311140 676350 311142
rect 676239 311137 676305 311140
rect 674170 310990 674176 311054
rect 674240 311052 674246 311054
rect 674240 310992 676320 311052
rect 674240 310990 674246 310992
rect 675514 310398 675520 310462
rect 675584 310460 675590 310462
rect 675584 310400 676320 310460
rect 675584 310398 675590 310400
rect 674170 309806 674176 309870
rect 674240 309868 674246 309870
rect 674240 309808 676320 309868
rect 674240 309806 674246 309808
rect 674554 309066 674560 309130
rect 674624 309128 674630 309130
rect 676290 309128 676350 309468
rect 674624 309068 676350 309128
rect 674624 309066 674630 309068
rect 674362 308918 674368 308982
rect 674432 308980 674438 308982
rect 674432 308920 676320 308980
rect 674432 308918 674438 308920
rect 674746 308326 674752 308390
rect 674816 308388 674822 308390
rect 674816 308328 676320 308388
rect 674816 308326 674822 308328
rect 676047 308018 676113 308021
rect 676047 308016 676320 308018
rect 676047 307960 676052 308016
rect 676108 307960 676320 308016
rect 676047 307958 676320 307960
rect 676047 307955 676113 307958
rect 676866 307207 676926 307470
rect 676815 307202 676926 307207
rect 676815 307146 676820 307202
rect 676876 307146 676926 307202
rect 676815 307144 676926 307146
rect 676815 307141 676881 307144
rect 676290 306763 676350 306878
rect 676239 306758 676350 306763
rect 676239 306702 676244 306758
rect 676300 306702 676350 306758
rect 676239 306700 676350 306702
rect 676239 306697 676305 306700
rect 675706 306402 675712 306466
rect 675776 306464 675782 306466
rect 675776 306404 676320 306464
rect 675776 306402 675782 306404
rect 675322 305958 675328 306022
rect 675392 306020 675398 306022
rect 675392 305960 676320 306020
rect 675392 305958 675398 305960
rect 674938 305366 674944 305430
rect 675008 305428 675014 305430
rect 675008 305368 676320 305428
rect 675008 305366 675014 305368
rect 676290 304839 676350 304954
rect 676239 304834 676350 304839
rect 676239 304778 676244 304834
rect 676300 304778 676350 304834
rect 676239 304776 676350 304778
rect 676239 304773 676305 304776
rect 676047 304466 676113 304469
rect 676047 304464 676320 304466
rect 676047 304408 676052 304464
rect 676108 304408 676320 304464
rect 676047 304406 676320 304408
rect 676047 304403 676113 304406
rect 675951 303948 676017 303951
rect 675951 303946 676320 303948
rect 675951 303890 675956 303946
rect 676012 303890 676320 303946
rect 675951 303888 676320 303890
rect 675951 303885 676017 303888
rect 675130 303442 675136 303506
rect 675200 303504 675206 303506
rect 675200 303444 676320 303504
rect 675200 303442 675206 303444
rect 654159 303356 654225 303359
rect 649986 303354 654225 303356
rect 649986 303298 654164 303354
rect 654220 303298 654225 303354
rect 649986 303296 654225 303298
rect 649986 302776 650046 303296
rect 654159 303293 654225 303296
rect 673978 302554 673984 302618
rect 674048 302616 674054 302618
rect 676290 302616 676350 302956
rect 674048 302556 676350 302616
rect 674048 302554 674054 302556
rect 675898 302406 675904 302470
rect 675968 302468 675974 302470
rect 675968 302408 676320 302468
rect 675968 302406 675974 302408
rect 654063 302172 654129 302175
rect 649986 302170 654129 302172
rect 649986 302114 654068 302170
rect 654124 302114 654129 302170
rect 649986 302112 654129 302114
rect 649986 301594 650046 302112
rect 654063 302109 654129 302112
rect 676047 302024 676113 302027
rect 676047 302022 676320 302024
rect 676047 301966 676052 302022
rect 676108 301966 676320 302022
rect 676047 301964 676320 301966
rect 676047 301961 676113 301964
rect 676290 301287 676350 301402
rect 676239 301282 676350 301287
rect 676239 301226 676244 301282
rect 676300 301226 676350 301282
rect 676239 301224 676350 301226
rect 676239 301221 676305 301224
rect 654255 300988 654321 300991
rect 649986 300986 654321 300988
rect 649986 300930 654260 300986
rect 654316 300930 654321 300986
rect 649986 300928 654321 300930
rect 649986 300412 650046 300928
rect 654255 300925 654321 300928
rect 679938 300695 679998 300958
rect 679938 300690 680049 300695
rect 679938 300634 679988 300690
rect 680044 300634 680049 300690
rect 679938 300632 680049 300634
rect 679983 300629 680049 300632
rect 679746 300251 679806 300514
rect 679746 300246 679857 300251
rect 679983 300248 680049 300251
rect 679746 300190 679796 300246
rect 679852 300190 679857 300246
rect 679746 300188 679857 300190
rect 679791 300185 679857 300188
rect 679938 300246 680049 300248
rect 679938 300190 679988 300246
rect 680044 300190 680049 300246
rect 679938 300185 680049 300190
rect 679938 299922 679998 300185
rect 679791 299804 679857 299807
rect 679746 299802 679857 299804
rect 679746 299746 679796 299802
rect 679852 299746 679857 299802
rect 679746 299741 679857 299746
rect 41775 299656 41841 299659
rect 41568 299654 41841 299656
rect 41568 299598 41780 299654
rect 41836 299598 41841 299654
rect 41568 299596 41841 299598
rect 41775 299593 41841 299596
rect 679746 299404 679806 299741
rect 41775 299212 41841 299215
rect 41568 299210 41841 299212
rect 41568 299154 41780 299210
rect 41836 299154 41841 299210
rect 41568 299152 41841 299154
rect 41775 299149 41841 299152
rect 39663 298768 39729 298771
rect 39618 298766 39729 298768
rect 39618 298710 39668 298766
rect 39724 298710 39729 298766
rect 39618 298705 39729 298710
rect 649986 298768 650046 299230
rect 676090 299150 676096 299214
rect 676160 299212 676166 299214
rect 676815 299212 676881 299215
rect 676160 299210 676881 299212
rect 676160 299154 676820 299210
rect 676876 299154 676881 299210
rect 676160 299152 676881 299154
rect 676160 299150 676166 299152
rect 676815 299149 676881 299152
rect 656559 298768 656625 298771
rect 649986 298766 656625 298768
rect 649986 298710 656564 298766
rect 656620 298710 656625 298766
rect 649986 298708 656625 298710
rect 656559 298705 656625 298708
rect 39618 298590 39678 298705
rect 41775 298176 41841 298179
rect 41568 298174 41841 298176
rect 41568 298118 41780 298174
rect 41836 298118 41841 298174
rect 41568 298116 41841 298118
rect 41775 298113 41841 298116
rect 41775 297658 41841 297661
rect 41568 297656 41841 297658
rect 41568 297600 41780 297656
rect 41836 297600 41841 297656
rect 41568 297598 41841 297600
rect 41775 297595 41841 297598
rect 649986 297584 650046 298048
rect 656079 297584 656145 297587
rect 649986 297582 656145 297584
rect 649986 297526 656084 297582
rect 656140 297526 656145 297582
rect 649986 297524 656145 297526
rect 656079 297521 656145 297524
rect 41775 297140 41841 297143
rect 41568 297138 41841 297140
rect 41568 297082 41780 297138
rect 41836 297082 41841 297138
rect 41568 297080 41841 297082
rect 41775 297077 41841 297080
rect 649986 296844 650046 296866
rect 656271 296844 656337 296847
rect 649986 296842 656337 296844
rect 649986 296786 656276 296842
rect 656332 296786 656337 296842
rect 649986 296784 656337 296786
rect 656271 296781 656337 296784
rect 39810 296551 39870 296670
rect 39759 296546 39870 296551
rect 39759 296490 39764 296546
rect 39820 296490 39870 296546
rect 39759 296488 39870 296490
rect 39759 296485 39825 296488
rect 41538 295959 41598 296074
rect 39951 295956 40017 295959
rect 39951 295954 40062 295956
rect 39951 295898 39956 295954
rect 40012 295898 40062 295954
rect 39951 295893 40062 295898
rect 41538 295954 41649 295959
rect 41538 295898 41588 295954
rect 41644 295898 41649 295954
rect 41538 295896 41649 295898
rect 41583 295893 41649 295896
rect 40002 295630 40062 295893
rect 59631 295216 59697 295219
rect 64578 295216 64638 295684
rect 59631 295214 64638 295216
rect 28674 294923 28734 295186
rect 59631 295158 59636 295214
rect 59692 295158 64638 295214
rect 59631 295156 64638 295158
rect 649986 295216 650046 295684
rect 656367 295216 656433 295219
rect 649986 295214 656433 295216
rect 649986 295158 656372 295214
rect 656428 295158 656433 295214
rect 649986 295156 656433 295158
rect 59631 295153 59697 295156
rect 656367 295153 656433 295156
rect 28674 294918 28785 294923
rect 28674 294862 28724 294918
rect 28780 294862 28785 294918
rect 28674 294860 28785 294862
rect 28719 294857 28785 294860
rect 41722 294624 41728 294626
rect 41568 294564 41728 294624
rect 41722 294562 41728 294564
rect 41792 294562 41798 294626
rect 41914 294180 41920 294182
rect 41568 294120 41920 294180
rect 41914 294118 41920 294120
rect 41984 294118 41990 294182
rect 60303 294032 60369 294035
rect 64578 294032 64638 294502
rect 60303 294030 64638 294032
rect 60303 293974 60308 294030
rect 60364 293974 64638 294030
rect 60303 293972 64638 293974
rect 649986 294032 650046 294502
rect 655887 294032 655953 294035
rect 649986 294030 655953 294032
rect 649986 293974 655892 294030
rect 655948 293974 655953 294030
rect 649986 293972 655953 293974
rect 60303 293969 60369 293972
rect 655887 293969 655953 293972
rect 41154 293442 41214 293706
rect 41146 293378 41152 293442
rect 41216 293378 41222 293442
rect 41538 292998 41598 293114
rect 41530 292934 41536 292998
rect 41600 292934 41606 292998
rect 58383 292848 58449 292851
rect 64578 292848 64638 293320
rect 58383 292846 64638 292848
rect 58383 292790 58388 292846
rect 58444 292790 64638 292846
rect 58383 292788 64638 292790
rect 649986 292848 650046 293320
rect 655791 292848 655857 292851
rect 649986 292846 655857 292848
rect 649986 292790 655796 292846
rect 655852 292790 655857 292846
rect 649986 292788 655857 292790
rect 58383 292785 58449 292788
rect 655791 292785 655857 292788
rect 675663 292850 675729 292851
rect 675663 292846 675712 292850
rect 675776 292848 675782 292850
rect 675663 292790 675668 292846
rect 675663 292786 675712 292790
rect 675776 292788 675820 292848
rect 675776 292786 675782 292788
rect 675663 292785 675729 292786
rect 58767 292700 58833 292703
rect 58767 292698 64638 292700
rect 58767 292642 58772 292698
rect 58828 292642 64638 292698
rect 58767 292640 64638 292642
rect 58767 292637 58833 292640
rect 41775 292626 41841 292629
rect 41568 292624 41841 292626
rect 41568 292568 41780 292624
rect 41836 292568 41841 292624
rect 41568 292566 41841 292568
rect 41775 292563 41841 292566
rect 40386 291962 40446 292226
rect 64578 292138 64638 292640
rect 40378 291898 40384 291962
rect 40448 291898 40454 291962
rect 649986 291664 650046 292138
rect 656175 291664 656241 291667
rect 649986 291662 656241 291664
rect 40962 291518 41022 291634
rect 649986 291606 656180 291662
rect 656236 291606 656241 291662
rect 649986 291604 656241 291606
rect 656175 291601 656241 291604
rect 40954 291454 40960 291518
rect 41024 291454 41030 291518
rect 60207 291516 60273 291519
rect 60207 291514 64638 291516
rect 60207 291458 60212 291514
rect 60268 291458 64638 291514
rect 60207 291456 64638 291458
rect 60207 291453 60273 291456
rect 41346 290926 41406 291042
rect 64578 290956 64638 291456
rect 41338 290862 41344 290926
rect 41408 290862 41414 290926
rect 649986 290924 650046 290956
rect 655983 290924 656049 290927
rect 649986 290922 656049 290924
rect 649986 290866 655988 290922
rect 656044 290866 656049 290922
rect 649986 290864 656049 290866
rect 655983 290861 656049 290864
rect 675759 290776 675825 290779
rect 675898 290776 675904 290778
rect 675759 290774 675904 290776
rect 41538 290483 41598 290746
rect 675759 290718 675764 290774
rect 675820 290718 675904 290774
rect 675759 290716 675904 290718
rect 675759 290713 675825 290716
rect 675898 290714 675904 290716
rect 675968 290714 675974 290778
rect 41487 290478 41598 290483
rect 41487 290422 41492 290478
rect 41548 290422 41598 290478
rect 41487 290420 41598 290422
rect 41487 290417 41553 290420
rect 42447 290184 42513 290187
rect 41568 290182 42513 290184
rect 41568 290126 42452 290182
rect 42508 290126 42513 290182
rect 41568 290124 42513 290126
rect 42447 290121 42513 290124
rect 57999 289592 58065 289595
rect 64578 289592 64638 289774
rect 57999 289590 64638 289592
rect 40578 289446 40638 289562
rect 57999 289534 58004 289590
rect 58060 289534 64638 289590
rect 57999 289532 64638 289534
rect 57999 289529 58065 289532
rect 40570 289382 40576 289446
rect 40640 289382 40646 289446
rect 649986 289296 650046 289774
rect 655599 289296 655665 289299
rect 649986 289294 655665 289296
rect 649986 289238 655604 289294
rect 655660 289238 655665 289294
rect 649986 289236 655665 289238
rect 655599 289233 655665 289236
rect 41538 288852 41598 289192
rect 41679 288852 41745 288855
rect 41538 288850 41745 288852
rect 41538 288794 41684 288850
rect 41740 288794 41745 288850
rect 41538 288792 41745 288794
rect 41679 288789 41745 288792
rect 41538 288411 41598 288674
rect 41538 288406 41649 288411
rect 41538 288350 41588 288406
rect 41644 288350 41649 288406
rect 41538 288348 41649 288350
rect 41583 288345 41649 288348
rect 59631 288112 59697 288115
rect 64578 288112 64638 288592
rect 59631 288110 64638 288112
rect 41538 287964 41598 288082
rect 59631 288054 59636 288110
rect 59692 288054 64638 288110
rect 59631 288052 64638 288054
rect 649986 288112 650046 288592
rect 675322 288494 675328 288558
rect 675392 288556 675398 288558
rect 675471 288556 675537 288559
rect 675392 288554 675537 288556
rect 675392 288498 675476 288554
rect 675532 288498 675537 288554
rect 675392 288496 675537 288498
rect 675392 288494 675398 288496
rect 675471 288493 675537 288496
rect 655407 288112 655473 288115
rect 649986 288110 655473 288112
rect 649986 288054 655412 288110
rect 655468 288054 655473 288110
rect 649986 288052 655473 288054
rect 59631 288049 59697 288052
rect 655407 288049 655473 288052
rect 41538 287904 41790 287964
rect 28866 287375 28926 287712
rect 41730 287520 41790 287904
rect 28815 287370 28926 287375
rect 28815 287314 28820 287370
rect 28876 287314 28926 287370
rect 28815 287312 28926 287314
rect 41538 287460 41790 287520
rect 28815 287309 28881 287312
rect 41538 287224 41598 287460
rect 41871 287224 41937 287227
rect 41538 287222 41937 287224
rect 41538 287194 41876 287222
rect 41568 287166 41876 287194
rect 41932 287166 41937 287222
rect 41568 287164 41937 287166
rect 41871 287161 41937 287164
rect 28815 286928 28881 286931
rect 58959 286928 59025 286931
rect 64578 286928 64638 287410
rect 28815 286926 28926 286928
rect 28815 286870 28820 286926
rect 28876 286870 28926 286926
rect 28815 286865 28926 286870
rect 58959 286926 64638 286928
rect 58959 286870 58964 286926
rect 59020 286870 64638 286926
rect 58959 286868 64638 286870
rect 649986 286928 650046 287410
rect 673978 287162 673984 287226
rect 674048 287224 674054 287226
rect 675471 287224 675537 287227
rect 674048 287222 675537 287224
rect 674048 287166 675476 287222
rect 675532 287166 675537 287222
rect 674048 287164 675537 287166
rect 674048 287162 674054 287164
rect 675471 287161 675537 287164
rect 655503 286928 655569 286931
rect 649986 286926 655569 286928
rect 649986 286870 655508 286926
rect 655564 286870 655569 286926
rect 649986 286868 655569 286870
rect 58959 286865 59025 286868
rect 655503 286865 655569 286868
rect 28866 286602 28926 286865
rect 59055 285744 59121 285747
rect 64578 285744 64638 286228
rect 59055 285742 64638 285744
rect 59055 285686 59060 285742
rect 59116 285686 64638 285742
rect 59055 285684 64638 285686
rect 649986 285744 650046 286228
rect 655695 285744 655761 285747
rect 649986 285742 655761 285744
rect 649986 285686 655700 285742
rect 655756 285686 655761 285742
rect 649986 285684 655761 285686
rect 59055 285681 59121 285684
rect 655695 285681 655761 285684
rect 675130 285238 675136 285302
rect 675200 285300 675206 285302
rect 675471 285300 675537 285303
rect 675200 285298 675537 285300
rect 675200 285242 675476 285298
rect 675532 285242 675537 285298
rect 675200 285240 675537 285242
rect 675200 285238 675206 285240
rect 675471 285237 675537 285240
rect 28719 285152 28785 285155
rect 42106 285152 42112 285154
rect 28719 285150 42112 285152
rect 28719 285094 28724 285150
rect 28780 285094 42112 285150
rect 28719 285092 42112 285094
rect 28719 285089 28785 285092
rect 42106 285090 42112 285092
rect 42176 285090 42182 285154
rect 57615 284560 57681 284563
rect 64578 284560 64638 285046
rect 57615 284558 64638 284560
rect 57615 284502 57620 284558
rect 57676 284502 64638 284558
rect 57615 284500 64638 284502
rect 649986 284560 650046 285046
rect 653775 284560 653841 284563
rect 649986 284558 653841 284560
rect 649986 284502 653780 284558
rect 653836 284502 653841 284558
rect 649986 284500 653841 284502
rect 57615 284497 57681 284500
rect 653775 284497 653841 284500
rect 59631 283376 59697 283379
rect 64578 283376 64638 283864
rect 59631 283374 64638 283376
rect 59631 283318 59636 283374
rect 59692 283318 64638 283374
rect 59631 283316 64638 283318
rect 649986 283376 650046 283864
rect 675759 283672 675825 283675
rect 676090 283672 676096 283674
rect 675759 283670 676096 283672
rect 675759 283614 675764 283670
rect 675820 283614 676096 283670
rect 675759 283612 676096 283614
rect 675759 283609 675825 283612
rect 676090 283610 676096 283612
rect 676160 283610 676166 283674
rect 655119 283376 655185 283379
rect 649986 283374 655185 283376
rect 649986 283318 655124 283374
rect 655180 283318 655185 283374
rect 649986 283316 655185 283318
rect 59631 283313 59697 283316
rect 655119 283313 655185 283316
rect 58959 282488 59025 282491
rect 64578 282488 64638 282682
rect 58959 282486 64638 282488
rect 58959 282430 58964 282486
rect 59020 282430 64638 282486
rect 58959 282428 64638 282430
rect 58959 282425 59025 282428
rect 649986 282340 650046 282682
rect 655311 282340 655377 282343
rect 649986 282338 655377 282340
rect 649986 282282 655316 282338
rect 655372 282282 655377 282338
rect 649986 282280 655377 282282
rect 655311 282277 655377 282280
rect 674938 281834 674944 281898
rect 675008 281896 675014 281898
rect 675375 281896 675441 281899
rect 675008 281894 675441 281896
rect 675008 281838 675380 281894
rect 675436 281838 675441 281894
rect 675008 281836 675441 281838
rect 675008 281834 675014 281836
rect 675375 281833 675441 281836
rect 41722 281686 41728 281750
rect 41792 281748 41798 281750
rect 41871 281748 41937 281751
rect 41792 281746 41937 281748
rect 41792 281690 41876 281746
rect 41932 281690 41937 281746
rect 41792 281688 41937 281690
rect 41792 281686 41798 281688
rect 41871 281685 41937 281688
rect 42447 281602 42513 281603
rect 42447 281598 42496 281602
rect 42560 281600 42566 281602
rect 42447 281542 42452 281598
rect 42447 281538 42496 281542
rect 42560 281540 42604 281600
rect 42560 281538 42566 281540
rect 42447 281537 42513 281538
rect 59535 281008 59601 281011
rect 64578 281008 64638 281500
rect 59535 281006 64638 281008
rect 59535 280950 59540 281006
rect 59596 280950 64638 281006
rect 59535 280948 64638 280950
rect 649986 281008 650046 281500
rect 655215 281008 655281 281011
rect 649986 281006 655281 281008
rect 649986 280950 655220 281006
rect 655276 280950 655281 281006
rect 649986 280948 655281 280950
rect 59535 280945 59601 280948
rect 655215 280945 655281 280948
rect 59343 279824 59409 279827
rect 64578 279824 64638 280318
rect 59343 279822 64638 279824
rect 59343 279766 59348 279822
rect 59404 279766 64638 279822
rect 59343 279764 64638 279766
rect 649986 279824 650046 280318
rect 654159 279824 654225 279827
rect 649986 279822 654225 279824
rect 649986 279766 654164 279822
rect 654220 279766 654225 279822
rect 649986 279764 654225 279766
rect 59343 279761 59409 279764
rect 654159 279761 654225 279764
rect 42298 278578 42304 278642
rect 42368 278640 42374 278642
rect 672303 278640 672369 278643
rect 42368 278638 672369 278640
rect 42368 278582 672308 278638
rect 672364 278582 672369 278638
rect 42368 278580 672369 278582
rect 42368 278578 42374 278580
rect 672303 278577 672369 278580
rect 43066 278430 43072 278494
rect 43136 278492 43142 278494
rect 674170 278492 674176 278494
rect 43136 278432 674176 278492
rect 43136 278430 43142 278432
rect 674170 278430 674176 278432
rect 674240 278430 674246 278494
rect 45135 278344 45201 278347
rect 672783 278344 672849 278347
rect 45135 278342 672849 278344
rect 45135 278286 45140 278342
rect 45196 278286 672788 278342
rect 672844 278286 672849 278342
rect 45135 278284 672849 278286
rect 45135 278281 45201 278284
rect 672783 278281 672849 278284
rect 61935 278196 62001 278199
rect 674746 278196 674752 278198
rect 61935 278194 674752 278196
rect 61935 278138 61940 278194
rect 61996 278138 674752 278194
rect 61935 278136 674752 278138
rect 61935 278133 62001 278136
rect 674746 278134 674752 278136
rect 674816 278196 674822 278198
rect 676527 278196 676593 278199
rect 674816 278194 676593 278196
rect 674816 278138 676532 278194
rect 676588 278138 676593 278194
rect 674816 278136 676593 278138
rect 674816 278134 674822 278136
rect 676527 278133 676593 278136
rect 42159 278048 42225 278051
rect 42490 278048 42496 278050
rect 42159 278046 42496 278048
rect 42159 277990 42164 278046
rect 42220 277990 42496 278046
rect 42159 277988 42496 277990
rect 42159 277985 42225 277988
rect 42490 277986 42496 277988
rect 42560 277986 42566 278050
rect 62607 278048 62673 278051
rect 672399 278048 672465 278051
rect 62607 278046 672465 278048
rect 62607 277990 62612 278046
rect 62668 277990 672404 278046
rect 672460 277990 672465 278046
rect 62607 277988 672465 277990
rect 62607 277985 62673 277988
rect 672399 277985 672465 277988
rect 62319 277900 62385 277903
rect 670479 277900 670545 277903
rect 62319 277898 670545 277900
rect 62319 277842 62324 277898
rect 62380 277842 670484 277898
rect 670540 277842 670545 277898
rect 62319 277840 670545 277842
rect 62319 277837 62385 277840
rect 670479 277837 670545 277840
rect 62799 277752 62865 277755
rect 670095 277752 670161 277755
rect 62799 277750 670161 277752
rect 62799 277694 62804 277750
rect 62860 277694 670100 277750
rect 670156 277694 670161 277750
rect 62799 277692 670161 277694
rect 62799 277689 62865 277692
rect 670095 277689 670161 277692
rect 62991 277604 63057 277607
rect 669903 277604 669969 277607
rect 62991 277602 669969 277604
rect 62991 277546 62996 277602
rect 63052 277546 669908 277602
rect 669964 277546 669969 277602
rect 62991 277544 669969 277546
rect 62991 277541 63057 277544
rect 669903 277541 669969 277544
rect 64719 277456 64785 277459
rect 670287 277456 670353 277459
rect 64719 277454 670353 277456
rect 64719 277398 64724 277454
rect 64780 277398 670292 277454
rect 670348 277398 670353 277454
rect 64719 277396 670353 277398
rect 64719 277393 64785 277396
rect 670287 277393 670353 277396
rect 405423 276864 405489 276867
rect 522543 276864 522609 276867
rect 405423 276862 522609 276864
rect 405423 276806 405428 276862
rect 405484 276806 522548 276862
rect 522604 276806 522609 276862
rect 405423 276804 522609 276806
rect 405423 276801 405489 276804
rect 522543 276801 522609 276804
rect 402543 276716 402609 276719
rect 529839 276716 529905 276719
rect 402543 276714 529905 276716
rect 402543 276658 402548 276714
rect 402604 276658 529844 276714
rect 529900 276658 529905 276714
rect 402543 276656 529905 276658
rect 402543 276653 402609 276656
rect 529839 276653 529905 276656
rect 41530 276506 41536 276570
rect 41600 276568 41606 276570
rect 41775 276568 41841 276571
rect 41600 276566 41841 276568
rect 41600 276510 41780 276566
rect 41836 276510 41841 276566
rect 41600 276508 41841 276510
rect 41600 276506 41606 276508
rect 41775 276505 41841 276508
rect 395151 276568 395217 276571
rect 607215 276568 607281 276571
rect 395151 276566 607281 276568
rect 395151 276510 395156 276566
rect 395212 276510 607220 276566
rect 607276 276510 607281 276566
rect 395151 276508 607281 276510
rect 395151 276505 395217 276508
rect 607215 276505 607281 276508
rect 674554 276506 674560 276570
rect 674624 276568 674630 276570
rect 679695 276568 679761 276571
rect 674624 276566 679761 276568
rect 674624 276510 679700 276566
rect 679756 276510 679761 276566
rect 674624 276508 679761 276510
rect 674624 276506 674630 276508
rect 45231 276272 45297 276275
rect 672495 276272 672561 276275
rect 45231 276270 672561 276272
rect 45231 276214 45236 276270
rect 45292 276214 672500 276270
rect 672556 276214 672561 276270
rect 45231 276212 672561 276214
rect 45231 276209 45297 276212
rect 672495 276209 672561 276212
rect 62127 276124 62193 276127
rect 674562 276124 674622 276506
rect 679695 276505 679761 276508
rect 62127 276122 674622 276124
rect 62127 276066 62132 276122
rect 62188 276066 674622 276122
rect 62127 276064 674622 276066
rect 62127 276061 62193 276064
rect 383439 275976 383505 275979
rect 577647 275976 577713 275979
rect 383439 275974 577713 275976
rect 383439 275918 383444 275974
rect 383500 275918 577652 275974
rect 577708 275918 577713 275974
rect 383439 275916 577713 275918
rect 383439 275913 383505 275916
rect 577647 275913 577713 275916
rect 390351 275828 390417 275831
rect 595407 275828 595473 275831
rect 390351 275826 595473 275828
rect 390351 275770 390356 275826
rect 390412 275770 595412 275826
rect 595468 275770 595473 275826
rect 390351 275768 595473 275770
rect 390351 275765 390417 275768
rect 595407 275765 595473 275768
rect 398895 275680 398961 275683
rect 616623 275680 616689 275683
rect 398895 275678 616689 275680
rect 398895 275622 398900 275678
rect 398956 275622 616628 275678
rect 616684 275622 616689 275678
rect 398895 275620 616689 275622
rect 398895 275617 398961 275620
rect 616623 275617 616689 275620
rect 407823 275532 407889 275535
rect 637935 275532 638001 275535
rect 407823 275530 638001 275532
rect 407823 275474 407828 275530
rect 407884 275474 637940 275530
rect 637996 275474 638001 275530
rect 407823 275472 638001 275474
rect 407823 275469 407889 275472
rect 637935 275469 638001 275472
rect 44751 275384 44817 275387
rect 646479 275384 646545 275387
rect 44751 275382 646545 275384
rect 44751 275326 44756 275382
rect 44812 275326 646484 275382
rect 646540 275326 646545 275382
rect 44751 275324 646545 275326
rect 44751 275321 44817 275324
rect 646479 275321 646545 275324
rect 50415 275236 50481 275239
rect 669519 275236 669585 275239
rect 50415 275234 669585 275236
rect 50415 275178 50420 275234
rect 50476 275178 669524 275234
rect 669580 275178 669585 275234
rect 50415 275176 669585 275178
rect 50415 275173 50481 275176
rect 669519 275173 669585 275176
rect 50607 275088 50673 275091
rect 669711 275088 669777 275091
rect 50607 275086 669777 275088
rect 50607 275030 50612 275086
rect 50668 275030 669716 275086
rect 669772 275030 669777 275086
rect 50607 275028 669777 275030
rect 50607 275025 50673 275028
rect 669711 275025 669777 275028
rect 379119 274940 379185 274943
rect 566991 274940 567057 274943
rect 379119 274938 567057 274940
rect 379119 274882 379124 274938
rect 379180 274882 566996 274938
rect 567052 274882 567057 274938
rect 379119 274880 567057 274882
rect 379119 274877 379185 274880
rect 566991 274877 567057 274880
rect 353391 274792 353457 274795
rect 503151 274792 503217 274795
rect 353391 274790 503217 274792
rect 353391 274734 353396 274790
rect 353452 274734 503156 274790
rect 503212 274734 503217 274790
rect 353391 274732 503217 274734
rect 353391 274729 353457 274732
rect 503151 274729 503217 274732
rect 350223 274644 350289 274647
rect 496047 274644 496113 274647
rect 350223 274642 496113 274644
rect 350223 274586 350228 274642
rect 350284 274586 496052 274642
rect 496108 274586 496113 274642
rect 350223 274584 496113 274586
rect 350223 274581 350289 274584
rect 496047 274581 496113 274584
rect 347631 274496 347697 274499
rect 489039 274496 489105 274499
rect 347631 274494 489105 274496
rect 347631 274438 347636 274494
rect 347692 274438 489044 274494
rect 489100 274438 489105 274494
rect 347631 274436 489105 274438
rect 347631 274433 347697 274436
rect 489039 274433 489105 274436
rect 341679 274348 341745 274351
rect 474831 274348 474897 274351
rect 341679 274346 474897 274348
rect 341679 274290 341684 274346
rect 341740 274290 474836 274346
rect 474892 274290 474897 274346
rect 341679 274288 474897 274290
rect 341679 274285 341745 274288
rect 474831 274285 474897 274288
rect 40570 274138 40576 274202
rect 40640 274200 40646 274202
rect 41775 274200 41841 274203
rect 40640 274198 41841 274200
rect 40640 274142 41780 274198
rect 41836 274142 41841 274198
rect 40640 274140 41841 274142
rect 40640 274138 40646 274140
rect 41775 274137 41841 274140
rect 45039 274200 45105 274203
rect 674362 274200 674368 274202
rect 45039 274198 674368 274200
rect 45039 274142 45044 274198
rect 45100 274142 674368 274198
rect 45039 274140 674368 274142
rect 45039 274137 45105 274140
rect 674362 274138 674368 274140
rect 674432 274138 674438 274202
rect 41338 273546 41344 273610
rect 41408 273608 41414 273610
rect 41775 273608 41841 273611
rect 41408 273606 41841 273608
rect 41408 273550 41780 273606
rect 41836 273550 41841 273606
rect 41408 273548 41841 273550
rect 41408 273546 41414 273548
rect 41775 273545 41841 273548
rect 45327 273608 45393 273611
rect 669999 273608 670065 273611
rect 45327 273606 670065 273608
rect 45327 273550 45332 273606
rect 45388 273550 670004 273606
rect 670060 273550 670065 273606
rect 45327 273548 670065 273550
rect 45327 273545 45393 273548
rect 669999 273545 670065 273548
rect 375567 273460 375633 273463
rect 558735 273460 558801 273463
rect 375567 273458 558801 273460
rect 375567 273402 375572 273458
rect 375628 273402 558740 273458
rect 558796 273402 558801 273458
rect 375567 273400 558801 273402
rect 375567 273397 375633 273400
rect 558735 273397 558801 273400
rect 378639 273312 378705 273315
rect 565839 273312 565905 273315
rect 378639 273310 565905 273312
rect 378639 273254 378644 273310
rect 378700 273254 565844 273310
rect 565900 273254 565905 273310
rect 378639 273252 565905 273254
rect 378639 273249 378705 273252
rect 565839 273249 565905 273252
rect 382959 273164 383025 273167
rect 576495 273164 576561 273167
rect 382959 273162 576561 273164
rect 382959 273106 382964 273162
rect 383020 273106 576500 273162
rect 576556 273106 576561 273162
rect 382959 273104 576561 273106
rect 382959 273101 383025 273104
rect 576495 273101 576561 273104
rect 390159 273016 390225 273019
rect 594159 273016 594225 273019
rect 390159 273014 594225 273016
rect 390159 272958 390164 273014
rect 390220 272958 594164 273014
rect 594220 272958 594225 273014
rect 390159 272956 594225 272958
rect 390159 272953 390225 272956
rect 594159 272953 594225 272956
rect 40954 272806 40960 272870
rect 41024 272868 41030 272870
rect 41775 272868 41841 272871
rect 41024 272866 41841 272868
rect 41024 272810 41780 272866
rect 41836 272810 41841 272866
rect 41024 272808 41841 272810
rect 41024 272806 41030 272808
rect 41775 272805 41841 272808
rect 392751 272868 392817 272871
rect 601263 272868 601329 272871
rect 392751 272866 601329 272868
rect 392751 272810 392756 272866
rect 392812 272810 601268 272866
rect 601324 272810 601329 272866
rect 392751 272808 601329 272810
rect 392751 272805 392817 272808
rect 601263 272805 601329 272808
rect 91887 272720 91953 272723
rect 200463 272720 200529 272723
rect 91887 272718 200529 272720
rect 91887 272662 91892 272718
rect 91948 272662 200468 272718
rect 200524 272662 200529 272718
rect 91887 272660 200529 272662
rect 91887 272657 91953 272660
rect 200463 272657 200529 272660
rect 398703 272720 398769 272723
rect 615471 272720 615537 272723
rect 398703 272718 615537 272720
rect 398703 272662 398708 272718
rect 398764 272662 615476 272718
rect 615532 272662 615537 272718
rect 398703 272660 615537 272662
rect 398703 272657 398769 272660
rect 615471 272657 615537 272660
rect 88335 272572 88401 272575
rect 199215 272572 199281 272575
rect 88335 272570 199281 272572
rect 88335 272514 88340 272570
rect 88396 272514 199220 272570
rect 199276 272514 199281 272570
rect 88335 272512 199281 272514
rect 88335 272509 88401 272512
rect 199215 272509 199281 272512
rect 404175 272572 404241 272575
rect 629679 272572 629745 272575
rect 404175 272570 629745 272572
rect 404175 272514 404180 272570
rect 404236 272514 629684 272570
rect 629740 272514 629745 272570
rect 404175 272512 629745 272514
rect 404175 272509 404241 272512
rect 629679 272509 629745 272512
rect 41146 272362 41152 272426
rect 41216 272424 41222 272426
rect 41775 272424 41841 272427
rect 41216 272422 41841 272424
rect 41216 272366 41780 272422
rect 41836 272366 41841 272422
rect 41216 272364 41841 272366
rect 41216 272362 41222 272364
rect 41775 272361 41841 272364
rect 78831 272424 78897 272427
rect 196623 272424 196689 272427
rect 78831 272422 196689 272424
rect 78831 272366 78836 272422
rect 78892 272366 196628 272422
rect 196684 272366 196689 272422
rect 78831 272364 196689 272366
rect 78831 272361 78897 272364
rect 196623 272361 196689 272364
rect 407247 272424 407313 272427
rect 636783 272424 636849 272427
rect 407247 272422 636849 272424
rect 407247 272366 407252 272422
rect 407308 272366 636788 272422
rect 636844 272366 636849 272422
rect 407247 272364 636849 272366
rect 407247 272361 407313 272364
rect 636783 272361 636849 272364
rect 72975 272276 73041 272279
rect 194415 272276 194481 272279
rect 72975 272274 194481 272276
rect 72975 272218 72980 272274
rect 73036 272218 194420 272274
rect 194476 272218 194481 272274
rect 72975 272216 194481 272218
rect 72975 272213 73041 272216
rect 194415 272213 194481 272216
rect 410895 272276 410961 272279
rect 646191 272276 646257 272279
rect 410895 272274 646257 272276
rect 410895 272218 410900 272274
rect 410956 272218 646196 272274
rect 646252 272218 646257 272274
rect 410895 272216 646257 272218
rect 410895 272213 410961 272216
rect 646191 272213 646257 272216
rect 70575 272128 70641 272131
rect 193743 272128 193809 272131
rect 70575 272126 193809 272128
rect 70575 272070 70580 272126
rect 70636 272070 193748 272126
rect 193804 272070 193809 272126
rect 70575 272068 193809 272070
rect 70575 272065 70641 272068
rect 193743 272065 193809 272068
rect 411759 272128 411825 272131
rect 648591 272128 648657 272131
rect 411759 272126 648657 272128
rect 411759 272070 411764 272126
rect 411820 272070 648596 272126
rect 648652 272070 648657 272126
rect 411759 272068 648657 272070
rect 411759 272065 411825 272068
rect 648591 272065 648657 272068
rect 370095 271980 370161 271983
rect 544527 271980 544593 271983
rect 370095 271978 544593 271980
rect 370095 271922 370100 271978
rect 370156 271922 544532 271978
rect 544588 271922 544593 271978
rect 370095 271920 544593 271922
rect 370095 271917 370161 271920
rect 544527 271917 544593 271920
rect 369615 271832 369681 271835
rect 543375 271832 543441 271835
rect 369615 271830 543441 271832
rect 369615 271774 369620 271830
rect 369676 271774 543380 271830
rect 543436 271774 543441 271830
rect 369615 271772 543441 271774
rect 369615 271769 369681 271772
rect 543375 271769 543441 271772
rect 42063 270650 42129 270651
rect 42063 270646 42112 270650
rect 42176 270648 42182 270650
rect 62511 270648 62577 270651
rect 670191 270648 670257 270651
rect 42063 270590 42068 270646
rect 42063 270586 42112 270590
rect 42176 270588 42220 270648
rect 62511 270646 670257 270648
rect 62511 270590 62516 270646
rect 62572 270590 670196 270646
rect 670252 270590 670257 270646
rect 62511 270588 670257 270590
rect 42176 270586 42182 270588
rect 42063 270585 42129 270586
rect 62511 270585 62577 270588
rect 670191 270585 670257 270588
rect 209679 270500 209745 270503
rect 214287 270500 214353 270503
rect 209679 270498 214353 270500
rect 209679 270442 209684 270498
rect 209740 270442 214292 270498
rect 214348 270442 214353 270498
rect 209679 270440 214353 270442
rect 209679 270437 209745 270440
rect 214287 270437 214353 270440
rect 374319 270500 374385 270503
rect 555183 270500 555249 270503
rect 374319 270498 555249 270500
rect 374319 270442 374324 270498
rect 374380 270442 555188 270498
rect 555244 270442 555249 270498
rect 374319 270440 555249 270442
rect 374319 270437 374385 270440
rect 555183 270437 555249 270440
rect 377007 270352 377073 270355
rect 562287 270352 562353 270355
rect 377007 270350 562353 270352
rect 377007 270294 377012 270350
rect 377068 270294 562292 270350
rect 562348 270294 562353 270350
rect 377007 270292 562353 270294
rect 377007 270289 377073 270292
rect 562287 270289 562353 270292
rect 385551 270204 385617 270207
rect 583599 270204 583665 270207
rect 385551 270202 583665 270204
rect 385551 270146 385556 270202
rect 385612 270146 583604 270202
rect 583660 270146 583665 270202
rect 385551 270144 583665 270146
rect 385551 270141 385617 270144
rect 583599 270141 583665 270144
rect 40378 269994 40384 270058
rect 40448 270056 40454 270058
rect 41775 270056 41841 270059
rect 40448 270054 41841 270056
rect 40448 269998 41780 270054
rect 41836 269998 41841 270054
rect 40448 269996 41841 269998
rect 40448 269994 40454 269996
rect 41775 269993 41841 269996
rect 388431 270056 388497 270059
rect 590607 270056 590673 270059
rect 388431 270054 590673 270056
rect 388431 269998 388436 270054
rect 388492 269998 590612 270054
rect 590668 269998 590673 270054
rect 388431 269996 590673 269998
rect 388431 269993 388497 269996
rect 590607 269993 590673 269996
rect 139119 269908 139185 269911
rect 213327 269908 213393 269911
rect 139119 269906 213393 269908
rect 139119 269850 139124 269906
rect 139180 269850 213332 269906
rect 213388 269850 213393 269906
rect 139119 269848 213393 269850
rect 139119 269845 139185 269848
rect 213327 269845 213393 269848
rect 391503 269908 391569 269911
rect 597711 269908 597777 269911
rect 391503 269906 597777 269908
rect 391503 269850 391508 269906
rect 391564 269850 597716 269906
rect 597772 269850 597777 269906
rect 391503 269848 597777 269850
rect 391503 269845 391569 269848
rect 597711 269845 597777 269848
rect 77583 269760 77649 269763
rect 196143 269760 196209 269763
rect 77583 269758 196209 269760
rect 77583 269702 77588 269758
rect 77644 269702 196148 269758
rect 196204 269702 196209 269758
rect 77583 269700 196209 269702
rect 77583 269697 77649 269700
rect 196143 269697 196209 269700
rect 403023 269760 403089 269763
rect 626127 269760 626193 269763
rect 403023 269758 626193 269760
rect 403023 269702 403028 269758
rect 403084 269702 626132 269758
rect 626188 269702 626193 269758
rect 403023 269700 626193 269702
rect 403023 269697 403089 269700
rect 626127 269697 626193 269700
rect 69423 269612 69489 269615
rect 193071 269612 193137 269615
rect 69423 269610 193137 269612
rect 69423 269554 69428 269610
rect 69484 269554 193076 269610
rect 193132 269554 193137 269610
rect 69423 269552 193137 269554
rect 69423 269549 69489 269552
rect 193071 269549 193137 269552
rect 405615 269612 405681 269615
rect 633231 269612 633297 269615
rect 405615 269610 633297 269612
rect 405615 269554 405620 269610
rect 405676 269554 633236 269610
rect 633292 269554 633297 269610
rect 405615 269552 633297 269554
rect 405615 269549 405681 269552
rect 633231 269549 633297 269552
rect 71727 269464 71793 269467
rect 194223 269464 194289 269467
rect 71727 269462 194289 269464
rect 71727 269406 71732 269462
rect 71788 269406 194228 269462
rect 194284 269406 194289 269462
rect 71727 269404 194289 269406
rect 71727 269401 71793 269404
rect 194223 269401 194289 269404
rect 410415 269464 410481 269467
rect 645039 269464 645105 269467
rect 410415 269462 645105 269464
rect 410415 269406 410420 269462
rect 410476 269406 645044 269462
rect 645100 269406 645105 269462
rect 410415 269404 645105 269406
rect 410415 269401 410481 269404
rect 645039 269401 645105 269404
rect 41871 269318 41937 269319
rect 41871 269314 41920 269318
rect 41984 269316 41990 269318
rect 65871 269316 65937 269319
rect 192399 269316 192465 269319
rect 41871 269258 41876 269314
rect 41871 269254 41920 269258
rect 41984 269256 42028 269316
rect 65871 269314 192465 269316
rect 65871 269258 65876 269314
rect 65932 269258 192404 269314
rect 192460 269258 192465 269314
rect 65871 269256 192465 269258
rect 41984 269254 41990 269256
rect 41871 269253 41937 269254
rect 65871 269253 65937 269256
rect 192399 269253 192465 269256
rect 411567 269316 411633 269319
rect 647343 269316 647409 269319
rect 411567 269314 647409 269316
rect 411567 269258 411572 269314
rect 411628 269258 647348 269314
rect 647404 269258 647409 269314
rect 411567 269256 647409 269258
rect 411567 269253 411633 269256
rect 647343 269253 647409 269256
rect 367887 269168 367953 269171
rect 539823 269168 539889 269171
rect 367887 269166 539889 269168
rect 367887 269110 367892 269166
rect 367948 269110 539828 269166
rect 539884 269110 539889 269166
rect 367887 269108 539889 269110
rect 367887 269105 367953 269108
rect 539823 269105 539889 269108
rect 368367 269020 368433 269023
rect 540975 269020 541041 269023
rect 368367 269018 541041 269020
rect 368367 268962 368372 269018
rect 368428 268962 540980 269018
rect 541036 268962 541041 269018
rect 368367 268960 541041 268962
rect 368367 268957 368433 268960
rect 540975 268957 541041 268960
rect 397071 268872 397137 268875
rect 523791 268872 523857 268875
rect 397071 268870 523857 268872
rect 397071 268814 397076 268870
rect 397132 268814 523796 268870
rect 523852 268814 523857 268870
rect 397071 268812 523857 268814
rect 397071 268809 397137 268812
rect 523791 268809 523857 268812
rect 44655 267096 44721 267099
rect 646575 267096 646641 267099
rect 44655 267094 646641 267096
rect 44655 267038 44660 267094
rect 44716 267038 646580 267094
rect 646636 267038 646641 267094
rect 44655 267036 646641 267038
rect 44655 267033 44721 267036
rect 646575 267033 646641 267036
rect 676290 266951 676350 267214
rect 43503 266948 43569 266951
rect 652239 266948 652305 266951
rect 43503 266946 652305 266948
rect 43503 266890 43508 266946
rect 43564 266890 652244 266946
rect 652300 266890 652305 266946
rect 43503 266888 652305 266890
rect 43503 266885 43569 266888
rect 652239 266885 652305 266888
rect 676239 266946 676350 266951
rect 676239 266890 676244 266946
rect 676300 266890 676350 266946
rect 676239 266888 676350 266890
rect 676239 266885 676305 266888
rect 62415 266800 62481 266803
rect 672783 266800 672849 266803
rect 62415 266798 672849 266800
rect 62415 266742 62420 266798
rect 62476 266742 672788 266798
rect 672844 266742 672849 266798
rect 62415 266740 672849 266742
rect 62415 266737 62481 266740
rect 672783 266737 672849 266740
rect 62031 266652 62097 266655
rect 672399 266652 672465 266655
rect 62031 266650 672465 266652
rect 62031 266594 62036 266650
rect 62092 266594 672404 266650
rect 672460 266594 672465 266650
rect 62031 266592 672465 266594
rect 62031 266589 62097 266592
rect 672399 266589 672465 266592
rect 62223 266504 62289 266507
rect 672975 266504 673041 266507
rect 62223 266502 673041 266504
rect 62223 266446 62228 266502
rect 62284 266446 672980 266502
rect 673036 266446 673041 266502
rect 62223 266444 673041 266446
rect 62223 266441 62289 266444
rect 672975 266441 673041 266444
rect 676143 266504 676209 266507
rect 676290 266504 676350 266770
rect 676143 266502 676350 266504
rect 676143 266446 676148 266502
rect 676204 266446 676350 266502
rect 676143 266444 676350 266446
rect 676143 266441 676209 266444
rect 61839 266356 61905 266359
rect 672591 266356 672657 266359
rect 61839 266354 672657 266356
rect 61839 266298 61844 266354
rect 61900 266298 672596 266354
rect 672652 266298 672657 266354
rect 61839 266296 672657 266298
rect 61839 266293 61905 266296
rect 672591 266293 672657 266296
rect 676047 266208 676113 266211
rect 676047 266206 676320 266208
rect 676047 266150 676052 266206
rect 676108 266150 676320 266206
rect 676047 266148 676320 266150
rect 676047 266145 676113 266148
rect 675514 265702 675520 265766
rect 675584 265764 675590 265766
rect 675584 265704 676320 265764
rect 675584 265702 675590 265704
rect 676047 265246 676113 265249
rect 676047 265244 676320 265246
rect 676047 265188 676052 265244
rect 676108 265188 676320 265244
rect 676047 265186 676320 265188
rect 676047 265183 676113 265186
rect 679695 264876 679761 264879
rect 679695 264874 679806 264876
rect 679695 264818 679700 264874
rect 679756 264818 679806 264874
rect 679695 264813 679806 264818
rect 679746 264698 679806 264813
rect 676047 264284 676113 264287
rect 676047 264282 676320 264284
rect 676047 264226 676052 264282
rect 676108 264226 676320 264282
rect 676047 264224 676320 264226
rect 676047 264221 676113 264224
rect 679791 264136 679857 264139
rect 679746 264134 679857 264136
rect 679746 264078 679796 264134
rect 679852 264078 679857 264134
rect 679746 264073 679857 264078
rect 679746 263736 679806 264073
rect 43311 263544 43377 263547
rect 649743 263544 649809 263547
rect 43311 263542 649809 263544
rect 43311 263486 43316 263542
rect 43372 263486 649748 263542
rect 649804 263486 649809 263542
rect 43311 263484 649809 263486
rect 43311 263481 43377 263484
rect 649743 263481 649809 263484
rect 673978 263248 673984 263250
rect 659490 263188 673984 263248
rect 44847 263100 44913 263103
rect 659490 263100 659550 263188
rect 673978 263186 673984 263188
rect 674048 263248 674054 263250
rect 674048 263188 676320 263248
rect 674048 263186 674054 263188
rect 44847 263098 659550 263100
rect 44847 263042 44852 263098
rect 44908 263042 659550 263098
rect 44847 263040 659550 263042
rect 44847 263037 44913 263040
rect 675514 262742 675520 262806
rect 675584 262804 675590 262806
rect 675584 262744 676320 262804
rect 675584 262742 675590 262744
rect 420399 262212 420465 262215
rect 412512 262210 420465 262212
rect 412512 262154 420404 262210
rect 420460 262154 420465 262210
rect 412512 262152 420465 262154
rect 420399 262149 420465 262152
rect 676866 262067 676926 262182
rect 676866 262062 676977 262067
rect 676866 262006 676916 262062
rect 676972 262006 676977 262062
rect 676866 262004 676977 262006
rect 676911 262001 676977 262004
rect 676290 261474 676350 261738
rect 676282 261410 676288 261474
rect 676352 261410 676358 261474
rect 676047 261324 676113 261327
rect 676047 261322 676320 261324
rect 676047 261266 676052 261322
rect 676108 261266 676320 261322
rect 676047 261264 676320 261266
rect 676047 261261 676113 261264
rect 675706 260670 675712 260734
rect 675776 260732 675782 260734
rect 675776 260672 676320 260732
rect 675776 260670 675782 260672
rect 676866 259995 676926 260184
rect 676815 259990 676926 259995
rect 676815 259934 676820 259990
rect 676876 259934 676926 259990
rect 676815 259932 676926 259934
rect 676815 259929 676881 259932
rect 420399 259844 420465 259847
rect 412512 259842 420465 259844
rect 412512 259786 420404 259842
rect 420460 259786 420465 259842
rect 412512 259784 420465 259786
rect 420399 259781 420465 259784
rect 675279 259844 675345 259847
rect 675279 259842 676320 259844
rect 675279 259786 675284 259842
rect 675340 259786 676320 259842
rect 675279 259784 676320 259786
rect 675279 259781 675345 259784
rect 191535 259400 191601 259403
rect 191535 259398 191904 259400
rect 191535 259342 191540 259398
rect 191596 259342 191904 259398
rect 191535 259340 191904 259342
rect 191535 259337 191601 259340
rect 675951 259252 676017 259255
rect 675951 259250 676320 259252
rect 675951 259194 675956 259250
rect 676012 259194 676320 259250
rect 675951 259192 676320 259194
rect 675951 259189 676017 259192
rect 676047 258734 676113 258737
rect 676047 258732 676320 258734
rect 676047 258676 676052 258732
rect 676108 258676 676320 258732
rect 676047 258674 676320 258676
rect 676047 258671 676113 258674
rect 674362 258302 674368 258366
rect 674432 258364 674438 258366
rect 674432 258304 676320 258364
rect 674432 258302 674438 258304
rect 674938 257710 674944 257774
rect 675008 257772 675014 257774
rect 675008 257712 676320 257772
rect 675008 257710 675014 257712
rect 412482 257032 412542 257520
rect 676290 257035 676350 257150
rect 420399 257032 420465 257035
rect 412482 257030 420465 257032
rect 412482 256974 420404 257030
rect 420460 256974 420465 257030
rect 412482 256972 420465 256974
rect 420399 256969 420465 256972
rect 676239 257030 676350 257035
rect 676239 256974 676244 257030
rect 676300 256974 676350 257030
rect 676239 256972 676350 256974
rect 676239 256969 676305 256972
rect 676047 256884 676113 256887
rect 676047 256882 676320 256884
rect 676047 256826 676052 256882
rect 676108 256826 676320 256882
rect 676047 256824 676320 256826
rect 676047 256821 676113 256824
rect 40194 256295 40254 256410
rect 40194 256290 40305 256295
rect 40194 256234 40244 256290
rect 40300 256234 40305 256290
rect 40194 256232 40305 256234
rect 40239 256229 40305 256232
rect 676047 256292 676113 256295
rect 676047 256290 676320 256292
rect 676047 256234 676052 256290
rect 676108 256234 676320 256290
rect 676047 256232 676320 256234
rect 676047 256229 676113 256232
rect 41538 255703 41598 255966
rect 41538 255698 41649 255703
rect 41538 255642 41588 255698
rect 41644 255642 41649 255698
rect 41538 255640 41649 255642
rect 41583 255637 41649 255640
rect 679746 255555 679806 255670
rect 679695 255550 679806 255555
rect 679695 255494 679700 255550
rect 679756 255494 679806 255550
rect 679695 255492 679806 255494
rect 679695 255489 679761 255492
rect 41775 255404 41841 255407
rect 41568 255402 41841 255404
rect 41568 255346 41780 255402
rect 41836 255346 41841 255402
rect 41568 255344 41841 255346
rect 41775 255341 41841 255344
rect 420399 255256 420465 255259
rect 412512 255254 420465 255256
rect 412512 255198 420404 255254
rect 420460 255198 420465 255254
rect 412512 255196 420465 255198
rect 420399 255193 420465 255196
rect 685506 254963 685566 255300
rect 41775 254960 41841 254963
rect 41568 254958 41841 254960
rect 41568 254902 41780 254958
rect 41836 254902 41841 254958
rect 41568 254900 41841 254902
rect 41775 254897 41841 254900
rect 679695 254960 679761 254963
rect 679695 254958 679806 254960
rect 679695 254902 679700 254958
rect 679756 254902 679806 254958
rect 679695 254897 679806 254902
rect 685455 254958 685566 254963
rect 685455 254902 685460 254958
rect 685516 254902 685566 254958
rect 685455 254900 685566 254902
rect 685455 254897 685521 254900
rect 679746 254782 679806 254897
rect 41775 254516 41841 254519
rect 41568 254514 41841 254516
rect 41568 254458 41780 254514
rect 41836 254458 41841 254514
rect 41568 254456 41841 254458
rect 41775 254453 41841 254456
rect 685455 254516 685521 254519
rect 685455 254514 685566 254516
rect 685455 254458 685460 254514
rect 685516 254458 685566 254514
rect 685455 254453 685566 254458
rect 23151 254220 23217 254223
rect 23106 254218 23217 254220
rect 23106 254162 23156 254218
rect 23212 254162 23217 254218
rect 685506 254190 685566 254453
rect 23106 254157 23217 254162
rect 23106 253894 23166 254157
rect 23298 253335 23358 253450
rect 23055 253332 23121 253335
rect 23055 253330 23166 253332
rect 23055 253274 23060 253330
rect 23116 253274 23166 253330
rect 23055 253269 23166 253274
rect 23298 253330 23409 253335
rect 23298 253274 23348 253330
rect 23404 253274 23409 253330
rect 23298 253272 23409 253274
rect 23343 253269 23409 253272
rect 675898 253270 675904 253334
rect 675968 253332 675974 253334
rect 676815 253332 676881 253335
rect 675968 253330 676881 253332
rect 675968 253274 676820 253330
rect 676876 253274 676881 253330
rect 675968 253272 676881 253274
rect 675968 253270 675974 253272
rect 676815 253269 676881 253272
rect 23106 252932 23166 253269
rect 676090 253122 676096 253186
rect 676160 253184 676166 253186
rect 676911 253184 676977 253187
rect 676160 253182 676977 253184
rect 676160 253126 676916 253182
rect 676972 253126 676977 253182
rect 676160 253124 676977 253126
rect 676160 253122 676166 253124
rect 676911 253121 676977 253124
rect 420399 252888 420465 252891
rect 412512 252886 420465 252888
rect 412512 252830 420404 252886
rect 420460 252830 420465 252886
rect 412512 252828 420465 252830
rect 420399 252825 420465 252828
rect 23247 252740 23313 252743
rect 23247 252738 23358 252740
rect 23247 252682 23252 252738
rect 23308 252682 23358 252738
rect 23247 252677 23358 252682
rect 23298 252414 23358 252677
rect 41914 252000 41920 252002
rect 41568 251940 41920 252000
rect 41914 251938 41920 251940
rect 41984 251938 41990 252002
rect 190191 251704 190257 251707
rect 190191 251702 191904 251704
rect 190191 251646 190196 251702
rect 190252 251646 191904 251702
rect 190191 251644 191904 251646
rect 190191 251641 190257 251644
rect 41538 251262 41598 251378
rect 41530 251198 41536 251262
rect 41600 251198 41606 251262
rect 42106 250964 42112 250966
rect 41568 250904 42112 250964
rect 42106 250902 42112 250904
rect 42176 250902 42182 250966
rect 675759 250816 675825 250819
rect 676282 250816 676288 250818
rect 675759 250814 676288 250816
rect 675759 250758 675764 250814
rect 675820 250758 676288 250814
rect 675759 250756 676288 250758
rect 675759 250753 675825 250756
rect 676282 250754 676288 250756
rect 676352 250754 676358 250818
rect 420303 250520 420369 250523
rect 412512 250518 420369 250520
rect 40962 250226 41022 250490
rect 412512 250462 420308 250518
rect 420364 250462 420369 250518
rect 412512 250460 420369 250462
rect 420303 250457 420369 250460
rect 40954 250162 40960 250226
rect 41024 250162 41030 250226
rect 40578 249782 40638 249898
rect 40570 249718 40576 249782
rect 40640 249718 40646 249782
rect 675567 249634 675633 249635
rect 675514 249570 675520 249634
rect 675584 249632 675633 249634
rect 675584 249630 675676 249632
rect 675628 249574 675676 249630
rect 675584 249572 675676 249574
rect 675584 249570 675633 249572
rect 675567 249569 675633 249570
rect 41871 249484 41937 249487
rect 41568 249482 41937 249484
rect 41568 249426 41876 249482
rect 41932 249426 41937 249482
rect 41568 249424 41937 249426
rect 41871 249421 41937 249424
rect 40770 248746 40830 249010
rect 40762 248682 40768 248746
rect 40832 248682 40838 248746
rect 41346 248302 41406 248418
rect 41338 248238 41344 248302
rect 41408 248238 41414 248302
rect 420399 248152 420465 248155
rect 412512 248150 420465 248152
rect 412512 248094 420404 248150
rect 420460 248094 420465 248150
rect 412512 248092 420465 248094
rect 420399 248089 420465 248092
rect 41154 247710 41214 247900
rect 41146 247646 41152 247710
rect 41216 247646 41222 247710
rect 41538 247264 41598 247530
rect 41679 247264 41745 247267
rect 41538 247262 41745 247264
rect 41538 247206 41684 247262
rect 41740 247206 41745 247262
rect 41538 247204 41745 247206
rect 41679 247201 41745 247204
rect 41346 246823 41406 246938
rect 41295 246818 41406 246823
rect 41295 246762 41300 246818
rect 41356 246762 41406 246818
rect 41295 246760 41406 246762
rect 41295 246757 41361 246760
rect 40386 246230 40446 246346
rect 40378 246166 40384 246230
rect 40448 246166 40454 246230
rect 41346 245639 41406 246050
rect 41346 245634 41457 245639
rect 41346 245578 41396 245634
rect 41452 245578 41457 245634
rect 41346 245576 41457 245578
rect 41391 245573 41457 245576
rect 41538 245195 41598 245458
rect 412482 245340 412542 245828
rect 420399 245340 420465 245343
rect 412482 245338 420465 245340
rect 412482 245282 420404 245338
rect 420460 245282 420465 245338
rect 412482 245280 420465 245282
rect 420399 245277 420465 245280
rect 41487 245190 41598 245195
rect 41487 245134 41492 245190
rect 41548 245134 41598 245190
rect 41487 245132 41598 245134
rect 41487 245129 41553 245132
rect 41775 244896 41841 244899
rect 41568 244894 41841 244896
rect 41568 244838 41780 244894
rect 41836 244838 41841 244894
rect 41568 244836 41841 244838
rect 41775 244833 41841 244836
rect 41583 244748 41649 244751
rect 41538 244746 41649 244748
rect 41538 244690 41588 244746
rect 41644 244690 41649 244746
rect 41538 244685 41649 244690
rect 41538 244496 41598 244685
rect 148335 244600 148401 244603
rect 143904 244598 148401 244600
rect 143904 244542 148340 244598
rect 148396 244542 148401 244598
rect 143904 244540 148401 244542
rect 148335 244537 148401 244540
rect 41538 243715 41598 243978
rect 41538 243710 41649 243715
rect 41538 243654 41588 243710
rect 41644 243654 41649 243710
rect 41538 243652 41649 243654
rect 41583 243649 41649 243652
rect 148719 243416 148785 243419
rect 143904 243414 148785 243416
rect 143904 243358 148724 243414
rect 148780 243358 148785 243414
rect 143904 243356 148785 243358
rect 148719 243353 148785 243356
rect 187119 243416 187185 243419
rect 191874 243416 191934 243904
rect 420303 243564 420369 243567
rect 412512 243562 420369 243564
rect 412512 243506 420308 243562
rect 420364 243506 420369 243562
rect 412512 243504 420369 243506
rect 420303 243501 420369 243504
rect 675663 243566 675729 243567
rect 675663 243562 675712 243566
rect 675776 243564 675782 243566
rect 675663 243506 675668 243562
rect 675663 243502 675712 243506
rect 675776 243504 675820 243564
rect 675776 243502 675782 243504
rect 675663 243501 675729 243502
rect 187119 243414 191934 243416
rect 187119 243358 187124 243414
rect 187180 243358 191934 243414
rect 187119 243356 191934 243358
rect 187119 243353 187185 243356
rect 143874 242084 143934 242128
rect 148527 242084 148593 242087
rect 143874 242082 148593 242084
rect 143874 242026 148532 242082
rect 148588 242026 148593 242082
rect 143874 242024 148593 242026
rect 148527 242021 148593 242024
rect 674938 242022 674944 242086
rect 675008 242084 675014 242086
rect 675375 242084 675441 242087
rect 675008 242082 675441 242084
rect 675008 242026 675380 242082
rect 675436 242026 675441 242082
rect 675008 242024 675441 242026
rect 675008 242022 675014 242024
rect 675375 242021 675441 242024
rect 420303 241196 420369 241199
rect 412512 241194 420369 241196
rect 412512 241138 420308 241194
rect 420364 241138 420369 241194
rect 412512 241136 420369 241138
rect 420303 241133 420369 241136
rect 149007 240900 149073 240903
rect 143904 240898 149073 240900
rect 143904 240842 149012 240898
rect 149068 240842 149073 240898
rect 143904 240840 149073 240842
rect 149007 240837 149073 240840
rect 674362 240542 674368 240606
rect 674432 240604 674438 240606
rect 675471 240604 675537 240607
rect 674432 240602 675537 240604
rect 674432 240546 675476 240602
rect 675532 240546 675537 240602
rect 674432 240544 675537 240546
rect 674432 240542 674438 240544
rect 675471 240541 675537 240544
rect 412239 240308 412305 240311
rect 581775 240308 581841 240311
rect 412239 240306 581841 240308
rect 412239 240250 412244 240306
rect 412300 240250 581780 240306
rect 581836 240250 581841 240306
rect 412239 240248 581841 240250
rect 412239 240245 412305 240248
rect 581775 240245 581841 240248
rect 412143 240160 412209 240163
rect 627183 240160 627249 240163
rect 412143 240158 627249 240160
rect 412143 240102 412148 240158
rect 412204 240102 627188 240158
rect 627244 240102 627249 240158
rect 412143 240100 627249 240102
rect 412143 240097 412209 240100
rect 627183 240097 627249 240100
rect 412047 240012 412113 240015
rect 567375 240012 567441 240015
rect 412047 240010 567441 240012
rect 412047 239954 412052 240010
rect 412108 239954 567380 240010
rect 567436 239954 567441 240010
rect 412047 239952 567441 239954
rect 412047 239949 412113 239952
rect 567375 239949 567441 239952
rect 148239 239716 148305 239719
rect 143904 239714 148305 239716
rect 143904 239658 148244 239714
rect 148300 239658 148305 239714
rect 143904 239656 148305 239658
rect 148239 239653 148305 239656
rect 413391 238976 413457 238979
rect 550191 238976 550257 238979
rect 413391 238974 550257 238976
rect 413391 238918 413396 238974
rect 413452 238918 550196 238974
rect 550252 238918 550257 238974
rect 413391 238916 550257 238918
rect 413391 238913 413457 238916
rect 550191 238913 550257 238916
rect 414639 238828 414705 238831
rect 573135 238828 573201 238831
rect 414639 238826 573201 238828
rect 414639 238770 414644 238826
rect 414700 238770 573140 238826
rect 573196 238770 573201 238826
rect 414639 238768 573201 238770
rect 414639 238765 414705 238768
rect 573135 238765 573201 238768
rect 413679 238680 413745 238683
rect 544335 238680 544401 238683
rect 413679 238678 544401 238680
rect 413679 238622 413684 238678
rect 413740 238622 544340 238678
rect 544396 238622 544401 238678
rect 413679 238620 544401 238622
rect 413679 238617 413745 238620
rect 544335 238617 544401 238620
rect 675759 238680 675825 238683
rect 676090 238680 676096 238682
rect 675759 238678 676096 238680
rect 675759 238622 675764 238678
rect 675820 238622 676096 238678
rect 675759 238620 676096 238622
rect 675759 238617 675825 238620
rect 676090 238618 676096 238620
rect 676160 238618 676166 238682
rect 148431 238532 148497 238535
rect 143904 238530 148497 238532
rect 143904 238474 148436 238530
rect 148492 238474 148497 238530
rect 143904 238472 148497 238474
rect 148431 238469 148497 238472
rect 413967 238384 414033 238387
rect 533487 238384 533553 238387
rect 413967 238382 533553 238384
rect 413967 238326 413972 238382
rect 414028 238326 533492 238382
rect 533548 238326 533553 238382
rect 413967 238324 533553 238326
rect 413967 238321 414033 238324
rect 533487 238321 533553 238324
rect 414255 238236 414321 238239
rect 559887 238236 559953 238239
rect 414255 238234 559953 238236
rect 414255 238178 414260 238234
rect 414316 238178 559892 238234
rect 559948 238178 559953 238234
rect 414255 238176 559953 238178
rect 414255 238173 414321 238176
rect 559887 238173 559953 238176
rect 414447 238088 414513 238091
rect 537999 238088 538065 238091
rect 414447 238086 538065 238088
rect 414447 238030 414452 238086
rect 414508 238030 538004 238086
rect 538060 238030 538065 238086
rect 414447 238028 538065 238030
rect 414447 238025 414513 238028
rect 537999 238025 538065 238028
rect 41530 237878 41536 237942
rect 41600 237940 41606 237942
rect 41775 237940 41841 237943
rect 41600 237938 41841 237940
rect 41600 237882 41780 237938
rect 41836 237882 41841 237938
rect 41600 237880 41841 237882
rect 41600 237878 41606 237880
rect 41775 237877 41841 237880
rect 143874 236756 143934 237244
rect 419151 237200 419217 237203
rect 414978 237198 419217 237200
rect 414978 237142 419156 237198
rect 419212 237142 419217 237198
rect 414978 237140 419217 237142
rect 361743 237052 361809 237055
rect 368943 237052 369009 237055
rect 377775 237052 377841 237055
rect 361743 237050 368670 237052
rect 361743 236994 361748 237050
rect 361804 236994 368670 237050
rect 361743 236992 368670 236994
rect 361743 236989 361809 236992
rect 148911 236756 148977 236759
rect 143874 236754 148977 236756
rect 143874 236698 148916 236754
rect 148972 236698 148977 236754
rect 143874 236696 148977 236698
rect 148911 236693 148977 236696
rect 368610 236460 368670 236992
rect 368943 237050 377841 237052
rect 368943 236994 368948 237050
rect 369004 236994 377780 237050
rect 377836 236994 377841 237050
rect 368943 236992 377841 236994
rect 368943 236989 369009 236992
rect 377775 236989 377841 236992
rect 377967 237052 378033 237055
rect 388431 237052 388497 237055
rect 377967 237050 388497 237052
rect 377967 236994 377972 237050
rect 378028 236994 388436 237050
rect 388492 236994 388497 237050
rect 377967 236992 388497 236994
rect 377967 236989 378033 236992
rect 388431 236989 388497 236992
rect 388719 237052 388785 237055
rect 397455 237052 397521 237055
rect 388719 237050 397521 237052
rect 388719 236994 388724 237050
rect 388780 236994 397460 237050
rect 397516 236994 397521 237050
rect 388719 236992 397521 236994
rect 388719 236989 388785 236992
rect 397455 236989 397521 236992
rect 397743 237052 397809 237055
rect 411375 237052 411441 237055
rect 397743 237050 411441 237052
rect 397743 236994 397748 237050
rect 397804 236994 411380 237050
rect 411436 236994 411441 237050
rect 397743 236992 411441 236994
rect 397743 236989 397809 236992
rect 411375 236989 411441 236992
rect 411567 237052 411633 237055
rect 414978 237052 415038 237140
rect 419151 237137 419217 237140
rect 565263 237052 565329 237055
rect 411567 237050 415038 237052
rect 411567 236994 411572 237050
rect 411628 236994 415038 237050
rect 411567 236992 415038 236994
rect 419010 237050 565329 237052
rect 419010 236994 565268 237050
rect 565324 236994 565329 237050
rect 419010 236992 565329 236994
rect 411567 236989 411633 236992
rect 370383 236904 370449 236907
rect 397551 236904 397617 236907
rect 370383 236902 397617 236904
rect 370383 236846 370388 236902
rect 370444 236846 397556 236902
rect 397612 236846 397617 236902
rect 370383 236844 397617 236846
rect 370383 236841 370449 236844
rect 397551 236841 397617 236844
rect 397743 236904 397809 236907
rect 419010 236904 419070 236992
rect 565263 236989 565329 236992
rect 397743 236902 419070 236904
rect 397743 236846 397748 236902
rect 397804 236846 419070 236902
rect 397743 236844 419070 236846
rect 419151 236904 419217 236907
rect 562191 236904 562257 236907
rect 419151 236902 562257 236904
rect 419151 236846 419156 236902
rect 419212 236846 562196 236902
rect 562252 236846 562257 236902
rect 419151 236844 562257 236846
rect 397743 236841 397809 236844
rect 419151 236841 419217 236844
rect 562191 236841 562257 236844
rect 675759 236904 675825 236907
rect 675898 236904 675904 236906
rect 675759 236902 675904 236904
rect 675759 236846 675764 236902
rect 675820 236846 675904 236902
rect 675759 236844 675904 236846
rect 675759 236841 675825 236844
rect 675898 236842 675904 236844
rect 675968 236842 675974 236906
rect 374895 236756 374961 236759
rect 559215 236756 559281 236759
rect 374895 236754 559281 236756
rect 374895 236698 374900 236754
rect 374956 236698 559220 236754
rect 559276 236698 559281 236754
rect 374895 236696 559281 236698
rect 374895 236693 374961 236696
rect 559215 236693 559281 236696
rect 373455 236608 373521 236611
rect 557007 236608 557073 236611
rect 373455 236606 557073 236608
rect 373455 236550 373460 236606
rect 373516 236550 557012 236606
rect 557068 236550 557073 236606
rect 373455 236548 557073 236550
rect 373455 236545 373521 236548
rect 557007 236545 557073 236548
rect 397071 236460 397137 236463
rect 368610 236458 397137 236460
rect 368610 236402 397076 236458
rect 397132 236402 397137 236458
rect 368610 236400 397137 236402
rect 397071 236397 397137 236400
rect 397359 236460 397425 236463
rect 553935 236460 554001 236463
rect 397359 236458 554001 236460
rect 397359 236402 397364 236458
rect 397420 236402 553940 236458
rect 553996 236402 554001 236458
rect 397359 236400 554001 236402
rect 397359 236397 397425 236400
rect 553935 236397 554001 236400
rect 372207 236312 372273 236315
rect 376527 236312 376593 236315
rect 372207 236310 376593 236312
rect 372207 236254 372212 236310
rect 372268 236254 376532 236310
rect 376588 236254 376593 236310
rect 372207 236252 376593 236254
rect 372207 236249 372273 236252
rect 376527 236249 376593 236252
rect 376719 236312 376785 236315
rect 411567 236312 411633 236315
rect 376719 236310 411633 236312
rect 376719 236254 376724 236310
rect 376780 236254 411572 236310
rect 411628 236254 411633 236310
rect 376719 236252 411633 236254
rect 376719 236249 376785 236252
rect 411567 236249 411633 236252
rect 411759 236312 411825 236315
rect 621135 236312 621201 236315
rect 411759 236310 621201 236312
rect 411759 236254 411764 236310
rect 411820 236254 621140 236310
rect 621196 236254 621201 236310
rect 411759 236252 621201 236254
rect 411759 236249 411825 236252
rect 621135 236249 621201 236252
rect 403983 236164 404049 236167
rect 587343 236164 587409 236167
rect 403983 236162 587409 236164
rect 403983 236106 403988 236162
rect 404044 236106 587348 236162
rect 587404 236106 587409 236162
rect 403983 236104 587409 236106
rect 403983 236101 404049 236104
rect 587343 236101 587409 236104
rect 149103 236016 149169 236019
rect 143904 236014 149169 236016
rect 143904 235958 149108 236014
rect 149164 235958 149169 236014
rect 143904 235956 149169 235958
rect 149103 235953 149169 235956
rect 367215 236016 367281 236019
rect 400431 236016 400497 236019
rect 367215 236014 400497 236016
rect 367215 235958 367220 236014
rect 367276 235958 400436 236014
rect 400492 235958 400497 236014
rect 367215 235956 400497 235958
rect 367215 235953 367281 235956
rect 400431 235953 400497 235956
rect 405423 236016 405489 236019
rect 588975 236016 589041 236019
rect 405423 236014 589041 236016
rect 405423 235958 405428 236014
rect 405484 235958 588980 236014
rect 589036 235958 589041 236014
rect 405423 235956 589041 235958
rect 405423 235953 405489 235956
rect 588975 235953 589041 235956
rect 393039 235868 393105 235871
rect 587823 235868 587889 235871
rect 393039 235866 587889 235868
rect 393039 235810 393044 235866
rect 393100 235810 587828 235866
rect 587884 235810 587889 235866
rect 393039 235808 587889 235810
rect 393039 235805 393105 235808
rect 587823 235805 587889 235808
rect 396783 235720 396849 235723
rect 602223 235720 602289 235723
rect 396783 235718 602289 235720
rect 396783 235662 396788 235718
rect 396844 235662 602228 235718
rect 602284 235662 602289 235718
rect 396783 235660 602289 235662
rect 396783 235657 396849 235660
rect 602223 235657 602289 235660
rect 399855 235572 399921 235575
rect 608271 235572 608337 235575
rect 399855 235570 608337 235572
rect 399855 235514 399860 235570
rect 399916 235514 608276 235570
rect 608332 235514 608337 235570
rect 399855 235512 608337 235514
rect 399855 235509 399921 235512
rect 608271 235509 608337 235512
rect 401391 235424 401457 235427
rect 611247 235424 611313 235427
rect 401391 235422 611313 235424
rect 401391 235366 401396 235422
rect 401452 235366 611252 235422
rect 611308 235366 611313 235422
rect 401391 235364 611313 235366
rect 401391 235361 401457 235364
rect 611247 235361 611313 235364
rect 356751 235276 356817 235279
rect 402543 235276 402609 235279
rect 356751 235274 402609 235276
rect 356751 235218 356756 235274
rect 356812 235218 402548 235274
rect 402604 235218 402609 235274
rect 356751 235216 402609 235218
rect 356751 235213 356817 235216
rect 402543 235213 402609 235216
rect 402735 235276 402801 235279
rect 614319 235276 614385 235279
rect 402735 235274 614385 235276
rect 402735 235218 402740 235274
rect 402796 235218 614324 235274
rect 614380 235218 614385 235274
rect 402735 235216 614385 235218
rect 402735 235213 402801 235216
rect 614319 235213 614385 235216
rect 344367 235128 344433 235131
rect 396975 235128 397041 235131
rect 344367 235126 397041 235128
rect 344367 235070 344372 235126
rect 344428 235070 396980 235126
rect 397036 235070 397041 235126
rect 344367 235068 397041 235070
rect 344367 235065 344433 235068
rect 396975 235065 397041 235068
rect 408111 235128 408177 235131
rect 624879 235128 624945 235131
rect 408111 235126 624945 235128
rect 408111 235070 408116 235126
rect 408172 235070 624884 235126
rect 624940 235070 624945 235126
rect 408111 235068 624945 235070
rect 408111 235065 408177 235068
rect 624879 235065 624945 235068
rect 299439 234980 299505 234983
rect 354351 234980 354417 234983
rect 299439 234978 354417 234980
rect 299439 234922 299444 234978
rect 299500 234922 354356 234978
rect 354412 234922 354417 234978
rect 299439 234920 354417 234922
rect 299439 234917 299505 234920
rect 354351 234917 354417 234920
rect 356847 234980 356913 234983
rect 403407 234980 403473 234983
rect 356847 234978 403473 234980
rect 356847 234922 356852 234978
rect 356908 234922 403412 234978
rect 403468 234922 403473 234978
rect 356847 234920 403473 234922
rect 356847 234917 356913 234920
rect 403407 234917 403473 234920
rect 408495 234980 408561 234983
rect 625551 234980 625617 234983
rect 408495 234978 625617 234980
rect 408495 234922 408500 234978
rect 408556 234922 625556 234978
rect 625612 234922 625617 234978
rect 408495 234920 625617 234922
rect 408495 234917 408561 234920
rect 625551 234917 625617 234920
rect 148815 234832 148881 234835
rect 143904 234830 148881 234832
rect 143904 234774 148820 234830
rect 148876 234774 148881 234830
rect 143904 234772 148881 234774
rect 148815 234769 148881 234772
rect 301647 234832 301713 234835
rect 345327 234832 345393 234835
rect 301647 234830 345393 234832
rect 301647 234774 301652 234830
rect 301708 234774 345332 234830
rect 345388 234774 345393 234830
rect 301647 234772 345393 234774
rect 301647 234769 301713 234772
rect 345327 234769 345393 234772
rect 347631 234832 347697 234835
rect 407439 234832 407505 234835
rect 347631 234830 407505 234832
rect 347631 234774 347636 234830
rect 347692 234774 407444 234830
rect 407500 234774 407505 234830
rect 347631 234772 407505 234774
rect 347631 234769 347697 234772
rect 407439 234769 407505 234772
rect 409935 234832 410001 234835
rect 627855 234832 627921 234835
rect 409935 234830 627921 234832
rect 409935 234774 409940 234830
rect 409996 234774 627860 234830
rect 627916 234774 627921 234830
rect 409935 234772 627921 234774
rect 409935 234769 410001 234772
rect 627855 234769 627921 234772
rect 299343 234684 299409 234687
rect 405327 234684 405393 234687
rect 299343 234682 405393 234684
rect 299343 234626 299348 234682
rect 299404 234626 405332 234682
rect 405388 234626 405393 234682
rect 299343 234624 405393 234626
rect 299343 234621 299409 234624
rect 405327 234621 405393 234624
rect 405519 234684 405585 234687
rect 411279 234684 411345 234687
rect 630927 234684 630993 234687
rect 405519 234682 406206 234684
rect 405519 234626 405524 234682
rect 405580 234626 406206 234682
rect 405519 234624 406206 234626
rect 405519 234621 405585 234624
rect 364047 234536 364113 234539
rect 405903 234536 405969 234539
rect 364047 234534 405969 234536
rect 364047 234478 364052 234534
rect 364108 234478 405908 234534
rect 405964 234478 405969 234534
rect 364047 234476 405969 234478
rect 406146 234536 406206 234624
rect 411279 234682 630993 234684
rect 411279 234626 411284 234682
rect 411340 234626 630932 234682
rect 630988 234626 630993 234682
rect 411279 234624 630993 234626
rect 411279 234621 411345 234624
rect 630927 234621 630993 234624
rect 587439 234536 587505 234539
rect 406146 234534 587505 234536
rect 406146 234478 587444 234534
rect 587500 234478 587505 234534
rect 406146 234476 587505 234478
rect 364047 234473 364113 234476
rect 405903 234473 405969 234476
rect 587439 234473 587505 234476
rect 341583 234388 341649 234391
rect 490479 234388 490545 234391
rect 341583 234386 490545 234388
rect 341583 234330 341588 234386
rect 341644 234330 490484 234386
rect 490540 234330 490545 234386
rect 341583 234328 490545 234330
rect 341583 234325 341649 234328
rect 490479 234325 490545 234328
rect 338607 234240 338673 234243
rect 466479 234240 466545 234243
rect 338607 234238 466545 234240
rect 338607 234182 338612 234238
rect 338668 234182 466484 234238
rect 466540 234182 466545 234238
rect 338607 234180 466545 234182
rect 338607 234177 338673 234180
rect 466479 234177 466545 234180
rect 407247 234092 407313 234095
rect 506799 234092 506865 234095
rect 407247 234090 506865 234092
rect 407247 234034 407252 234090
rect 407308 234034 506804 234090
rect 506860 234034 506865 234090
rect 407247 234032 506865 234034
rect 407247 234029 407313 234032
rect 506799 234029 506865 234032
rect 379119 233944 379185 233947
rect 411471 233944 411537 233947
rect 379119 233942 411537 233944
rect 379119 233886 379124 233942
rect 379180 233886 411476 233942
rect 411532 233886 411537 233942
rect 379119 233884 411537 233886
rect 379119 233881 379185 233884
rect 411471 233881 411537 233884
rect 382095 233796 382161 233799
rect 411759 233796 411825 233799
rect 382095 233794 411825 233796
rect 382095 233738 382100 233794
rect 382156 233738 411764 233794
rect 411820 233738 411825 233794
rect 382095 233736 411825 233738
rect 382095 233733 382161 233736
rect 411759 233733 411825 233736
rect 148623 233648 148689 233651
rect 143904 233646 148689 233648
rect 143904 233590 148628 233646
rect 148684 233590 148689 233646
rect 143904 233588 148689 233590
rect 148623 233585 148689 233588
rect 376335 233648 376401 233651
rect 408783 233648 408849 233651
rect 376335 233646 408849 233648
rect 376335 233590 376340 233646
rect 376396 233590 408788 233646
rect 408844 233590 408849 233646
rect 376335 233588 408849 233590
rect 376335 233585 376401 233588
rect 408783 233585 408849 233588
rect 40570 233290 40576 233354
rect 40640 233352 40646 233354
rect 41775 233352 41841 233355
rect 40640 233350 41841 233352
rect 40640 233294 41780 233350
rect 41836 233294 41841 233350
rect 40640 233292 41841 233294
rect 40640 233290 40646 233292
rect 41775 233289 41841 233292
rect 365679 233352 365745 233355
rect 377199 233352 377265 233355
rect 365679 233350 377265 233352
rect 365679 233294 365684 233350
rect 365740 233294 377204 233350
rect 377260 233294 377265 233350
rect 365679 233292 377265 233294
rect 365679 233289 365745 233292
rect 377199 233289 377265 233292
rect 334863 233204 334929 233207
rect 479055 233204 479121 233207
rect 334863 233202 479121 233204
rect 334863 233146 334868 233202
rect 334924 233146 479060 233202
rect 479116 233146 479121 233202
rect 334863 233144 479121 233146
rect 334863 233141 334929 233144
rect 479055 233141 479121 233144
rect 359055 233056 359121 233059
rect 525231 233056 525297 233059
rect 359055 233054 525297 233056
rect 359055 232998 359060 233054
rect 359116 232998 525236 233054
rect 525292 232998 525297 233054
rect 359055 232996 525297 232998
rect 359055 232993 359121 232996
rect 525231 232993 525297 232996
rect 370767 232908 370833 232911
rect 551631 232908 551697 232911
rect 370767 232906 551697 232908
rect 370767 232850 370772 232906
rect 370828 232850 551636 232906
rect 551692 232850 551697 232906
rect 370767 232848 551697 232850
rect 370767 232845 370833 232848
rect 551631 232845 551697 232848
rect 375375 232760 375441 232763
rect 560751 232760 560817 232763
rect 375375 232758 560817 232760
rect 375375 232702 375380 232758
rect 375436 232702 560756 232758
rect 560812 232702 560817 232758
rect 375375 232700 560817 232702
rect 375375 232697 375441 232700
rect 560751 232697 560817 232700
rect 378735 232612 378801 232615
rect 564495 232612 564561 232615
rect 378735 232610 564561 232612
rect 378735 232554 378740 232610
rect 378796 232554 564500 232610
rect 564556 232554 564561 232610
rect 378735 232552 564561 232554
rect 378735 232549 378801 232552
rect 564495 232549 564561 232552
rect 381711 232464 381777 232467
rect 570447 232464 570513 232467
rect 381711 232462 570513 232464
rect 381711 232406 381716 232462
rect 381772 232406 570452 232462
rect 570508 232406 570513 232462
rect 381711 232404 570513 232406
rect 381711 232401 381777 232404
rect 570447 232401 570513 232404
rect 147855 232316 147921 232319
rect 143904 232314 147921 232316
rect 143904 232258 147860 232314
rect 147916 232258 147921 232314
rect 143904 232256 147921 232258
rect 147855 232253 147921 232256
rect 384975 232316 385041 232319
rect 576591 232316 576657 232319
rect 384975 232314 576657 232316
rect 384975 232258 384980 232314
rect 385036 232258 576596 232314
rect 576652 232258 576657 232314
rect 384975 232256 576657 232258
rect 384975 232253 385041 232256
rect 576591 232253 576657 232256
rect 385359 232168 385425 232171
rect 578031 232168 578097 232171
rect 385359 232166 578097 232168
rect 385359 232110 385364 232166
rect 385420 232110 578036 232166
rect 578092 232110 578097 232166
rect 385359 232108 578097 232110
rect 385359 232105 385425 232108
rect 578031 232105 578097 232108
rect 382959 232020 383025 232023
rect 575823 232020 575889 232023
rect 382959 232018 575889 232020
rect 382959 231962 382964 232018
rect 383020 231962 575828 232018
rect 575884 231962 575889 232018
rect 382959 231960 575889 231962
rect 382959 231957 383025 231960
rect 575823 231957 575889 231960
rect 298959 231872 299025 231875
rect 385839 231872 385905 231875
rect 298959 231870 385905 231872
rect 298959 231814 298964 231870
rect 299020 231814 385844 231870
rect 385900 231814 385905 231870
rect 298959 231812 385905 231814
rect 298959 231809 299025 231812
rect 385839 231809 385905 231812
rect 405231 231872 405297 231875
rect 604527 231872 604593 231875
rect 405231 231870 604593 231872
rect 405231 231814 405236 231870
rect 405292 231814 604532 231870
rect 604588 231814 604593 231870
rect 405231 231812 604593 231814
rect 405231 231809 405297 231812
rect 604527 231809 604593 231812
rect 330255 231724 330321 231727
rect 470127 231724 470193 231727
rect 330255 231722 470193 231724
rect 330255 231666 330260 231722
rect 330316 231666 470132 231722
rect 470188 231666 470193 231722
rect 330255 231664 470193 231666
rect 330255 231661 330321 231664
rect 470127 231661 470193 231664
rect 327087 231576 327153 231579
rect 464079 231576 464145 231579
rect 327087 231574 464145 231576
rect 327087 231518 327092 231574
rect 327148 231518 464084 231574
rect 464140 231518 464145 231574
rect 327087 231516 464145 231518
rect 327087 231513 327153 231516
rect 464079 231513 464145 231516
rect 322479 231428 322545 231431
rect 455151 231428 455217 231431
rect 322479 231426 455217 231428
rect 322479 231370 322484 231426
rect 322540 231370 455156 231426
rect 455212 231370 455217 231426
rect 322479 231368 455217 231370
rect 322479 231365 322545 231368
rect 455151 231365 455217 231368
rect 316719 231280 316785 231283
rect 442863 231280 442929 231283
rect 316719 231278 442929 231280
rect 316719 231222 316724 231278
rect 316780 231222 442868 231278
rect 442924 231222 442929 231278
rect 316719 231220 442929 231222
rect 316719 231217 316785 231220
rect 442863 231217 442929 231220
rect 40378 231070 40384 231134
rect 40448 231132 40454 231134
rect 41775 231132 41841 231135
rect 149391 231132 149457 231135
rect 40448 231130 41841 231132
rect 40448 231074 41780 231130
rect 41836 231074 41841 231130
rect 40448 231072 41841 231074
rect 143904 231130 149457 231132
rect 143904 231074 149396 231130
rect 149452 231074 149457 231130
rect 143904 231072 149457 231074
rect 40448 231070 40454 231072
rect 41775 231069 41841 231072
rect 149391 231069 149457 231072
rect 307599 231132 307665 231135
rect 424719 231132 424785 231135
rect 307599 231130 424785 231132
rect 307599 231074 307604 231130
rect 307660 231074 424724 231130
rect 424780 231074 424785 231130
rect 307599 231072 424785 231074
rect 307599 231069 307665 231072
rect 424719 231069 424785 231072
rect 352719 230836 352785 230839
rect 359055 230836 359121 230839
rect 352719 230834 359121 230836
rect 352719 230778 352724 230834
rect 352780 230778 359060 230834
rect 359116 230778 359121 230834
rect 352719 230776 359121 230778
rect 352719 230773 352785 230776
rect 359055 230773 359121 230776
rect 41146 230330 41152 230394
rect 41216 230392 41222 230394
rect 41775 230392 41841 230395
rect 41216 230390 41841 230392
rect 41216 230334 41780 230390
rect 41836 230334 41841 230390
rect 41216 230332 41841 230334
rect 41216 230330 41222 230332
rect 41775 230329 41841 230332
rect 339855 230392 339921 230395
rect 354255 230392 354321 230395
rect 339855 230390 354321 230392
rect 339855 230334 339860 230390
rect 339916 230334 354260 230390
rect 354316 230334 354321 230390
rect 339855 230332 354321 230334
rect 339855 230329 339921 230332
rect 354255 230329 354321 230332
rect 360879 230392 360945 230395
rect 528303 230392 528369 230395
rect 360879 230390 528369 230392
rect 360879 230334 360884 230390
rect 360940 230334 528308 230390
rect 528364 230334 528369 230390
rect 360879 230332 528369 230334
rect 360879 230329 360945 230332
rect 528303 230329 528369 230332
rect 407631 230244 407697 230247
rect 575055 230244 575121 230247
rect 407631 230242 575121 230244
rect 407631 230186 407636 230242
rect 407692 230186 575060 230242
rect 575116 230186 575121 230242
rect 407631 230184 575121 230186
rect 407631 230181 407697 230184
rect 575055 230181 575121 230184
rect 363567 230096 363633 230099
rect 534255 230096 534321 230099
rect 363567 230094 534321 230096
rect 363567 230038 363572 230094
rect 363628 230038 534260 230094
rect 534316 230038 534321 230094
rect 363567 230036 534321 230038
rect 363567 230033 363633 230036
rect 534255 230033 534321 230036
rect 146895 229948 146961 229951
rect 143904 229946 146961 229948
rect 143904 229890 146900 229946
rect 146956 229890 146961 229946
rect 143904 229888 146961 229890
rect 146895 229885 146961 229888
rect 358959 229948 359025 229951
rect 527535 229948 527601 229951
rect 358959 229946 527601 229948
rect 358959 229890 358964 229946
rect 359020 229890 527540 229946
rect 527596 229890 527601 229946
rect 358959 229888 527601 229890
rect 358959 229885 359025 229888
rect 527535 229885 527601 229888
rect 41338 229738 41344 229802
rect 41408 229800 41414 229802
rect 41775 229800 41841 229803
rect 41408 229798 41841 229800
rect 41408 229742 41780 229798
rect 41836 229742 41841 229798
rect 41408 229740 41841 229742
rect 41408 229738 41414 229740
rect 41775 229737 41841 229740
rect 373071 229800 373137 229803
rect 553935 229800 554001 229803
rect 373071 229798 554001 229800
rect 373071 229742 373076 229798
rect 373132 229742 553940 229798
rect 553996 229742 554001 229798
rect 373071 229740 554001 229742
rect 373071 229737 373137 229740
rect 553935 229737 554001 229740
rect 376815 229652 376881 229655
rect 563631 229652 563697 229655
rect 376815 229650 563697 229652
rect 376815 229594 376820 229650
rect 376876 229594 563636 229650
rect 563692 229594 563697 229650
rect 376815 229592 563697 229594
rect 376815 229589 376881 229592
rect 563631 229589 563697 229592
rect 381327 229504 381393 229507
rect 572751 229504 572817 229507
rect 381327 229502 572817 229504
rect 381327 229446 381332 229502
rect 381388 229446 572756 229502
rect 572812 229446 572817 229502
rect 381327 229444 572817 229446
rect 381327 229441 381393 229444
rect 572751 229441 572817 229444
rect 383535 229356 383601 229359
rect 573519 229356 573585 229359
rect 383535 229354 573585 229356
rect 383535 229298 383540 229354
rect 383596 229298 573524 229354
rect 573580 229298 573585 229354
rect 383535 229296 573585 229298
rect 383535 229293 383601 229296
rect 573519 229293 573585 229296
rect 384399 229208 384465 229211
rect 578895 229208 578961 229211
rect 384399 229206 578961 229208
rect 384399 229150 384404 229206
rect 384460 229150 578900 229206
rect 578956 229150 578961 229206
rect 384399 229148 578961 229150
rect 384399 229145 384465 229148
rect 578895 229145 578961 229148
rect 40954 228998 40960 229062
rect 41024 229060 41030 229062
rect 41775 229060 41841 229063
rect 41024 229058 41841 229060
rect 41024 229002 41780 229058
rect 41836 229002 41841 229058
rect 41024 229000 41841 229002
rect 41024 228998 41030 229000
rect 41775 228997 41841 229000
rect 398127 229060 398193 229063
rect 599919 229060 599985 229063
rect 398127 229058 599985 229060
rect 398127 229002 398132 229058
rect 398188 229002 599924 229058
rect 599980 229002 599985 229058
rect 398127 229000 599985 229002
rect 398127 228997 398193 229000
rect 599919 228997 599985 229000
rect 292143 228912 292209 228915
rect 359823 228912 359889 228915
rect 292143 228910 359889 228912
rect 292143 228854 292148 228910
rect 292204 228854 359828 228910
rect 359884 228854 359889 228910
rect 292143 228852 359889 228854
rect 292143 228849 292209 228852
rect 359823 228849 359889 228852
rect 399471 228912 399537 228915
rect 607503 228912 607569 228915
rect 399471 228910 607569 228912
rect 399471 228854 399476 228910
rect 399532 228854 607508 228910
rect 607564 228854 607569 228910
rect 399471 228852 607569 228854
rect 399471 228849 399537 228852
rect 607503 228849 607569 228852
rect 342159 228764 342225 228767
rect 494223 228764 494289 228767
rect 342159 228762 494289 228764
rect 342159 228706 342164 228762
rect 342220 228706 494228 228762
rect 494284 228706 494289 228762
rect 342159 228704 494289 228706
rect 342159 228701 342225 228704
rect 494223 228701 494289 228704
rect 143874 228172 143934 228660
rect 345423 228616 345489 228619
rect 497967 228616 498033 228619
rect 345423 228614 498033 228616
rect 345423 228558 345428 228614
rect 345484 228558 497972 228614
rect 498028 228558 498033 228614
rect 345423 228556 498033 228558
rect 345423 228553 345489 228556
rect 497967 228553 498033 228556
rect 339375 228468 339441 228471
rect 488271 228468 488337 228471
rect 339375 228466 488337 228468
rect 339375 228410 339380 228466
rect 339436 228410 488276 228466
rect 488332 228410 488337 228466
rect 339375 228408 488337 228410
rect 339375 228405 339441 228408
rect 488271 228405 488337 228408
rect 333039 228320 333105 228323
rect 476175 228320 476241 228323
rect 333039 228318 476241 228320
rect 333039 228262 333044 228318
rect 333100 228262 476180 228318
rect 476236 228262 476241 228318
rect 333039 228260 476241 228262
rect 333039 228257 333105 228260
rect 476175 228257 476241 228260
rect 149391 228172 149457 228175
rect 143874 228170 149457 228172
rect 143874 228114 149396 228170
rect 149452 228114 149457 228170
rect 143874 228112 149457 228114
rect 149391 228109 149457 228112
rect 313455 228172 313521 228175
rect 436911 228172 436977 228175
rect 313455 228170 436977 228172
rect 313455 228114 313460 228170
rect 313516 228114 436916 228170
rect 436972 228114 436977 228170
rect 313455 228112 436977 228114
rect 313455 228109 313521 228112
rect 436911 228109 436977 228112
rect 41530 227370 41536 227434
rect 41600 227432 41606 227434
rect 41775 227432 41841 227435
rect 149391 227432 149457 227435
rect 41600 227430 41841 227432
rect 41600 227374 41780 227430
rect 41836 227374 41841 227430
rect 41600 227372 41841 227374
rect 143904 227430 149457 227432
rect 143904 227374 149396 227430
rect 149452 227374 149457 227430
rect 143904 227372 149457 227374
rect 41600 227370 41606 227372
rect 41775 227369 41841 227372
rect 149391 227369 149457 227372
rect 336879 227432 336945 227435
rect 481455 227432 481521 227435
rect 336879 227430 481521 227432
rect 336879 227374 336884 227430
rect 336940 227374 481460 227430
rect 481516 227374 481521 227430
rect 336879 227372 481521 227374
rect 336879 227369 336945 227372
rect 481455 227369 481521 227372
rect 343119 227284 343185 227287
rect 493455 227284 493521 227287
rect 343119 227282 493521 227284
rect 343119 227226 343124 227282
rect 343180 227226 493460 227282
rect 493516 227226 493521 227282
rect 343119 227224 493521 227226
rect 343119 227221 343185 227224
rect 493455 227221 493521 227224
rect 344751 227136 344817 227139
rect 498831 227136 498897 227139
rect 344751 227134 498897 227136
rect 344751 227078 344756 227134
rect 344812 227078 498836 227134
rect 498892 227078 498897 227134
rect 344751 227076 498897 227078
rect 344751 227073 344817 227076
rect 498831 227073 498897 227076
rect 391215 226988 391281 226991
rect 590895 226988 590961 226991
rect 391215 226986 590961 226988
rect 391215 226930 391220 226986
rect 391276 226930 590900 226986
rect 590956 226930 590961 226986
rect 391215 226928 590961 226930
rect 391215 226925 391281 226928
rect 590895 226925 590961 226928
rect 391599 226840 391665 226843
rect 591663 226840 591729 226843
rect 391599 226838 591729 226840
rect 391599 226782 391604 226838
rect 391660 226782 591668 226838
rect 591724 226782 591729 226838
rect 391599 226780 591729 226782
rect 391599 226777 391665 226780
rect 591663 226777 591729 226780
rect 40762 226630 40768 226694
rect 40832 226692 40838 226694
rect 41775 226692 41841 226695
rect 40832 226690 41841 226692
rect 40832 226634 41780 226690
rect 41836 226634 41841 226690
rect 40832 226632 41841 226634
rect 40832 226630 40838 226632
rect 41775 226629 41841 226632
rect 394479 226692 394545 226695
rect 596943 226692 597009 226695
rect 394479 226690 597009 226692
rect 394479 226634 394484 226690
rect 394540 226634 596948 226690
rect 597004 226634 597009 226690
rect 394479 226632 597009 226634
rect 394479 226629 394545 226632
rect 596943 226629 597009 226632
rect 394095 226544 394161 226547
rect 596175 226544 596241 226547
rect 394095 226542 596241 226544
rect 394095 226486 394100 226542
rect 394156 226486 596180 226542
rect 596236 226486 596241 226542
rect 394095 226484 596241 226486
rect 394095 226481 394161 226484
rect 596175 226481 596241 226484
rect 147087 226396 147153 226399
rect 143904 226394 147153 226396
rect 143904 226338 147092 226394
rect 147148 226338 147153 226394
rect 143904 226336 147153 226338
rect 147087 226333 147153 226336
rect 402639 226396 402705 226399
rect 613551 226396 613617 226399
rect 402639 226394 613617 226396
rect 402639 226338 402644 226394
rect 402700 226338 613556 226394
rect 613612 226338 613617 226394
rect 402639 226336 613617 226338
rect 402639 226333 402705 226336
rect 613551 226333 613617 226336
rect 42063 226250 42129 226251
rect 42063 226246 42112 226250
rect 42176 226248 42182 226250
rect 407535 226248 407601 226251
rect 623343 226248 623409 226251
rect 42063 226190 42068 226246
rect 42063 226186 42112 226190
rect 42176 226188 42220 226248
rect 407535 226246 623409 226248
rect 407535 226190 407540 226246
rect 407596 226190 623348 226246
rect 623404 226190 623409 226246
rect 407535 226188 623409 226190
rect 42176 226186 42182 226188
rect 42063 226185 42129 226186
rect 407535 226185 407601 226188
rect 623343 226185 623409 226188
rect 405807 226100 405873 226103
rect 620367 226100 620433 226103
rect 405807 226098 620433 226100
rect 405807 226042 405812 226098
rect 405868 226042 620372 226098
rect 620428 226042 620433 226098
rect 405807 226040 620433 226042
rect 405807 226037 405873 226040
rect 620367 226037 620433 226040
rect 333807 225952 333873 225955
rect 475311 225952 475377 225955
rect 333807 225950 475377 225952
rect 333807 225894 333812 225950
rect 333868 225894 475316 225950
rect 475372 225894 475377 225950
rect 333807 225892 475377 225894
rect 333807 225889 333873 225892
rect 475311 225889 475377 225892
rect 331023 225804 331089 225807
rect 469359 225804 469425 225807
rect 331023 225802 469425 225804
rect 331023 225746 331028 225802
rect 331084 225746 469364 225802
rect 469420 225746 469425 225802
rect 331023 225744 469425 225746
rect 331023 225741 331089 225744
rect 469359 225741 469425 225744
rect 327951 225656 328017 225659
rect 463311 225656 463377 225659
rect 327951 225654 463377 225656
rect 327951 225598 327956 225654
rect 328012 225598 463316 225654
rect 463372 225598 463377 225654
rect 327951 225596 463377 225598
rect 327951 225593 328017 225596
rect 463311 225593 463377 225596
rect 354255 225508 354321 225511
rect 487503 225508 487569 225511
rect 354255 225506 487569 225508
rect 354255 225450 354260 225506
rect 354316 225450 487508 225506
rect 487564 225450 487569 225506
rect 354255 225448 487569 225450
rect 354255 225445 354321 225448
rect 487503 225445 487569 225448
rect 325935 225360 326001 225363
rect 457263 225360 457329 225363
rect 325935 225358 457329 225360
rect 325935 225302 325940 225358
rect 325996 225302 457268 225358
rect 457324 225302 457329 225358
rect 325935 225300 457329 225302
rect 325935 225297 326001 225300
rect 457263 225297 457329 225300
rect 149487 225212 149553 225215
rect 143904 225210 149553 225212
rect 143904 225154 149492 225210
rect 149548 225154 149553 225210
rect 143904 225152 149553 225154
rect 149487 225149 149553 225152
rect 318927 225212 318993 225215
rect 445167 225212 445233 225215
rect 318927 225210 445233 225212
rect 318927 225154 318932 225210
rect 318988 225154 445172 225210
rect 445228 225154 445233 225210
rect 318927 225152 445233 225154
rect 318927 225149 318993 225152
rect 445167 225149 445233 225152
rect 359439 224620 359505 224623
rect 526671 224620 526737 224623
rect 359439 224618 526737 224620
rect 359439 224562 359444 224618
rect 359500 224562 526676 224618
rect 526732 224562 526737 224618
rect 359439 224560 526737 224562
rect 359439 224557 359505 224560
rect 526671 224557 526737 224560
rect 354159 224472 354225 224475
rect 518415 224472 518481 224475
rect 354159 224470 518481 224472
rect 354159 224414 354164 224470
rect 354220 224414 518420 224470
rect 518476 224414 518481 224470
rect 354159 224412 518481 224414
rect 354159 224409 354225 224412
rect 518415 224409 518481 224412
rect 360975 224324 361041 224327
rect 530511 224324 530577 224327
rect 360975 224322 530577 224324
rect 360975 224266 360980 224322
rect 361036 224266 530516 224322
rect 530572 224266 530577 224322
rect 360975 224264 530577 224266
rect 360975 224261 361041 224264
rect 530511 224261 530577 224264
rect 359727 224176 359793 224179
rect 528975 224176 529041 224179
rect 359727 224174 529041 224176
rect 359727 224118 359732 224174
rect 359788 224118 528980 224174
rect 529036 224118 529041 224174
rect 359727 224116 529041 224118
rect 359727 224113 359793 224116
rect 528975 224113 529041 224116
rect 363471 224028 363537 224031
rect 536559 224028 536625 224031
rect 363471 224026 536625 224028
rect 363471 223970 363476 224026
rect 363532 223970 536564 224026
rect 536620 223970 536625 224026
rect 363471 223968 536625 223970
rect 363471 223965 363537 223968
rect 536559 223965 536625 223968
rect 149487 223880 149553 223883
rect 143904 223878 149553 223880
rect 143904 223822 149492 223878
rect 149548 223822 149553 223878
rect 143904 223820 149553 223822
rect 149487 223817 149553 223820
rect 366159 223880 366225 223883
rect 541071 223880 541137 223883
rect 366159 223878 541137 223880
rect 366159 223822 366164 223878
rect 366220 223822 541076 223878
rect 541132 223822 541137 223878
rect 366159 223820 541137 223822
rect 366159 223817 366225 223820
rect 541071 223817 541137 223820
rect 367599 223732 367665 223735
rect 544047 223732 544113 223735
rect 367599 223730 544113 223732
rect 367599 223674 367604 223730
rect 367660 223674 544052 223730
rect 544108 223674 544113 223730
rect 367599 223672 544113 223674
rect 367599 223669 367665 223672
rect 544047 223669 544113 223672
rect 377583 223584 377649 223587
rect 562959 223584 563025 223587
rect 377583 223582 563025 223584
rect 377583 223526 377588 223582
rect 377644 223526 562964 223582
rect 563020 223526 563025 223582
rect 377583 223524 563025 223526
rect 377583 223521 377649 223524
rect 562959 223521 563025 223524
rect 379791 223436 379857 223439
rect 568239 223436 568305 223439
rect 379791 223434 568305 223436
rect 379791 223378 379796 223434
rect 379852 223378 568244 223434
rect 568300 223378 568305 223434
rect 379791 223376 568305 223378
rect 379791 223373 379857 223376
rect 568239 223373 568305 223376
rect 381231 223288 381297 223291
rect 571311 223288 571377 223291
rect 381231 223286 571377 223288
rect 381231 223230 381236 223286
rect 381292 223230 571316 223286
rect 571372 223230 571377 223286
rect 381231 223228 571377 223230
rect 381231 223225 381297 223228
rect 571311 223225 571377 223228
rect 384303 223140 384369 223143
rect 577263 223140 577329 223143
rect 384303 223138 577329 223140
rect 384303 223082 384308 223138
rect 384364 223082 577268 223138
rect 577324 223082 577329 223138
rect 384303 223080 577329 223082
rect 384303 223077 384369 223080
rect 577263 223077 577329 223080
rect 357423 222992 357489 222995
rect 524463 222992 524529 222995
rect 357423 222990 524529 222992
rect 357423 222934 357428 222990
rect 357484 222934 524468 222990
rect 524524 222934 524529 222990
rect 357423 222932 524529 222934
rect 357423 222929 357489 222932
rect 524463 222929 524529 222932
rect 385743 222844 385809 222847
rect 532047 222844 532113 222847
rect 385743 222842 532113 222844
rect 385743 222786 385748 222842
rect 385804 222786 532052 222842
rect 532108 222786 532113 222842
rect 385743 222784 532113 222786
rect 385743 222781 385809 222784
rect 532047 222781 532113 222784
rect 149391 222696 149457 222699
rect 143904 222694 149457 222696
rect 143904 222638 149396 222694
rect 149452 222638 149457 222694
rect 143904 222636 149457 222638
rect 149391 222633 149457 222636
rect 400047 222696 400113 222699
rect 523791 222696 523857 222699
rect 400047 222694 523857 222696
rect 400047 222638 400052 222694
rect 400108 222638 523796 222694
rect 523852 222638 523857 222694
rect 400047 222636 523857 222638
rect 400047 222633 400113 222636
rect 523791 222633 523857 222636
rect 403407 222548 403473 222551
rect 522927 222548 522993 222551
rect 403407 222546 522993 222548
rect 403407 222490 403412 222546
rect 403468 222490 522932 222546
rect 522988 222490 522993 222546
rect 403407 222488 522993 222490
rect 403407 222485 403473 222488
rect 522927 222485 522993 222488
rect 676290 221811 676350 222074
rect 676239 221806 676350 221811
rect 513999 221790 514065 221793
rect 513999 221788 514110 221790
rect 513999 221732 514004 221788
rect 514060 221732 514110 221788
rect 676239 221750 676244 221806
rect 676300 221750 676350 221806
rect 676239 221748 676350 221750
rect 676239 221745 676305 221748
rect 513999 221727 514110 221732
rect 513903 221660 513969 221663
rect 514050 221660 514110 221727
rect 513903 221658 514110 221660
rect 513903 221602 513908 221658
rect 513964 221602 514110 221658
rect 513903 221600 514110 221602
rect 513903 221597 513969 221600
rect 147279 221512 147345 221515
rect 143904 221510 147345 221512
rect 143904 221454 147284 221510
rect 147340 221454 147345 221510
rect 143904 221452 147345 221454
rect 147279 221449 147345 221452
rect 676143 221216 676209 221219
rect 676290 221216 676350 221482
rect 676143 221214 676350 221216
rect 676143 221158 676148 221214
rect 676204 221158 676350 221214
rect 676143 221156 676350 221158
rect 676143 221153 676209 221156
rect 186927 221068 186993 221071
rect 186927 221066 190560 221068
rect 186927 221010 186932 221066
rect 186988 221010 190560 221066
rect 186927 221008 190560 221010
rect 186927 221005 186993 221008
rect 676290 220775 676350 221038
rect 676239 220770 676350 220775
rect 676239 220714 676244 220770
rect 676300 220714 676350 220770
rect 676239 220712 676350 220714
rect 676239 220709 676305 220712
rect 676047 220624 676113 220627
rect 676047 220622 676320 220624
rect 185583 220328 185649 220331
rect 185583 220326 190560 220328
rect 185583 220270 185588 220326
rect 185644 220270 190560 220326
rect 185583 220268 190560 220270
rect 185583 220265 185649 220268
rect 143874 219736 143934 220224
rect 149487 219736 149553 219739
rect 143874 219734 149553 219736
rect 143874 219678 149492 219734
rect 149548 219678 149553 219734
rect 143874 219676 149553 219678
rect 149487 219673 149553 219676
rect 184335 219588 184401 219591
rect 184335 219586 190560 219588
rect 184335 219530 184340 219586
rect 184396 219530 190560 219586
rect 184335 219528 190560 219530
rect 184335 219525 184401 219528
rect 149391 218996 149457 218999
rect 143904 218994 149457 218996
rect 143904 218938 149396 218994
rect 149452 218938 149457 218994
rect 143904 218936 149457 218938
rect 149391 218933 149457 218936
rect 184335 218848 184401 218851
rect 184335 218846 190560 218848
rect 184335 218790 184340 218846
rect 184396 218790 190560 218846
rect 184335 218788 190560 218790
rect 184335 218785 184401 218788
rect 639810 218670 639870 220594
rect 676047 220566 676052 220622
rect 676108 220566 676320 220622
rect 676047 220564 676320 220566
rect 676047 220561 676113 220564
rect 674170 219970 674176 220034
rect 674240 220032 674246 220034
rect 674240 219972 676320 220032
rect 674240 219970 674246 219972
rect 676047 219514 676113 219517
rect 676047 219512 676320 219514
rect 676047 219456 676052 219512
rect 676108 219456 676320 219512
rect 676047 219454 676320 219456
rect 676047 219451 676113 219454
rect 672975 219144 673041 219147
rect 675322 219144 675328 219146
rect 672975 219142 675328 219144
rect 672975 219086 672980 219142
rect 673036 219086 675328 219142
rect 672975 219084 675328 219086
rect 672975 219081 673041 219084
rect 675322 219082 675328 219084
rect 675392 219144 675398 219146
rect 675392 219084 676320 219144
rect 675392 219082 675398 219084
rect 673978 218490 673984 218554
rect 674048 218552 674054 218554
rect 674048 218492 676320 218552
rect 674048 218490 674054 218492
rect 187023 218108 187089 218111
rect 187023 218106 190560 218108
rect 187023 218050 187028 218106
rect 187084 218050 190560 218106
rect 187023 218048 190560 218050
rect 187023 218045 187089 218048
rect 149391 217812 149457 217815
rect 143904 217810 149457 217812
rect 143904 217754 149396 217810
rect 149452 217754 149457 217810
rect 143904 217752 149457 217754
rect 149391 217749 149457 217752
rect 190146 217294 190206 218048
rect 672783 217960 672849 217963
rect 674362 217960 674368 217962
rect 672783 217958 674368 217960
rect 672783 217902 672788 217958
rect 672844 217902 674368 217958
rect 672783 217900 674368 217902
rect 672783 217897 672849 217900
rect 674362 217898 674368 217900
rect 674432 217960 674438 217962
rect 674432 217900 676320 217960
rect 674432 217898 674438 217900
rect 675898 217602 675904 217666
rect 675968 217664 675974 217666
rect 675968 217604 676320 217664
rect 675968 217602 675974 217604
rect 190146 217234 190560 217294
rect 676866 216779 676926 217042
rect 676866 216774 676977 216779
rect 149487 216628 149553 216631
rect 143904 216626 149553 216628
rect 143904 216570 149492 216626
rect 149548 216570 149553 216626
rect 143904 216568 149553 216570
rect 149487 216565 149553 216568
rect 186831 216480 186897 216483
rect 186831 216478 190560 216480
rect 186831 216422 186836 216478
rect 186892 216422 190560 216478
rect 186831 216420 190560 216422
rect 186831 216417 186897 216420
rect 190146 215814 190206 216420
rect 190146 215754 190560 215814
rect 143874 215000 143934 215340
rect 149391 215000 149457 215003
rect 143874 214998 149457 215000
rect 143874 214942 149396 214998
rect 149452 214942 149457 214998
rect 143874 214940 149457 214942
rect 149391 214937 149457 214940
rect 186735 215000 186801 215003
rect 186735 214998 190560 215000
rect 186735 214942 186740 214998
rect 186796 214942 190560 214998
rect 186735 214940 190560 214942
rect 186735 214937 186801 214940
rect 190146 214334 190206 214940
rect 640386 214822 640446 216746
rect 676866 216718 676916 216774
rect 676972 216718 676977 216774
rect 676866 216716 676977 216718
rect 676911 216713 676977 216716
rect 675759 216480 675825 216483
rect 675759 216478 676320 216480
rect 675759 216422 675764 216478
rect 675820 216422 676320 216478
rect 675759 216420 676320 216422
rect 675759 216417 675825 216420
rect 675706 216048 675712 216112
rect 675776 216110 675782 216112
rect 675776 216050 676320 216110
rect 675776 216048 675782 216050
rect 676090 215234 676096 215298
rect 676160 215296 676166 215298
rect 676290 215296 676350 215562
rect 676160 215236 676350 215296
rect 676160 215234 676166 215236
rect 676866 214855 676926 214970
rect 676815 214850 676926 214855
rect 676815 214794 676820 214850
rect 676876 214794 676926 214850
rect 676815 214792 676926 214794
rect 676815 214789 676881 214792
rect 676047 214630 676113 214633
rect 676047 214628 676320 214630
rect 676047 214572 676052 214628
rect 676108 214572 676320 214628
rect 676047 214570 676320 214572
rect 676047 214567 676113 214570
rect 190146 214274 190560 214334
rect 147279 214112 147345 214115
rect 143904 214110 147345 214112
rect 143904 214054 147284 214110
rect 147340 214054 147345 214110
rect 143904 214052 147345 214054
rect 147279 214049 147345 214052
rect 675951 214112 676017 214115
rect 675951 214110 676320 214112
rect 675951 214054 675956 214110
rect 676012 214054 676320 214110
rect 675951 214052 676320 214054
rect 675951 214049 676017 214052
rect 186543 213520 186609 213523
rect 186543 213518 190560 213520
rect 186543 213462 186548 213518
rect 186604 213462 190560 213518
rect 186543 213460 190560 213462
rect 186543 213457 186609 213460
rect 41775 213298 41841 213301
rect 41568 213296 41841 213298
rect 41568 213240 41780 213296
rect 41836 213240 41841 213296
rect 41568 213238 41841 213240
rect 41775 213235 41841 213238
rect 41583 212928 41649 212931
rect 146895 212928 146961 212931
rect 41538 212926 41649 212928
rect 41538 212870 41588 212926
rect 41644 212870 41649 212926
rect 41538 212865 41649 212870
rect 143904 212926 146961 212928
rect 143904 212870 146900 212926
rect 146956 212870 146961 212926
rect 143904 212868 146961 212870
rect 146895 212865 146961 212868
rect 41538 212750 41598 212865
rect 190146 212706 190206 213460
rect 675514 213458 675520 213522
rect 675584 213520 675590 213522
rect 675584 213460 676320 213520
rect 675584 213458 675590 213460
rect 674554 213014 674560 213078
rect 674624 213076 674630 213078
rect 674624 213016 676320 213076
rect 674624 213014 674630 213016
rect 190146 212646 190560 212706
rect 640194 212339 640254 212898
rect 676047 212632 676113 212635
rect 676047 212630 676320 212632
rect 676047 212574 676052 212630
rect 676108 212574 676320 212630
rect 676047 212572 676320 212574
rect 676047 212569 676113 212572
rect 640143 212334 640254 212339
rect 640143 212278 640148 212334
rect 640204 212278 640254 212334
rect 640143 212276 640254 212278
rect 640143 212273 640209 212276
rect 41775 212188 41841 212191
rect 41568 212186 41841 212188
rect 41568 212130 41780 212186
rect 41836 212130 41841 212186
rect 41568 212128 41841 212130
rect 41775 212125 41841 212128
rect 186063 212040 186129 212043
rect 676047 212040 676113 212043
rect 186063 212038 190560 212040
rect 186063 211982 186068 212038
rect 186124 211982 190560 212038
rect 186063 211980 190560 211982
rect 676047 212038 676320 212040
rect 676047 211982 676052 212038
rect 676108 211982 676320 212038
rect 676047 211980 676320 211982
rect 186063 211977 186129 211980
rect 41775 211744 41841 211747
rect 147087 211744 147153 211747
rect 41568 211742 41841 211744
rect 41568 211686 41780 211742
rect 41836 211686 41841 211742
rect 41568 211684 41841 211686
rect 143904 211742 147153 211744
rect 143904 211686 147092 211742
rect 147148 211686 147153 211742
rect 143904 211684 147153 211686
rect 41775 211681 41841 211684
rect 147087 211681 147153 211684
rect 41583 211448 41649 211451
rect 41538 211446 41649 211448
rect 41538 211390 41588 211446
rect 41644 211390 41649 211446
rect 41538 211385 41649 211390
rect 41538 211270 41598 211385
rect 190146 211152 190206 211980
rect 676047 211977 676113 211980
rect 640143 211596 640209 211599
rect 640143 211594 640254 211596
rect 640143 211538 640148 211594
rect 640204 211538 640254 211594
rect 640143 211533 640254 211538
rect 190146 211092 190560 211152
rect 640194 210974 640254 211533
rect 676290 211451 676350 211566
rect 676239 211446 676350 211451
rect 676239 211390 676244 211446
rect 676300 211390 676350 211446
rect 676239 211388 676350 211390
rect 676239 211385 676305 211388
rect 675951 211078 676017 211081
rect 675951 211076 676320 211078
rect 675951 211020 675956 211076
rect 676012 211020 676320 211076
rect 675951 211018 676320 211020
rect 675951 211015 676017 211018
rect 41775 210708 41841 210711
rect 679791 210708 679857 210711
rect 41568 210706 41841 210708
rect 41568 210650 41780 210706
rect 41836 210650 41841 210706
rect 41568 210648 41841 210650
rect 41775 210645 41841 210648
rect 679746 210706 679857 210708
rect 679746 210650 679796 210706
rect 679852 210650 679857 210706
rect 679746 210645 679857 210650
rect 186351 210560 186417 210563
rect 186351 210558 190206 210560
rect 186351 210502 186356 210558
rect 186412 210502 190206 210558
rect 679746 210530 679806 210645
rect 186351 210500 190206 210502
rect 186351 210497 186417 210500
rect 190146 210486 190206 210500
rect 190146 210426 190560 210486
rect 147471 210412 147537 210415
rect 143904 210410 147537 210412
rect 143904 210354 147476 210410
rect 147532 210354 147537 210410
rect 143904 210352 147537 210354
rect 147471 210349 147537 210352
rect 41775 210264 41841 210267
rect 41568 210262 41841 210264
rect 41568 210206 41780 210262
rect 41836 210206 41841 210262
rect 41568 210204 41841 210206
rect 41775 210201 41841 210204
rect 41583 209968 41649 209971
rect 41538 209966 41649 209968
rect 41538 209910 41588 209966
rect 41644 209910 41649 209966
rect 41538 209905 41649 209910
rect 41538 209790 41598 209905
rect 190146 209672 190206 210426
rect 685506 209823 685566 210086
rect 679791 209820 679857 209823
rect 679746 209818 679857 209820
rect 679746 209762 679796 209818
rect 679852 209762 679857 209818
rect 679746 209757 679857 209762
rect 685455 209818 685566 209823
rect 685455 209762 685460 209818
rect 685516 209762 685566 209818
rect 685455 209760 685566 209762
rect 685455 209757 685521 209760
rect 190146 209612 190560 209672
rect 679746 209568 679806 209757
rect 41583 209376 41649 209379
rect 41538 209374 41649 209376
rect 41538 209318 41588 209374
rect 41644 209318 41649 209374
rect 41538 209313 41649 209318
rect 685455 209376 685521 209379
rect 685455 209374 685566 209376
rect 685455 209318 685460 209374
rect 685516 209318 685566 209374
rect 685455 209313 685566 209318
rect 41538 209198 41598 209313
rect 146895 209228 146961 209231
rect 143904 209226 146961 209228
rect 143904 209170 146900 209226
rect 146956 209170 146961 209226
rect 143904 209168 146961 209170
rect 146895 209165 146961 209168
rect 186639 209080 186705 209083
rect 186639 209078 190206 209080
rect 186639 209022 186644 209078
rect 186700 209022 190206 209078
rect 186639 209020 190206 209022
rect 186639 209017 186705 209020
rect 190146 209006 190206 209020
rect 190146 208946 190560 209006
rect 25602 208491 25662 208754
rect 25551 208486 25662 208491
rect 25551 208430 25556 208486
rect 25612 208430 25662 208486
rect 25551 208428 25662 208430
rect 25551 208425 25617 208428
rect 25794 208047 25854 208236
rect 190146 208192 190206 208946
rect 190146 208132 190560 208192
rect 25743 208042 25854 208047
rect 147183 208044 147249 208047
rect 25743 207986 25748 208042
rect 25804 207986 25854 208042
rect 25743 207984 25854 207986
rect 143904 208042 147249 208044
rect 143904 207986 147188 208042
rect 147244 207986 147249 208042
rect 143904 207984 147249 207986
rect 25743 207981 25809 207984
rect 147183 207981 147249 207984
rect 25839 207896 25905 207899
rect 25794 207894 25905 207896
rect 25794 207838 25844 207894
rect 25900 207838 25905 207894
rect 25794 207833 25905 207838
rect 25794 207718 25854 207833
rect 190146 207318 190560 207378
rect 186255 207304 186321 207307
rect 190146 207304 190206 207318
rect 186255 207302 190206 207304
rect 40770 207158 40830 207274
rect 186255 207246 186260 207302
rect 186316 207246 190206 207302
rect 639810 207274 639870 209124
rect 685506 209050 685566 209313
rect 676666 207538 676672 207602
rect 676736 207600 676742 207602
rect 676815 207600 676881 207603
rect 676736 207598 676881 207600
rect 676736 207542 676820 207598
rect 676876 207542 676881 207598
rect 676736 207540 676881 207542
rect 676736 207538 676742 207540
rect 676815 207537 676881 207540
rect 676474 207390 676480 207454
rect 676544 207452 676550 207454
rect 676911 207452 676977 207455
rect 676544 207450 676977 207452
rect 676544 207394 676916 207450
rect 676972 207394 676977 207450
rect 676544 207392 676977 207394
rect 676544 207390 676550 207392
rect 676911 207389 676977 207392
rect 186255 207244 190206 207246
rect 186255 207241 186321 207244
rect 40762 207094 40768 207158
rect 40832 207094 40838 207158
rect 25602 206419 25662 206682
rect 25602 206414 25713 206419
rect 25602 206358 25652 206414
rect 25708 206358 25713 206414
rect 25602 206356 25713 206358
rect 143874 206416 143934 206904
rect 190146 206712 190206 207244
rect 190146 206652 190560 206712
rect 147087 206416 147153 206419
rect 143874 206414 147153 206416
rect 143874 206358 147092 206414
rect 147148 206358 147153 206414
rect 143874 206356 147153 206358
rect 25647 206353 25713 206356
rect 147087 206353 147153 206356
rect 41967 206268 42033 206271
rect 41568 206266 42033 206268
rect 41568 206210 41972 206266
rect 42028 206210 42033 206266
rect 41568 206208 42033 206210
rect 41967 206205 42033 206208
rect 186447 205972 186513 205975
rect 186447 205970 190206 205972
rect 186447 205914 186452 205970
rect 186508 205914 190206 205970
rect 186447 205912 190206 205914
rect 186447 205909 186513 205912
rect 190146 205898 190206 205912
rect 190146 205838 190560 205898
rect 41154 205530 41214 205794
rect 149391 205676 149457 205679
rect 143904 205674 149457 205676
rect 143904 205618 149396 205674
rect 149452 205618 149457 205674
rect 143904 205616 149457 205618
rect 149391 205613 149457 205616
rect 41146 205466 41152 205530
rect 41216 205466 41222 205530
rect 190146 205232 190206 205838
rect 40962 205086 41022 205202
rect 190146 205172 190560 205232
rect 40954 205022 40960 205086
rect 41024 205022 41030 205086
rect 42106 204788 42112 204790
rect 41568 204728 42112 204788
rect 42106 204726 42112 204728
rect 42176 204726 42182 204790
rect 149295 204492 149361 204495
rect 143904 204490 149361 204492
rect 143904 204434 149300 204490
rect 149356 204434 149361 204490
rect 143904 204432 149361 204434
rect 149295 204429 149361 204432
rect 185967 204344 186033 204347
rect 185967 204342 190560 204344
rect 41538 204048 41598 204314
rect 185967 204286 185972 204342
rect 186028 204286 190560 204342
rect 185967 204284 190560 204286
rect 185967 204281 186033 204284
rect 41679 204048 41745 204051
rect 41538 204046 41745 204048
rect 41538 203990 41684 204046
rect 41740 203990 41745 204046
rect 41538 203988 41745 203990
rect 41679 203985 41745 203988
rect 41775 203752 41841 203755
rect 41568 203750 41841 203752
rect 41568 203694 41780 203750
rect 41836 203694 41841 203750
rect 41568 203692 41841 203694
rect 41775 203689 41841 203692
rect 190146 203604 190206 204284
rect 190146 203544 190560 203604
rect 639810 203426 639870 205350
rect 675759 204492 675825 204495
rect 675898 204492 675904 204494
rect 675759 204490 675904 204492
rect 675759 204434 675764 204490
rect 675820 204434 675904 204490
rect 675759 204432 675904 204434
rect 675759 204429 675825 204432
rect 675898 204430 675904 204432
rect 675968 204430 675974 204494
rect 149487 203308 149553 203311
rect 143904 203306 149553 203308
rect 143904 203250 149492 203306
rect 149548 203250 149553 203306
rect 143904 203248 149553 203250
rect 149487 203245 149553 203248
rect 41914 203234 41920 203236
rect 41568 203174 41920 203234
rect 41914 203172 41920 203174
rect 41984 203172 41990 203236
rect 186159 202864 186225 202867
rect 186159 202862 190560 202864
rect 41538 202571 41598 202834
rect 186159 202806 186164 202862
rect 186220 202806 190560 202862
rect 186159 202804 190560 202806
rect 186159 202801 186225 202804
rect 41487 202566 41598 202571
rect 41487 202510 41492 202566
rect 41548 202510 41598 202566
rect 41487 202508 41598 202510
rect 41487 202505 41553 202508
rect 41538 202127 41598 202242
rect 41538 202122 41649 202127
rect 41538 202066 41588 202122
rect 41644 202066 41649 202122
rect 41538 202064 41649 202066
rect 190146 202124 190206 202804
rect 675663 202718 675729 202719
rect 675663 202714 675712 202718
rect 675776 202716 675782 202718
rect 675663 202658 675668 202714
rect 675663 202654 675712 202658
rect 675776 202656 675820 202716
rect 675776 202654 675782 202656
rect 675663 202653 675729 202654
rect 190146 202064 190560 202124
rect 41583 202061 41649 202064
rect 143874 201976 143934 202020
rect 149391 201976 149457 201979
rect 143874 201974 149457 201976
rect 143874 201918 149396 201974
rect 149452 201918 149457 201974
rect 143874 201916 149457 201918
rect 149391 201913 149457 201916
rect 41871 201680 41937 201683
rect 41568 201678 41937 201680
rect 41568 201622 41876 201678
rect 41932 201622 41937 201678
rect 41568 201620 41937 201622
rect 41871 201617 41937 201620
rect 41871 201384 41937 201387
rect 41568 201382 41937 201384
rect 41568 201326 41876 201382
rect 41932 201326 41937 201382
rect 41568 201324 41937 201326
rect 41871 201321 41937 201324
rect 190287 201384 190353 201387
rect 190287 201382 190560 201384
rect 190287 201326 190292 201382
rect 190348 201326 190560 201382
rect 190287 201324 190560 201326
rect 190287 201321 190353 201324
rect 42298 201088 42304 201090
rect 25890 201028 42304 201088
rect 25890 200943 25950 201028
rect 42298 201026 42304 201028
rect 42368 201026 42374 201090
rect 640194 200943 640254 201502
rect 675567 201386 675633 201387
rect 675514 201322 675520 201386
rect 675584 201384 675633 201386
rect 675584 201382 675676 201384
rect 675628 201326 675676 201382
rect 675584 201324 675676 201326
rect 675584 201322 675633 201324
rect 675567 201321 675633 201322
rect 25839 200938 25950 200943
rect 25839 200882 25844 200938
rect 25900 200882 25950 200938
rect 25839 200880 25950 200882
rect 41487 200940 41553 200943
rect 41487 200938 41598 200940
rect 41487 200882 41492 200938
rect 41548 200882 41598 200938
rect 25839 200877 25905 200880
rect 41487 200877 41598 200882
rect 640143 200938 640254 200943
rect 640143 200882 640148 200938
rect 640204 200882 640254 200938
rect 640143 200880 640254 200882
rect 640143 200877 640209 200880
rect 41538 200762 41598 200877
rect 149391 200792 149457 200795
rect 143904 200790 149457 200792
rect 143904 200734 149396 200790
rect 149452 200734 149457 200790
rect 143904 200732 149457 200734
rect 149391 200729 149457 200732
rect 190287 200570 190353 200573
rect 190287 200568 190560 200570
rect 190287 200512 190292 200568
rect 190348 200512 190560 200568
rect 190287 200510 190560 200512
rect 190287 200507 190353 200510
rect 25743 200496 25809 200499
rect 41722 200496 41728 200498
rect 25743 200494 41728 200496
rect 25743 200438 25748 200494
rect 25804 200438 41728 200494
rect 25743 200436 41728 200438
rect 25743 200433 25809 200436
rect 41722 200434 41728 200436
rect 41792 200434 41798 200498
rect 640143 200200 640209 200203
rect 640143 200198 640254 200200
rect 640143 200142 640148 200198
rect 640204 200142 640254 200198
rect 640143 200137 640254 200142
rect 25551 200052 25617 200055
rect 41338 200052 41344 200054
rect 25551 200050 41344 200052
rect 25551 199994 25556 200050
rect 25612 199994 41344 200050
rect 25551 199992 41344 199994
rect 25551 199989 25617 199992
rect 41338 199990 41344 199992
rect 41408 199990 41414 200054
rect 184335 199756 184401 199759
rect 184335 199754 190560 199756
rect 184335 199698 184340 199754
rect 184396 199698 190560 199754
rect 184335 199696 190560 199698
rect 184335 199693 184401 199696
rect 25647 199608 25713 199611
rect 41530 199608 41536 199610
rect 25647 199606 41536 199608
rect 25647 199550 25652 199606
rect 25708 199550 41536 199606
rect 25647 199548 41536 199550
rect 25647 199545 25713 199548
rect 41530 199546 41536 199548
rect 41600 199546 41606 199610
rect 147471 199608 147537 199611
rect 143904 199606 147537 199608
rect 143904 199550 147476 199606
rect 147532 199550 147537 199606
rect 640194 199578 640254 200137
rect 143904 199548 147537 199550
rect 147471 199545 147537 199548
rect 187215 199164 187281 199167
rect 187215 199162 190014 199164
rect 187215 199106 187220 199162
rect 187276 199106 190014 199162
rect 187215 199104 190014 199106
rect 187215 199101 187281 199104
rect 189954 199090 190014 199104
rect 189954 199030 190560 199090
rect 149487 198424 149553 198427
rect 143904 198422 149553 198424
rect 143904 198366 149492 198422
rect 149548 198366 149553 198422
rect 143904 198364 149553 198366
rect 149487 198361 149553 198364
rect 675759 198424 675825 198427
rect 676090 198424 676096 198426
rect 675759 198422 676096 198424
rect 675759 198366 675764 198422
rect 675820 198366 676096 198422
rect 675759 198364 676096 198366
rect 675759 198361 675825 198364
rect 676090 198362 676096 198364
rect 676160 198362 676166 198426
rect 185487 198276 185553 198279
rect 185487 198274 190560 198276
rect 185487 198218 185492 198274
rect 185548 198218 190560 198274
rect 185487 198216 190560 198218
rect 185487 198213 185553 198216
rect 184239 197684 184305 197687
rect 184239 197682 190014 197684
rect 184239 197626 184244 197682
rect 184300 197626 190014 197682
rect 184239 197624 190014 197626
rect 184239 197621 184305 197624
rect 189954 197610 190014 197624
rect 189954 197550 190560 197610
rect 149391 197092 149457 197095
rect 143904 197090 149457 197092
rect 143904 197034 149396 197090
rect 149452 197034 149457 197090
rect 143904 197032 149457 197034
rect 149391 197029 149457 197032
rect 184431 196796 184497 196799
rect 184431 196794 190560 196796
rect 184431 196738 184436 196794
rect 184492 196738 190560 196794
rect 184431 196736 190560 196738
rect 184431 196733 184497 196736
rect 184335 196056 184401 196059
rect 184335 196054 190560 196056
rect 184335 195998 184340 196054
rect 184396 195998 190560 196054
rect 184335 195996 190560 195998
rect 184335 195993 184401 195996
rect 149391 195908 149457 195911
rect 143904 195906 149457 195908
rect 143904 195850 149396 195906
rect 149452 195850 149457 195906
rect 143904 195848 149457 195850
rect 149391 195845 149457 195848
rect 639810 195730 639870 197654
rect 41775 195318 41841 195319
rect 41722 195316 41728 195318
rect 41684 195256 41728 195316
rect 41792 195314 41841 195318
rect 41836 195258 41841 195314
rect 41722 195254 41728 195256
rect 41792 195254 41841 195258
rect 41775 195253 41841 195254
rect 184335 195316 184401 195319
rect 184335 195314 190560 195316
rect 184335 195258 184340 195314
rect 184396 195258 190560 195314
rect 184335 195256 190560 195258
rect 184335 195253 184401 195256
rect 674554 195254 674560 195318
rect 674624 195316 674630 195318
rect 675471 195316 675537 195319
rect 674624 195314 675537 195316
rect 674624 195258 675476 195314
rect 675532 195258 675537 195314
rect 674624 195256 675537 195258
rect 674624 195254 674630 195256
rect 675471 195253 675537 195256
rect 149487 194724 149553 194727
rect 143904 194722 149553 194724
rect 143904 194666 149492 194722
rect 149548 194666 149553 194722
rect 143904 194664 149553 194666
rect 149487 194661 149553 194664
rect 184431 194428 184497 194431
rect 184431 194426 190560 194428
rect 184431 194370 184436 194426
rect 184492 194370 190560 194426
rect 184431 194368 190560 194370
rect 184431 194365 184497 194368
rect 184527 193836 184593 193839
rect 184527 193834 190014 193836
rect 184527 193778 184532 193834
rect 184588 193778 190014 193834
rect 184527 193776 190014 193778
rect 184527 193773 184593 193776
rect 189954 193762 190014 193776
rect 189954 193702 190560 193762
rect 143874 193392 143934 193436
rect 149391 193392 149457 193395
rect 143874 193390 149457 193392
rect 143874 193334 149396 193390
rect 149452 193334 149457 193390
rect 143874 193332 149457 193334
rect 149391 193329 149457 193332
rect 184431 192948 184497 192951
rect 184431 192946 190560 192948
rect 184431 192890 184436 192946
rect 184492 192890 190560 192946
rect 184431 192888 190560 192890
rect 184431 192885 184497 192888
rect 184335 192356 184401 192359
rect 184335 192354 190014 192356
rect 184335 192298 184340 192354
rect 184396 192298 190014 192354
rect 184335 192296 190014 192298
rect 184335 192293 184401 192296
rect 189954 192282 190014 192296
rect 189954 192222 190560 192282
rect 149391 192208 149457 192211
rect 143904 192206 149457 192208
rect 143904 192150 149396 192206
rect 149452 192150 149457 192206
rect 143904 192148 149457 192150
rect 149391 192145 149457 192148
rect 639810 192030 639870 193880
rect 675759 193540 675825 193543
rect 676474 193540 676480 193542
rect 675759 193538 676480 193540
rect 675759 193482 675764 193538
rect 675820 193482 676480 193538
rect 675759 193480 676480 193482
rect 675759 193477 675825 193480
rect 676474 193478 676480 193480
rect 676544 193478 676550 193542
rect 675759 191616 675825 191619
rect 676666 191616 676672 191618
rect 675759 191614 676672 191616
rect 675759 191558 675764 191614
rect 675820 191558 676672 191614
rect 675759 191556 676672 191558
rect 675759 191553 675825 191556
rect 676666 191554 676672 191556
rect 676736 191554 676742 191618
rect 184527 191468 184593 191471
rect 184527 191466 190560 191468
rect 184527 191410 184532 191466
rect 184588 191410 190560 191466
rect 184527 191408 190560 191410
rect 184527 191405 184593 191408
rect 147375 191024 147441 191027
rect 143904 191022 147441 191024
rect 143904 190966 147380 191022
rect 147436 190966 147441 191022
rect 143904 190964 147441 190966
rect 147375 190961 147441 190964
rect 184623 190728 184689 190731
rect 184623 190726 190014 190728
rect 184623 190670 184628 190726
rect 184684 190670 190014 190726
rect 184623 190668 190014 190670
rect 184623 190665 184689 190668
rect 189954 190654 190014 190668
rect 189954 190594 190560 190654
rect 41530 190074 41536 190138
rect 41600 190136 41606 190138
rect 41775 190136 41841 190139
rect 41600 190134 41841 190136
rect 41600 190078 41780 190134
rect 41836 190078 41841 190134
rect 41600 190076 41841 190078
rect 41600 190074 41606 190076
rect 41775 190073 41841 190076
rect 184335 189988 184401 189991
rect 184335 189986 190560 189988
rect 184335 189930 184340 189986
rect 184396 189930 190560 189986
rect 184335 189928 190560 189930
rect 184335 189925 184401 189928
rect 149391 189840 149457 189843
rect 143904 189838 149457 189840
rect 143904 189782 149396 189838
rect 149452 189782 149457 189838
rect 143904 189780 149457 189782
rect 149391 189777 149457 189780
rect 184527 189248 184593 189251
rect 184527 189246 190014 189248
rect 184527 189190 184532 189246
rect 184588 189190 190014 189246
rect 184527 189188 190014 189190
rect 184527 189185 184593 189188
rect 189954 189174 190014 189188
rect 189954 189114 190560 189174
rect 143874 188064 143934 188552
rect 184335 188508 184401 188511
rect 184335 188506 190560 188508
rect 184335 188450 184340 188506
rect 184396 188450 190560 188506
rect 184335 188448 190560 188450
rect 184335 188445 184401 188448
rect 639810 188182 639870 190106
rect 149487 188064 149553 188067
rect 143874 188062 149553 188064
rect 143874 188006 149492 188062
rect 149548 188006 149553 188062
rect 143874 188004 149553 188006
rect 149487 188001 149553 188004
rect 41871 187918 41937 187919
rect 41871 187914 41920 187918
rect 41984 187916 41990 187918
rect 41871 187858 41876 187914
rect 41871 187854 41920 187858
rect 41984 187856 42028 187916
rect 41984 187854 41990 187856
rect 41871 187853 41937 187854
rect 184431 187620 184497 187623
rect 184431 187618 190560 187620
rect 184431 187562 184436 187618
rect 184492 187562 190560 187618
rect 184431 187560 190560 187562
rect 184431 187557 184497 187560
rect 149295 187472 149361 187475
rect 143904 187470 149361 187472
rect 143904 187414 149300 187470
rect 149356 187414 149361 187470
rect 143904 187412 149361 187414
rect 149295 187409 149361 187412
rect 42159 187178 42225 187179
rect 42106 187176 42112 187178
rect 42068 187116 42112 187176
rect 42176 187174 42225 187178
rect 42220 187118 42225 187174
rect 42106 187114 42112 187116
rect 42176 187114 42225 187118
rect 42159 187113 42225 187114
rect 184335 186880 184401 186883
rect 184335 186878 190560 186880
rect 184335 186822 184340 186878
rect 184396 186822 190560 186878
rect 184335 186820 190560 186822
rect 184335 186817 184401 186820
rect 40954 186374 40960 186438
rect 41024 186436 41030 186438
rect 41775 186436 41841 186439
rect 41024 186434 41841 186436
rect 41024 186378 41780 186434
rect 41836 186378 41841 186434
rect 41024 186376 41841 186378
rect 41024 186374 41030 186376
rect 41775 186373 41841 186376
rect 149199 186288 149265 186291
rect 143904 186286 149265 186288
rect 143904 186230 149204 186286
rect 149260 186230 149265 186286
rect 143904 186228 149265 186230
rect 149199 186225 149265 186228
rect 184431 186140 184497 186143
rect 184431 186138 190560 186140
rect 184431 186082 184436 186138
rect 184492 186082 190560 186138
rect 184431 186080 190560 186082
rect 184431 186077 184497 186080
rect 40762 185782 40768 185846
rect 40832 185844 40838 185846
rect 41775 185844 41841 185847
rect 40832 185842 41841 185844
rect 40832 185786 41780 185842
rect 41836 185786 41841 185842
rect 40832 185784 41841 185786
rect 40832 185782 40838 185784
rect 41775 185781 41841 185784
rect 640194 185699 640254 186258
rect 640194 185694 640305 185699
rect 640194 185638 640244 185694
rect 640300 185638 640305 185694
rect 640194 185636 640305 185638
rect 640239 185633 640305 185636
rect 184623 185400 184689 185403
rect 184623 185398 190014 185400
rect 184623 185342 184628 185398
rect 184684 185342 190014 185398
rect 184623 185340 190014 185342
rect 184623 185337 184689 185340
rect 189954 185326 190014 185340
rect 189954 185266 190560 185326
rect 143874 184512 143934 185000
rect 640239 184956 640305 184959
rect 640194 184954 640305 184956
rect 640194 184898 640244 184954
rect 640300 184898 640305 184954
rect 640194 184893 640305 184898
rect 184527 184660 184593 184663
rect 184527 184658 190560 184660
rect 184527 184602 184532 184658
rect 184588 184602 190560 184658
rect 184527 184600 190560 184602
rect 184527 184597 184593 184600
rect 149583 184512 149649 184515
rect 143874 184510 149649 184512
rect 143874 184454 149588 184510
rect 149644 184454 149649 184510
rect 143874 184452 149649 184454
rect 149583 184449 149649 184452
rect 640194 184334 640254 184893
rect 41338 184154 41344 184218
rect 41408 184216 41414 184218
rect 41775 184216 41841 184219
rect 41408 184214 41841 184216
rect 41408 184158 41780 184214
rect 41836 184158 41841 184214
rect 41408 184156 41841 184158
rect 41408 184154 41414 184156
rect 41775 184153 41841 184156
rect 184335 183920 184401 183923
rect 184335 183918 190014 183920
rect 184335 183862 184340 183918
rect 184396 183862 190014 183918
rect 184335 183860 190014 183862
rect 184335 183857 184401 183860
rect 189954 183846 190014 183860
rect 189954 183786 190560 183846
rect 149391 183772 149457 183775
rect 143904 183770 149457 183772
rect 143904 183714 149396 183770
rect 149452 183714 149457 183770
rect 143904 183712 149457 183714
rect 149391 183709 149457 183712
rect 41146 183414 41152 183478
rect 41216 183476 41222 183478
rect 41775 183476 41841 183479
rect 41216 183474 41841 183476
rect 41216 183418 41780 183474
rect 41836 183418 41841 183474
rect 41216 183416 41841 183418
rect 41216 183414 41222 183416
rect 41775 183413 41841 183416
rect 186735 183180 186801 183183
rect 186735 183178 190560 183180
rect 186735 183122 186740 183178
rect 186796 183122 190560 183178
rect 186735 183120 190560 183122
rect 186735 183117 186801 183120
rect 42063 183032 42129 183035
rect 42298 183032 42304 183034
rect 42063 183030 42304 183032
rect 42063 182974 42068 183030
rect 42124 182974 42304 183030
rect 42063 182972 42304 182974
rect 42063 182969 42129 182972
rect 42298 182970 42304 182972
rect 42368 182970 42374 183034
rect 645135 183032 645201 183035
rect 640386 183030 645201 183032
rect 640386 182974 645140 183030
rect 645196 182974 645201 183030
rect 640386 182972 645201 182974
rect 149487 182588 149553 182591
rect 143904 182586 149553 182588
rect 143904 182530 149492 182586
rect 149548 182530 149553 182586
rect 143904 182528 149553 182530
rect 149487 182525 149553 182528
rect 185775 182440 185841 182443
rect 640386 182440 640446 182972
rect 645135 182969 645201 182972
rect 185775 182438 190014 182440
rect 185775 182382 185780 182438
rect 185836 182382 190014 182438
rect 640224 182410 640446 182440
rect 185775 182380 190014 182382
rect 185775 182377 185841 182380
rect 189954 182366 190014 182380
rect 640194 182380 640416 182410
rect 189954 182306 190560 182366
rect 184431 181552 184497 181555
rect 184431 181550 190560 181552
rect 184431 181494 184436 181550
rect 184492 181494 190560 181550
rect 184431 181492 190560 181494
rect 184431 181489 184497 181492
rect 149295 181404 149361 181407
rect 143904 181402 149361 181404
rect 143904 181346 149300 181402
rect 149356 181346 149361 181402
rect 143904 181344 149361 181346
rect 149295 181341 149361 181344
rect 184335 180812 184401 180815
rect 184335 180810 190560 180812
rect 184335 180754 184340 180810
rect 184396 180754 190560 180810
rect 184335 180752 190560 180754
rect 184335 180749 184401 180752
rect 640194 180560 640254 182380
rect 143874 179628 143934 180116
rect 184431 180072 184497 180075
rect 184431 180070 190560 180072
rect 184431 180014 184436 180070
rect 184492 180014 190560 180070
rect 184431 180012 190560 180014
rect 184431 180009 184497 180012
rect 149487 179628 149553 179631
rect 143874 179626 149553 179628
rect 143874 179570 149492 179626
rect 149548 179570 149553 179626
rect 143874 179568 149553 179570
rect 149487 179565 149553 179568
rect 184623 179332 184689 179335
rect 645135 179332 645201 179335
rect 184623 179330 190560 179332
rect 184623 179274 184628 179330
rect 184684 179274 190560 179330
rect 184623 179272 190560 179274
rect 640194 179330 645201 179332
rect 640194 179274 645140 179330
rect 645196 179274 645201 179330
rect 640194 179272 645201 179274
rect 184623 179269 184689 179272
rect 149391 178888 149457 178891
rect 143904 178886 149457 178888
rect 143904 178830 149396 178886
rect 149452 178830 149457 178886
rect 143904 178828 149457 178830
rect 149391 178825 149457 178828
rect 184527 178592 184593 178595
rect 184527 178590 190560 178592
rect 184527 178534 184532 178590
rect 184588 178534 190560 178590
rect 184527 178532 190560 178534
rect 184527 178529 184593 178532
rect 149391 177704 149457 177707
rect 143904 177702 149457 177704
rect 143904 177646 149396 177702
rect 149452 177646 149457 177702
rect 143904 177644 149457 177646
rect 149391 177641 149457 177644
rect 184431 177704 184497 177707
rect 184431 177702 190560 177704
rect 184431 177646 184436 177702
rect 184492 177646 190560 177702
rect 184431 177644 190560 177646
rect 184431 177641 184497 177644
rect 184335 177112 184401 177115
rect 184335 177110 190014 177112
rect 184335 177054 184340 177110
rect 184396 177054 190014 177110
rect 184335 177052 190014 177054
rect 184335 177049 184401 177052
rect 189954 177038 190014 177052
rect 189954 176978 190560 177038
rect 640194 176786 640254 179272
rect 645135 179269 645201 179272
rect 676290 177411 676350 177674
rect 676290 177406 676401 177411
rect 676290 177350 676340 177406
rect 676396 177350 676401 177406
rect 676290 177348 676401 177350
rect 676335 177345 676401 177348
rect 676143 176816 676209 176819
rect 676290 176816 676350 177082
rect 676143 176814 676350 176816
rect 676143 176758 676148 176814
rect 676204 176758 676350 176814
rect 676143 176756 676350 176758
rect 676143 176753 676209 176756
rect 147759 176520 147825 176523
rect 143904 176518 147825 176520
rect 143904 176462 147764 176518
rect 147820 176462 147825 176518
rect 143904 176460 147825 176462
rect 147759 176457 147825 176460
rect 676290 176375 676350 176638
rect 676239 176370 676350 176375
rect 676239 176314 676244 176370
rect 676300 176314 676350 176370
rect 676239 176312 676350 176314
rect 676239 176309 676305 176312
rect 184527 176224 184593 176227
rect 184527 176222 190560 176224
rect 184527 176166 184532 176222
rect 184588 176166 190560 176222
rect 184527 176164 190560 176166
rect 184527 176161 184593 176164
rect 674170 176162 674176 176226
rect 674240 176224 674246 176226
rect 674240 176164 676320 176224
rect 674240 176162 674246 176164
rect 184335 175632 184401 175635
rect 184335 175630 190014 175632
rect 184335 175574 184340 175630
rect 184396 175574 190014 175630
rect 184335 175572 190014 175574
rect 184335 175569 184401 175572
rect 189954 175558 190014 175572
rect 674554 175570 674560 175634
rect 674624 175632 674630 175634
rect 674624 175572 676320 175632
rect 674624 175570 674630 175572
rect 189954 175498 190560 175558
rect 675322 175422 675328 175486
rect 675392 175484 675398 175486
rect 675392 175424 676350 175484
rect 675392 175422 675398 175424
rect 149391 175188 149457 175191
rect 143904 175186 149457 175188
rect 143904 175130 149396 175186
rect 149452 175130 149457 175186
rect 143904 175128 149457 175130
rect 149391 175125 149457 175128
rect 676290 175084 676350 175424
rect 645135 174892 645201 174895
rect 640416 174890 645201 174892
rect 640416 174862 645140 174890
rect 640386 174834 645140 174862
rect 645196 174834 645201 174890
rect 640386 174832 645201 174834
rect 185679 174744 185745 174747
rect 185679 174742 190560 174744
rect 185679 174686 185684 174742
rect 185740 174686 190560 174742
rect 185679 174684 190560 174686
rect 185679 174681 185745 174684
rect 149103 174004 149169 174007
rect 143904 174002 149169 174004
rect 143904 173946 149108 174002
rect 149164 173946 149169 174002
rect 143904 173944 149169 173946
rect 149103 173941 149169 173944
rect 184431 174004 184497 174007
rect 184431 174002 190014 174004
rect 184431 173946 184436 174002
rect 184492 173946 190014 174002
rect 184431 173944 190014 173946
rect 184431 173941 184497 173944
rect 189954 173930 190014 173944
rect 189954 173870 190560 173930
rect 186351 173264 186417 173267
rect 186351 173262 190560 173264
rect 186351 173206 186356 173262
rect 186412 173206 190560 173262
rect 186351 173204 190560 173206
rect 186351 173201 186417 173204
rect 640386 172938 640446 174832
rect 645135 174829 645201 174832
rect 672399 174744 672465 174747
rect 673978 174744 673984 174746
rect 672399 174742 673984 174744
rect 672399 174686 672404 174742
rect 672460 174686 673984 174742
rect 672399 174684 673984 174686
rect 672399 174681 672465 174684
rect 673978 174682 673984 174684
rect 674048 174744 674054 174746
rect 674048 174684 676320 174744
rect 674048 174682 674054 174684
rect 674362 174090 674368 174154
rect 674432 174152 674438 174154
rect 674432 174092 676320 174152
rect 674432 174090 674438 174092
rect 672591 173560 672657 173563
rect 674170 173560 674176 173562
rect 672591 173558 674176 173560
rect 672591 173502 672596 173558
rect 672652 173502 674176 173558
rect 672591 173500 674176 173502
rect 672591 173497 672657 173500
rect 674170 173498 674176 173500
rect 674240 173560 674246 173562
rect 674240 173500 676320 173560
rect 674240 173498 674246 173500
rect 676290 172970 676350 173234
rect 676282 172906 676288 172970
rect 676352 172906 676358 172970
rect 149583 172820 149649 172823
rect 143904 172818 149649 172820
rect 143904 172762 149588 172818
rect 149644 172762 149649 172818
rect 143904 172760 149649 172762
rect 149583 172757 149649 172760
rect 674746 172610 674752 172674
rect 674816 172672 674822 172674
rect 674816 172612 676320 172672
rect 674816 172610 674822 172612
rect 184527 172524 184593 172527
rect 184527 172522 190014 172524
rect 184527 172466 184532 172522
rect 184588 172466 190014 172522
rect 184527 172464 190014 172466
rect 184527 172461 184593 172464
rect 189954 172450 190014 172464
rect 189954 172390 190560 172450
rect 676290 171935 676350 172050
rect 676239 171930 676350 171935
rect 676239 171874 676244 171930
rect 676300 171874 676350 171930
rect 676239 171872 676350 171874
rect 676239 171869 676305 171872
rect 184335 171784 184401 171787
rect 184335 171782 190560 171784
rect 184335 171726 184340 171782
rect 184396 171726 190560 171782
rect 184335 171724 190560 171726
rect 184335 171721 184401 171724
rect 675706 171648 675712 171712
rect 675776 171710 675782 171712
rect 675776 171650 676320 171710
rect 675776 171648 675782 171650
rect 143874 171044 143934 171532
rect 675322 171130 675328 171194
rect 675392 171192 675398 171194
rect 675392 171132 676320 171192
rect 675392 171130 675398 171132
rect 149487 171044 149553 171047
rect 645135 171044 645201 171047
rect 143874 171042 149553 171044
rect 143874 170986 149492 171042
rect 149548 170986 149553 171042
rect 640416 171042 645201 171044
rect 640416 171014 645140 171042
rect 143874 170984 149553 170986
rect 149487 170981 149553 170984
rect 640386 170986 645140 171014
rect 645196 170986 645201 171042
rect 640386 170984 645201 170986
rect 184431 170896 184497 170899
rect 184431 170894 190560 170896
rect 184431 170838 184436 170894
rect 184492 170838 190560 170894
rect 184431 170836 190560 170838
rect 184431 170833 184497 170836
rect 149007 170304 149073 170307
rect 143904 170302 149073 170304
rect 143904 170246 149012 170302
rect 149068 170246 149073 170302
rect 143904 170244 149073 170246
rect 149007 170241 149073 170244
rect 184623 170304 184689 170307
rect 184623 170302 190014 170304
rect 184623 170246 184628 170302
rect 184684 170246 190014 170302
rect 184623 170244 190014 170246
rect 184623 170241 184689 170244
rect 189954 170230 190014 170244
rect 189954 170170 190560 170230
rect 184335 169416 184401 169419
rect 184335 169414 190560 169416
rect 184335 169358 184340 169414
rect 184396 169358 190560 169414
rect 184335 169356 190560 169358
rect 184335 169353 184401 169356
rect 148527 169120 148593 169123
rect 143904 169118 148593 169120
rect 143904 169062 148532 169118
rect 148588 169062 148593 169118
rect 640386 169090 640446 170984
rect 645135 170981 645201 170984
rect 676090 170390 676096 170454
rect 676160 170452 676166 170454
rect 676290 170452 676350 170570
rect 676160 170392 676350 170452
rect 676160 170390 676166 170392
rect 676047 170230 676113 170233
rect 676047 170228 676320 170230
rect 676047 170172 676052 170228
rect 676108 170172 676320 170228
rect 676047 170170 676320 170172
rect 676047 170167 676113 170170
rect 676047 169712 676113 169715
rect 676047 169710 676320 169712
rect 676047 169654 676052 169710
rect 676108 169654 676320 169710
rect 676047 169652 676320 169654
rect 676047 169649 676113 169652
rect 143904 169060 148593 169062
rect 148527 169057 148593 169060
rect 676290 168975 676350 169090
rect 676239 168970 676350 168975
rect 676239 168914 676244 168970
rect 676300 168914 676350 168970
rect 676239 168912 676350 168914
rect 676239 168909 676305 168912
rect 184527 168676 184593 168679
rect 184527 168674 190014 168676
rect 184527 168618 184532 168674
rect 184588 168618 190014 168674
rect 184527 168616 190014 168618
rect 184527 168613 184593 168616
rect 189954 168602 190014 168616
rect 674938 168614 674944 168678
rect 675008 168676 675014 168678
rect 675008 168616 676320 168676
rect 675008 168614 675014 168616
rect 189954 168542 190560 168602
rect 675514 168170 675520 168234
rect 675584 168232 675590 168234
rect 675584 168172 676320 168232
rect 675584 168170 675590 168172
rect 148335 168084 148401 168087
rect 143904 168082 148401 168084
rect 143904 168026 148340 168082
rect 148396 168026 148401 168082
rect 143904 168024 148401 168026
rect 148335 168021 148401 168024
rect 184431 167936 184497 167939
rect 184431 167934 190560 167936
rect 184431 167878 184436 167934
rect 184492 167878 190560 167934
rect 184431 167876 190560 167878
rect 184431 167873 184497 167876
rect 645135 167788 645201 167791
rect 640386 167786 645201 167788
rect 640386 167730 645140 167786
rect 645196 167730 645201 167786
rect 640386 167728 645201 167730
rect 184623 167196 184689 167199
rect 184623 167194 190014 167196
rect 184623 167138 184628 167194
rect 184684 167138 190014 167194
rect 184623 167136 190014 167138
rect 184623 167133 184689 167136
rect 189954 167122 190014 167136
rect 189954 167062 190560 167122
rect 143874 166308 143934 166796
rect 184335 166456 184401 166459
rect 184335 166454 190560 166456
rect 184335 166398 184340 166454
rect 184396 166398 190560 166454
rect 184335 166396 190560 166398
rect 184335 166393 184401 166396
rect 148431 166308 148497 166311
rect 143874 166306 148497 166308
rect 143874 166250 148436 166306
rect 148492 166250 148497 166306
rect 143874 166248 148497 166250
rect 148431 166245 148497 166248
rect 640386 166012 640446 167728
rect 645135 167725 645201 167728
rect 675898 167578 675904 167642
rect 675968 167640 675974 167642
rect 675968 167580 676320 167640
rect 675968 167578 675974 167580
rect 675130 167134 675136 167198
rect 675200 167196 675206 167198
rect 675200 167136 676320 167196
rect 675200 167134 675206 167136
rect 676047 166678 676113 166681
rect 676047 166676 676320 166678
rect 676047 166620 676052 166676
rect 676108 166620 676320 166676
rect 676047 166618 676320 166620
rect 676047 166615 676113 166618
rect 676047 166160 676113 166163
rect 676047 166158 676320 166160
rect 676047 166102 676052 166158
rect 676108 166102 676320 166158
rect 676047 166100 676320 166102
rect 676047 166097 676113 166100
rect 640194 165952 640446 166012
rect 184431 165716 184497 165719
rect 184431 165714 190014 165716
rect 184431 165658 184436 165714
rect 184492 165658 190014 165714
rect 184431 165656 190014 165658
rect 184431 165653 184497 165656
rect 189954 165642 190014 165656
rect 189954 165582 190560 165642
rect 148719 165568 148785 165571
rect 143904 165566 148785 165568
rect 143904 165510 148724 165566
rect 148780 165510 148785 165566
rect 143904 165508 148785 165510
rect 148719 165505 148785 165508
rect 640194 165242 640254 165952
rect 676143 165568 676209 165571
rect 676290 165568 676350 165686
rect 676143 165566 676350 165568
rect 676143 165510 676148 165566
rect 676204 165510 676350 165566
rect 676143 165508 676350 165510
rect 676143 165505 676209 165508
rect 676290 164979 676350 165168
rect 676239 164974 676350 164979
rect 676239 164918 676244 164974
rect 676300 164918 676350 164974
rect 676239 164916 676350 164918
rect 676239 164913 676305 164916
rect 184527 164828 184593 164831
rect 184527 164826 190560 164828
rect 184527 164770 184532 164826
rect 184588 164770 190560 164826
rect 184527 164768 190560 164770
rect 184527 164765 184593 164768
rect 148239 164384 148305 164387
rect 143904 164382 148305 164384
rect 143904 164326 148244 164382
rect 148300 164326 148305 164382
rect 143904 164324 148305 164326
rect 148239 164321 148305 164324
rect 184335 164088 184401 164091
rect 184335 164086 190560 164088
rect 184335 164030 184340 164086
rect 184396 164030 190560 164086
rect 184335 164028 190560 164030
rect 184335 164025 184401 164028
rect 184527 163348 184593 163351
rect 645135 163348 645201 163351
rect 184527 163346 190560 163348
rect 184527 163290 184532 163346
rect 184588 163290 190560 163346
rect 640416 163346 645201 163348
rect 640416 163318 645140 163346
rect 184527 163288 190560 163290
rect 640386 163290 645140 163318
rect 645196 163290 645201 163346
rect 640386 163288 645201 163290
rect 184527 163285 184593 163288
rect 148911 163200 148977 163203
rect 143904 163198 148977 163200
rect 143904 163142 148916 163198
rect 148972 163142 148977 163198
rect 143904 163140 148977 163142
rect 148911 163137 148977 163140
rect 184335 162608 184401 162611
rect 184335 162606 190560 162608
rect 184335 162550 184340 162606
rect 184396 162550 190560 162606
rect 184335 162548 190560 162550
rect 184335 162545 184401 162548
rect 148623 161868 148689 161871
rect 143904 161866 148689 161868
rect 143904 161810 148628 161866
rect 148684 161810 148689 161866
rect 143904 161808 148689 161810
rect 148623 161805 148689 161808
rect 184431 161868 184497 161871
rect 184431 161866 190560 161868
rect 184431 161810 184436 161866
rect 184492 161810 190560 161866
rect 184431 161808 190560 161810
rect 184431 161805 184497 161808
rect 640386 161394 640446 163288
rect 645135 163285 645201 163288
rect 184431 160980 184497 160983
rect 184431 160978 190560 160980
rect 184431 160922 184436 160978
rect 184492 160922 190560 160978
rect 184431 160920 190560 160922
rect 184431 160917 184497 160920
rect 148815 160684 148881 160687
rect 143904 160682 148881 160684
rect 143904 160626 148820 160682
rect 148876 160626 148881 160682
rect 143904 160624 148881 160626
rect 148815 160621 148881 160624
rect 184527 160388 184593 160391
rect 184527 160386 190014 160388
rect 184527 160330 184532 160386
rect 184588 160330 190014 160386
rect 184527 160328 190014 160330
rect 184527 160325 184593 160328
rect 189954 160314 190014 160328
rect 189954 160254 190560 160314
rect 147471 159500 147537 159503
rect 143904 159498 147537 159500
rect 143904 159442 147476 159498
rect 147532 159442 147537 159498
rect 143904 159440 147537 159442
rect 147471 159437 147537 159440
rect 184335 159500 184401 159503
rect 645135 159500 645201 159503
rect 184335 159498 190560 159500
rect 184335 159442 184340 159498
rect 184396 159442 190560 159498
rect 640416 159498 645201 159500
rect 640416 159470 645140 159498
rect 184335 159440 190560 159442
rect 640386 159442 645140 159470
rect 645196 159442 645201 159498
rect 640386 159440 645201 159442
rect 184335 159437 184401 159440
rect 184623 158908 184689 158911
rect 184623 158906 190014 158908
rect 184623 158850 184628 158906
rect 184684 158850 190014 158906
rect 184623 158848 190014 158850
rect 184623 158845 184689 158848
rect 189954 158834 190014 158848
rect 189954 158774 190560 158834
rect 143874 157724 143934 158212
rect 184335 158020 184401 158023
rect 184335 158018 190560 158020
rect 184335 157962 184340 158018
rect 184396 157962 190560 158018
rect 184335 157960 190560 157962
rect 184335 157957 184401 157960
rect 149295 157724 149361 157727
rect 143874 157722 149361 157724
rect 143874 157666 149300 157722
rect 149356 157666 149361 157722
rect 143874 157664 149361 157666
rect 149295 157661 149361 157664
rect 640386 157546 640446 159440
rect 645135 159437 645201 159440
rect 675759 159352 675825 159355
rect 676282 159352 676288 159354
rect 675759 159350 676288 159352
rect 675759 159294 675764 159350
rect 675820 159294 676288 159350
rect 675759 159292 676288 159294
rect 675759 159289 675825 159292
rect 676282 159290 676288 159292
rect 676352 159290 676358 159354
rect 675759 157726 675825 157727
rect 675706 157662 675712 157726
rect 675776 157724 675825 157726
rect 675776 157722 675868 157724
rect 675820 157666 675868 157722
rect 675776 157664 675868 157666
rect 675776 157662 675825 157664
rect 675759 157661 675825 157662
rect 184431 157428 184497 157431
rect 184431 157426 190014 157428
rect 184431 157370 184436 157426
rect 184492 157370 190014 157426
rect 184431 157368 190014 157370
rect 184431 157365 184497 157368
rect 189954 157354 190014 157368
rect 189954 157294 190560 157354
rect 146895 156984 146961 156987
rect 143904 156982 146961 156984
rect 143904 156926 146900 156982
rect 146956 156926 146961 156982
rect 143904 156924 146961 156926
rect 146895 156921 146961 156924
rect 184527 156540 184593 156543
rect 184527 156538 190560 156540
rect 184527 156482 184532 156538
rect 184588 156482 190560 156538
rect 184527 156480 190560 156482
rect 184527 156477 184593 156480
rect 149391 155800 149457 155803
rect 143904 155798 149457 155800
rect 143904 155742 149396 155798
rect 149452 155742 149457 155798
rect 143904 155740 149457 155742
rect 149391 155737 149457 155740
rect 184623 155652 184689 155655
rect 184623 155650 190560 155652
rect 184623 155594 184628 155650
rect 184684 155594 190560 155650
rect 184623 155592 190560 155594
rect 184623 155589 184689 155592
rect 640194 155504 640254 155622
rect 645135 155504 645201 155507
rect 640194 155502 645201 155504
rect 640194 155446 645140 155502
rect 645196 155446 645201 155502
rect 640194 155444 645201 155446
rect 184335 155060 184401 155063
rect 184335 155058 190560 155060
rect 184335 155002 184340 155058
rect 184396 155002 190560 155058
rect 184335 155000 190560 155002
rect 184335 154997 184401 155000
rect 149295 154616 149361 154619
rect 143904 154614 149361 154616
rect 143904 154558 149300 154614
rect 149356 154558 149361 154614
rect 143904 154556 149361 154558
rect 149295 154553 149361 154556
rect 184431 154172 184497 154175
rect 184431 154170 190560 154172
rect 184431 154114 184436 154170
rect 184492 154114 190560 154170
rect 184431 154112 190560 154114
rect 184431 154109 184497 154112
rect 640386 153772 640446 155444
rect 645135 155441 645201 155444
rect 675759 155504 675825 155507
rect 675898 155504 675904 155506
rect 675759 155502 675904 155504
rect 675759 155446 675764 155502
rect 675820 155446 675904 155502
rect 675759 155444 675904 155446
rect 675759 155441 675825 155444
rect 675898 155442 675904 155444
rect 675968 155442 675974 155506
rect 184527 153580 184593 153583
rect 184527 153578 190014 153580
rect 184527 153522 184532 153578
rect 184588 153522 190014 153578
rect 184527 153520 190014 153522
rect 184527 153517 184593 153520
rect 189954 153506 190014 153520
rect 189954 153446 190560 153506
rect 675322 153370 675328 153434
rect 675392 153432 675398 153434
rect 675471 153432 675537 153435
rect 675392 153430 675537 153432
rect 675392 153374 675476 153430
rect 675532 153374 675537 153430
rect 675392 153372 675537 153374
rect 675392 153370 675398 153372
rect 675471 153369 675537 153372
rect 143874 153136 143934 153328
rect 149391 153136 149457 153139
rect 143874 153134 149457 153136
rect 143874 153078 149396 153134
rect 149452 153078 149457 153134
rect 143874 153076 149457 153078
rect 149391 153073 149457 153076
rect 184623 152692 184689 152695
rect 184623 152690 190560 152692
rect 184623 152634 184628 152690
rect 184684 152634 190560 152690
rect 184623 152632 190560 152634
rect 184623 152629 184689 152632
rect 645135 152544 645201 152547
rect 640194 152542 645201 152544
rect 640194 152486 645140 152542
rect 645196 152486 645201 152542
rect 640194 152484 645201 152486
rect 149199 152100 149265 152103
rect 143904 152098 149265 152100
rect 143904 152042 149204 152098
rect 149260 152042 149265 152098
rect 143904 152040 149265 152042
rect 149199 152037 149265 152040
rect 184335 151952 184401 151955
rect 184335 151950 190014 151952
rect 184335 151894 184340 151950
rect 184396 151894 190014 151950
rect 184335 151892 190014 151894
rect 184335 151889 184401 151892
rect 189954 151878 190014 151892
rect 189954 151818 190560 151878
rect 184431 151212 184497 151215
rect 184431 151210 190560 151212
rect 184431 151154 184436 151210
rect 184492 151154 190560 151210
rect 184431 151152 190560 151154
rect 184431 151149 184497 151152
rect 149391 150916 149457 150919
rect 143904 150914 149457 150916
rect 143904 150858 149396 150914
rect 149452 150858 149457 150914
rect 143904 150856 149457 150858
rect 149391 150853 149457 150856
rect 184527 150472 184593 150475
rect 184527 150470 190014 150472
rect 184527 150414 184532 150470
rect 184588 150414 190014 150470
rect 184527 150412 190014 150414
rect 184527 150409 184593 150412
rect 189954 150398 190014 150412
rect 189954 150338 190560 150398
rect 640194 149998 640254 152484
rect 645135 152481 645201 152484
rect 675130 152482 675136 152546
rect 675200 152544 675206 152546
rect 675375 152544 675441 152547
rect 675200 152542 675441 152544
rect 675200 152486 675380 152542
rect 675436 152486 675441 152542
rect 675200 152484 675441 152486
rect 675200 152482 675206 152484
rect 675375 152481 675441 152484
rect 675471 152250 675537 152251
rect 675471 152246 675520 152250
rect 675584 152248 675590 152250
rect 675471 152190 675476 152246
rect 675471 152186 675520 152190
rect 675584 152188 675628 152248
rect 675584 152186 675590 152188
rect 675471 152185 675537 152186
rect 674938 150262 674944 150326
rect 675008 150324 675014 150326
rect 675471 150324 675537 150327
rect 675008 150322 675537 150324
rect 675008 150266 675476 150322
rect 675532 150266 675537 150322
rect 675008 150264 675537 150266
rect 675008 150262 675014 150264
rect 675471 150261 675537 150264
rect 149295 149880 149361 149883
rect 143874 149878 149361 149880
rect 143874 149822 149300 149878
rect 149356 149822 149361 149878
rect 143874 149820 149361 149822
rect 143874 149776 143934 149820
rect 149295 149817 149361 149820
rect 184335 149732 184401 149735
rect 184335 149730 190560 149732
rect 184335 149674 184340 149730
rect 184396 149674 190560 149730
rect 184335 149672 190560 149674
rect 184335 149669 184401 149672
rect 184431 148992 184497 148995
rect 184431 148990 190014 148992
rect 184431 148934 184436 148990
rect 184492 148934 190014 148990
rect 184431 148932 190014 148934
rect 184431 148929 184497 148932
rect 189954 148918 190014 148932
rect 189954 148858 190560 148918
rect 149295 148548 149361 148551
rect 143904 148546 149361 148548
rect 143904 148490 149300 148546
rect 149356 148490 149361 148546
rect 143904 148488 149361 148490
rect 149295 148485 149361 148488
rect 674746 148486 674752 148550
rect 674816 148548 674822 148550
rect 675471 148548 675537 148551
rect 674816 148546 675537 148548
rect 674816 148490 675476 148546
rect 675532 148490 675537 148546
rect 674816 148488 675537 148490
rect 674816 148486 674822 148488
rect 675471 148485 675537 148488
rect 184719 148104 184785 148107
rect 645135 148104 645201 148107
rect 184719 148102 190560 148104
rect 184719 148046 184724 148102
rect 184780 148046 190560 148102
rect 640416 148102 645201 148104
rect 640416 148074 645140 148102
rect 184719 148044 190560 148046
rect 640386 148046 645140 148074
rect 645196 148046 645201 148102
rect 640386 148044 645201 148046
rect 184719 148041 184785 148044
rect 149391 147364 149457 147367
rect 143904 147362 149457 147364
rect 143904 147306 149396 147362
rect 149452 147306 149457 147362
rect 143904 147304 149457 147306
rect 149391 147301 149457 147304
rect 184527 147364 184593 147367
rect 184527 147362 190560 147364
rect 184527 147306 184532 147362
rect 184588 147306 190560 147362
rect 184527 147304 190560 147306
rect 184527 147301 184593 147304
rect 184623 146624 184689 146627
rect 184623 146622 190560 146624
rect 184623 146566 184628 146622
rect 184684 146566 190560 146622
rect 184623 146564 190560 146566
rect 184623 146561 184689 146564
rect 147663 146180 147729 146183
rect 143904 146178 147729 146180
rect 143904 146122 147668 146178
rect 147724 146122 147729 146178
rect 640386 146150 640446 148044
rect 645135 148041 645201 148044
rect 675759 146624 675825 146627
rect 676090 146624 676096 146626
rect 675759 146622 676096 146624
rect 675759 146566 675764 146622
rect 675820 146566 676096 146622
rect 675759 146564 676096 146566
rect 675759 146561 675825 146564
rect 676090 146562 676096 146564
rect 676160 146562 676166 146626
rect 143904 146120 147729 146122
rect 147663 146117 147729 146120
rect 184335 145884 184401 145887
rect 184335 145882 190560 145884
rect 184335 145826 184340 145882
rect 184396 145826 190560 145882
rect 184335 145824 190560 145826
rect 184335 145821 184401 145824
rect 184431 145144 184497 145147
rect 184431 145142 190014 145144
rect 184431 145086 184436 145142
rect 184492 145086 190014 145142
rect 184431 145084 190014 145086
rect 184431 145081 184497 145084
rect 189954 145070 190014 145084
rect 189954 145010 190560 145070
rect 143874 144552 143934 144892
rect 147471 144552 147537 144555
rect 143874 144550 147537 144552
rect 143874 144494 147476 144550
rect 147532 144494 147537 144550
rect 143874 144492 147537 144494
rect 147471 144489 147537 144492
rect 184527 144404 184593 144407
rect 184527 144402 190560 144404
rect 184527 144346 184532 144402
rect 184588 144346 190560 144402
rect 184527 144344 190560 144346
rect 184527 144341 184593 144344
rect 646671 144256 646737 144259
rect 640416 144254 646737 144256
rect 640416 144226 646676 144254
rect 640386 144198 646676 144226
rect 646732 144198 646737 144254
rect 640386 144196 646737 144198
rect 147471 143664 147537 143667
rect 143904 143662 147537 143664
rect 143904 143606 147476 143662
rect 147532 143606 147537 143662
rect 143904 143604 147537 143606
rect 147471 143601 147537 143604
rect 184335 143664 184401 143667
rect 184335 143662 190014 143664
rect 184335 143606 184340 143662
rect 184396 143606 190014 143662
rect 184335 143604 190014 143606
rect 184335 143601 184401 143604
rect 189954 143590 190014 143604
rect 189954 143530 190560 143590
rect 184431 142776 184497 142779
rect 184431 142774 190560 142776
rect 184431 142718 184436 142774
rect 184492 142718 190560 142774
rect 184431 142716 190560 142718
rect 184431 142713 184497 142716
rect 147663 142480 147729 142483
rect 143904 142478 147729 142480
rect 143904 142422 147668 142478
rect 147724 142422 147729 142478
rect 143904 142420 147729 142422
rect 147663 142417 147729 142420
rect 640386 142302 640446 144196
rect 646671 144193 646737 144196
rect 184623 142184 184689 142187
rect 184623 142182 190014 142184
rect 184623 142126 184628 142182
rect 184684 142126 190014 142182
rect 184623 142124 190014 142126
rect 184623 142121 184689 142124
rect 189954 142110 190014 142124
rect 189954 142050 190560 142110
rect 149679 141296 149745 141299
rect 143904 141294 149745 141296
rect 143904 141238 149684 141294
rect 149740 141238 149745 141294
rect 143904 141236 149745 141238
rect 149679 141233 149745 141236
rect 184527 141296 184593 141299
rect 184527 141294 190560 141296
rect 184527 141238 184532 141294
rect 184588 141238 190560 141294
rect 184527 141236 190560 141238
rect 184527 141233 184593 141236
rect 646767 141000 646833 141003
rect 640386 140998 646833 141000
rect 640386 140942 646772 140998
rect 646828 140942 646833 140998
rect 640386 140940 646833 140942
rect 184335 140556 184401 140559
rect 184335 140554 190560 140556
rect 184335 140498 184340 140554
rect 184396 140498 190560 140554
rect 184335 140496 190560 140498
rect 184335 140493 184401 140496
rect 640386 140408 640446 140940
rect 646767 140937 646833 140940
rect 640224 140378 640446 140408
rect 640194 140348 640416 140378
rect 147471 139964 147537 139967
rect 143904 139962 147537 139964
rect 143904 139906 147476 139962
rect 147532 139906 147537 139962
rect 143904 139904 147537 139906
rect 147471 139901 147537 139904
rect 184431 139816 184497 139819
rect 184431 139814 190560 139816
rect 184431 139758 184436 139814
rect 184492 139758 190560 139814
rect 184431 139756 190560 139758
rect 184431 139753 184497 139756
rect 184527 138928 184593 138931
rect 184527 138926 190560 138928
rect 184527 138870 184532 138926
rect 184588 138870 190560 138926
rect 184527 138868 190560 138870
rect 184527 138865 184593 138868
rect 147471 138780 147537 138783
rect 143904 138778 147537 138780
rect 143904 138722 147476 138778
rect 147532 138722 147537 138778
rect 143904 138720 147537 138722
rect 147471 138717 147537 138720
rect 640194 138528 640254 140348
rect 185967 138336 186033 138339
rect 185967 138334 190560 138336
rect 185967 138278 185972 138334
rect 186028 138278 190560 138334
rect 185967 138276 190560 138278
rect 185967 138273 186033 138276
rect 149583 137596 149649 137599
rect 143904 137594 149649 137596
rect 143904 137538 149588 137594
rect 149644 137538 149649 137594
rect 143904 137536 149649 137538
rect 149583 137533 149649 137536
rect 186063 137448 186129 137451
rect 186063 137446 190560 137448
rect 186063 137390 186068 137446
rect 186124 137390 190560 137446
rect 186063 137388 190560 137390
rect 186063 137385 186129 137388
rect 186255 136856 186321 136859
rect 186255 136854 190014 136856
rect 186255 136798 186260 136854
rect 186316 136798 190014 136854
rect 186255 136796 190014 136798
rect 186255 136793 186321 136796
rect 189954 136782 190014 136796
rect 189954 136722 190560 136782
rect 143874 135968 143934 136308
rect 149679 135968 149745 135971
rect 143874 135966 149745 135968
rect 143874 135910 149684 135966
rect 149740 135910 149745 135966
rect 143874 135908 149745 135910
rect 149679 135905 149745 135908
rect 186447 135968 186513 135971
rect 186447 135966 190560 135968
rect 186447 135910 186452 135966
rect 186508 135910 190560 135966
rect 186447 135908 190560 135910
rect 186447 135905 186513 135908
rect 185775 135228 185841 135231
rect 185775 135226 190014 135228
rect 185775 135170 185780 135226
rect 185836 135170 190014 135226
rect 185775 135168 190014 135170
rect 185775 135165 185841 135168
rect 189954 135154 190014 135168
rect 189954 135094 190560 135154
rect 149679 135080 149745 135083
rect 143904 135078 149745 135080
rect 143904 135022 149684 135078
rect 149740 135022 149745 135078
rect 143904 135020 149745 135022
rect 149679 135017 149745 135020
rect 647055 134784 647121 134787
rect 640416 134782 647121 134784
rect 640416 134726 647060 134782
rect 647116 134726 647121 134782
rect 640416 134724 647121 134726
rect 647055 134721 647121 134724
rect 184335 134488 184401 134491
rect 184335 134486 190560 134488
rect 184335 134430 184340 134486
rect 184396 134430 190560 134486
rect 184335 134428 190560 134430
rect 184335 134425 184401 134428
rect 148815 133896 148881 133899
rect 143904 133894 148881 133896
rect 143904 133838 148820 133894
rect 148876 133838 148881 133894
rect 143904 133836 148881 133838
rect 148815 133833 148881 133836
rect 186159 133748 186225 133751
rect 186159 133746 190014 133748
rect 186159 133690 186164 133746
rect 186220 133690 190014 133746
rect 186159 133688 190014 133690
rect 186159 133685 186225 133688
rect 189954 133674 190014 133688
rect 189954 133614 190560 133674
rect 184431 133008 184497 133011
rect 184431 133006 190560 133008
rect 184431 132950 184436 133006
rect 184492 132950 190560 133006
rect 184431 132948 190560 132950
rect 184431 132945 184497 132948
rect 149007 132712 149073 132715
rect 143904 132710 149073 132712
rect 143904 132654 149012 132710
rect 149068 132654 149073 132710
rect 143904 132652 149073 132654
rect 149007 132649 149073 132652
rect 184335 132268 184401 132271
rect 184335 132266 190014 132268
rect 184335 132210 184340 132266
rect 184396 132210 190014 132266
rect 184335 132208 190014 132210
rect 184335 132205 184401 132208
rect 189954 132194 190014 132208
rect 189954 132134 190560 132194
rect 676143 131824 676209 131827
rect 676290 131824 676350 132090
rect 676143 131822 676350 131824
rect 676143 131766 676148 131822
rect 676204 131766 676350 131822
rect 676143 131764 676350 131766
rect 676143 131761 676209 131764
rect 184431 131528 184497 131531
rect 184431 131526 190560 131528
rect 184431 131470 184436 131526
rect 184492 131470 190560 131526
rect 184431 131468 190560 131470
rect 184431 131465 184497 131468
rect 143874 130936 143934 131424
rect 676290 131235 676350 131498
rect 676290 131230 676401 131235
rect 676290 131174 676340 131230
rect 676396 131174 676401 131230
rect 676290 131172 676401 131174
rect 676335 131169 676401 131172
rect 149679 130936 149745 130939
rect 647823 130936 647889 130939
rect 143874 130934 149745 130936
rect 143874 130878 149684 130934
rect 149740 130878 149745 130934
rect 143874 130876 149745 130878
rect 640416 130934 647889 130936
rect 640416 130878 647828 130934
rect 647884 130878 647889 130934
rect 640416 130876 647889 130878
rect 149679 130873 149745 130876
rect 647823 130873 647889 130876
rect 676290 130791 676350 130980
rect 676239 130786 676350 130791
rect 676239 130730 676244 130786
rect 676300 130730 676350 130786
rect 676239 130728 676350 130730
rect 676239 130725 676305 130728
rect 184527 130640 184593 130643
rect 184527 130638 190560 130640
rect 184527 130582 184532 130638
rect 184588 130582 190560 130638
rect 184527 130580 190560 130582
rect 184527 130577 184593 130580
rect 674362 130578 674368 130642
rect 674432 130640 674438 130642
rect 674432 130580 676320 130640
rect 674432 130578 674438 130580
rect 147471 130344 147537 130347
rect 143904 130342 147537 130344
rect 143904 130286 147476 130342
rect 147532 130286 147537 130342
rect 143904 130284 147537 130286
rect 147471 130281 147537 130284
rect 184623 129900 184689 129903
rect 184623 129898 190560 129900
rect 184623 129842 184628 129898
rect 184684 129842 190560 129898
rect 184623 129840 190560 129842
rect 184623 129837 184689 129840
rect 676290 129755 676350 130018
rect 676239 129750 676350 129755
rect 676239 129694 676244 129750
rect 676300 129694 676350 129750
rect 676239 129692 676350 129694
rect 676239 129689 676305 129692
rect 673978 129394 673984 129458
rect 674048 129456 674054 129458
rect 674048 129396 676320 129456
rect 674048 129394 674054 129396
rect 149103 129160 149169 129163
rect 143904 129158 149169 129160
rect 143904 129102 149108 129158
rect 149164 129102 149169 129158
rect 143904 129100 149169 129102
rect 149103 129097 149169 129100
rect 186735 129160 186801 129163
rect 186735 129158 190560 129160
rect 186735 129102 186740 129158
rect 186796 129102 190560 129158
rect 186735 129100 190560 129102
rect 186735 129097 186801 129100
rect 645711 129012 645777 129015
rect 640416 129010 645777 129012
rect 640416 128954 645716 129010
rect 645772 128954 645777 129010
rect 640416 128952 645777 128954
rect 645711 128949 645777 128952
rect 676143 128864 676209 128867
rect 676290 128864 676350 129130
rect 676143 128862 676350 128864
rect 676143 128806 676148 128862
rect 676204 128806 676350 128862
rect 676143 128804 676350 128806
rect 676143 128801 676209 128804
rect 674170 128506 674176 128570
rect 674240 128568 674246 128570
rect 674240 128508 676320 128568
rect 674240 128506 674246 128508
rect 184335 128420 184401 128423
rect 184335 128418 190014 128420
rect 184335 128362 184340 128418
rect 184396 128362 190014 128418
rect 184335 128360 190014 128362
rect 184335 128357 184401 128360
rect 189954 128346 190014 128360
rect 189954 128286 190560 128346
rect 147471 127976 147537 127979
rect 143904 127974 147537 127976
rect 143904 127918 147476 127974
rect 147532 127918 147537 127974
rect 143904 127916 147537 127918
rect 147471 127913 147537 127916
rect 676290 127831 676350 127946
rect 676239 127826 676350 127831
rect 676239 127770 676244 127826
rect 676300 127770 676350 127826
rect 676239 127768 676350 127770
rect 676239 127765 676305 127768
rect 184431 127680 184497 127683
rect 646959 127680 647025 127683
rect 184431 127678 190560 127680
rect 184431 127622 184436 127678
rect 184492 127622 190560 127678
rect 184431 127620 190560 127622
rect 640386 127678 647025 127680
rect 640386 127622 646964 127678
rect 647020 127622 647025 127678
rect 640386 127620 647025 127622
rect 184431 127617 184497 127620
rect 640386 127058 640446 127620
rect 646959 127617 647025 127620
rect 676047 127606 676113 127609
rect 676047 127604 676320 127606
rect 676047 127548 676052 127604
rect 676108 127548 676320 127604
rect 676047 127546 676320 127548
rect 676047 127543 676113 127546
rect 184527 126940 184593 126943
rect 184527 126938 190014 126940
rect 184527 126882 184532 126938
rect 184588 126882 190014 126938
rect 184527 126880 190014 126882
rect 184527 126877 184593 126880
rect 189954 126866 190014 126880
rect 189954 126806 190560 126866
rect 676866 126795 676926 127058
rect 676866 126790 676977 126795
rect 676866 126734 676916 126790
rect 676972 126734 676977 126790
rect 676866 126732 676977 126734
rect 676911 126729 676977 126732
rect 149295 126644 149361 126647
rect 143904 126642 149361 126644
rect 143904 126586 149300 126642
rect 149356 126586 149361 126642
rect 143904 126584 149361 126586
rect 149295 126581 149361 126584
rect 675567 126496 675633 126499
rect 675567 126494 676320 126496
rect 675567 126438 675572 126494
rect 675628 126438 676320 126494
rect 675567 126436 676320 126438
rect 675567 126433 675633 126436
rect 676047 126126 676113 126129
rect 676047 126124 676320 126126
rect 676047 126068 676052 126124
rect 676108 126068 676320 126124
rect 676047 126066 676320 126068
rect 676047 126063 676113 126066
rect 184335 126052 184401 126055
rect 184335 126050 190560 126052
rect 184335 125994 184340 126050
rect 184396 125994 190560 126050
rect 184335 125992 190560 125994
rect 184335 125989 184401 125992
rect 646863 125756 646929 125759
rect 640386 125754 646929 125756
rect 640386 125698 646868 125754
rect 646924 125698 646929 125754
rect 640386 125696 646929 125698
rect 149583 125460 149649 125463
rect 143904 125458 149649 125460
rect 143904 125402 149588 125458
rect 149644 125402 149649 125458
rect 143904 125400 149649 125402
rect 149583 125397 149649 125400
rect 184431 125460 184497 125463
rect 184431 125458 190014 125460
rect 184431 125402 184436 125458
rect 184492 125402 190014 125458
rect 184431 125400 190014 125402
rect 184431 125397 184497 125400
rect 189954 125386 190014 125400
rect 189954 125326 190560 125386
rect 640386 125208 640446 125696
rect 646863 125693 646929 125696
rect 675706 125546 675712 125610
rect 675776 125608 675782 125610
rect 675776 125548 676320 125608
rect 675776 125546 675782 125548
rect 676866 124871 676926 124986
rect 676815 124866 676926 124871
rect 676815 124810 676820 124866
rect 676876 124810 676926 124866
rect 676815 124808 676926 124810
rect 676815 124805 676881 124808
rect 184527 124572 184593 124575
rect 184527 124570 190560 124572
rect 184527 124514 184532 124570
rect 184588 124514 190560 124570
rect 184527 124512 190560 124514
rect 184527 124509 184593 124512
rect 676290 124427 676350 124542
rect 676239 124422 676350 124427
rect 676239 124366 676244 124422
rect 676300 124366 676350 124422
rect 676239 124364 676350 124366
rect 676239 124361 676305 124364
rect 149391 124276 149457 124279
rect 143904 124274 149457 124276
rect 143904 124218 149396 124274
rect 149452 124218 149457 124274
rect 143904 124216 149457 124218
rect 149391 124213 149457 124216
rect 676047 124128 676113 124131
rect 676047 124126 676320 124128
rect 676047 124070 676052 124126
rect 676108 124070 676320 124126
rect 676047 124068 676320 124070
rect 676047 124065 676113 124068
rect 184431 123832 184497 123835
rect 646575 123832 646641 123835
rect 184431 123830 190560 123832
rect 184431 123774 184436 123830
rect 184492 123774 190560 123830
rect 184431 123772 190560 123774
rect 640194 123830 646641 123832
rect 640194 123774 646580 123830
rect 646636 123774 646641 123830
rect 640194 123772 646641 123774
rect 184431 123769 184497 123772
rect 640194 123358 640254 123772
rect 646575 123769 646641 123772
rect 676047 123536 676113 123539
rect 676047 123534 676320 123536
rect 676047 123478 676052 123534
rect 676108 123478 676320 123534
rect 676047 123476 676320 123478
rect 676047 123473 676113 123476
rect 184335 123092 184401 123095
rect 184335 123090 190560 123092
rect 184335 123034 184340 123090
rect 184396 123034 190560 123090
rect 184335 123032 190560 123034
rect 184335 123029 184401 123032
rect 673978 123030 673984 123094
rect 674048 123092 674054 123094
rect 674048 123032 676320 123092
rect 674048 123030 674054 123032
rect 143874 122500 143934 122988
rect 148335 122500 148401 122503
rect 143874 122498 148401 122500
rect 143874 122442 148340 122498
rect 148396 122442 148401 122498
rect 143874 122440 148401 122442
rect 148335 122437 148401 122440
rect 184623 122204 184689 122207
rect 184623 122202 190560 122204
rect 184623 122146 184628 122202
rect 184684 122146 190560 122202
rect 184623 122144 190560 122146
rect 184623 122141 184689 122144
rect 675514 122142 675520 122206
rect 675584 122204 675590 122206
rect 676290 122204 676350 122544
rect 675584 122144 676350 122204
rect 675584 122142 675590 122144
rect 646479 122056 646545 122059
rect 640194 122054 646545 122056
rect 640194 121998 646484 122054
rect 646540 121998 646545 122054
rect 640194 121996 646545 121998
rect 148527 121760 148593 121763
rect 143904 121758 148593 121760
rect 143904 121702 148532 121758
rect 148588 121702 148593 121758
rect 143904 121700 148593 121702
rect 148527 121697 148593 121700
rect 184527 121612 184593 121615
rect 184527 121610 190560 121612
rect 184527 121554 184532 121610
rect 184588 121554 190560 121610
rect 184527 121552 190560 121554
rect 184527 121549 184593 121552
rect 640194 121434 640254 121996
rect 646479 121993 646545 121996
rect 676047 122056 676113 122059
rect 676047 122054 676320 122056
rect 676047 121998 676052 122054
rect 676108 121998 676320 122054
rect 676047 121996 676320 121998
rect 676047 121993 676113 121996
rect 676290 121467 676350 121582
rect 676239 121462 676350 121467
rect 676239 121406 676244 121462
rect 676300 121406 676350 121462
rect 676239 121404 676350 121406
rect 676239 121401 676305 121404
rect 675951 121094 676017 121097
rect 675951 121092 676320 121094
rect 675951 121036 675956 121092
rect 676012 121036 676320 121092
rect 675951 121034 676320 121036
rect 675951 121031 676017 121034
rect 184335 120724 184401 120727
rect 184335 120722 190560 120724
rect 184335 120666 184340 120722
rect 184396 120666 190560 120722
rect 184335 120664 190560 120666
rect 184335 120661 184401 120664
rect 147855 120576 147921 120579
rect 143904 120574 147921 120576
rect 143904 120518 147860 120574
rect 147916 120518 147921 120574
rect 143904 120516 147921 120518
rect 147855 120513 147921 120516
rect 676047 120576 676113 120579
rect 676047 120574 676320 120576
rect 676047 120518 676052 120574
rect 676108 120518 676320 120574
rect 676047 120516 676320 120518
rect 676047 120513 676113 120516
rect 184527 120132 184593 120135
rect 184527 120130 190014 120132
rect 184527 120074 184532 120130
rect 184588 120074 190014 120130
rect 184527 120072 190014 120074
rect 184527 120069 184593 120072
rect 189954 120058 190014 120072
rect 189954 119998 190560 120058
rect 676143 119836 676209 119839
rect 676290 119836 676350 120102
rect 676143 119834 676350 119836
rect 676143 119778 676148 119834
rect 676204 119778 676350 119834
rect 676143 119776 676350 119778
rect 676143 119773 676209 119776
rect 647919 119540 647985 119543
rect 640416 119538 647985 119540
rect 640416 119482 647924 119538
rect 647980 119482 647985 119538
rect 640416 119480 647985 119482
rect 647919 119477 647985 119480
rect 676290 119395 676350 119510
rect 149487 119392 149553 119395
rect 143904 119390 149553 119392
rect 143904 119334 149492 119390
rect 149548 119334 149553 119390
rect 143904 119332 149553 119334
rect 149487 119329 149553 119332
rect 676239 119390 676350 119395
rect 676239 119334 676244 119390
rect 676300 119334 676350 119390
rect 676239 119332 676350 119334
rect 676239 119329 676305 119332
rect 184431 119244 184497 119247
rect 184431 119242 190560 119244
rect 184431 119186 184436 119242
rect 184492 119186 190560 119242
rect 184431 119184 190560 119186
rect 184431 119181 184497 119184
rect 184719 118652 184785 118655
rect 184719 118650 190014 118652
rect 184719 118594 184724 118650
rect 184780 118594 190014 118650
rect 184719 118592 190014 118594
rect 184719 118589 184785 118592
rect 189954 118578 190014 118592
rect 189954 118518 190560 118578
rect 149391 118208 149457 118211
rect 143874 118206 149457 118208
rect 143874 118150 149396 118206
rect 149452 118150 149457 118206
rect 143874 118148 149457 118150
rect 143874 118104 143934 118148
rect 149391 118145 149457 118148
rect 184335 117764 184401 117767
rect 184335 117762 190560 117764
rect 184335 117706 184340 117762
rect 184396 117706 190560 117762
rect 184335 117704 190560 117706
rect 184335 117701 184401 117704
rect 645231 117616 645297 117619
rect 640416 117614 645297 117616
rect 640416 117558 645236 117614
rect 645292 117558 645297 117614
rect 640416 117556 645297 117558
rect 645231 117553 645297 117556
rect 184431 117024 184497 117027
rect 184431 117022 190014 117024
rect 184431 116966 184436 117022
rect 184492 116966 190014 117022
rect 184431 116964 190014 116966
rect 184431 116961 184497 116964
rect 189954 116950 190014 116964
rect 189954 116890 190560 116950
rect 149487 116876 149553 116879
rect 143904 116874 149553 116876
rect 143904 116818 149492 116874
rect 149548 116818 149553 116874
rect 143904 116816 149553 116818
rect 149487 116813 149553 116816
rect 675898 116666 675904 116730
rect 675968 116728 675974 116730
rect 676911 116728 676977 116731
rect 675968 116726 676977 116728
rect 675968 116670 676916 116726
rect 676972 116670 676977 116726
rect 675968 116668 676977 116670
rect 675968 116666 675974 116668
rect 676911 116665 676977 116668
rect 184527 116284 184593 116287
rect 184527 116282 190560 116284
rect 184527 116226 184532 116282
rect 184588 116226 190560 116282
rect 184527 116224 190560 116226
rect 184527 116221 184593 116224
rect 676666 116074 676672 116138
rect 676736 116136 676742 116138
rect 676815 116136 676881 116139
rect 676736 116134 676881 116136
rect 676736 116078 676820 116134
rect 676876 116078 676881 116134
rect 676736 116076 676881 116078
rect 676736 116074 676742 116076
rect 676815 116073 676881 116076
rect 149391 115692 149457 115695
rect 647919 115692 647985 115695
rect 143904 115690 149457 115692
rect 143904 115634 149396 115690
rect 149452 115634 149457 115690
rect 143904 115632 149457 115634
rect 640416 115690 647985 115692
rect 640416 115634 647924 115690
rect 647980 115634 647985 115690
rect 640416 115632 647985 115634
rect 149391 115629 149457 115632
rect 647919 115629 647985 115632
rect 184623 115396 184689 115399
rect 184623 115394 190560 115396
rect 184623 115338 184628 115394
rect 184684 115338 190560 115394
rect 184623 115336 190560 115338
rect 184623 115333 184689 115336
rect 148815 115248 148881 115251
rect 149391 115248 149457 115251
rect 148815 115246 149457 115248
rect 148815 115190 148820 115246
rect 148876 115190 149396 115246
rect 149452 115190 149457 115246
rect 148815 115188 149457 115190
rect 148815 115185 148881 115188
rect 149391 115185 149457 115188
rect 184335 114804 184401 114807
rect 184335 114802 190560 114804
rect 184335 114746 184340 114802
rect 184396 114746 190560 114802
rect 184335 114744 190560 114746
rect 184335 114741 184401 114744
rect 149391 114508 149457 114511
rect 143904 114506 149457 114508
rect 143904 114450 149396 114506
rect 149452 114450 149457 114506
rect 143904 114448 149457 114450
rect 149391 114445 149457 114448
rect 184431 113916 184497 113919
rect 184431 113914 190560 113916
rect 184431 113858 184436 113914
rect 184492 113858 190560 113914
rect 184431 113856 190560 113858
rect 184431 113853 184497 113856
rect 149391 113176 149457 113179
rect 143904 113174 149457 113176
rect 143904 113118 149396 113174
rect 149452 113118 149457 113174
rect 143904 113116 149457 113118
rect 149391 113113 149457 113116
rect 184527 113176 184593 113179
rect 640194 113176 640254 113738
rect 646575 113176 646641 113179
rect 184527 113174 190560 113176
rect 184527 113118 184532 113174
rect 184588 113118 190560 113174
rect 184527 113116 190560 113118
rect 640194 113174 646641 113176
rect 640194 113118 646580 113174
rect 646636 113118 646641 113174
rect 640194 113116 646641 113118
rect 184527 113113 184593 113116
rect 646575 113113 646641 113116
rect 184623 112436 184689 112439
rect 184623 112434 190560 112436
rect 184623 112378 184628 112434
rect 184684 112378 190560 112434
rect 184623 112376 190560 112378
rect 184623 112373 184689 112376
rect 148239 111992 148305 111995
rect 143904 111990 148305 111992
rect 143904 111934 148244 111990
rect 148300 111934 148305 111990
rect 143904 111932 148305 111934
rect 148239 111929 148305 111932
rect 184335 111696 184401 111699
rect 184335 111694 190014 111696
rect 184335 111638 184340 111694
rect 184396 111638 190014 111694
rect 184335 111636 190014 111638
rect 184335 111633 184401 111636
rect 189954 111622 190014 111636
rect 189954 111562 190560 111622
rect 640386 111400 640446 111888
rect 647055 111400 647121 111403
rect 640386 111398 647121 111400
rect 640386 111342 647060 111398
rect 647116 111342 647121 111398
rect 640386 111340 647121 111342
rect 647055 111337 647121 111340
rect 149391 110956 149457 110959
rect 143904 110954 149457 110956
rect 143904 110898 149396 110954
rect 149452 110898 149457 110954
rect 143904 110896 149457 110898
rect 149391 110893 149457 110896
rect 184431 110956 184497 110959
rect 184431 110954 190560 110956
rect 184431 110898 184436 110954
rect 184492 110898 190560 110954
rect 184431 110896 190560 110898
rect 184431 110893 184497 110896
rect 184527 110216 184593 110219
rect 184527 110214 190014 110216
rect 184527 110158 184532 110214
rect 184588 110158 190014 110214
rect 184527 110156 190014 110158
rect 184527 110153 184593 110156
rect 189954 110142 190014 110156
rect 189954 110082 190560 110142
rect 143874 109624 143934 109668
rect 148623 109624 148689 109627
rect 143874 109622 148689 109624
rect 143874 109566 148628 109622
rect 148684 109566 148689 109622
rect 143874 109564 148689 109566
rect 148623 109561 148689 109564
rect 640386 109476 640446 109890
rect 646671 109476 646737 109479
rect 640386 109474 646737 109476
rect 640386 109418 646676 109474
rect 646732 109418 646737 109474
rect 640386 109416 646737 109418
rect 646671 109413 646737 109416
rect 184335 109328 184401 109331
rect 184335 109326 190560 109328
rect 184335 109270 184340 109326
rect 184396 109270 190560 109326
rect 184335 109268 190560 109270
rect 184335 109265 184401 109268
rect 185583 108736 185649 108739
rect 185583 108734 190014 108736
rect 185583 108678 185588 108734
rect 185644 108678 190014 108734
rect 185583 108676 190014 108678
rect 185583 108673 185649 108676
rect 189954 108662 190014 108676
rect 189954 108602 190560 108662
rect 147183 108440 147249 108443
rect 143904 108438 147249 108440
rect 143904 108382 147188 108438
rect 147244 108382 147249 108438
rect 143904 108380 147249 108382
rect 147183 108377 147249 108380
rect 675759 108146 675825 108147
rect 675706 108082 675712 108146
rect 675776 108144 675825 108146
rect 675776 108142 675868 108144
rect 675820 108086 675868 108142
rect 675776 108084 675868 108086
rect 675776 108082 675825 108084
rect 675759 108081 675825 108082
rect 646767 107996 646833 107999
rect 640416 107994 646833 107996
rect 640416 107938 646772 107994
rect 646828 107938 646833 107994
rect 640416 107936 646833 107938
rect 646767 107933 646833 107936
rect 186159 107848 186225 107851
rect 186159 107846 190560 107848
rect 186159 107790 186164 107846
rect 186220 107790 190560 107846
rect 186159 107788 190560 107790
rect 186159 107785 186225 107788
rect 148431 107256 148497 107259
rect 143904 107254 148497 107256
rect 143904 107198 148436 107254
rect 148492 107198 148497 107254
rect 143904 107196 148497 107198
rect 148431 107193 148497 107196
rect 184431 107108 184497 107111
rect 184431 107106 190560 107108
rect 184431 107050 184436 107106
rect 184492 107050 190560 107106
rect 184431 107048 190560 107050
rect 184431 107045 184497 107048
rect 675471 106666 675537 106667
rect 675471 106664 675520 106666
rect 675428 106662 675520 106664
rect 675428 106606 675476 106662
rect 675428 106604 675520 106606
rect 675471 106602 675520 106604
rect 675584 106602 675590 106666
rect 675471 106601 675537 106602
rect 185295 106368 185361 106371
rect 185295 106366 190560 106368
rect 185295 106310 185300 106366
rect 185356 106310 190560 106366
rect 185295 106308 190560 106310
rect 185295 106305 185361 106308
rect 148815 106072 148881 106075
rect 645903 106072 645969 106075
rect 143904 106070 148881 106072
rect 143904 106014 148820 106070
rect 148876 106014 148881 106070
rect 143904 106012 148881 106014
rect 640416 106070 645969 106072
rect 640416 106014 645908 106070
rect 645964 106014 645969 106070
rect 665472 106072 665982 106112
rect 668271 106072 668337 106075
rect 665472 106070 668337 106072
rect 665472 106052 668276 106070
rect 640416 106012 645969 106014
rect 665922 106014 668276 106052
rect 668332 106014 668337 106070
rect 665922 106012 668337 106014
rect 148815 106009 148881 106012
rect 645903 106009 645969 106012
rect 668271 106009 668337 106012
rect 184335 105628 184401 105631
rect 665199 105628 665265 105631
rect 184335 105626 190560 105628
rect 184335 105570 184340 105626
rect 184396 105570 190560 105626
rect 184335 105568 190560 105570
rect 665154 105626 665265 105628
rect 665154 105570 665204 105626
rect 665260 105570 665265 105626
rect 184335 105565 184401 105568
rect 665154 105565 665265 105570
rect 665154 105361 665214 105565
rect 665295 105184 665361 105187
rect 665295 105182 665406 105184
rect 665295 105126 665300 105182
rect 665356 105126 665406 105182
rect 665295 105121 665406 105126
rect 673978 105122 673984 105186
rect 674048 105184 674054 105186
rect 675375 105184 675441 105187
rect 674048 105182 675441 105184
rect 674048 105126 675380 105182
rect 675436 105126 675441 105182
rect 674048 105124 675441 105126
rect 674048 105122 674054 105124
rect 675375 105121 675441 105124
rect 665346 104996 665406 105121
rect 184527 104888 184593 104891
rect 184527 104886 190014 104888
rect 184527 104830 184532 104886
rect 184588 104830 190014 104886
rect 184527 104828 190014 104830
rect 184527 104825 184593 104828
rect 189954 104814 190014 104828
rect 189954 104754 190560 104814
rect 148623 104740 148689 104743
rect 143904 104738 148689 104740
rect 143904 104682 148628 104738
rect 148684 104682 148689 104738
rect 143904 104680 148689 104682
rect 148623 104677 148689 104680
rect 647919 104148 647985 104151
rect 640416 104146 647985 104148
rect 640416 104090 647924 104146
rect 647980 104090 647985 104146
rect 640416 104088 647985 104090
rect 647919 104085 647985 104088
rect 184431 104000 184497 104003
rect 184431 103998 190560 104000
rect 184431 103942 184436 103998
rect 184492 103942 190560 103998
rect 184431 103940 190560 103942
rect 184431 103937 184497 103940
rect 148719 103556 148785 103559
rect 143904 103554 148785 103556
rect 143904 103498 148724 103554
rect 148780 103498 148785 103554
rect 143904 103496 148785 103498
rect 148719 103493 148785 103496
rect 184431 103408 184497 103411
rect 184431 103406 190014 103408
rect 184431 103350 184436 103406
rect 184492 103350 190014 103406
rect 184431 103348 190014 103350
rect 184431 103345 184497 103348
rect 189954 103334 190014 103348
rect 189954 103274 190560 103334
rect 675759 103260 675825 103263
rect 675898 103260 675904 103262
rect 675759 103258 675904 103260
rect 675759 103202 675764 103258
rect 675820 103202 675904 103258
rect 675759 103200 675904 103202
rect 675759 103197 675825 103200
rect 675898 103198 675904 103200
rect 675968 103198 675974 103262
rect 184335 102520 184401 102523
rect 184335 102518 190560 102520
rect 184335 102462 184340 102518
rect 184396 102462 190560 102518
rect 184335 102460 190560 102462
rect 184335 102457 184401 102460
rect 148911 102372 148977 102375
rect 143904 102370 148977 102372
rect 143904 102314 148916 102370
rect 148972 102314 148977 102370
rect 143904 102312 148977 102314
rect 148911 102309 148977 102312
rect 645135 102224 645201 102227
rect 640416 102222 645201 102224
rect 640416 102166 645140 102222
rect 645196 102166 645201 102222
rect 640416 102164 645201 102166
rect 645135 102161 645201 102164
rect 184527 101928 184593 101931
rect 184527 101926 190014 101928
rect 184527 101870 184532 101926
rect 184588 101870 190014 101926
rect 184527 101868 190014 101870
rect 184527 101865 184593 101868
rect 189954 101854 190014 101868
rect 189954 101794 190560 101854
rect 675759 101484 675825 101487
rect 676666 101484 676672 101486
rect 675759 101482 676672 101484
rect 675759 101426 675764 101482
rect 675820 101426 676672 101482
rect 675759 101424 676672 101426
rect 675759 101421 675825 101424
rect 676666 101422 676672 101424
rect 676736 101422 676742 101486
rect 143874 100892 143934 101084
rect 184623 101040 184689 101043
rect 184623 101038 190560 101040
rect 184623 100982 184628 101038
rect 184684 100982 190560 101038
rect 184623 100980 190560 100982
rect 184623 100977 184689 100980
rect 149391 100892 149457 100895
rect 143874 100890 149457 100892
rect 143874 100834 149396 100890
rect 149452 100834 149457 100890
rect 143874 100832 149457 100834
rect 149391 100829 149457 100832
rect 184335 100300 184401 100303
rect 184335 100298 190014 100300
rect 184335 100242 184340 100298
rect 184396 100242 190014 100298
rect 184335 100240 190014 100242
rect 184335 100237 184401 100240
rect 189954 100226 190014 100240
rect 189954 100166 190560 100226
rect 149487 99856 149553 99859
rect 143904 99854 149553 99856
rect 143904 99798 149492 99854
rect 149548 99798 149553 99854
rect 143904 99796 149553 99798
rect 149487 99793 149553 99796
rect 640194 99708 640254 100270
rect 647919 99708 647985 99711
rect 640194 99706 647985 99708
rect 640194 99650 647924 99706
rect 647980 99650 647985 99706
rect 640194 99648 647985 99650
rect 647919 99645 647985 99648
rect 184431 99560 184497 99563
rect 184431 99558 190560 99560
rect 184431 99502 184436 99558
rect 184492 99502 190560 99558
rect 184431 99500 190560 99502
rect 184431 99497 184497 99500
rect 149391 98672 149457 98675
rect 143904 98670 149457 98672
rect 143904 98614 149396 98670
rect 149452 98614 149457 98670
rect 143904 98612 149457 98614
rect 149391 98609 149457 98612
rect 184623 98672 184689 98675
rect 184623 98670 190560 98672
rect 184623 98614 184628 98670
rect 184684 98614 190560 98670
rect 184623 98612 190560 98614
rect 184623 98609 184689 98612
rect 184527 98080 184593 98083
rect 640386 98080 640446 98420
rect 647151 98080 647217 98083
rect 184527 98078 190560 98080
rect 184527 98022 184532 98078
rect 184588 98022 190560 98078
rect 184527 98020 190560 98022
rect 640386 98078 647217 98080
rect 640386 98022 647156 98078
rect 647212 98022 647217 98078
rect 640386 98020 647217 98022
rect 184527 98017 184593 98020
rect 647151 98017 647217 98020
rect 149487 97488 149553 97491
rect 143904 97486 149553 97488
rect 143904 97430 149492 97486
rect 149548 97430 149553 97486
rect 143904 97428 149553 97430
rect 149487 97425 149553 97428
rect 184335 97192 184401 97195
rect 184335 97190 190560 97192
rect 184335 97134 184340 97190
rect 184396 97134 190560 97190
rect 184335 97132 190560 97134
rect 184335 97129 184401 97132
rect 184431 96452 184497 96455
rect 184431 96450 190560 96452
rect 184431 96394 184436 96450
rect 184492 96394 190560 96450
rect 184431 96392 190560 96394
rect 184431 96389 184497 96392
rect 143874 95712 143934 96200
rect 640386 96008 640446 96570
rect 645423 96008 645489 96011
rect 640386 96006 645489 96008
rect 640386 95950 645428 96006
rect 645484 95950 645489 96006
rect 640386 95948 645489 95950
rect 645423 95945 645489 95948
rect 149391 95712 149457 95715
rect 143874 95710 149457 95712
rect 143874 95654 149396 95710
rect 149452 95654 149457 95710
rect 143874 95652 149457 95654
rect 149391 95649 149457 95652
rect 184719 95712 184785 95715
rect 184719 95710 190560 95712
rect 184719 95654 184724 95710
rect 184780 95654 190560 95710
rect 184719 95652 190560 95654
rect 184719 95649 184785 95652
rect 149583 94972 149649 94975
rect 143904 94970 149649 94972
rect 143904 94914 149588 94970
rect 149644 94914 149649 94970
rect 143904 94912 149649 94914
rect 149583 94909 149649 94912
rect 189954 94838 190560 94898
rect 184335 94824 184401 94827
rect 189954 94824 190014 94838
rect 184335 94822 190014 94824
rect 184335 94766 184340 94822
rect 184396 94766 190014 94822
rect 184335 94764 190014 94766
rect 184335 94761 184401 94764
rect 184431 94232 184497 94235
rect 184431 94230 190560 94232
rect 184431 94174 184436 94230
rect 184492 94174 190560 94230
rect 184431 94172 190560 94174
rect 184431 94169 184497 94172
rect 640386 94084 640446 94646
rect 647727 94084 647793 94087
rect 640386 94082 647793 94084
rect 640386 94026 647732 94082
rect 647788 94026 647793 94082
rect 640386 94024 647793 94026
rect 647727 94021 647793 94024
rect 149487 93788 149553 93791
rect 143904 93786 149553 93788
rect 143904 93730 149492 93786
rect 149548 93730 149553 93786
rect 143904 93728 149553 93730
rect 149487 93725 149553 93728
rect 184527 93492 184593 93495
rect 184527 93490 190014 93492
rect 184527 93434 184532 93490
rect 184588 93434 190014 93490
rect 184527 93432 190014 93434
rect 184527 93429 184593 93432
rect 189954 93418 190014 93432
rect 189954 93358 190560 93418
rect 184623 92752 184689 92755
rect 647823 92752 647889 92755
rect 184623 92750 190560 92752
rect 184623 92694 184628 92750
rect 184684 92694 190560 92750
rect 184623 92692 190560 92694
rect 640416 92750 647889 92752
rect 640416 92694 647828 92750
rect 647884 92694 647889 92750
rect 640416 92692 647889 92694
rect 184623 92689 184689 92692
rect 647823 92689 647889 92692
rect 149391 92604 149457 92607
rect 143904 92602 149457 92604
rect 143904 92546 149396 92602
rect 149452 92546 149457 92602
rect 143904 92544 149457 92546
rect 149391 92541 149457 92544
rect 184335 92012 184401 92015
rect 184335 92010 190014 92012
rect 184335 91954 184340 92010
rect 184396 91954 190014 92010
rect 184335 91952 190014 91954
rect 184335 91949 184401 91952
rect 189954 91938 190014 91952
rect 189954 91878 190560 91938
rect 149295 91420 149361 91423
rect 143904 91418 149361 91420
rect 143904 91362 149300 91418
rect 149356 91362 149361 91418
rect 143904 91360 149361 91362
rect 149295 91357 149361 91360
rect 184623 91124 184689 91127
rect 184623 91122 190560 91124
rect 184623 91066 184628 91122
rect 184684 91066 190560 91122
rect 184623 91064 190560 91066
rect 184623 91061 184689 91064
rect 659343 90828 659409 90831
rect 640416 90826 659409 90828
rect 640416 90770 659348 90826
rect 659404 90770 659409 90826
rect 640416 90768 659409 90770
rect 659343 90765 659409 90768
rect 184431 90384 184497 90387
rect 184431 90382 190560 90384
rect 184431 90326 184436 90382
rect 184492 90326 190560 90382
rect 184431 90324 190560 90326
rect 184431 90321 184497 90324
rect 149391 90236 149457 90239
rect 143904 90234 149457 90236
rect 143904 90178 149396 90234
rect 149452 90178 149457 90234
rect 143904 90176 149457 90178
rect 149391 90173 149457 90176
rect 184527 89644 184593 89647
rect 184527 89642 190560 89644
rect 184527 89586 184532 89642
rect 184588 89586 190560 89642
rect 184527 89584 190560 89586
rect 184527 89581 184593 89584
rect 149391 89052 149457 89055
rect 143904 89050 149457 89052
rect 143904 88994 149396 89050
rect 149452 88994 149457 89050
rect 143904 88992 149457 88994
rect 149391 88989 149457 88992
rect 184335 88904 184401 88907
rect 645903 88904 645969 88907
rect 184335 88902 190560 88904
rect 184335 88846 184340 88902
rect 184396 88846 190560 88902
rect 184335 88844 190560 88846
rect 640416 88902 645969 88904
rect 640416 88846 645908 88902
rect 645964 88846 645969 88902
rect 640416 88844 645969 88846
rect 184335 88841 184401 88844
rect 645903 88841 645969 88844
rect 184431 88164 184497 88167
rect 184431 88162 190014 88164
rect 184431 88106 184436 88162
rect 184492 88106 190014 88162
rect 184431 88104 190014 88106
rect 184431 88101 184497 88104
rect 189954 88090 190014 88104
rect 189954 88030 190560 88090
rect 143874 87276 143934 87764
rect 149487 87276 149553 87279
rect 143874 87274 149553 87276
rect 143874 87218 149492 87274
rect 149548 87218 149553 87274
rect 143874 87216 149553 87218
rect 149487 87213 149553 87216
rect 184527 87276 184593 87279
rect 184527 87274 190560 87276
rect 184527 87218 184532 87274
rect 184588 87218 190560 87274
rect 184527 87216 190560 87218
rect 184527 87213 184593 87216
rect 647919 87128 647985 87131
rect 640386 87126 647985 87128
rect 640386 87070 647924 87126
rect 647980 87070 647985 87126
rect 640386 87068 647985 87070
rect 640386 86950 640446 87068
rect 647919 87065 647985 87068
rect 653679 86980 653745 86983
rect 653679 86978 656736 86980
rect 653679 86922 653684 86978
rect 653740 86922 656736 86978
rect 653679 86920 656736 86922
rect 653679 86917 653745 86920
rect 184623 86684 184689 86687
rect 184623 86682 190014 86684
rect 184623 86626 184628 86682
rect 184684 86626 190014 86682
rect 184623 86624 190014 86626
rect 184623 86621 184689 86624
rect 189954 86610 190014 86624
rect 189954 86550 190560 86610
rect 148815 86536 148881 86539
rect 143904 86534 148881 86536
rect 143904 86478 148820 86534
rect 148876 86478 148881 86534
rect 143904 86476 148881 86478
rect 148815 86473 148881 86476
rect 663279 86388 663345 86391
rect 663234 86386 663345 86388
rect 663234 86330 663284 86386
rect 663340 86330 663345 86386
rect 663234 86325 663345 86330
rect 650895 86240 650961 86243
rect 650895 86238 656736 86240
rect 650895 86182 650900 86238
rect 650956 86182 656736 86238
rect 663234 86210 663294 86325
rect 650895 86180 656736 86182
rect 650895 86177 650961 86180
rect 184335 85796 184401 85799
rect 184335 85794 190560 85796
rect 184335 85738 184340 85794
rect 184396 85738 190560 85794
rect 184335 85736 190560 85738
rect 184335 85733 184401 85736
rect 148815 85352 148881 85355
rect 143904 85350 148881 85352
rect 143904 85294 148820 85350
rect 148876 85294 148881 85350
rect 143904 85292 148881 85294
rect 148815 85289 148881 85292
rect 652335 85352 652401 85355
rect 652335 85350 656736 85352
rect 652335 85294 652340 85350
rect 652396 85294 656736 85350
rect 652335 85292 656736 85294
rect 652335 85289 652401 85292
rect 184431 85204 184497 85207
rect 184431 85202 190014 85204
rect 184431 85146 184436 85202
rect 184492 85146 190014 85202
rect 184431 85144 190014 85146
rect 184431 85141 184497 85144
rect 189954 85130 190014 85144
rect 189954 85070 190560 85130
rect 640194 84464 640254 85026
rect 663234 84763 663294 85322
rect 663234 84758 663345 84763
rect 663234 84702 663284 84758
rect 663340 84702 663345 84758
rect 663234 84700 663345 84702
rect 663279 84697 663345 84700
rect 645903 84464 645969 84467
rect 640194 84462 645969 84464
rect 640194 84406 645908 84462
rect 645964 84406 645969 84462
rect 640194 84404 645969 84406
rect 645903 84401 645969 84404
rect 184527 84316 184593 84319
rect 651759 84316 651825 84319
rect 184527 84314 190560 84316
rect 184527 84258 184532 84314
rect 184588 84258 190560 84314
rect 184527 84256 190560 84258
rect 651759 84314 656736 84316
rect 651759 84258 651764 84314
rect 651820 84258 656736 84314
rect 651759 84256 656736 84258
rect 184527 84253 184593 84256
rect 651759 84253 651825 84256
rect 147087 84168 147153 84171
rect 143904 84166 147153 84168
rect 143904 84110 147092 84166
rect 147148 84110 147153 84166
rect 143904 84108 147153 84110
rect 147087 84105 147153 84108
rect 663426 84023 663486 84582
rect 663426 84018 663537 84023
rect 663426 83962 663476 84018
rect 663532 83962 663537 84018
rect 663426 83960 663537 83962
rect 663471 83957 663537 83960
rect 189954 83442 190560 83502
rect 184335 83428 184401 83431
rect 189954 83428 190014 83442
rect 184335 83426 190014 83428
rect 184335 83370 184340 83426
rect 184396 83370 190014 83426
rect 184335 83368 190014 83370
rect 652239 83428 652305 83431
rect 652239 83426 656736 83428
rect 652239 83370 652244 83426
rect 652300 83370 656736 83426
rect 652239 83368 656736 83370
rect 184335 83365 184401 83368
rect 652239 83365 652305 83368
rect 143874 82392 143934 82880
rect 186159 82836 186225 82839
rect 186159 82834 190560 82836
rect 186159 82778 186164 82834
rect 186220 82778 190560 82834
rect 186159 82776 190560 82778
rect 186159 82773 186225 82776
rect 640386 82688 640446 83176
rect 663426 82839 663486 83398
rect 663375 82834 663486 82839
rect 663375 82778 663380 82834
rect 663436 82778 663486 82834
rect 663375 82776 663486 82778
rect 663375 82773 663441 82776
rect 647919 82688 647985 82691
rect 640386 82686 647985 82688
rect 640386 82630 647924 82686
rect 647980 82630 647985 82686
rect 640386 82628 647985 82630
rect 647919 82625 647985 82628
rect 652431 82688 652497 82691
rect 652431 82686 656736 82688
rect 652431 82630 652436 82686
rect 652492 82630 656736 82686
rect 652431 82628 656736 82630
rect 652431 82625 652497 82628
rect 149103 82392 149169 82395
rect 143874 82390 149169 82392
rect 143874 82334 149108 82390
rect 149164 82334 149169 82390
rect 143874 82332 149169 82334
rect 149103 82329 149169 82332
rect 663234 82099 663294 82658
rect 663234 82094 663345 82099
rect 663234 82038 663284 82094
rect 663340 82038 663345 82094
rect 663234 82036 663345 82038
rect 663279 82033 663345 82036
rect 184239 81948 184305 81951
rect 184239 81946 190560 81948
rect 184239 81890 184244 81946
rect 184300 81890 190560 81946
rect 184239 81888 190560 81890
rect 184239 81885 184305 81888
rect 148431 81652 148497 81655
rect 143904 81650 148497 81652
rect 143904 81594 148436 81650
rect 148492 81594 148497 81650
rect 143904 81592 148497 81594
rect 148431 81589 148497 81592
rect 662415 81652 662481 81655
rect 663042 81652 663102 81770
rect 662415 81650 663102 81652
rect 662415 81594 662420 81650
rect 662476 81594 663102 81650
rect 662415 81592 663102 81594
rect 662415 81589 662481 81592
rect 184431 81356 184497 81359
rect 184431 81354 190560 81356
rect 184431 81298 184436 81354
rect 184492 81298 190560 81354
rect 184431 81296 190560 81298
rect 184431 81293 184497 81296
rect 640386 81060 640446 81326
rect 647919 81060 647985 81063
rect 640386 81058 647985 81060
rect 640386 81002 647924 81058
rect 647980 81002 647985 81058
rect 640386 81000 647985 81002
rect 647919 80997 647985 81000
rect 149583 80468 149649 80471
rect 143904 80466 149649 80468
rect 143904 80410 149588 80466
rect 149644 80410 149649 80466
rect 143904 80408 149649 80410
rect 149583 80405 149649 80408
rect 184623 80468 184689 80471
rect 184623 80466 190560 80468
rect 184623 80410 184628 80466
rect 184684 80410 190560 80466
rect 184623 80408 190560 80410
rect 184623 80405 184689 80408
rect 184431 79876 184497 79879
rect 184431 79874 190014 79876
rect 184431 79818 184436 79874
rect 184492 79818 190014 79874
rect 184431 79816 190014 79818
rect 184431 79813 184497 79816
rect 189954 79802 190014 79816
rect 189954 79742 190560 79802
rect 645519 79432 645585 79435
rect 640416 79430 645585 79432
rect 640416 79374 645524 79430
rect 645580 79374 645585 79430
rect 640416 79372 645585 79374
rect 645519 79369 645585 79372
rect 149679 79284 149745 79287
rect 143904 79282 149745 79284
rect 143904 79226 149684 79282
rect 149740 79226 149745 79282
rect 143904 79224 149745 79226
rect 149679 79221 149745 79224
rect 184335 78988 184401 78991
rect 184335 78986 190560 78988
rect 184335 78930 184340 78986
rect 184396 78930 190560 78986
rect 184335 78928 190560 78930
rect 184335 78925 184401 78928
rect 184527 78248 184593 78251
rect 184527 78246 190014 78248
rect 184527 78190 184532 78246
rect 184588 78190 190014 78246
rect 184527 78188 190014 78190
rect 184527 78185 184593 78188
rect 189954 78174 190014 78188
rect 189954 78114 190560 78174
rect 148911 77952 148977 77955
rect 143904 77950 148977 77952
rect 143904 77894 148916 77950
rect 148972 77894 148977 77950
rect 143904 77892 148977 77894
rect 148911 77889 148977 77892
rect 184431 77508 184497 77511
rect 647919 77508 647985 77511
rect 184431 77506 190560 77508
rect 184431 77450 184436 77506
rect 184492 77450 190560 77506
rect 184431 77448 190560 77450
rect 640416 77506 647985 77508
rect 640416 77450 647924 77506
rect 647980 77450 647985 77506
rect 640416 77448 647985 77450
rect 184431 77445 184497 77448
rect 647919 77445 647985 77448
rect 149391 76768 149457 76771
rect 143904 76766 149457 76768
rect 143904 76710 149396 76766
rect 149452 76710 149457 76766
rect 143904 76708 149457 76710
rect 149391 76705 149457 76708
rect 184335 76768 184401 76771
rect 184335 76766 190014 76768
rect 184335 76710 184340 76766
rect 184396 76710 190014 76766
rect 184335 76708 190014 76710
rect 184335 76705 184401 76708
rect 189954 76694 190014 76708
rect 189954 76634 190560 76694
rect 184527 76028 184593 76031
rect 184527 76026 190560 76028
rect 184527 75970 184532 76026
rect 184588 75970 190560 76026
rect 184527 75968 190560 75970
rect 184527 75965 184593 75968
rect 149199 75584 149265 75587
rect 645999 75584 646065 75587
rect 143904 75582 149265 75584
rect 143904 75526 149204 75582
rect 149260 75526 149265 75582
rect 143904 75524 149265 75526
rect 640416 75582 646065 75584
rect 640416 75526 646004 75582
rect 646060 75526 646065 75582
rect 640416 75524 646065 75526
rect 149199 75521 149265 75524
rect 645999 75521 646065 75524
rect 184623 75140 184689 75143
rect 184623 75138 190560 75140
rect 184623 75082 184628 75138
rect 184684 75082 190560 75138
rect 184623 75080 190560 75082
rect 184623 75077 184689 75080
rect 184335 74400 184401 74403
rect 184335 74398 190560 74400
rect 184335 74342 184340 74398
rect 184396 74342 190560 74398
rect 184335 74340 190560 74342
rect 184335 74337 184401 74340
rect 143874 73808 143934 74296
rect 149295 73808 149361 73811
rect 143874 73806 149361 73808
rect 143874 73750 149300 73806
rect 149356 73750 149361 73806
rect 143874 73748 149361 73750
rect 149295 73745 149361 73748
rect 184527 73660 184593 73663
rect 647919 73660 647985 73663
rect 184527 73658 190560 73660
rect 184527 73602 184532 73658
rect 184588 73602 190560 73658
rect 184527 73600 190560 73602
rect 640416 73658 647985 73660
rect 640416 73602 647924 73658
rect 647980 73602 647985 73658
rect 640416 73600 647985 73602
rect 184527 73597 184593 73600
rect 647919 73597 647985 73600
rect 149007 73068 149073 73071
rect 143904 73066 149073 73068
rect 143904 73010 149012 73066
rect 149068 73010 149073 73066
rect 143904 73008 149073 73010
rect 149007 73005 149073 73008
rect 184431 72920 184497 72923
rect 184431 72918 190560 72920
rect 184431 72862 184436 72918
rect 184492 72862 190560 72918
rect 184431 72860 190560 72862
rect 184431 72857 184497 72860
rect 184623 72180 184689 72183
rect 184623 72178 190560 72180
rect 184623 72122 184628 72178
rect 184684 72122 190560 72178
rect 184623 72120 190560 72122
rect 184623 72117 184689 72120
rect 149103 72032 149169 72035
rect 143904 72030 149169 72032
rect 143904 71974 149108 72030
rect 149164 71974 149169 72030
rect 143904 71972 149169 71974
rect 149103 71969 149169 71972
rect 646959 71884 647025 71887
rect 640386 71882 647025 71884
rect 640386 71826 646964 71882
rect 647020 71826 647025 71882
rect 640386 71824 647025 71826
rect 640386 71706 640446 71824
rect 646959 71821 647025 71824
rect 184431 71440 184497 71443
rect 184431 71438 190014 71440
rect 184431 71382 184436 71438
rect 184492 71382 190014 71438
rect 184431 71380 190014 71382
rect 184431 71377 184497 71380
rect 189954 71366 190014 71380
rect 189954 71306 190560 71366
rect 149487 70848 149553 70851
rect 143904 70846 149553 70848
rect 143904 70790 149492 70846
rect 149548 70790 149553 70846
rect 143904 70788 149553 70790
rect 149487 70785 149553 70788
rect 184335 70552 184401 70555
rect 184335 70550 190560 70552
rect 184335 70494 184340 70550
rect 184396 70494 190560 70550
rect 184335 70492 190560 70494
rect 184335 70489 184401 70492
rect 184527 69960 184593 69963
rect 184527 69958 190014 69960
rect 184527 69902 184532 69958
rect 184588 69902 190014 69958
rect 184527 69900 190014 69902
rect 184527 69897 184593 69900
rect 189954 69886 190014 69900
rect 189954 69826 190560 69886
rect 640386 69664 640446 69856
rect 647919 69664 647985 69667
rect 640386 69662 647985 69664
rect 640386 69606 647924 69662
rect 647980 69606 647985 69662
rect 640386 69604 647985 69606
rect 647919 69601 647985 69604
rect 149391 69516 149457 69519
rect 143904 69514 149457 69516
rect 143904 69458 149396 69514
rect 149452 69458 149457 69514
rect 143904 69456 149457 69458
rect 149391 69453 149457 69456
rect 184335 69072 184401 69075
rect 184335 69070 190560 69072
rect 184335 69014 184340 69070
rect 184396 69014 190560 69070
rect 184335 69012 190560 69014
rect 184335 69009 184401 69012
rect 646863 68628 646929 68631
rect 640194 68626 646929 68628
rect 640194 68570 646868 68626
rect 646924 68570 646929 68626
rect 640194 68568 646929 68570
rect 184527 68480 184593 68483
rect 184527 68478 190014 68480
rect 184527 68422 184532 68478
rect 184588 68422 190014 68478
rect 184527 68420 190014 68422
rect 184527 68417 184593 68420
rect 189954 68406 190014 68420
rect 189954 68346 190560 68406
rect 149199 68332 149265 68335
rect 143904 68330 149265 68332
rect 143904 68274 149204 68330
rect 149260 68274 149265 68330
rect 143904 68272 149265 68274
rect 149199 68269 149265 68272
rect 640194 68006 640254 68568
rect 646863 68565 646929 68568
rect 184431 67592 184497 67595
rect 184431 67590 190560 67592
rect 184431 67534 184436 67590
rect 184492 67534 190560 67590
rect 184431 67532 190560 67534
rect 184431 67529 184497 67532
rect 149583 67148 149649 67151
rect 143904 67146 149649 67148
rect 143904 67090 149588 67146
rect 149644 67090 149649 67146
rect 143904 67088 149649 67090
rect 149583 67085 149649 67088
rect 184335 66852 184401 66855
rect 184335 66850 190560 66852
rect 184335 66794 184340 66850
rect 184396 66794 190560 66850
rect 184335 66792 190560 66794
rect 184335 66789 184401 66792
rect 645999 66260 646065 66263
rect 640194 66258 646065 66260
rect 640194 66202 646004 66258
rect 646060 66202 646065 66258
rect 640194 66200 646065 66202
rect 184335 66112 184401 66115
rect 184335 66110 190560 66112
rect 184335 66054 184340 66110
rect 184396 66054 190560 66110
rect 640194 66082 640254 66200
rect 645999 66197 646065 66200
rect 184335 66052 190560 66054
rect 184335 66049 184401 66052
rect 143874 65372 143934 65860
rect 149487 65372 149553 65375
rect 143874 65370 149553 65372
rect 143874 65314 149492 65370
rect 149548 65314 149553 65370
rect 143874 65312 149553 65314
rect 149487 65309 149553 65312
rect 184527 65224 184593 65227
rect 184527 65222 190560 65224
rect 184527 65166 184532 65222
rect 184588 65166 190560 65222
rect 184527 65164 190560 65166
rect 184527 65161 184593 65164
rect 149391 64632 149457 64635
rect 143904 64630 149457 64632
rect 143904 64574 149396 64630
rect 149452 64574 149457 64630
rect 143904 64572 149457 64574
rect 149391 64569 149457 64572
rect 184431 64632 184497 64635
rect 184431 64630 190014 64632
rect 184431 64574 184436 64630
rect 184492 64574 190014 64630
rect 184431 64572 190014 64574
rect 184431 64569 184497 64572
rect 189954 64558 190014 64572
rect 189954 64498 190560 64558
rect 647919 64188 647985 64191
rect 640416 64186 647985 64188
rect 640416 64130 647924 64186
rect 647980 64130 647985 64186
rect 640416 64128 647985 64130
rect 647919 64125 647985 64128
rect 184623 63744 184689 63747
rect 184623 63742 190560 63744
rect 184623 63686 184628 63742
rect 184684 63686 190560 63742
rect 184623 63684 190560 63686
rect 184623 63681 184689 63684
rect 149295 63448 149361 63451
rect 143904 63446 149361 63448
rect 143904 63390 149300 63446
rect 149356 63390 149361 63446
rect 143904 63388 149361 63390
rect 149295 63385 149361 63388
rect 184431 63152 184497 63155
rect 184431 63150 190014 63152
rect 184431 63094 184436 63150
rect 184492 63094 190014 63150
rect 184431 63092 190014 63094
rect 184431 63089 184497 63092
rect 189954 63078 190014 63092
rect 189954 63018 190560 63078
rect 149391 62264 149457 62267
rect 143904 62262 149457 62264
rect 143904 62206 149396 62262
rect 149452 62206 149457 62262
rect 143904 62204 149457 62206
rect 149391 62201 149457 62204
rect 184335 62264 184401 62267
rect 647919 62264 647985 62267
rect 184335 62262 190560 62264
rect 184335 62206 184340 62262
rect 184396 62206 190560 62262
rect 184335 62204 190560 62206
rect 640416 62262 647985 62264
rect 640416 62206 647924 62262
rect 647980 62206 647985 62262
rect 640416 62204 647985 62206
rect 184335 62201 184401 62204
rect 647919 62201 647985 62204
rect 184527 61524 184593 61527
rect 184527 61522 190014 61524
rect 184527 61466 184532 61522
rect 184588 61466 190014 61522
rect 184527 61464 190014 61466
rect 184527 61461 184593 61464
rect 189954 61450 190014 61464
rect 189954 61390 190560 61450
rect 143874 60636 143934 60976
rect 184623 60784 184689 60787
rect 184623 60782 190560 60784
rect 184623 60726 184628 60782
rect 184684 60726 190560 60782
rect 184623 60724 190560 60726
rect 184623 60721 184689 60724
rect 149487 60636 149553 60639
rect 143874 60634 149553 60636
rect 143874 60578 149492 60634
rect 149548 60578 149553 60634
rect 143874 60576 149553 60578
rect 149487 60573 149553 60576
rect 647055 60340 647121 60343
rect 640416 60338 647121 60340
rect 640416 60282 647060 60338
rect 647116 60282 647121 60338
rect 640416 60280 647121 60282
rect 647055 60277 647121 60280
rect 184431 60044 184497 60047
rect 184431 60042 190014 60044
rect 184431 59986 184436 60042
rect 184492 59986 190014 60042
rect 184431 59984 190014 59986
rect 184431 59981 184497 59984
rect 189954 59970 190014 59984
rect 189954 59910 190560 59970
rect 149391 59748 149457 59751
rect 143904 59746 149457 59748
rect 143904 59690 149396 59746
rect 149452 59690 149457 59746
rect 143904 59688 149457 59690
rect 149391 59685 149457 59688
rect 184335 59304 184401 59307
rect 184335 59302 190560 59304
rect 184335 59246 184340 59302
rect 184396 59246 190560 59302
rect 184335 59244 190560 59246
rect 184335 59241 184401 59244
rect 645999 59008 646065 59011
rect 640386 59006 646065 59008
rect 640386 58950 646004 59006
rect 646060 58950 646065 59006
rect 640386 58948 646065 58950
rect 149391 58564 149457 58567
rect 143904 58562 149457 58564
rect 143904 58506 149396 58562
rect 149452 58506 149457 58562
rect 143904 58504 149457 58506
rect 149391 58501 149457 58504
rect 184527 58416 184593 58419
rect 184527 58414 190560 58416
rect 184527 58358 184532 58414
rect 184588 58358 190560 58414
rect 640386 58386 640446 58948
rect 645999 58945 646065 58948
rect 184527 58356 190560 58358
rect 184527 58353 184593 58356
rect 184335 57676 184401 57679
rect 184335 57674 190560 57676
rect 184335 57618 184340 57674
rect 184396 57618 190560 57674
rect 184335 57616 190560 57618
rect 184335 57613 184401 57616
rect 149487 57380 149553 57383
rect 143904 57378 149553 57380
rect 143904 57322 149492 57378
rect 149548 57322 149553 57378
rect 143904 57320 149553 57322
rect 149487 57317 149553 57320
rect 646767 57084 646833 57087
rect 640386 57082 646833 57084
rect 640386 57026 646772 57082
rect 646828 57026 646833 57082
rect 640386 57024 646833 57026
rect 184335 56936 184401 56939
rect 184335 56934 190560 56936
rect 184335 56878 184340 56934
rect 184396 56878 190560 56934
rect 184335 56876 190560 56878
rect 184335 56873 184401 56876
rect 640386 56536 640446 57024
rect 646767 57021 646833 57024
rect 149391 56196 149457 56199
rect 143874 56194 149457 56196
rect 143874 56138 149396 56194
rect 149452 56138 149457 56194
rect 143874 56136 149457 56138
rect 143874 56092 143934 56136
rect 149391 56133 149457 56136
rect 184335 56196 184401 56199
rect 184335 56194 190560 56196
rect 184335 56138 184340 56194
rect 184396 56138 190560 56194
rect 184335 56136 190560 56138
rect 184335 56133 184401 56136
rect 184431 55456 184497 55459
rect 184431 55454 190560 55456
rect 184431 55398 184436 55454
rect 184492 55398 190560 55454
rect 184431 55396 190560 55398
rect 184431 55393 184497 55396
rect 149679 54864 149745 54867
rect 143904 54862 149745 54864
rect 143904 54806 149684 54862
rect 149740 54806 149745 54862
rect 143904 54804 149745 54806
rect 149679 54801 149745 54804
rect 184335 54716 184401 54719
rect 646479 54716 646545 54719
rect 184335 54714 190014 54716
rect 184335 54658 184340 54714
rect 184396 54658 190014 54714
rect 184335 54656 190014 54658
rect 184335 54653 184401 54656
rect 189954 54642 190014 54656
rect 640386 54714 646545 54716
rect 640386 54658 646484 54714
rect 646540 54658 646545 54714
rect 640386 54656 646545 54658
rect 189954 54582 190560 54642
rect 640386 54612 640446 54656
rect 646479 54653 646545 54656
rect 184335 53976 184401 53979
rect 184335 53974 190560 53976
rect 184335 53918 184340 53974
rect 184396 53918 190560 53974
rect 184335 53916 190560 53918
rect 184335 53913 184401 53916
rect 149391 53828 149457 53831
rect 143904 53826 149457 53828
rect 143904 53770 149396 53826
rect 149452 53770 149457 53826
rect 143904 53768 149457 53770
rect 149391 53765 149457 53768
rect 417519 44948 417585 44951
rect 472239 44948 472305 44951
rect 417474 44946 417585 44948
rect 417474 44890 417524 44946
rect 417580 44890 417585 44946
rect 417474 44885 417585 44890
rect 472194 44946 472305 44948
rect 472194 44890 472244 44946
rect 472300 44890 472305 44946
rect 472194 44885 472305 44890
rect 417474 44404 417534 44885
rect 472194 44404 472254 44885
rect 415215 41988 415281 41991
rect 415215 41986 417630 41988
rect 415215 41930 415220 41986
rect 415276 41930 417630 41986
rect 415215 41928 417630 41930
rect 415215 41925 415281 41928
rect 416847 41840 416913 41843
rect 416847 41838 416958 41840
rect 416847 41782 416852 41838
rect 416908 41782 416958 41838
rect 416847 41777 416958 41782
rect 416898 40508 416958 41777
rect 417570 40656 417630 41928
rect 464847 41840 464913 41843
rect 457890 41838 464913 41840
rect 457890 41782 464852 41838
rect 464908 41782 464913 41838
rect 457890 41780 464913 41782
rect 457890 40656 457950 41780
rect 464847 41777 464913 41780
rect 470319 41840 470385 41843
rect 512175 41840 512241 41843
rect 525903 41840 525969 41843
rect 470319 41838 478110 41840
rect 470319 41782 470324 41838
rect 470380 41782 478110 41838
rect 470319 41780 478110 41782
rect 470319 41777 470385 41780
rect 417570 40596 457950 40656
rect 417466 40508 417472 40510
rect 416898 40448 417472 40508
rect 417466 40446 417472 40448
rect 417536 40446 417542 40510
rect 417658 40446 417664 40510
rect 417728 40508 417734 40510
rect 420783 40508 420849 40511
rect 417728 40506 420849 40508
rect 417728 40450 420788 40506
rect 420844 40450 420849 40506
rect 417728 40448 420849 40450
rect 478050 40508 478110 41780
rect 512175 41838 525969 41840
rect 512175 41782 512180 41838
rect 512236 41782 525908 41838
rect 525964 41782 525969 41838
rect 512175 41780 525969 41782
rect 512175 41777 512241 41780
rect 525903 41777 525969 41780
rect 539727 40508 539793 40511
rect 478050 40506 539793 40508
rect 478050 40450 539732 40506
rect 539788 40450 539793 40506
rect 478050 40448 539793 40450
rect 417728 40446 417734 40448
rect 420783 40445 420849 40448
rect 539727 40445 539793 40448
rect 142095 40212 142161 40215
rect 141762 40210 142161 40212
rect 141762 40154 142100 40210
rect 142156 40154 142161 40210
rect 141762 40152 142161 40154
rect 141762 39886 141822 40152
rect 142095 40149 142161 40152
rect 311055 37252 311121 37255
rect 331215 37252 331281 37255
rect 311055 37250 331281 37252
rect 311055 37194 311060 37250
rect 311116 37194 331220 37250
rect 331276 37194 331281 37250
rect 311055 37192 331281 37194
rect 311055 37189 311121 37192
rect 331215 37189 331281 37192
rect 311151 31628 311217 31631
rect 328335 31628 328401 31631
rect 311151 31626 328401 31628
rect 311151 31570 311156 31626
rect 311212 31570 328340 31626
rect 328396 31570 328401 31626
rect 311151 31568 328401 31570
rect 311151 31565 311217 31568
rect 328335 31565 328401 31568
<< via3 >>
rect 40384 815078 40448 815142
rect 40576 814042 40640 814106
rect 41536 810194 41600 810258
rect 41344 802054 41408 802118
rect 42688 800930 42752 800934
rect 42688 800874 42740 800930
rect 42740 800874 42752 800930
rect 42688 800870 42752 800874
rect 41728 800486 41792 800490
rect 41728 800430 41740 800486
rect 41740 800430 41792 800486
rect 41728 800426 41792 800430
rect 42112 800486 42176 800490
rect 42112 800430 42124 800486
rect 42124 800430 42176 800486
rect 42112 800426 42176 800430
rect 41920 800338 41984 800342
rect 41920 800282 41972 800338
rect 41972 800282 41984 800338
rect 41920 800278 41984 800282
rect 41728 794270 41792 794274
rect 41728 794214 41780 794270
rect 41780 794214 41792 794270
rect 41728 794210 41792 794214
rect 42688 793530 42752 793534
rect 42688 793474 42740 793530
rect 42740 793474 42752 793530
rect 42688 793470 42752 793474
rect 41920 792938 41984 792942
rect 41920 792882 41972 792938
rect 41972 792882 41984 792938
rect 41920 792878 41984 792882
rect 42112 790126 42176 790130
rect 42112 790070 42164 790126
rect 42164 790070 42176 790126
rect 42112 790066 42176 790070
rect 41344 789326 41408 789390
rect 41536 789178 41600 789242
rect 674752 787994 674816 788058
rect 676096 787402 676160 787466
rect 675520 786722 675584 786726
rect 675520 786666 675532 786722
rect 675532 786666 675584 786722
rect 675520 786662 675584 786666
rect 675136 784738 675200 784802
rect 674368 784146 674432 784210
rect 673984 783406 674048 783470
rect 676480 782962 676544 783026
rect 675712 780654 675776 780658
rect 675712 780598 675724 780654
rect 675724 780598 675776 780654
rect 675712 780594 675776 780598
rect 676288 779854 676352 779918
rect 676672 779114 676736 779178
rect 675328 777634 675392 777698
rect 675904 775414 675968 775478
rect 40576 772898 40640 772962
rect 676096 772010 676160 772074
rect 40384 771808 40448 771872
rect 40576 771862 40640 771926
rect 675520 771862 675584 771926
rect 40576 770826 40640 770890
rect 40768 766978 40832 767042
rect 41728 764610 41792 764674
rect 40960 759874 41024 759938
rect 42880 757862 42944 757866
rect 42880 757806 42892 757862
rect 42892 757806 42944 757862
rect 42880 757802 42944 757806
rect 42112 757358 42176 757422
rect 42304 757210 42368 757274
rect 41920 757122 41984 757126
rect 41920 757066 41972 757122
rect 41972 757066 41984 757122
rect 41920 757062 41984 757066
rect 41920 754902 41984 754906
rect 41920 754846 41972 754902
rect 41972 754846 41984 754902
rect 41920 754842 41984 754846
rect 42880 751350 42944 751354
rect 42880 751294 42932 751350
rect 42932 751294 42944 751350
rect 42880 751290 42944 751294
rect 42112 747738 42176 747802
rect 41728 747502 41792 747506
rect 41728 747446 41780 747502
rect 41780 747446 41792 747502
rect 41728 747442 41792 747446
rect 40768 747146 40832 747210
rect 42304 746850 42368 746914
rect 40960 746554 41024 746618
rect 676288 745814 676352 745878
rect 677248 745814 677312 745878
rect 676480 743002 676544 743066
rect 676864 743002 676928 743066
rect 674176 742410 674240 742474
rect 674944 741078 675008 741142
rect 674560 740338 674624 740402
rect 675520 739214 675584 739218
rect 675520 739158 675532 739214
rect 675532 739158 675584 739214
rect 675520 739154 675584 739158
rect 676288 735454 676352 735518
rect 676096 730570 676160 730634
rect 676864 729830 676928 729894
rect 677056 729386 677120 729450
rect 40576 729238 40640 729302
rect 40384 728706 40448 728710
rect 40384 728650 40436 728706
rect 40436 728650 40448 728706
rect 40384 728646 40448 728650
rect 676672 728054 676736 728118
rect 677248 728054 677312 728118
rect 40576 727610 40640 727674
rect 41920 721394 41984 721458
rect 41728 720950 41792 721014
rect 40576 716658 40640 716722
rect 40384 716066 40448 716130
rect 43072 714142 43136 714206
rect 42880 713994 42944 714058
rect 42112 713906 42176 713910
rect 42112 713850 42124 713906
rect 42124 713850 42176 713906
rect 42112 713846 42176 713850
rect 42496 712278 42560 712282
rect 42496 712222 42508 712278
rect 42508 712222 42560 712278
rect 42496 712218 42560 712222
rect 42112 711686 42176 711690
rect 42112 711630 42124 711686
rect 42124 711630 42176 711686
rect 42112 711626 42176 711630
rect 42688 711626 42752 711690
rect 42304 711478 42368 711542
rect 42688 711182 42752 711246
rect 42304 711034 42368 711098
rect 675904 710590 675968 710654
rect 674752 710442 674816 710506
rect 675136 709702 675200 709766
rect 675712 709110 675776 709174
rect 41920 708814 41984 708878
rect 42880 707986 42944 707990
rect 42880 707930 42932 707986
rect 42932 707930 42944 707986
rect 42880 707926 42944 707930
rect 674368 707630 674432 707694
rect 41728 707394 41792 707398
rect 41728 707338 41780 707394
rect 41780 707338 41792 707394
rect 41728 707334 41792 707338
rect 673984 707038 674048 707102
rect 675328 706890 675392 706954
rect 677248 706446 677312 706510
rect 677056 705854 677120 705918
rect 676864 705410 676928 705474
rect 40576 705114 40640 705178
rect 42496 704818 42560 704882
rect 43072 703546 43136 703550
rect 43072 703490 43084 703546
rect 43084 703490 43136 703546
rect 43072 703486 43136 703490
rect 40384 699934 40448 699998
rect 675136 697862 675200 697926
rect 674368 697122 674432 697186
rect 674752 696974 674816 697038
rect 675712 694962 675776 694966
rect 675712 694906 675724 694962
rect 675724 694906 675776 694962
rect 675712 694902 675776 694906
rect 675328 694666 675392 694670
rect 675328 694610 675340 694666
rect 675340 694610 675392 694666
rect 675328 694606 675392 694610
rect 40384 685430 40448 685494
rect 40576 684394 40640 684458
rect 40576 672406 40640 672470
rect 41152 671074 41216 671138
rect 42304 670630 42368 670694
rect 674944 666190 675008 666254
rect 42304 665006 42368 665070
rect 676096 664858 676160 664922
rect 674560 664710 674624 664774
rect 676288 664414 676352 664478
rect 674176 663378 674240 663442
rect 675520 662638 675584 662702
rect 41152 662342 41216 662406
rect 40576 660714 40640 660778
rect 673984 652722 674048 652786
rect 674176 652130 674240 652194
rect 674944 651390 675008 651454
rect 674560 649614 674624 649678
rect 675520 645382 675584 645386
rect 675520 645326 675532 645382
rect 675532 645326 675584 645382
rect 675520 645322 675584 645326
rect 40768 644730 40832 644794
rect 40384 642214 40448 642278
rect 40576 642214 40640 642278
rect 42880 642214 42944 642278
rect 676096 640290 676160 640354
rect 675904 638514 675968 638578
rect 40768 629190 40832 629254
rect 40576 628302 40640 628366
rect 43072 627562 43136 627626
rect 41920 627414 41984 627478
rect 42304 627414 42368 627478
rect 41920 625194 41984 625258
rect 42304 622086 42368 622150
rect 674752 620902 674816 620966
rect 675136 619866 675200 619930
rect 675712 619422 675776 619486
rect 43072 619126 43136 619190
rect 674368 617942 674432 618006
rect 675328 617794 675392 617858
rect 40576 616462 40640 616526
rect 40768 616314 40832 616378
rect 674368 607730 674432 607794
rect 675136 606014 675200 606018
rect 675136 605958 675188 606014
rect 675188 605958 675200 606014
rect 675136 605954 675200 605958
rect 674752 604770 674816 604834
rect 40384 601722 40448 601726
rect 40384 601666 40396 601722
rect 40396 601666 40448 601722
rect 40384 601662 40448 601666
rect 675328 600182 675392 600246
rect 43072 599442 43136 599506
rect 676288 595298 676352 595362
rect 675712 593434 675776 593438
rect 675712 593378 675724 593434
rect 675724 593378 675776 593434
rect 675712 593374 675776 593378
rect 40384 585678 40448 585742
rect 40576 585234 40640 585298
rect 42688 584790 42752 584854
rect 41920 584258 41984 584262
rect 41920 584202 41932 584258
rect 41932 584202 41984 584258
rect 41920 584198 41984 584202
rect 42304 584258 42368 584262
rect 42304 584202 42316 584258
rect 42316 584202 42368 584258
rect 42304 584198 42368 584202
rect 42688 578722 42752 578786
rect 42304 578278 42368 578342
rect 40576 575318 40640 575382
rect 40384 573986 40448 574050
rect 674944 573986 675008 574050
rect 676096 573690 676160 573754
rect 673984 572802 674048 572866
rect 41920 572714 41984 572718
rect 41920 572658 41932 572714
rect 41932 572658 41984 572714
rect 41920 572654 41984 572658
rect 674560 572506 674624 572570
rect 675520 571914 675584 571978
rect 675904 571322 675968 571386
rect 674176 571174 674240 571238
rect 675520 562502 675584 562506
rect 675520 562446 675532 562502
rect 675532 562446 675584 562502
rect 675520 562442 675584 562446
rect 674176 561702 674240 561766
rect 674944 561406 675008 561470
rect 674560 558890 674624 558954
rect 40384 539798 40448 539862
rect 41152 538022 41216 538086
rect 42880 536986 42944 537050
rect 40960 536246 41024 536310
rect 40768 535062 40832 535126
rect 41536 534174 41600 534238
rect 40576 533878 40640 533942
rect 41728 533198 41792 533202
rect 41728 533142 41780 533198
rect 41780 533142 41792 533198
rect 41728 533138 41792 533142
rect 41344 530770 41408 530834
rect 675136 530770 675200 530834
rect 41920 530090 41984 530094
rect 41920 530034 41932 530090
rect 41932 530034 41984 530090
rect 41920 530030 41984 530034
rect 676288 530474 676352 530538
rect 674368 529882 674432 529946
rect 42112 529350 42176 529354
rect 42112 529294 42124 529350
rect 42124 529294 42176 529350
rect 42112 529290 42176 529294
rect 674752 529290 674816 529354
rect 42304 528698 42368 528762
rect 675328 528698 675392 528762
rect 675712 528106 675776 528170
rect 42496 527070 42560 527134
rect 674944 486370 675008 486434
rect 675520 485630 675584 485694
rect 674176 483410 674240 483474
rect 674560 482818 674624 482882
rect 42496 471570 42560 471634
rect 41152 471274 41216 471338
rect 42304 470090 42368 470154
rect 41728 469498 41792 469562
rect 40384 469350 40448 469414
rect 42112 468018 42176 468082
rect 41920 467426 41984 467490
rect 40960 467278 41024 467342
rect 41536 466834 41600 466898
rect 41344 466242 41408 466306
rect 40576 465798 40640 465862
rect 40768 465354 40832 465418
rect 41536 422286 41600 422350
rect 40384 421842 40448 421906
rect 42496 421694 42560 421758
rect 40576 421250 40640 421314
rect 40960 417698 41024 417762
rect 41920 417254 41984 417318
rect 41728 416958 41792 417022
rect 42112 416810 42176 416874
rect 41152 416366 41216 416430
rect 42304 416218 42368 416282
rect 41344 414886 41408 414950
rect 40384 411186 40448 411250
rect 40960 407634 41024 407698
rect 42112 406066 42176 406070
rect 42112 406010 42124 406066
rect 42124 406010 42176 406066
rect 42112 406006 42176 406010
rect 41728 403846 41792 403850
rect 41728 403790 41780 403846
rect 41780 403790 41792 403846
rect 41728 403786 41792 403790
rect 42304 403046 42368 403110
rect 41920 402662 41984 402666
rect 41920 402606 41932 402662
rect 41932 402606 41984 402662
rect 41920 402602 41984 402606
rect 41344 401862 41408 401926
rect 41536 400086 41600 400150
rect 41152 399346 41216 399410
rect 40576 398754 40640 398818
rect 676672 397866 676736 397930
rect 673984 397570 674048 397634
rect 675136 396830 675200 396894
rect 676672 396386 676736 396450
rect 674752 396090 674816 396154
rect 675904 395202 675968 395266
rect 675328 394610 675392 394674
rect 676480 393870 676544 393934
rect 676096 393278 676160 393342
rect 674368 393130 674432 393194
rect 675712 392538 675776 392602
rect 675520 391798 675584 391862
rect 676288 391354 676352 391418
rect 42496 388690 42560 388754
rect 675136 385938 675200 385942
rect 675136 385882 675188 385938
rect 675188 385882 675200 385938
rect 675136 385878 675200 385882
rect 675904 385582 675968 385646
rect 674944 384398 675008 384462
rect 676672 382918 676736 382982
rect 675328 382326 675392 382390
rect 676480 381734 676544 381798
rect 675712 381202 675776 381206
rect 675712 381146 675764 381202
rect 675764 381146 675776 381202
rect 675712 381142 675776 381146
rect 39808 380254 39872 380318
rect 40576 379810 40640 379874
rect 40000 379218 40064 379282
rect 42304 378774 42368 378838
rect 674752 378774 674816 378838
rect 675520 378094 675584 378098
rect 675520 378038 675572 378094
rect 675572 378038 675584 378094
rect 675520 378034 675584 378038
rect 674368 377146 674432 377210
rect 676288 376702 676352 376766
rect 41344 375814 41408 375878
rect 676096 375666 676160 375730
rect 40960 373890 41024 373954
rect 673984 373890 674048 373954
rect 41728 373742 41792 373806
rect 41920 373298 41984 373362
rect 42112 373150 42176 373214
rect 39808 372410 39872 372474
rect 42496 372410 42560 372474
rect 40768 372262 40832 372326
rect 41728 368178 41792 368182
rect 41728 368122 41780 368178
rect 41780 368122 41792 368178
rect 41728 368118 41792 368122
rect 40384 362790 40448 362854
rect 41344 360570 41408 360634
rect 41920 359890 41984 359894
rect 41920 359834 41972 359890
rect 41972 359834 41984 359890
rect 41920 359830 41984 359834
rect 42112 359298 42176 359302
rect 42112 359242 42124 359298
rect 42124 359242 42176 359298
rect 42112 359238 42176 359242
rect 40576 358794 40640 358858
rect 40768 357166 40832 357230
rect 41920 357166 41984 357230
rect 41920 356930 41984 356934
rect 41920 356874 41932 356930
rect 41932 356874 41984 356930
rect 41920 356870 41984 356874
rect 40960 356130 41024 356194
rect 42496 355538 42560 355602
rect 674176 355834 674240 355898
rect 673984 355242 674048 355306
rect 674368 354206 674432 354270
rect 675904 353762 675968 353826
rect 674560 353170 674624 353234
rect 674752 351690 674816 351754
rect 674944 348730 675008 348794
rect 41728 343166 41792 343170
rect 41728 343110 41740 343166
rect 41740 343110 41792 343166
rect 41728 343106 41792 343110
rect 675712 342958 675776 343022
rect 676672 342810 676736 342874
rect 675904 339554 675968 339618
rect 41920 338814 41984 338878
rect 40384 336594 40448 336658
rect 40768 336002 40832 336066
rect 40960 335114 41024 335178
rect 41344 334522 41408 334586
rect 41152 334078 41216 334142
rect 674752 333486 674816 333550
rect 41536 332598 41600 332662
rect 674944 332302 675008 332366
rect 40576 332006 40640 332070
rect 41728 331118 41792 331182
rect 42304 330674 42368 330738
rect 675712 330586 675776 330590
rect 675712 330530 675764 330586
rect 675764 330530 675776 330586
rect 675712 330526 675776 330530
rect 42112 329046 42176 329110
rect 674560 328306 674624 328370
rect 676672 326826 676736 326890
rect 41728 324962 41792 324966
rect 41728 324906 41780 324962
rect 41780 324906 41792 324962
rect 41728 324902 41792 324906
rect 40576 320462 40640 320526
rect 40768 319722 40832 319786
rect 41536 317354 41600 317418
rect 41152 316614 41216 316678
rect 41344 316170 41408 316234
rect 40384 315430 40448 315494
rect 42112 313714 42176 313718
rect 42112 313658 42124 313714
rect 42124 313658 42176 313714
rect 42112 313654 42176 313658
rect 40960 313062 41024 313126
rect 42304 312470 42368 312534
rect 674176 310990 674240 311054
rect 675520 310398 675584 310462
rect 674176 309806 674240 309870
rect 674560 309066 674624 309130
rect 674368 308918 674432 308982
rect 674752 308326 674816 308390
rect 675712 306402 675776 306466
rect 675328 305958 675392 306022
rect 674944 305366 675008 305430
rect 675136 303442 675200 303506
rect 673984 302554 674048 302618
rect 675904 302406 675968 302470
rect 676096 299150 676160 299214
rect 41728 294562 41792 294626
rect 41920 294118 41984 294182
rect 41152 293378 41216 293442
rect 41536 292934 41600 292998
rect 675712 292846 675776 292850
rect 675712 292790 675724 292846
rect 675724 292790 675776 292846
rect 675712 292786 675776 292790
rect 40384 291898 40448 291962
rect 40960 291454 41024 291518
rect 41344 290862 41408 290926
rect 675904 290714 675968 290778
rect 40576 289382 40640 289446
rect 675328 288494 675392 288558
rect 673984 287162 674048 287226
rect 675136 285238 675200 285302
rect 42112 285090 42176 285154
rect 676096 283610 676160 283674
rect 674944 281834 675008 281898
rect 41728 281686 41792 281750
rect 42496 281598 42560 281602
rect 42496 281542 42508 281598
rect 42508 281542 42560 281598
rect 42496 281538 42560 281542
rect 42304 278578 42368 278642
rect 43072 278430 43136 278494
rect 674176 278430 674240 278494
rect 674752 278134 674816 278198
rect 42496 277986 42560 278050
rect 41536 276506 41600 276570
rect 674560 276506 674624 276570
rect 40576 274138 40640 274202
rect 674368 274138 674432 274202
rect 41344 273546 41408 273610
rect 40960 272806 41024 272870
rect 41152 272362 41216 272426
rect 42112 270646 42176 270650
rect 42112 270590 42124 270646
rect 42124 270590 42176 270646
rect 42112 270586 42176 270590
rect 40384 269994 40448 270058
rect 41920 269314 41984 269318
rect 41920 269258 41932 269314
rect 41932 269258 41984 269314
rect 41920 269254 41984 269258
rect 675520 265702 675584 265766
rect 673984 263186 674048 263250
rect 675520 262742 675584 262806
rect 676288 261410 676352 261474
rect 675712 260670 675776 260734
rect 674368 258302 674432 258366
rect 674944 257710 675008 257774
rect 675904 253270 675968 253334
rect 676096 253122 676160 253186
rect 41920 251938 41984 252002
rect 41536 251198 41600 251262
rect 42112 250902 42176 250966
rect 676288 250754 676352 250818
rect 40960 250162 41024 250226
rect 40576 249718 40640 249782
rect 675520 249630 675584 249634
rect 675520 249574 675572 249630
rect 675572 249574 675584 249630
rect 675520 249570 675584 249574
rect 40768 248682 40832 248746
rect 41344 248238 41408 248302
rect 41152 247646 41216 247710
rect 40384 246166 40448 246230
rect 675712 243562 675776 243566
rect 675712 243506 675724 243562
rect 675724 243506 675776 243562
rect 675712 243502 675776 243506
rect 674944 242022 675008 242086
rect 674368 240542 674432 240606
rect 676096 238618 676160 238682
rect 41536 237878 41600 237942
rect 675904 236842 675968 236906
rect 40576 233290 40640 233354
rect 40384 231070 40448 231134
rect 41152 230330 41216 230394
rect 41344 229738 41408 229802
rect 40960 228998 41024 229062
rect 41536 227370 41600 227434
rect 40768 226630 40832 226694
rect 42112 226246 42176 226250
rect 42112 226190 42124 226246
rect 42124 226190 42176 226246
rect 42112 226186 42176 226190
rect 674176 219970 674240 220034
rect 675328 219082 675392 219146
rect 673984 218490 674048 218554
rect 674368 217898 674432 217962
rect 675904 217602 675968 217666
rect 675712 216048 675776 216112
rect 676096 215234 676160 215298
rect 675520 213458 675584 213522
rect 674560 213014 674624 213078
rect 676672 207538 676736 207602
rect 676480 207390 676544 207454
rect 40768 207094 40832 207158
rect 41152 205466 41216 205530
rect 40960 205022 41024 205086
rect 42112 204726 42176 204790
rect 675904 204430 675968 204494
rect 41920 203172 41984 203236
rect 675712 202714 675776 202718
rect 675712 202658 675724 202714
rect 675724 202658 675776 202714
rect 675712 202654 675776 202658
rect 42304 201026 42368 201090
rect 675520 201382 675584 201386
rect 675520 201326 675572 201382
rect 675572 201326 675584 201382
rect 675520 201322 675584 201326
rect 41728 200434 41792 200498
rect 41344 199990 41408 200054
rect 41536 199546 41600 199610
rect 676096 198362 676160 198426
rect 41728 195314 41792 195318
rect 41728 195258 41780 195314
rect 41780 195258 41792 195314
rect 41728 195254 41792 195258
rect 674560 195254 674624 195318
rect 676480 193478 676544 193542
rect 676672 191554 676736 191618
rect 41536 190074 41600 190138
rect 41920 187914 41984 187918
rect 41920 187858 41932 187914
rect 41932 187858 41984 187914
rect 41920 187854 41984 187858
rect 42112 187174 42176 187178
rect 42112 187118 42164 187174
rect 42164 187118 42176 187174
rect 42112 187114 42176 187118
rect 40960 186374 41024 186438
rect 40768 185782 40832 185846
rect 41344 184154 41408 184218
rect 41152 183414 41216 183478
rect 42304 182970 42368 183034
rect 674176 176162 674240 176226
rect 674560 175570 674624 175634
rect 675328 175422 675392 175486
rect 673984 174682 674048 174746
rect 674368 174090 674432 174154
rect 674176 173498 674240 173562
rect 676288 172906 676352 172970
rect 674752 172610 674816 172674
rect 675712 171648 675776 171712
rect 675328 171130 675392 171194
rect 676096 170390 676160 170454
rect 674944 168614 675008 168678
rect 675520 168170 675584 168234
rect 675904 167578 675968 167642
rect 675136 167134 675200 167198
rect 676288 159290 676352 159354
rect 675712 157722 675776 157726
rect 675712 157666 675764 157722
rect 675764 157666 675776 157722
rect 675712 157662 675776 157666
rect 675904 155442 675968 155506
rect 675328 153370 675392 153434
rect 675136 152482 675200 152546
rect 675520 152246 675584 152250
rect 675520 152190 675532 152246
rect 675532 152190 675584 152246
rect 675520 152186 675584 152190
rect 674944 150262 675008 150326
rect 674752 148486 674816 148550
rect 676096 146562 676160 146626
rect 674368 130578 674432 130642
rect 673984 129394 674048 129458
rect 674176 128506 674240 128570
rect 675712 125546 675776 125610
rect 673984 123030 674048 123094
rect 675520 122142 675584 122206
rect 675904 116666 675968 116730
rect 676672 116074 676736 116138
rect 675712 108142 675776 108146
rect 675712 108086 675764 108142
rect 675764 108086 675776 108142
rect 675712 108082 675776 108086
rect 675520 106662 675584 106666
rect 675520 106606 675532 106662
rect 675532 106606 675584 106662
rect 675520 106602 675584 106606
rect 673984 105122 674048 105186
rect 675904 103198 675968 103262
rect 676672 101422 676736 101486
rect 417472 40446 417536 40510
rect 417664 40446 417728 40510
<< metal4 >>
rect 40383 815142 40449 815143
rect 40383 815078 40384 815142
rect 40448 815078 40449 815142
rect 40383 815077 40449 815078
rect 40386 772257 40446 815077
rect 40575 814106 40641 814107
rect 40575 814042 40576 814106
rect 40640 814042 40641 814106
rect 40575 814041 40641 814042
rect 40578 772963 40638 814041
rect 41535 810258 41601 810259
rect 41535 810194 41536 810258
rect 41600 810194 41601 810258
rect 41535 810193 41601 810194
rect 41343 802118 41409 802119
rect 41343 802054 41344 802118
rect 41408 802054 41409 802118
rect 41343 802053 41409 802054
rect 41346 789391 41406 802053
rect 41343 789390 41409 789391
rect 41343 789326 41344 789390
rect 41408 789326 41409 789390
rect 41343 789325 41409 789326
rect 41538 789243 41598 810193
rect 42687 800934 42753 800935
rect 42687 800870 42688 800934
rect 42752 800870 42753 800934
rect 42687 800869 42753 800870
rect 41727 800490 41793 800491
rect 41727 800426 41728 800490
rect 41792 800426 41793 800490
rect 41727 800425 41793 800426
rect 42111 800490 42177 800491
rect 42111 800426 42112 800490
rect 42176 800426 42177 800490
rect 42111 800425 42177 800426
rect 41730 794275 41790 800425
rect 41919 800342 41985 800343
rect 41919 800278 41920 800342
rect 41984 800278 41985 800342
rect 41919 800277 41985 800278
rect 41727 794274 41793 794275
rect 41727 794210 41728 794274
rect 41792 794210 41793 794274
rect 41727 794209 41793 794210
rect 41922 792943 41982 800277
rect 41919 792942 41985 792943
rect 41919 792878 41920 792942
rect 41984 792878 41985 792942
rect 41919 792877 41985 792878
rect 42114 790131 42174 800425
rect 42690 793535 42750 800869
rect 42687 793534 42753 793535
rect 42687 793470 42688 793534
rect 42752 793470 42753 793534
rect 42687 793469 42753 793470
rect 42111 790130 42177 790131
rect 42111 790066 42112 790130
rect 42176 790066 42177 790130
rect 42111 790065 42177 790066
rect 41535 789242 41601 789243
rect 41535 789178 41536 789242
rect 41600 789178 41601 789242
rect 41535 789177 41601 789178
rect 674751 788058 674817 788059
rect 674751 787994 674752 788058
rect 674816 787994 674817 788058
rect 674751 787993 674817 787994
rect 674367 784210 674433 784211
rect 674367 784146 674368 784210
rect 674432 784146 674433 784210
rect 674367 784145 674433 784146
rect 673983 783470 674049 783471
rect 673983 783406 673984 783470
rect 674048 783406 674049 783470
rect 673983 783405 674049 783406
rect 40575 772962 40641 772963
rect 40575 772898 40576 772962
rect 40640 772898 40641 772962
rect 40575 772897 40641 772898
rect 40386 772197 40638 772257
rect 40578 771927 40638 772197
rect 40575 771926 40641 771927
rect 40383 771872 40449 771873
rect 40383 771870 40384 771872
rect 40194 771810 40384 771870
rect 40194 771591 40254 771810
rect 40383 771808 40384 771810
rect 40448 771808 40449 771872
rect 40575 771862 40576 771926
rect 40640 771862 40641 771926
rect 40575 771861 40641 771862
rect 40383 771807 40449 771808
rect 40194 771531 40446 771591
rect 40386 728711 40446 771531
rect 40575 770890 40641 770891
rect 40575 770826 40576 770890
rect 40640 770826 40641 770890
rect 40575 770825 40641 770826
rect 40578 729303 40638 770825
rect 40767 767042 40833 767043
rect 40767 766978 40768 767042
rect 40832 766978 40833 767042
rect 40767 766977 40833 766978
rect 40770 747211 40830 766977
rect 41727 764674 41793 764675
rect 41727 764610 41728 764674
rect 41792 764610 41793 764674
rect 41727 764609 41793 764610
rect 40959 759938 41025 759939
rect 40959 759874 40960 759938
rect 41024 759874 41025 759938
rect 40959 759873 41025 759874
rect 40767 747210 40833 747211
rect 40767 747146 40768 747210
rect 40832 747146 40833 747210
rect 40767 747145 40833 747146
rect 40962 746619 41022 759873
rect 41730 747507 41790 764609
rect 42879 757866 42945 757867
rect 42879 757802 42880 757866
rect 42944 757802 42945 757866
rect 42879 757801 42945 757802
rect 42111 757422 42177 757423
rect 42111 757358 42112 757422
rect 42176 757358 42177 757422
rect 42111 757357 42177 757358
rect 41919 757126 41985 757127
rect 41919 757062 41920 757126
rect 41984 757062 41985 757126
rect 41919 757061 41985 757062
rect 41922 754907 41982 757061
rect 41919 754906 41985 754907
rect 41919 754842 41920 754906
rect 41984 754842 41985 754906
rect 41919 754841 41985 754842
rect 42114 747803 42174 757357
rect 42303 757274 42369 757275
rect 42303 757210 42304 757274
rect 42368 757210 42369 757274
rect 42303 757209 42369 757210
rect 42111 747802 42177 747803
rect 42111 747738 42112 747802
rect 42176 747738 42177 747802
rect 42111 747737 42177 747738
rect 41727 747506 41793 747507
rect 41727 747442 41728 747506
rect 41792 747442 41793 747506
rect 41727 747441 41793 747442
rect 42306 746915 42366 757209
rect 42882 751355 42942 757801
rect 42879 751354 42945 751355
rect 42879 751290 42880 751354
rect 42944 751290 42945 751354
rect 42879 751289 42945 751290
rect 42303 746914 42369 746915
rect 42303 746850 42304 746914
rect 42368 746850 42369 746914
rect 42303 746849 42369 746850
rect 40959 746618 41025 746619
rect 40959 746554 40960 746618
rect 41024 746554 41025 746618
rect 40959 746553 41025 746554
rect 40575 729302 40641 729303
rect 40575 729238 40576 729302
rect 40640 729238 40641 729302
rect 40575 729237 40641 729238
rect 40383 728710 40449 728711
rect 40383 728646 40384 728710
rect 40448 728646 40449 728710
rect 40383 728645 40449 728646
rect 40578 727675 40638 729237
rect 40575 727674 40641 727675
rect 40575 727610 40576 727674
rect 40640 727610 40641 727674
rect 40575 727609 40641 727610
rect 41919 721458 41985 721459
rect 41919 721394 41920 721458
rect 41984 721394 41985 721458
rect 41919 721393 41985 721394
rect 41727 721014 41793 721015
rect 41727 720950 41728 721014
rect 41792 720950 41793 721014
rect 41727 720949 41793 720950
rect 40575 716722 40641 716723
rect 40575 716658 40576 716722
rect 40640 716658 40641 716722
rect 40575 716657 40641 716658
rect 40383 716130 40449 716131
rect 40383 716066 40384 716130
rect 40448 716066 40449 716130
rect 40383 716065 40449 716066
rect 40386 699999 40446 716065
rect 40578 705179 40638 716657
rect 41730 707399 41790 720949
rect 41922 708879 41982 721393
rect 43071 714206 43137 714207
rect 43071 714142 43072 714206
rect 43136 714142 43137 714206
rect 43071 714141 43137 714142
rect 42879 714058 42945 714059
rect 42879 713994 42880 714058
rect 42944 713994 42945 714058
rect 42879 713993 42945 713994
rect 42111 713910 42177 713911
rect 42111 713846 42112 713910
rect 42176 713846 42177 713910
rect 42111 713845 42177 713846
rect 42114 711691 42174 713845
rect 42495 712282 42561 712283
rect 42495 712218 42496 712282
rect 42560 712218 42561 712282
rect 42495 712217 42561 712218
rect 42111 711690 42177 711691
rect 42111 711626 42112 711690
rect 42176 711626 42177 711690
rect 42111 711625 42177 711626
rect 42303 711542 42369 711543
rect 42303 711478 42304 711542
rect 42368 711478 42369 711542
rect 42303 711477 42369 711478
rect 42306 711099 42366 711477
rect 42303 711098 42369 711099
rect 42303 711034 42304 711098
rect 42368 711034 42369 711098
rect 42303 711033 42369 711034
rect 41919 708878 41985 708879
rect 41919 708814 41920 708878
rect 41984 708814 41985 708878
rect 41919 708813 41985 708814
rect 41727 707398 41793 707399
rect 41727 707334 41728 707398
rect 41792 707334 41793 707398
rect 41727 707333 41793 707334
rect 40575 705178 40641 705179
rect 40575 705114 40576 705178
rect 40640 705114 40641 705178
rect 40575 705113 40641 705114
rect 42498 704883 42558 712217
rect 42687 711690 42753 711691
rect 42687 711626 42688 711690
rect 42752 711626 42753 711690
rect 42687 711625 42753 711626
rect 42690 711247 42750 711625
rect 42687 711246 42753 711247
rect 42687 711182 42688 711246
rect 42752 711182 42753 711246
rect 42687 711181 42753 711182
rect 42882 707991 42942 713993
rect 42879 707990 42945 707991
rect 42879 707926 42880 707990
rect 42944 707926 42945 707990
rect 42879 707925 42945 707926
rect 42495 704882 42561 704883
rect 42495 704818 42496 704882
rect 42560 704818 42561 704882
rect 42495 704817 42561 704818
rect 43074 703551 43134 714141
rect 673986 707103 674046 783405
rect 674175 742474 674241 742475
rect 674175 742410 674176 742474
rect 674240 742410 674241 742474
rect 674175 742409 674241 742410
rect 673983 707102 674049 707103
rect 673983 707038 673984 707102
rect 674048 707038 674049 707102
rect 673983 707037 674049 707038
rect 43071 703550 43137 703551
rect 43071 703486 43072 703550
rect 43136 703486 43137 703550
rect 43071 703485 43137 703486
rect 40383 699998 40449 699999
rect 40383 699934 40384 699998
rect 40448 699934 40449 699998
rect 40383 699933 40449 699934
rect 40383 685494 40449 685495
rect 40383 685430 40384 685494
rect 40448 685430 40449 685494
rect 40383 685429 40449 685430
rect 40386 647049 40446 685429
rect 40575 684458 40641 684459
rect 40575 684394 40576 684458
rect 40640 684394 40641 684458
rect 40575 684393 40641 684394
rect 40578 679710 40638 684393
rect 40578 679650 40830 679710
rect 40575 672470 40641 672471
rect 40575 672406 40576 672470
rect 40640 672406 40641 672470
rect 40575 672405 40641 672406
rect 40578 660779 40638 672405
rect 40575 660778 40641 660779
rect 40575 660714 40576 660778
rect 40640 660714 40641 660778
rect 40575 660713 40641 660714
rect 40386 646989 40638 647049
rect 40578 642279 40638 646989
rect 40770 644795 40830 679650
rect 41151 671138 41217 671139
rect 41151 671074 41152 671138
rect 41216 671074 41217 671138
rect 41151 671073 41217 671074
rect 41154 662407 41214 671073
rect 42303 670694 42369 670695
rect 42303 670630 42304 670694
rect 42368 670630 42369 670694
rect 42303 670629 42369 670630
rect 42306 665071 42366 670629
rect 42303 665070 42369 665071
rect 42303 665006 42304 665070
rect 42368 665006 42369 665070
rect 42303 665005 42369 665006
rect 674178 663443 674238 742409
rect 674370 707695 674430 784145
rect 674559 740402 674625 740403
rect 674559 740338 674560 740402
rect 674624 740338 674625 740402
rect 674559 740337 674625 740338
rect 674367 707694 674433 707695
rect 674367 707630 674368 707694
rect 674432 707630 674433 707694
rect 674367 707629 674433 707630
rect 674367 697186 674433 697187
rect 674367 697122 674368 697186
rect 674432 697122 674433 697186
rect 674367 697121 674433 697122
rect 674175 663442 674241 663443
rect 674175 663378 674176 663442
rect 674240 663378 674241 663442
rect 674175 663377 674241 663378
rect 41151 662406 41217 662407
rect 41151 662342 41152 662406
rect 41216 662342 41217 662406
rect 41151 662341 41217 662342
rect 673983 652786 674049 652787
rect 673983 652722 673984 652786
rect 674048 652722 674049 652786
rect 673983 652721 674049 652722
rect 40767 644794 40833 644795
rect 40767 644730 40768 644794
rect 40832 644730 40833 644794
rect 40767 644729 40833 644730
rect 40383 642278 40449 642279
rect 40383 642214 40384 642278
rect 40448 642214 40449 642278
rect 40383 642213 40449 642214
rect 40575 642278 40641 642279
rect 40575 642214 40576 642278
rect 40640 642214 40641 642278
rect 40575 642213 40641 642214
rect 42879 642278 42945 642279
rect 42879 642214 42880 642278
rect 42944 642214 42945 642278
rect 42879 642213 42945 642214
rect 40386 601727 40446 642213
rect 40767 629254 40833 629255
rect 40767 629190 40768 629254
rect 40832 629190 40833 629254
rect 40767 629189 40833 629190
rect 40575 628366 40641 628367
rect 40575 628302 40576 628366
rect 40640 628302 40641 628366
rect 40575 628301 40641 628302
rect 40578 616527 40638 628301
rect 40575 616526 40641 616527
rect 40575 616462 40576 616526
rect 40640 616462 40641 616526
rect 40575 616461 40641 616462
rect 40770 616379 40830 629189
rect 41919 627478 41985 627479
rect 41919 627414 41920 627478
rect 41984 627414 41985 627478
rect 41919 627413 41985 627414
rect 42303 627478 42369 627479
rect 42303 627414 42304 627478
rect 42368 627414 42369 627478
rect 42303 627413 42369 627414
rect 41922 625259 41982 627413
rect 41919 625258 41985 625259
rect 41919 625194 41920 625258
rect 41984 625194 41985 625258
rect 41919 625193 41985 625194
rect 42306 622151 42366 627413
rect 42303 622150 42369 622151
rect 42303 622086 42304 622150
rect 42368 622086 42369 622150
rect 42303 622085 42369 622086
rect 40767 616378 40833 616379
rect 40767 616314 40768 616378
rect 40832 616314 40833 616378
rect 40767 616313 40833 616314
rect 40383 601726 40449 601727
rect 40383 601662 40384 601726
rect 40448 601662 40449 601726
rect 40383 601661 40449 601662
rect 40383 585742 40449 585743
rect 40383 585678 40384 585742
rect 40448 585678 40449 585742
rect 40383 585677 40449 585678
rect 40386 574051 40446 585677
rect 40575 585298 40641 585299
rect 40575 585234 40576 585298
rect 40640 585234 40641 585298
rect 40575 585233 40641 585234
rect 40578 575383 40638 585233
rect 42687 584854 42753 584855
rect 42687 584790 42688 584854
rect 42752 584790 42753 584854
rect 42687 584789 42753 584790
rect 41919 584262 41985 584263
rect 41919 584198 41920 584262
rect 41984 584198 41985 584262
rect 41919 584197 41985 584198
rect 42303 584262 42369 584263
rect 42303 584198 42304 584262
rect 42368 584198 42369 584262
rect 42303 584197 42369 584198
rect 40575 575382 40641 575383
rect 40575 575318 40576 575382
rect 40640 575318 40641 575382
rect 40575 575317 40641 575318
rect 40383 574050 40449 574051
rect 40383 573986 40384 574050
rect 40448 573986 40449 574050
rect 40383 573985 40449 573986
rect 41922 572719 41982 584197
rect 42306 578343 42366 584197
rect 42690 578787 42750 584789
rect 42687 578786 42753 578787
rect 42687 578722 42688 578786
rect 42752 578722 42753 578786
rect 42687 578721 42753 578722
rect 42303 578342 42369 578343
rect 42303 578278 42304 578342
rect 42368 578278 42369 578342
rect 42303 578277 42369 578278
rect 41919 572718 41985 572719
rect 41919 572654 41920 572718
rect 41984 572654 41985 572718
rect 41919 572653 41985 572654
rect 40383 539862 40449 539863
rect 40383 539798 40384 539862
rect 40448 539798 40449 539862
rect 40383 539797 40449 539798
rect 40386 469415 40446 539797
rect 41151 538086 41217 538087
rect 41151 538022 41152 538086
rect 41216 538022 41217 538086
rect 41151 538021 41217 538022
rect 40959 536310 41025 536311
rect 40959 536246 40960 536310
rect 41024 536246 41025 536310
rect 40959 536245 41025 536246
rect 40767 535126 40833 535127
rect 40767 535062 40768 535126
rect 40832 535062 40833 535126
rect 40767 535061 40833 535062
rect 40575 533942 40641 533943
rect 40575 533878 40576 533942
rect 40640 533878 40641 533942
rect 40575 533877 40641 533878
rect 40383 469414 40449 469415
rect 40383 469350 40384 469414
rect 40448 469350 40449 469414
rect 40383 469349 40449 469350
rect 40578 465863 40638 533877
rect 40575 465862 40641 465863
rect 40575 465798 40576 465862
rect 40640 465798 40641 465862
rect 40575 465797 40641 465798
rect 40770 465419 40830 535061
rect 40962 467343 41022 536245
rect 41154 471339 41214 538021
rect 42882 537051 42942 642213
rect 43071 627626 43137 627627
rect 43071 627562 43072 627626
rect 43136 627562 43137 627626
rect 43071 627561 43137 627562
rect 43074 619191 43134 627561
rect 43071 619190 43137 619191
rect 43071 619126 43072 619190
rect 43136 619126 43137 619190
rect 43071 619125 43137 619126
rect 43071 599506 43137 599507
rect 43071 599442 43072 599506
rect 43136 599442 43137 599506
rect 43071 599441 43137 599442
rect 42879 537050 42945 537051
rect 42879 536986 42880 537050
rect 42944 536986 42945 537050
rect 42879 536985 42945 536986
rect 41535 534238 41601 534239
rect 41535 534174 41536 534238
rect 41600 534174 41601 534238
rect 41535 534173 41601 534174
rect 41343 530834 41409 530835
rect 41343 530770 41344 530834
rect 41408 530770 41409 530834
rect 41343 530769 41409 530770
rect 41151 471338 41217 471339
rect 41151 471274 41152 471338
rect 41216 471274 41217 471338
rect 41151 471273 41217 471274
rect 40959 467342 41025 467343
rect 40959 467278 40960 467342
rect 41024 467278 41025 467342
rect 40959 467277 41025 467278
rect 41346 466307 41406 530769
rect 41538 466899 41598 534173
rect 41727 533202 41793 533203
rect 41727 533138 41728 533202
rect 41792 533138 41793 533202
rect 41727 533137 41793 533138
rect 41730 469563 41790 533137
rect 41919 530094 41985 530095
rect 41919 530030 41920 530094
rect 41984 530030 41985 530094
rect 41919 530029 41985 530030
rect 41727 469562 41793 469563
rect 41727 469498 41728 469562
rect 41792 469498 41793 469562
rect 41727 469497 41793 469498
rect 41922 467491 41982 530029
rect 42111 529354 42177 529355
rect 42111 529290 42112 529354
rect 42176 529290 42177 529354
rect 42111 529289 42177 529290
rect 42114 468083 42174 529289
rect 42303 528762 42369 528763
rect 42303 528698 42304 528762
rect 42368 528698 42369 528762
rect 42303 528697 42369 528698
rect 42306 470155 42366 528697
rect 42495 527134 42561 527135
rect 42495 527070 42496 527134
rect 42560 527070 42561 527134
rect 42495 527069 42561 527070
rect 42498 471635 42558 527069
rect 42495 471634 42561 471635
rect 42495 471570 42496 471634
rect 42560 471570 42561 471634
rect 42495 471569 42561 471570
rect 42303 470154 42369 470155
rect 42303 470090 42304 470154
rect 42368 470090 42369 470154
rect 42303 470089 42369 470090
rect 42111 468082 42177 468083
rect 42111 468018 42112 468082
rect 42176 468018 42177 468082
rect 42111 468017 42177 468018
rect 41919 467490 41985 467491
rect 41919 467426 41920 467490
rect 41984 467426 41985 467490
rect 41919 467425 41985 467426
rect 41535 466898 41601 466899
rect 41535 466834 41536 466898
rect 41600 466834 41601 466898
rect 41535 466833 41601 466834
rect 41343 466306 41409 466307
rect 41343 466242 41344 466306
rect 41408 466242 41409 466306
rect 41343 466241 41409 466242
rect 40767 465418 40833 465419
rect 40767 465354 40768 465418
rect 40832 465354 40833 465418
rect 40767 465353 40833 465354
rect 41535 422350 41601 422351
rect 41535 422286 41536 422350
rect 41600 422286 41601 422350
rect 41535 422285 41601 422286
rect 40383 421906 40449 421907
rect 40383 421842 40384 421906
rect 40448 421842 40449 421906
rect 40383 421841 40449 421842
rect 40386 411251 40446 421841
rect 40575 421314 40641 421315
rect 40575 421250 40576 421314
rect 40640 421250 40641 421314
rect 40575 421249 40641 421250
rect 40383 411250 40449 411251
rect 40383 411186 40384 411250
rect 40448 411186 40449 411250
rect 40383 411185 40449 411186
rect 40578 398819 40638 421249
rect 40959 417762 41025 417763
rect 40959 417698 40960 417762
rect 41024 417698 41025 417762
rect 40959 417697 41025 417698
rect 40962 407699 41022 417697
rect 41151 416430 41217 416431
rect 41151 416366 41152 416430
rect 41216 416366 41217 416430
rect 41151 416365 41217 416366
rect 40959 407698 41025 407699
rect 40959 407634 40960 407698
rect 41024 407634 41025 407698
rect 40959 407633 41025 407634
rect 41154 399411 41214 416365
rect 41343 414950 41409 414951
rect 41343 414886 41344 414950
rect 41408 414886 41409 414950
rect 41343 414885 41409 414886
rect 41346 401927 41406 414885
rect 41343 401926 41409 401927
rect 41343 401862 41344 401926
rect 41408 401862 41409 401926
rect 41343 401861 41409 401862
rect 41538 400151 41598 422285
rect 42495 421758 42561 421759
rect 42495 421694 42496 421758
rect 42560 421694 42561 421758
rect 42495 421693 42561 421694
rect 41919 417318 41985 417319
rect 41919 417254 41920 417318
rect 41984 417254 41985 417318
rect 41919 417253 41985 417254
rect 41727 417022 41793 417023
rect 41727 416958 41728 417022
rect 41792 416958 41793 417022
rect 41727 416957 41793 416958
rect 41730 403851 41790 416957
rect 41727 403850 41793 403851
rect 41727 403786 41728 403850
rect 41792 403786 41793 403850
rect 41727 403785 41793 403786
rect 41922 402667 41982 417253
rect 42111 416874 42177 416875
rect 42111 416810 42112 416874
rect 42176 416810 42177 416874
rect 42111 416809 42177 416810
rect 42114 406071 42174 416809
rect 42303 416282 42369 416283
rect 42303 416218 42304 416282
rect 42368 416218 42369 416282
rect 42303 416217 42369 416218
rect 42111 406070 42177 406071
rect 42111 406006 42112 406070
rect 42176 406006 42177 406070
rect 42111 406005 42177 406006
rect 42306 403111 42366 416217
rect 42303 403110 42369 403111
rect 42303 403046 42304 403110
rect 42368 403046 42369 403110
rect 42303 403045 42369 403046
rect 41919 402666 41985 402667
rect 41919 402602 41920 402666
rect 41984 402602 41985 402666
rect 41919 402601 41985 402602
rect 41535 400150 41601 400151
rect 41535 400086 41536 400150
rect 41600 400086 41601 400150
rect 41535 400085 41601 400086
rect 41151 399410 41217 399411
rect 41151 399346 41152 399410
rect 41216 399346 41217 399410
rect 41151 399345 41217 399346
rect 40575 398818 40641 398819
rect 40575 398754 40576 398818
rect 40640 398754 40641 398818
rect 40575 398753 40641 398754
rect 42498 388755 42558 421693
rect 42495 388754 42561 388755
rect 42495 388690 42496 388754
rect 42560 388690 42561 388754
rect 42495 388689 42561 388690
rect 39807 380318 39873 380319
rect 39807 380254 39808 380318
rect 39872 380254 39873 380318
rect 39807 380253 39873 380254
rect 39810 372475 39870 380253
rect 40575 379874 40641 379875
rect 40575 379810 40576 379874
rect 40640 379810 40641 379874
rect 40575 379809 40641 379810
rect 39999 379282 40065 379283
rect 39999 379218 40000 379282
rect 40064 379218 40065 379282
rect 39999 379217 40065 379218
rect 40002 374655 40062 379217
rect 40002 374595 40446 374655
rect 39807 372474 39873 372475
rect 39807 372410 39808 372474
rect 39872 372410 39873 372474
rect 39807 372409 39873 372410
rect 40386 362855 40446 374595
rect 40383 362854 40449 362855
rect 40383 362790 40384 362854
rect 40448 362790 40449 362854
rect 40383 362789 40449 362790
rect 40578 358859 40638 379809
rect 42303 378838 42369 378839
rect 42303 378774 42304 378838
rect 42368 378774 42369 378838
rect 42303 378773 42369 378774
rect 41343 375878 41409 375879
rect 41343 375814 41344 375878
rect 41408 375814 41409 375878
rect 41343 375813 41409 375814
rect 40959 373954 41025 373955
rect 40959 373890 40960 373954
rect 41024 373890 41025 373954
rect 40959 373889 41025 373890
rect 40767 372326 40833 372327
rect 40767 372262 40768 372326
rect 40832 372262 40833 372326
rect 40767 372261 40833 372262
rect 40575 358858 40641 358859
rect 40575 358794 40576 358858
rect 40640 358794 40641 358858
rect 40575 358793 40641 358794
rect 40770 357231 40830 372261
rect 40767 357230 40833 357231
rect 40767 357166 40768 357230
rect 40832 357166 40833 357230
rect 40767 357165 40833 357166
rect 40962 356195 41022 373889
rect 41346 360635 41406 375813
rect 41727 373806 41793 373807
rect 41727 373742 41728 373806
rect 41792 373742 41793 373806
rect 41727 373741 41793 373742
rect 41730 368183 41790 373741
rect 41919 373362 41985 373363
rect 41919 373298 41920 373362
rect 41984 373298 41985 373362
rect 41919 373297 41985 373298
rect 41727 368182 41793 368183
rect 41727 368118 41728 368182
rect 41792 368118 41793 368182
rect 41727 368117 41793 368118
rect 41343 360634 41409 360635
rect 41343 360570 41344 360634
rect 41408 360570 41409 360634
rect 41343 360569 41409 360570
rect 41922 359895 41982 373297
rect 42111 373214 42177 373215
rect 42111 373150 42112 373214
rect 42176 373150 42177 373214
rect 42111 373149 42177 373150
rect 41919 359894 41985 359895
rect 41919 359830 41920 359894
rect 41984 359830 41985 359894
rect 41919 359829 41985 359830
rect 42114 359303 42174 373149
rect 42111 359302 42177 359303
rect 42111 359238 42112 359302
rect 42176 359238 42177 359302
rect 42111 359237 42177 359238
rect 42306 358671 42366 378773
rect 42495 372474 42561 372475
rect 42495 372410 42496 372474
rect 42560 372410 42561 372474
rect 42495 372409 42561 372410
rect 41730 358611 42366 358671
rect 40959 356194 41025 356195
rect 40959 356130 40960 356194
rect 41024 356130 41025 356194
rect 40959 356129 41025 356130
rect 41730 343171 41790 358611
rect 41919 357230 41985 357231
rect 41919 357166 41920 357230
rect 41984 357166 41985 357230
rect 41919 357165 41985 357166
rect 41922 356935 41982 357165
rect 41919 356934 41985 356935
rect 41919 356870 41920 356934
rect 41984 356870 41985 356934
rect 41919 356869 41985 356870
rect 42498 355603 42558 372409
rect 42495 355602 42561 355603
rect 42495 355538 42496 355602
rect 42560 355538 42561 355602
rect 42495 355537 42561 355538
rect 41727 343170 41793 343171
rect 41727 343106 41728 343170
rect 41792 343106 41793 343170
rect 41727 343105 41793 343106
rect 41919 338878 41985 338879
rect 41919 338814 41920 338878
rect 41984 338814 41985 338878
rect 41919 338813 41985 338814
rect 40383 336658 40449 336659
rect 40383 336594 40384 336658
rect 40448 336594 40449 336658
rect 40383 336593 40449 336594
rect 40386 315495 40446 336593
rect 40767 336066 40833 336067
rect 40767 336002 40768 336066
rect 40832 336002 40833 336066
rect 40767 336001 40833 336002
rect 40575 332070 40641 332071
rect 40575 332006 40576 332070
rect 40640 332006 40641 332070
rect 40575 332005 40641 332006
rect 40578 320527 40638 332005
rect 40575 320526 40641 320527
rect 40575 320462 40576 320526
rect 40640 320462 40641 320526
rect 40575 320461 40641 320462
rect 40770 319787 40830 336001
rect 40959 335178 41025 335179
rect 40959 335114 40960 335178
rect 41024 335114 41025 335178
rect 40959 335113 41025 335114
rect 40767 319786 40833 319787
rect 40767 319722 40768 319786
rect 40832 319722 40833 319786
rect 40767 319721 40833 319722
rect 40383 315494 40449 315495
rect 40383 315430 40384 315494
rect 40448 315430 40449 315494
rect 40383 315429 40449 315430
rect 40962 313127 41022 335113
rect 41343 334586 41409 334587
rect 41343 334522 41344 334586
rect 41408 334522 41409 334586
rect 41343 334521 41409 334522
rect 41151 334142 41217 334143
rect 41151 334078 41152 334142
rect 41216 334078 41217 334142
rect 41151 334077 41217 334078
rect 41154 316679 41214 334077
rect 41151 316678 41217 316679
rect 41151 316614 41152 316678
rect 41216 316614 41217 316678
rect 41151 316613 41217 316614
rect 41346 316235 41406 334521
rect 41535 332662 41601 332663
rect 41535 332598 41536 332662
rect 41600 332598 41601 332662
rect 41535 332597 41601 332598
rect 41538 317419 41598 332597
rect 41727 331182 41793 331183
rect 41727 331118 41728 331182
rect 41792 331118 41793 331182
rect 41727 331117 41793 331118
rect 41730 324967 41790 331117
rect 41727 324966 41793 324967
rect 41727 324902 41728 324966
rect 41792 324902 41793 324966
rect 41727 324901 41793 324902
rect 41535 317418 41601 317419
rect 41535 317354 41536 317418
rect 41600 317354 41601 317418
rect 41535 317353 41601 317354
rect 41343 316234 41409 316235
rect 41343 316170 41344 316234
rect 41408 316170 41409 316234
rect 41343 316169 41409 316170
rect 40959 313126 41025 313127
rect 40959 313062 40960 313126
rect 41024 313062 41025 313126
rect 40959 313061 41025 313062
rect 41922 308190 41982 338813
rect 42303 330738 42369 330739
rect 42303 330674 42304 330738
rect 42368 330674 42369 330738
rect 42303 330673 42369 330674
rect 42111 329110 42177 329111
rect 42111 329046 42112 329110
rect 42176 329046 42177 329110
rect 42111 329045 42177 329046
rect 42114 313719 42174 329045
rect 42111 313718 42177 313719
rect 42111 313654 42112 313718
rect 42176 313654 42177 313718
rect 42111 313653 42177 313654
rect 42306 312535 42366 330673
rect 42303 312534 42369 312535
rect 42303 312470 42304 312534
rect 42368 312470 42369 312534
rect 42303 312469 42369 312470
rect 41730 308130 41982 308190
rect 41730 296670 41790 308130
rect 41730 296610 42366 296670
rect 41727 294626 41793 294627
rect 41727 294562 41728 294626
rect 41792 294562 41793 294626
rect 41727 294561 41793 294562
rect 41151 293442 41217 293443
rect 41151 293378 41152 293442
rect 41216 293378 41217 293442
rect 41151 293377 41217 293378
rect 40383 291962 40449 291963
rect 40383 291898 40384 291962
rect 40448 291898 40449 291962
rect 40383 291897 40449 291898
rect 40386 270059 40446 291897
rect 40959 291518 41025 291519
rect 40959 291454 40960 291518
rect 41024 291454 41025 291518
rect 40959 291453 41025 291454
rect 40575 289446 40641 289447
rect 40575 289382 40576 289446
rect 40640 289382 40641 289446
rect 40575 289381 40641 289382
rect 40578 274203 40638 289381
rect 40575 274202 40641 274203
rect 40575 274138 40576 274202
rect 40640 274138 40641 274202
rect 40575 274137 40641 274138
rect 40962 272871 41022 291453
rect 40959 272870 41025 272871
rect 40959 272806 40960 272870
rect 41024 272806 41025 272870
rect 40959 272805 41025 272806
rect 41154 272427 41214 293377
rect 41535 292998 41601 292999
rect 41535 292934 41536 292998
rect 41600 292934 41601 292998
rect 41535 292933 41601 292934
rect 41343 290926 41409 290927
rect 41343 290862 41344 290926
rect 41408 290862 41409 290926
rect 41343 290861 41409 290862
rect 41346 273611 41406 290861
rect 41538 276571 41598 292933
rect 41730 281751 41790 294561
rect 41919 294182 41985 294183
rect 41919 294118 41920 294182
rect 41984 294118 41985 294182
rect 41919 294117 41985 294118
rect 41727 281750 41793 281751
rect 41727 281686 41728 281750
rect 41792 281686 41793 281750
rect 41727 281685 41793 281686
rect 41535 276570 41601 276571
rect 41535 276506 41536 276570
rect 41600 276506 41601 276570
rect 41535 276505 41601 276506
rect 41343 273610 41409 273611
rect 41343 273546 41344 273610
rect 41408 273546 41409 273610
rect 41343 273545 41409 273546
rect 41151 272426 41217 272427
rect 41151 272362 41152 272426
rect 41216 272362 41217 272426
rect 41151 272361 41217 272362
rect 40383 270058 40449 270059
rect 40383 269994 40384 270058
rect 40448 269994 40449 270058
rect 40383 269993 40449 269994
rect 41922 269319 41982 294117
rect 42111 285154 42177 285155
rect 42111 285090 42112 285154
rect 42176 285090 42177 285154
rect 42111 285089 42177 285090
rect 42114 270651 42174 285089
rect 42306 278643 42366 296610
rect 42495 281602 42561 281603
rect 42495 281538 42496 281602
rect 42560 281538 42561 281602
rect 42495 281537 42561 281538
rect 42303 278642 42369 278643
rect 42303 278578 42304 278642
rect 42368 278578 42369 278642
rect 42303 278577 42369 278578
rect 42498 278051 42558 281537
rect 43074 278495 43134 599441
rect 673986 572867 674046 652721
rect 674175 652194 674241 652195
rect 674175 652130 674176 652194
rect 674240 652130 674241 652194
rect 674175 652129 674241 652130
rect 673983 572866 674049 572867
rect 673983 572802 673984 572866
rect 674048 572802 674049 572866
rect 673983 572801 674049 572802
rect 674178 571239 674238 652129
rect 674370 618007 674430 697121
rect 674562 664775 674622 740337
rect 674754 710507 674814 787993
rect 676095 787466 676161 787467
rect 676095 787402 676096 787466
rect 676160 787402 676161 787466
rect 676095 787401 676161 787402
rect 675519 786726 675585 786727
rect 675519 786662 675520 786726
rect 675584 786662 675585 786726
rect 675519 786661 675585 786662
rect 675135 784802 675201 784803
rect 675135 784738 675136 784802
rect 675200 784738 675201 784802
rect 675135 784737 675201 784738
rect 674943 741142 675009 741143
rect 674943 741078 674944 741142
rect 675008 741078 675009 741142
rect 674943 741077 675009 741078
rect 674751 710506 674817 710507
rect 674751 710442 674752 710506
rect 674816 710442 674817 710506
rect 674751 710441 674817 710442
rect 674751 697038 674817 697039
rect 674751 696974 674752 697038
rect 674816 696974 674817 697038
rect 674751 696973 674817 696974
rect 674559 664774 674625 664775
rect 674559 664710 674560 664774
rect 674624 664710 674625 664774
rect 674559 664709 674625 664710
rect 674559 649678 674625 649679
rect 674559 649614 674560 649678
rect 674624 649614 674625 649678
rect 674559 649613 674625 649614
rect 674367 618006 674433 618007
rect 674367 617942 674368 618006
rect 674432 617942 674433 618006
rect 674367 617941 674433 617942
rect 674367 607794 674433 607795
rect 674367 607730 674368 607794
rect 674432 607730 674433 607794
rect 674367 607729 674433 607730
rect 674175 571238 674241 571239
rect 674175 571174 674176 571238
rect 674240 571174 674241 571238
rect 674175 571173 674241 571174
rect 674175 561766 674241 561767
rect 674175 561702 674176 561766
rect 674240 561702 674241 561766
rect 674175 561701 674241 561702
rect 674178 483475 674238 561701
rect 674370 529947 674430 607729
rect 674562 572571 674622 649613
rect 674754 620967 674814 696973
rect 674946 666255 675006 741077
rect 675138 709767 675198 784737
rect 675327 777698 675393 777699
rect 675327 777634 675328 777698
rect 675392 777634 675393 777698
rect 675327 777633 675393 777634
rect 675135 709766 675201 709767
rect 675135 709702 675136 709766
rect 675200 709702 675201 709766
rect 675135 709701 675201 709702
rect 675330 706955 675390 777633
rect 675522 771927 675582 786661
rect 675711 780658 675777 780659
rect 675711 780594 675712 780658
rect 675776 780594 675777 780658
rect 675711 780593 675777 780594
rect 675519 771926 675585 771927
rect 675519 771862 675520 771926
rect 675584 771862 675585 771926
rect 675519 771861 675585 771862
rect 675519 739218 675585 739219
rect 675519 739154 675520 739218
rect 675584 739154 675585 739218
rect 675519 739153 675585 739154
rect 675327 706954 675393 706955
rect 675327 706890 675328 706954
rect 675392 706890 675393 706954
rect 675327 706889 675393 706890
rect 675135 697926 675201 697927
rect 675135 697862 675136 697926
rect 675200 697862 675201 697926
rect 675135 697861 675201 697862
rect 674943 666254 675009 666255
rect 674943 666190 674944 666254
rect 675008 666190 675009 666254
rect 674943 666189 675009 666190
rect 674943 651454 675009 651455
rect 674943 651390 674944 651454
rect 675008 651390 675009 651454
rect 674943 651389 675009 651390
rect 674751 620966 674817 620967
rect 674751 620902 674752 620966
rect 674816 620902 674817 620966
rect 674751 620901 674817 620902
rect 674751 604834 674817 604835
rect 674751 604770 674752 604834
rect 674816 604770 674817 604834
rect 674751 604769 674817 604770
rect 674559 572570 674625 572571
rect 674559 572506 674560 572570
rect 674624 572506 674625 572570
rect 674559 572505 674625 572506
rect 674559 558954 674625 558955
rect 674559 558890 674560 558954
rect 674624 558890 674625 558954
rect 674559 558889 674625 558890
rect 674367 529946 674433 529947
rect 674367 529882 674368 529946
rect 674432 529882 674433 529946
rect 674367 529881 674433 529882
rect 674175 483474 674241 483475
rect 674175 483410 674176 483474
rect 674240 483410 674241 483474
rect 674175 483409 674241 483410
rect 674562 482883 674622 558889
rect 674754 529355 674814 604769
rect 674946 574051 675006 651389
rect 675138 619931 675198 697861
rect 675327 694670 675393 694671
rect 675327 694606 675328 694670
rect 675392 694606 675393 694670
rect 675327 694605 675393 694606
rect 675135 619930 675201 619931
rect 675135 619866 675136 619930
rect 675200 619866 675201 619930
rect 675135 619865 675201 619866
rect 675330 617859 675390 694605
rect 675522 662703 675582 739153
rect 675714 709175 675774 780593
rect 675903 775478 675969 775479
rect 675903 775414 675904 775478
rect 675968 775414 675969 775478
rect 675903 775413 675969 775414
rect 675906 710655 675966 775413
rect 676098 772075 676158 787401
rect 676479 783026 676545 783027
rect 676479 782962 676480 783026
rect 676544 782962 676545 783026
rect 676479 782961 676545 782962
rect 676287 779918 676353 779919
rect 676287 779854 676288 779918
rect 676352 779854 676353 779918
rect 676287 779853 676353 779854
rect 676095 772074 676161 772075
rect 676095 772010 676096 772074
rect 676160 772010 676161 772074
rect 676095 772009 676161 772010
rect 676290 745879 676350 779853
rect 676287 745878 676353 745879
rect 676287 745814 676288 745878
rect 676352 745814 676353 745878
rect 676287 745813 676353 745814
rect 676482 743067 676542 782961
rect 676671 779178 676737 779179
rect 676671 779114 676672 779178
rect 676736 779114 676737 779178
rect 676671 779113 676737 779114
rect 676479 743066 676545 743067
rect 676479 743002 676480 743066
rect 676544 743002 676545 743066
rect 676479 743001 676545 743002
rect 676287 735518 676353 735519
rect 676287 735454 676288 735518
rect 676352 735454 676353 735518
rect 676287 735453 676353 735454
rect 676095 730634 676161 730635
rect 676095 730570 676096 730634
rect 676160 730570 676161 730634
rect 676095 730569 676161 730570
rect 675903 710654 675969 710655
rect 675903 710590 675904 710654
rect 675968 710590 675969 710654
rect 675903 710589 675969 710590
rect 675711 709174 675777 709175
rect 675711 709110 675712 709174
rect 675776 709110 675777 709174
rect 675711 709109 675777 709110
rect 675711 694966 675777 694967
rect 675711 694902 675712 694966
rect 675776 694902 675777 694966
rect 675711 694901 675777 694902
rect 675519 662702 675585 662703
rect 675519 662638 675520 662702
rect 675584 662638 675585 662702
rect 675519 662637 675585 662638
rect 675519 645386 675585 645387
rect 675519 645322 675520 645386
rect 675584 645322 675585 645386
rect 675519 645321 675585 645322
rect 675327 617858 675393 617859
rect 675327 617794 675328 617858
rect 675392 617794 675393 617858
rect 675327 617793 675393 617794
rect 675135 606018 675201 606019
rect 675135 605954 675136 606018
rect 675200 605954 675201 606018
rect 675135 605953 675201 605954
rect 674943 574050 675009 574051
rect 674943 573986 674944 574050
rect 675008 573986 675009 574050
rect 674943 573985 675009 573986
rect 674943 561470 675009 561471
rect 674943 561406 674944 561470
rect 675008 561406 675009 561470
rect 674943 561405 675009 561406
rect 674751 529354 674817 529355
rect 674751 529290 674752 529354
rect 674816 529290 674817 529354
rect 674751 529289 674817 529290
rect 674946 486435 675006 561405
rect 675138 530835 675198 605953
rect 675327 600246 675393 600247
rect 675327 600182 675328 600246
rect 675392 600182 675393 600246
rect 675327 600181 675393 600182
rect 675135 530834 675201 530835
rect 675135 530770 675136 530834
rect 675200 530770 675201 530834
rect 675135 530769 675201 530770
rect 675330 528763 675390 600181
rect 675522 571979 675582 645321
rect 675714 619487 675774 694901
rect 676098 664923 676158 730569
rect 676095 664922 676161 664923
rect 676095 664858 676096 664922
rect 676160 664858 676161 664922
rect 676095 664857 676161 664858
rect 676290 664479 676350 735453
rect 676674 728119 676734 779113
rect 677247 745878 677313 745879
rect 677247 745814 677248 745878
rect 677312 745814 677313 745878
rect 677247 745813 677313 745814
rect 676863 743066 676929 743067
rect 676863 743002 676864 743066
rect 676928 743002 676929 743066
rect 676863 743001 676929 743002
rect 676866 729895 676926 743001
rect 676863 729894 676929 729895
rect 676863 729830 676864 729894
rect 676928 729830 676929 729894
rect 676863 729829 676929 729830
rect 677250 729633 677310 745813
rect 676866 729573 677310 729633
rect 676671 728118 676737 728119
rect 676671 728054 676672 728118
rect 676736 728054 676737 728118
rect 676671 728053 676737 728054
rect 676866 705475 676926 729573
rect 677055 729450 677121 729451
rect 677055 729386 677056 729450
rect 677120 729386 677121 729450
rect 677055 729385 677121 729386
rect 677058 705919 677118 729385
rect 677247 728118 677313 728119
rect 677247 728054 677248 728118
rect 677312 728054 677313 728118
rect 677247 728053 677313 728054
rect 677250 706511 677310 728053
rect 677247 706510 677313 706511
rect 677247 706446 677248 706510
rect 677312 706446 677313 706510
rect 677247 706445 677313 706446
rect 677055 705918 677121 705919
rect 677055 705854 677056 705918
rect 677120 705854 677121 705918
rect 677055 705853 677121 705854
rect 676863 705474 676929 705475
rect 676863 705410 676864 705474
rect 676928 705410 676929 705474
rect 676863 705409 676929 705410
rect 676287 664478 676353 664479
rect 676287 664414 676288 664478
rect 676352 664414 676353 664478
rect 676287 664413 676353 664414
rect 676095 640354 676161 640355
rect 676095 640290 676096 640354
rect 676160 640290 676161 640354
rect 676095 640289 676161 640290
rect 675903 638578 675969 638579
rect 675903 638514 675904 638578
rect 675968 638514 675969 638578
rect 675903 638513 675969 638514
rect 675711 619486 675777 619487
rect 675711 619422 675712 619486
rect 675776 619422 675777 619486
rect 675711 619421 675777 619422
rect 675711 593438 675777 593439
rect 675711 593374 675712 593438
rect 675776 593374 675777 593438
rect 675711 593373 675777 593374
rect 675519 571978 675585 571979
rect 675519 571914 675520 571978
rect 675584 571914 675585 571978
rect 675519 571913 675585 571914
rect 675519 562506 675585 562507
rect 675519 562442 675520 562506
rect 675584 562442 675585 562506
rect 675519 562441 675585 562442
rect 675327 528762 675393 528763
rect 675327 528698 675328 528762
rect 675392 528698 675393 528762
rect 675327 528697 675393 528698
rect 674943 486434 675009 486435
rect 674943 486370 674944 486434
rect 675008 486370 675009 486434
rect 674943 486369 675009 486370
rect 675522 485695 675582 562441
rect 675714 528171 675774 593373
rect 675906 571387 675966 638513
rect 676098 573755 676158 640289
rect 676287 595362 676353 595363
rect 676287 595298 676288 595362
rect 676352 595298 676353 595362
rect 676287 595297 676353 595298
rect 676095 573754 676161 573755
rect 676095 573690 676096 573754
rect 676160 573690 676161 573754
rect 676095 573689 676161 573690
rect 675903 571386 675969 571387
rect 675903 571322 675904 571386
rect 675968 571322 675969 571386
rect 675903 571321 675969 571322
rect 676290 530539 676350 595297
rect 676287 530538 676353 530539
rect 676287 530474 676288 530538
rect 676352 530474 676353 530538
rect 676287 530473 676353 530474
rect 675711 528170 675777 528171
rect 675711 528106 675712 528170
rect 675776 528106 675777 528170
rect 675711 528105 675777 528106
rect 675519 485694 675585 485695
rect 675519 485630 675520 485694
rect 675584 485630 675585 485694
rect 675519 485629 675585 485630
rect 674559 482882 674625 482883
rect 674559 482818 674560 482882
rect 674624 482818 674625 482882
rect 674559 482817 674625 482818
rect 676671 397930 676737 397931
rect 676671 397866 676672 397930
rect 676736 397866 676737 397930
rect 676671 397865 676737 397866
rect 673983 397634 674049 397635
rect 673983 397570 673984 397634
rect 674048 397570 674049 397634
rect 673983 397569 674049 397570
rect 673986 373955 674046 397569
rect 676674 397470 676734 397865
rect 674946 397410 676734 397470
rect 674751 396154 674817 396155
rect 674751 396090 674752 396154
rect 674816 396090 674817 396154
rect 674751 396089 674817 396090
rect 674367 393194 674433 393195
rect 674367 393130 674368 393194
rect 674432 393130 674433 393194
rect 674367 393129 674433 393130
rect 674370 377211 674430 393129
rect 674754 378839 674814 396089
rect 674946 384463 675006 397410
rect 675135 396894 675201 396895
rect 675135 396830 675136 396894
rect 675200 396830 675201 396894
rect 675135 396829 675201 396830
rect 675138 385943 675198 396829
rect 676671 396450 676737 396451
rect 676671 396386 676672 396450
rect 676736 396386 676737 396450
rect 676671 396385 676737 396386
rect 675903 395266 675969 395267
rect 675903 395202 675904 395266
rect 675968 395202 675969 395266
rect 675903 395201 675969 395202
rect 675327 394674 675393 394675
rect 675327 394610 675328 394674
rect 675392 394610 675393 394674
rect 675327 394609 675393 394610
rect 675135 385942 675201 385943
rect 675135 385878 675136 385942
rect 675200 385878 675201 385942
rect 675135 385877 675201 385878
rect 674943 384462 675009 384463
rect 674943 384398 674944 384462
rect 675008 384398 675009 384462
rect 674943 384397 675009 384398
rect 675330 382391 675390 394609
rect 675711 392602 675777 392603
rect 675711 392538 675712 392602
rect 675776 392538 675777 392602
rect 675711 392537 675777 392538
rect 675519 391862 675585 391863
rect 675519 391798 675520 391862
rect 675584 391798 675585 391862
rect 675519 391797 675585 391798
rect 675327 382390 675393 382391
rect 675327 382326 675328 382390
rect 675392 382326 675393 382390
rect 675327 382325 675393 382326
rect 674751 378838 674817 378839
rect 674751 378774 674752 378838
rect 674816 378774 674817 378838
rect 674751 378773 674817 378774
rect 675522 378099 675582 391797
rect 675714 381207 675774 392537
rect 675906 385647 675966 395201
rect 676479 393934 676545 393935
rect 676479 393870 676480 393934
rect 676544 393870 676545 393934
rect 676479 393869 676545 393870
rect 676095 393342 676161 393343
rect 676095 393278 676096 393342
rect 676160 393278 676161 393342
rect 676095 393277 676161 393278
rect 675903 385646 675969 385647
rect 675903 385582 675904 385646
rect 675968 385582 675969 385646
rect 675903 385581 675969 385582
rect 675711 381206 675777 381207
rect 675711 381142 675712 381206
rect 675776 381142 675777 381206
rect 675711 381141 675777 381142
rect 675519 378098 675585 378099
rect 675519 378034 675520 378098
rect 675584 378034 675585 378098
rect 675519 378033 675585 378034
rect 674367 377210 674433 377211
rect 674367 377146 674368 377210
rect 674432 377146 674433 377210
rect 674367 377145 674433 377146
rect 676098 375731 676158 393277
rect 676287 391418 676353 391419
rect 676287 391354 676288 391418
rect 676352 391354 676353 391418
rect 676287 391353 676353 391354
rect 676290 376767 676350 391353
rect 676482 381799 676542 393869
rect 676674 382983 676734 396385
rect 676671 382982 676737 382983
rect 676671 382918 676672 382982
rect 676736 382918 676737 382982
rect 676671 382917 676737 382918
rect 676479 381798 676545 381799
rect 676479 381734 676480 381798
rect 676544 381734 676545 381798
rect 676479 381733 676545 381734
rect 676287 376766 676353 376767
rect 676287 376702 676288 376766
rect 676352 376702 676353 376766
rect 676287 376701 676353 376702
rect 676095 375730 676161 375731
rect 676095 375666 676096 375730
rect 676160 375666 676161 375730
rect 676095 375665 676161 375666
rect 673983 373954 674049 373955
rect 673983 373890 673984 373954
rect 674048 373890 674049 373954
rect 673983 373889 674049 373890
rect 674175 355898 674241 355899
rect 674175 355834 674176 355898
rect 674240 355834 674241 355898
rect 674175 355833 674241 355834
rect 673983 355306 674049 355307
rect 673983 355242 673984 355306
rect 674048 355242 674049 355306
rect 673983 355241 674049 355242
rect 673986 310053 674046 355241
rect 674178 311055 674238 355833
rect 674367 354270 674433 354271
rect 674367 354206 674368 354270
rect 674432 354206 674433 354270
rect 674367 354205 674433 354206
rect 674175 311054 674241 311055
rect 674175 310990 674176 311054
rect 674240 310990 674241 311054
rect 674175 310989 674241 310990
rect 673986 309993 674238 310053
rect 674178 309871 674238 309993
rect 674175 309870 674241 309871
rect 674175 309806 674176 309870
rect 674240 309806 674241 309870
rect 674175 309805 674241 309806
rect 673983 302618 674049 302619
rect 673983 302554 673984 302618
rect 674048 302554 674049 302618
rect 673983 302553 674049 302554
rect 673986 287227 674046 302553
rect 673983 287226 674049 287227
rect 673983 287162 673984 287226
rect 674048 287162 674049 287226
rect 673983 287161 674049 287162
rect 674178 278495 674238 309805
rect 674370 308983 674430 354205
rect 675903 353826 675969 353827
rect 675903 353762 675904 353826
rect 675968 353762 675969 353826
rect 675903 353761 675969 353762
rect 674559 353234 674625 353235
rect 674559 353170 674560 353234
rect 674624 353170 674625 353234
rect 674559 353169 674625 353170
rect 674562 328371 674622 353169
rect 674751 351754 674817 351755
rect 674751 351690 674752 351754
rect 674816 351690 674817 351754
rect 674751 351689 674817 351690
rect 674754 333551 674814 351689
rect 674943 348794 675009 348795
rect 674943 348730 674944 348794
rect 675008 348730 675009 348794
rect 674943 348729 675009 348730
rect 674751 333550 674817 333551
rect 674751 333486 674752 333550
rect 674816 333486 674817 333550
rect 674751 333485 674817 333486
rect 674946 332367 675006 348729
rect 675711 343022 675777 343023
rect 675711 342958 675712 343022
rect 675776 342958 675777 343022
rect 675711 342957 675777 342958
rect 674943 332366 675009 332367
rect 674943 332302 674944 332366
rect 675008 332302 675009 332366
rect 674943 332301 675009 332302
rect 675714 330591 675774 342957
rect 675906 339619 675966 353761
rect 676671 342874 676737 342875
rect 676671 342810 676672 342874
rect 676736 342810 676737 342874
rect 676671 342809 676737 342810
rect 675903 339618 675969 339619
rect 675903 339554 675904 339618
rect 675968 339554 675969 339618
rect 675903 339553 675969 339554
rect 675711 330590 675777 330591
rect 675711 330526 675712 330590
rect 675776 330526 675777 330590
rect 675711 330525 675777 330526
rect 674559 328370 674625 328371
rect 674559 328306 674560 328370
rect 674624 328306 674625 328370
rect 674559 328305 674625 328306
rect 676674 326891 676734 342809
rect 676671 326890 676737 326891
rect 676671 326826 676672 326890
rect 676736 326826 676737 326890
rect 676671 326825 676737 326826
rect 675519 310462 675585 310463
rect 675519 310398 675520 310462
rect 675584 310398 675585 310462
rect 675519 310397 675585 310398
rect 674559 309130 674625 309131
rect 674559 309066 674560 309130
rect 674624 309066 674625 309130
rect 674559 309065 674625 309066
rect 674367 308982 674433 308983
rect 674367 308918 674368 308982
rect 674432 308918 674433 308982
rect 674367 308917 674433 308918
rect 43071 278494 43137 278495
rect 43071 278430 43072 278494
rect 43136 278430 43137 278494
rect 43071 278429 43137 278430
rect 674175 278494 674241 278495
rect 674175 278430 674176 278494
rect 674240 278430 674241 278494
rect 674175 278429 674241 278430
rect 42495 278050 42561 278051
rect 42495 277986 42496 278050
rect 42560 277986 42561 278050
rect 42495 277985 42561 277986
rect 674370 274203 674430 308917
rect 674562 276571 674622 309065
rect 674751 308390 674817 308391
rect 674751 308326 674752 308390
rect 674816 308326 674817 308390
rect 674751 308325 674817 308326
rect 674754 278199 674814 308325
rect 675327 306022 675393 306023
rect 675327 305958 675328 306022
rect 675392 305958 675393 306022
rect 675327 305957 675393 305958
rect 674943 305430 675009 305431
rect 674943 305366 674944 305430
rect 675008 305366 675009 305430
rect 674943 305365 675009 305366
rect 674946 281899 675006 305365
rect 675135 303506 675201 303507
rect 675135 303442 675136 303506
rect 675200 303442 675201 303506
rect 675135 303441 675201 303442
rect 675138 285303 675198 303441
rect 675330 288559 675390 305957
rect 675327 288558 675393 288559
rect 675327 288494 675328 288558
rect 675392 288494 675393 288558
rect 675327 288493 675393 288494
rect 675135 285302 675201 285303
rect 675135 285238 675136 285302
rect 675200 285238 675201 285302
rect 675135 285237 675201 285238
rect 674943 281898 675009 281899
rect 674943 281834 674944 281898
rect 675008 281834 675009 281898
rect 674943 281833 675009 281834
rect 674751 278198 674817 278199
rect 674751 278134 674752 278198
rect 674816 278134 674817 278198
rect 674751 278133 674817 278134
rect 674559 276570 674625 276571
rect 674559 276506 674560 276570
rect 674624 276506 674625 276570
rect 674559 276505 674625 276506
rect 674367 274202 674433 274203
rect 674367 274138 674368 274202
rect 674432 274138 674433 274202
rect 674367 274137 674433 274138
rect 42111 270650 42177 270651
rect 42111 270586 42112 270650
rect 42176 270586 42177 270650
rect 42111 270585 42177 270586
rect 41919 269318 41985 269319
rect 41919 269254 41920 269318
rect 41984 269254 41985 269318
rect 41919 269253 41985 269254
rect 675522 265767 675582 310397
rect 675711 306466 675777 306467
rect 675711 306402 675712 306466
rect 675776 306402 675777 306466
rect 675711 306401 675777 306402
rect 675714 292851 675774 306401
rect 675903 302470 675969 302471
rect 675903 302406 675904 302470
rect 675968 302406 675969 302470
rect 675903 302405 675969 302406
rect 675711 292850 675777 292851
rect 675711 292786 675712 292850
rect 675776 292786 675777 292850
rect 675711 292785 675777 292786
rect 675906 290779 675966 302405
rect 676095 299214 676161 299215
rect 676095 299150 676096 299214
rect 676160 299150 676161 299214
rect 676095 299149 676161 299150
rect 675903 290778 675969 290779
rect 675903 290714 675904 290778
rect 675968 290714 675969 290778
rect 675903 290713 675969 290714
rect 676098 283675 676158 299149
rect 676095 283674 676161 283675
rect 676095 283610 676096 283674
rect 676160 283610 676161 283674
rect 676095 283609 676161 283610
rect 675519 265766 675585 265767
rect 675519 265702 675520 265766
rect 675584 265702 675585 265766
rect 675519 265701 675585 265702
rect 673983 263250 674049 263251
rect 673983 263186 673984 263250
rect 674048 263186 674049 263250
rect 673983 263185 674049 263186
rect 41919 252002 41985 252003
rect 41919 251938 41920 252002
rect 41984 251938 41985 252002
rect 41919 251937 41985 251938
rect 41535 251262 41601 251263
rect 41535 251198 41536 251262
rect 41600 251198 41601 251262
rect 41535 251197 41601 251198
rect 40959 250226 41025 250227
rect 40959 250162 40960 250226
rect 41024 250162 41025 250226
rect 40959 250161 41025 250162
rect 40575 249782 40641 249783
rect 40575 249718 40576 249782
rect 40640 249718 40641 249782
rect 40575 249717 40641 249718
rect 40383 246230 40449 246231
rect 40383 246166 40384 246230
rect 40448 246166 40449 246230
rect 40383 246165 40449 246166
rect 40386 231135 40446 246165
rect 40578 233355 40638 249717
rect 40767 248746 40833 248747
rect 40767 248682 40768 248746
rect 40832 248682 40833 248746
rect 40767 248681 40833 248682
rect 40575 233354 40641 233355
rect 40575 233290 40576 233354
rect 40640 233290 40641 233354
rect 40575 233289 40641 233290
rect 40383 231134 40449 231135
rect 40383 231070 40384 231134
rect 40448 231070 40449 231134
rect 40383 231069 40449 231070
rect 40770 226695 40830 248681
rect 40962 229063 41022 250161
rect 41343 248302 41409 248303
rect 41343 248238 41344 248302
rect 41408 248238 41409 248302
rect 41343 248237 41409 248238
rect 41151 247710 41217 247711
rect 41151 247646 41152 247710
rect 41216 247646 41217 247710
rect 41151 247645 41217 247646
rect 41154 230395 41214 247645
rect 41151 230394 41217 230395
rect 41151 230330 41152 230394
rect 41216 230330 41217 230394
rect 41151 230329 41217 230330
rect 41346 229803 41406 248237
rect 41538 237943 41598 251197
rect 41535 237942 41601 237943
rect 41535 237878 41536 237942
rect 41600 237878 41601 237942
rect 41535 237877 41601 237878
rect 41922 236793 41982 251937
rect 42111 250966 42177 250967
rect 42111 250902 42112 250966
rect 42176 250902 42177 250966
rect 42111 250901 42177 250902
rect 41538 236733 41982 236793
rect 41343 229802 41409 229803
rect 41343 229738 41344 229802
rect 41408 229738 41409 229802
rect 41343 229737 41409 229738
rect 40959 229062 41025 229063
rect 40959 228998 40960 229062
rect 41024 228998 41025 229062
rect 40959 228997 41025 228998
rect 41538 227435 41598 236733
rect 41535 227434 41601 227435
rect 41535 227370 41536 227434
rect 41600 227370 41601 227434
rect 41535 227369 41601 227370
rect 40767 226694 40833 226695
rect 40767 226630 40768 226694
rect 40832 226630 40833 226694
rect 40767 226629 40833 226630
rect 42114 226251 42174 250901
rect 42111 226250 42177 226251
rect 42111 226186 42112 226250
rect 42176 226186 42177 226250
rect 42111 226185 42177 226186
rect 673986 218555 674046 263185
rect 675519 262806 675585 262807
rect 675519 262742 675520 262806
rect 675584 262742 675585 262806
rect 675519 262741 675585 262742
rect 674367 258366 674433 258367
rect 674367 258302 674368 258366
rect 674432 258302 674433 258366
rect 674367 258301 674433 258302
rect 674370 240607 674430 258301
rect 674943 257774 675009 257775
rect 674943 257710 674944 257774
rect 675008 257710 675009 257774
rect 674943 257709 675009 257710
rect 674946 242087 675006 257709
rect 675522 249635 675582 262741
rect 676287 261474 676353 261475
rect 676287 261410 676288 261474
rect 676352 261410 676353 261474
rect 676287 261409 676353 261410
rect 675711 260734 675777 260735
rect 675711 260670 675712 260734
rect 675776 260670 675777 260734
rect 675711 260669 675777 260670
rect 675519 249634 675585 249635
rect 675519 249570 675520 249634
rect 675584 249570 675585 249634
rect 675519 249569 675585 249570
rect 675714 243567 675774 260669
rect 675903 253334 675969 253335
rect 675903 253270 675904 253334
rect 675968 253270 675969 253334
rect 675903 253269 675969 253270
rect 675711 243566 675777 243567
rect 675711 243502 675712 243566
rect 675776 243502 675777 243566
rect 675711 243501 675777 243502
rect 674943 242086 675009 242087
rect 674943 242022 674944 242086
rect 675008 242022 675009 242086
rect 674943 242021 675009 242022
rect 674367 240606 674433 240607
rect 674367 240542 674368 240606
rect 674432 240542 674433 240606
rect 674367 240541 674433 240542
rect 675906 236907 675966 253269
rect 676095 253186 676161 253187
rect 676095 253122 676096 253186
rect 676160 253122 676161 253186
rect 676095 253121 676161 253122
rect 676098 238683 676158 253121
rect 676290 250819 676350 261409
rect 676287 250818 676353 250819
rect 676287 250754 676288 250818
rect 676352 250754 676353 250818
rect 676287 250753 676353 250754
rect 676095 238682 676161 238683
rect 676095 238618 676096 238682
rect 676160 238618 676161 238682
rect 676095 238617 676161 238618
rect 675903 236906 675969 236907
rect 675903 236842 675904 236906
rect 675968 236842 675969 236906
rect 675903 236841 675969 236842
rect 674175 220034 674241 220035
rect 674175 219970 674176 220034
rect 674240 219970 674241 220034
rect 674175 219969 674241 219970
rect 673983 218554 674049 218555
rect 673983 218490 673984 218554
rect 674048 218490 674049 218554
rect 673983 218489 674049 218490
rect 40767 207158 40833 207159
rect 40767 207094 40768 207158
rect 40832 207094 40833 207158
rect 40767 207093 40833 207094
rect 40770 185847 40830 207093
rect 41151 205530 41217 205531
rect 41151 205466 41152 205530
rect 41216 205466 41217 205530
rect 41151 205465 41217 205466
rect 40959 205086 41025 205087
rect 40959 205022 40960 205086
rect 41024 205022 41025 205086
rect 40959 205021 41025 205022
rect 40962 186439 41022 205021
rect 40959 186438 41025 186439
rect 40959 186374 40960 186438
rect 41024 186374 41025 186438
rect 40959 186373 41025 186374
rect 40767 185846 40833 185847
rect 40767 185782 40768 185846
rect 40832 185782 40833 185846
rect 40767 185781 40833 185782
rect 41154 183479 41214 205465
rect 42111 204790 42177 204791
rect 42111 204726 42112 204790
rect 42176 204726 42177 204790
rect 42111 204725 42177 204726
rect 41919 203236 41985 203237
rect 41919 203172 41920 203236
rect 41984 203172 41985 203236
rect 41919 203171 41985 203172
rect 41727 200498 41793 200499
rect 41727 200434 41728 200498
rect 41792 200434 41793 200498
rect 41727 200433 41793 200434
rect 41343 200054 41409 200055
rect 41343 199990 41344 200054
rect 41408 199990 41409 200054
rect 41343 199989 41409 199990
rect 41346 184219 41406 199989
rect 41535 199610 41601 199611
rect 41535 199546 41536 199610
rect 41600 199546 41601 199610
rect 41535 199545 41601 199546
rect 41538 190139 41598 199545
rect 41730 195319 41790 200433
rect 41727 195318 41793 195319
rect 41727 195254 41728 195318
rect 41792 195254 41793 195318
rect 41727 195253 41793 195254
rect 41535 190138 41601 190139
rect 41535 190074 41536 190138
rect 41600 190074 41601 190138
rect 41535 190073 41601 190074
rect 41922 187919 41982 203171
rect 41919 187918 41985 187919
rect 41919 187854 41920 187918
rect 41984 187854 41985 187918
rect 41919 187853 41985 187854
rect 42114 187179 42174 204725
rect 42303 201090 42369 201091
rect 42303 201026 42304 201090
rect 42368 201026 42369 201090
rect 42303 201025 42369 201026
rect 42111 187178 42177 187179
rect 42111 187114 42112 187178
rect 42176 187114 42177 187178
rect 42111 187113 42177 187114
rect 41343 184218 41409 184219
rect 41343 184154 41344 184218
rect 41408 184154 41409 184218
rect 41343 184153 41409 184154
rect 41151 183478 41217 183479
rect 41151 183414 41152 183478
rect 41216 183414 41217 183478
rect 41151 183413 41217 183414
rect 42306 183035 42366 201025
rect 42303 183034 42369 183035
rect 42303 182970 42304 183034
rect 42368 182970 42369 183034
rect 42303 182969 42369 182970
rect 674178 176227 674238 219969
rect 675327 219146 675393 219147
rect 675327 219082 675328 219146
rect 675392 219082 675393 219146
rect 675327 219081 675393 219082
rect 674367 217962 674433 217963
rect 674367 217898 674368 217962
rect 674432 217898 674433 217962
rect 674367 217897 674433 217898
rect 674175 176226 674241 176227
rect 674175 176162 674176 176226
rect 674240 176162 674241 176226
rect 674175 176161 674241 176162
rect 673983 174746 674049 174747
rect 673983 174682 673984 174746
rect 674048 174682 674049 174746
rect 673983 174681 674049 174682
rect 673986 129459 674046 174681
rect 674370 174155 674430 217897
rect 674559 213078 674625 213079
rect 674559 213014 674560 213078
rect 674624 213014 674625 213078
rect 674559 213013 674625 213014
rect 674562 195319 674622 213013
rect 674559 195318 674625 195319
rect 674559 195254 674560 195318
rect 674624 195254 674625 195318
rect 674559 195253 674625 195254
rect 674559 175634 674625 175635
rect 674559 175570 674560 175634
rect 674624 175570 674625 175634
rect 674559 175569 674625 175570
rect 674367 174154 674433 174155
rect 674367 174090 674368 174154
rect 674432 174090 674433 174154
rect 674367 174089 674433 174090
rect 674175 173562 674241 173563
rect 674175 173498 674176 173562
rect 674240 173498 674241 173562
rect 674175 173497 674241 173498
rect 673983 129458 674049 129459
rect 673983 129394 673984 129458
rect 674048 129394 674049 129458
rect 673983 129393 674049 129394
rect 674178 128571 674238 173497
rect 674562 135390 674622 175569
rect 675330 175487 675390 219081
rect 675903 217666 675969 217667
rect 675903 217602 675904 217666
rect 675968 217602 675969 217666
rect 675903 217601 675969 217602
rect 675711 216112 675777 216113
rect 675711 216048 675712 216112
rect 675776 216048 675777 216112
rect 675711 216047 675777 216048
rect 675519 213522 675585 213523
rect 675519 213458 675520 213522
rect 675584 213458 675585 213522
rect 675519 213457 675585 213458
rect 675522 201387 675582 213457
rect 675714 202719 675774 216047
rect 675906 204495 675966 217601
rect 676095 215298 676161 215299
rect 676095 215234 676096 215298
rect 676160 215234 676161 215298
rect 676095 215233 676161 215234
rect 675903 204494 675969 204495
rect 675903 204430 675904 204494
rect 675968 204430 675969 204494
rect 675903 204429 675969 204430
rect 675711 202718 675777 202719
rect 675711 202654 675712 202718
rect 675776 202654 675777 202718
rect 675711 202653 675777 202654
rect 675519 201386 675585 201387
rect 675519 201322 675520 201386
rect 675584 201322 675585 201386
rect 675519 201321 675585 201322
rect 676098 198427 676158 215233
rect 676671 207602 676737 207603
rect 676671 207538 676672 207602
rect 676736 207538 676737 207602
rect 676671 207537 676737 207538
rect 676479 207454 676545 207455
rect 676479 207390 676480 207454
rect 676544 207390 676545 207454
rect 676479 207389 676545 207390
rect 676095 198426 676161 198427
rect 676095 198362 676096 198426
rect 676160 198362 676161 198426
rect 676095 198361 676161 198362
rect 676482 193543 676542 207389
rect 676479 193542 676545 193543
rect 676479 193478 676480 193542
rect 676544 193478 676545 193542
rect 676479 193477 676545 193478
rect 676674 191619 676734 207537
rect 676671 191618 676737 191619
rect 676671 191554 676672 191618
rect 676736 191554 676737 191618
rect 676671 191553 676737 191554
rect 675327 175486 675393 175487
rect 675327 175422 675328 175486
rect 675392 175422 675393 175486
rect 675327 175421 675393 175422
rect 676287 172970 676353 172971
rect 676287 172906 676288 172970
rect 676352 172906 676353 172970
rect 676287 172905 676353 172906
rect 674751 172674 674817 172675
rect 674751 172610 674752 172674
rect 674816 172610 674817 172674
rect 674751 172609 674817 172610
rect 674754 148551 674814 172609
rect 675711 171712 675777 171713
rect 675711 171648 675712 171712
rect 675776 171648 675777 171712
rect 675711 171647 675777 171648
rect 675327 171194 675393 171195
rect 675327 171130 675328 171194
rect 675392 171130 675393 171194
rect 675327 171129 675393 171130
rect 674943 168678 675009 168679
rect 674943 168614 674944 168678
rect 675008 168614 675009 168678
rect 674943 168613 675009 168614
rect 674946 150327 675006 168613
rect 675135 167198 675201 167199
rect 675135 167134 675136 167198
rect 675200 167134 675201 167198
rect 675135 167133 675201 167134
rect 675138 152547 675198 167133
rect 675330 153435 675390 171129
rect 675519 168234 675585 168235
rect 675519 168170 675520 168234
rect 675584 168170 675585 168234
rect 675519 168169 675585 168170
rect 675327 153434 675393 153435
rect 675327 153370 675328 153434
rect 675392 153370 675393 153434
rect 675327 153369 675393 153370
rect 675135 152546 675201 152547
rect 675135 152482 675136 152546
rect 675200 152482 675201 152546
rect 675135 152481 675201 152482
rect 675522 152251 675582 168169
rect 675714 157727 675774 171647
rect 676095 170454 676161 170455
rect 676095 170390 676096 170454
rect 676160 170390 676161 170454
rect 676095 170389 676161 170390
rect 675903 167642 675969 167643
rect 675903 167578 675904 167642
rect 675968 167578 675969 167642
rect 675903 167577 675969 167578
rect 675711 157726 675777 157727
rect 675711 157662 675712 157726
rect 675776 157662 675777 157726
rect 675711 157661 675777 157662
rect 675906 155507 675966 167577
rect 675903 155506 675969 155507
rect 675903 155442 675904 155506
rect 675968 155442 675969 155506
rect 675903 155441 675969 155442
rect 675519 152250 675585 152251
rect 675519 152186 675520 152250
rect 675584 152186 675585 152250
rect 675519 152185 675585 152186
rect 674943 150326 675009 150327
rect 674943 150262 674944 150326
rect 675008 150262 675009 150326
rect 674943 150261 675009 150262
rect 674751 148550 674817 148551
rect 674751 148486 674752 148550
rect 674816 148486 674817 148550
rect 674751 148485 674817 148486
rect 676098 146627 676158 170389
rect 676290 159355 676350 172905
rect 676287 159354 676353 159355
rect 676287 159290 676288 159354
rect 676352 159290 676353 159354
rect 676287 159289 676353 159290
rect 676095 146626 676161 146627
rect 676095 146562 676096 146626
rect 676160 146562 676161 146626
rect 676095 146561 676161 146562
rect 674370 135330 674622 135390
rect 674370 130643 674430 135330
rect 674367 130642 674433 130643
rect 674367 130578 674368 130642
rect 674432 130578 674433 130642
rect 674367 130577 674433 130578
rect 674175 128570 674241 128571
rect 674175 128506 674176 128570
rect 674240 128506 674241 128570
rect 674175 128505 674241 128506
rect 675711 125610 675777 125611
rect 675711 125546 675712 125610
rect 675776 125546 675777 125610
rect 675711 125545 675777 125546
rect 673983 123094 674049 123095
rect 673983 123030 673984 123094
rect 674048 123030 674049 123094
rect 673983 123029 674049 123030
rect 673986 105187 674046 123029
rect 675519 122206 675585 122207
rect 675519 122142 675520 122206
rect 675584 122142 675585 122206
rect 675519 122141 675585 122142
rect 675522 106667 675582 122141
rect 675714 108147 675774 125545
rect 675903 116730 675969 116731
rect 675903 116666 675904 116730
rect 675968 116666 675969 116730
rect 675903 116665 675969 116666
rect 675711 108146 675777 108147
rect 675711 108082 675712 108146
rect 675776 108082 675777 108146
rect 675711 108081 675777 108082
rect 675519 106666 675585 106667
rect 675519 106602 675520 106666
rect 675584 106602 675585 106666
rect 675519 106601 675585 106602
rect 673983 105186 674049 105187
rect 673983 105122 673984 105186
rect 674048 105122 674049 105186
rect 673983 105121 674049 105122
rect 675906 103263 675966 116665
rect 676671 116138 676737 116139
rect 676671 116074 676672 116138
rect 676736 116074 676737 116138
rect 676671 116073 676737 116074
rect 675903 103262 675969 103263
rect 675903 103198 675904 103262
rect 675968 103198 675969 103262
rect 675903 103197 675969 103198
rect 676674 101487 676734 116073
rect 676671 101486 676737 101487
rect 676671 101422 676672 101486
rect 676736 101422 676737 101486
rect 676671 101421 676737 101422
rect 417471 40510 417537 40511
rect 417471 40446 417472 40510
rect 417536 40446 417537 40510
rect 417471 40445 417537 40446
rect 417663 40510 417729 40511
rect 417663 40446 417664 40510
rect 417728 40446 417729 40510
rect 417663 40445 417729 40446
rect 417474 40323 417534 40445
rect 417666 40323 417726 40445
rect 417474 40263 417726 40323
<< metal5 >>
rect 77610 1018624 89778 1030788
rect 129010 1018624 141178 1030788
rect 180410 1018624 192578 1030788
rect 231810 1018624 243978 1030788
rect 283410 1018624 295578 1030788
rect 334810 1018624 346978 1030788
rect 385210 1018624 397378 1030788
rect 474210 1018624 486378 1030788
rect 525610 1018624 537778 1030788
rect 577010 1018624 589178 1030788
rect 627410 1018624 639578 1030788
rect 6811 955610 18975 967778
rect 698624 954022 710788 966190
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876180
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786620 19088 799160
rect 698512 774440 711002 786980
rect 6598 743420 19088 755960
rect 698512 729440 711002 741980
rect 6598 700220 19088 712760
rect 698512 684440 711002 696980
rect 6598 657020 19088 669560
rect 698512 639240 711002 651780
rect 6598 613820 19088 626360
rect 698512 594240 711002 606780
rect 6598 570620 19088 583160
rect 698512 549040 711002 561580
rect 6598 527420 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399820 19088 412360
rect 698512 371840 711002 384380
rect 6598 356620 19088 369160
rect 698512 326640 711002 339180
rect 6598 313420 19088 325960
rect 6598 270220 19088 282760
rect 698512 281640 711002 294180
rect 6598 227020 19088 239560
rect 698512 236640 711002 249180
rect 6598 183820 19088 196360
rect 698512 191440 711002 203980
rect 698512 146440 711002 158980
rect 6811 111610 18975 123778
rect 698512 101240 711002 113780
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200180 19088
rect 243266 6167 254146 19619
rect 296240 6598 308780 19088
rect 351040 6598 363580 19088
rect 405840 6598 418380 19088
rect 460640 6598 473180 19088
rect 515440 6598 527980 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use user_id_programming  user_id_value
timestamp 1625094921
transform 1 0 656624 0 1 80926
box 0 0 7109 7077
use storage  storage
timestamp 1625094921
transform 1 0 52032 0 1 53156
box 1066 70 92000 191480
use mgmt_core  soc
timestamp 1625094921
transform 1 0 190434 0 1 53602
box 0 0 450000 168026
use sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped  rstb_level
timestamp 1625094921
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use simple_por  por
timestamp 1625094921
transform 1 0 654146 0 -1 112882
box 25 11 11344 8291
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1625094921
transform -1 0 710203 0 1 164000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1625094921
transform -1 0 710203 0 1 118400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1625094921
transform 1 0 7631 0 1 242800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1625094921
transform 1 0 7631 0 1 199600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1625094921
transform 1 0 7631 0 1 286000
box -1620 -364 34000 13964
use mgmt_protect  mgmt_buffers
timestamp 1625094921
transform 1 0 192180 0 1 240036
box -2762 -2778 222734 26170
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1625094921
transform -1 0 710203 0 1 208400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1625094921
transform -1 0 710203 0 1 253600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1625094921
transform 1 0 7631 0 1 372400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1625094921
transform 1 0 7631 0 1 329200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1625094921
transform -1 0 710203 0 1 298800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1625094921
transform -1 0 710203 0 1 344600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1625094921
transform 1 0 7631 0 1 413400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1625094921
transform 1 0 7631 0 1 462400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1625094921
transform -1 0 710203 0 1 477200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1625094921
transform -1 0 710203 0 1 389000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1625094921
transform 1 0 7631 0 1 588224
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1625094921
transform 1 0 7631 0 1 631400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1625094921
transform 1 0 7631 0 1 674600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1625094921
transform -1 0 710203 0 1 657000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1625094921
transform -1 0 710203 0 1 611800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1625094921
transform -1 0 710203 0 1 564800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1625094921
transform -1 0 710203 0 1 521600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1625094921
transform 1 0 7631 0 1 717800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1625094921
transform 1 0 7631 0 1 761000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1625094921
transform 1 0 7631 0 1 804200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1625094921
transform -1 0 710203 0 1 702000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[11\]
timestamp 1625094921
transform -1 0 710203 0 1 880800
box -1620 -364 34000 13964
use user_analog_project_wrapper  mprj
timestamp 1625094921
transform 1 0 65308 0 1 278718
box -800 -800 584800 704000
use chip_io_alt  padframe
timestamp 1625094921
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< labels >>
rlabel metal5 s 187640 6598 200180 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363580 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308780 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418380 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473180 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527980 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113780 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696980 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741980 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786980 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876180 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698624 954022 710788 966190 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 627410 1018624 639578 1030788 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 525610 1018624 537778 1030788 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 474210 1018624 486378 1030788 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 385210 1018624 397378 1030788 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 283410 1018624 295578 1030788 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158980 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 231810 1018624 243978 1030788 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 180410 1018624 192578 1030788 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 129010 1018624 141178 1030788 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 77610 1018624 89778 1030788 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6811 955610 18975 967778 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786620 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743420 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700220 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657020 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613820 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203980 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570620 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527420 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399820 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356620 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313420 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270220 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227020 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183820 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249180 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294180 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339180 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384380 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561580 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606780 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651780 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144149 18309 6 resetb
port 44 nsew signal input
rlabel metal5 s 697980 909666 711432 920546 6 vccd1
port 45 nsew signal bidirectional
rlabel metal5 s 6167 914054 19619 924934 6 vccd2
port 46 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18975 6 vdda
port 47 nsew signal bidirectional
rlabel metal5 s 698624 819822 710788 831990 6 vdda1
port 48 nsew signal bidirectional
rlabel metal5 s 698624 505222 710788 517390 6 vdda1_2
port 49 nsew signal bidirectional
rlabel metal5 s 6811 484410 18975 496578 6 vdda2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 871210 18975 883378 6 vddio_2
port 51 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030788 6 vssa1
port 52 nsew signal bidirectional
rlabel metal5 s 698624 417022 710788 429190 6 vssa1_2
port 53 nsew signal bidirectional
rlabel metal5 s 6811 829010 18975 841178 6 vssa2
port 54 nsew signal bidirectional
rlabel metal5 s 697980 461866 711432 472746 6 vssd1
port 55 nsew signal bidirectional
rlabel metal5 s 6167 442854 19619 453734 6 vssd2
port 56 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030788 6 vssio_2
port 57 nsew signal bidirectional
rlabel metal5 s 6811 111610 18975 123778 6 vddio
port 58 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18975 6 vssio
port 59 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18975 6 vssa
port 60 nsew signal bidirectional
rlabel metal5 s 6167 70054 19619 80934 6 vccd
port 61 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19619 6 vssd
port 62 nsew signal bidirectional
rlabel metal2 s 579796 53602 579852 54402 6 pwr_ctrl_out[0]
port 63 nsew signal tristate
rlabel metal2 s 597092 53602 597148 54402 6 pwr_ctrl_out[1]
port 64 nsew signal tristate
rlabel metal2 s 614388 53602 614444 54402 6 pwr_ctrl_out[2]
port 65 nsew signal tristate
rlabel metal2 s 631684 53602 631740 54402 6 pwr_ctrl_out[3]
port 66 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
