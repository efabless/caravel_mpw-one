magic
tech sky130A
magscale 1 2
timestamp 1605994897
<< pwell >>
rect -962 -458 962 458
<< mvnmos >>
rect -734 -200 -574 200
rect -516 -200 -356 200
rect -298 -200 -138 200
rect -80 -200 80 200
rect 138 -200 298 200
rect 356 -200 516 200
rect 574 -200 734 200
<< mvndiff >>
rect -792 188 -734 200
rect -792 -188 -780 188
rect -746 -188 -734 188
rect -792 -200 -734 -188
rect -574 188 -516 200
rect -574 -188 -562 188
rect -528 -188 -516 188
rect -574 -200 -516 -188
rect -356 188 -298 200
rect -356 -188 -344 188
rect -310 -188 -298 188
rect -356 -200 -298 -188
rect -138 188 -80 200
rect -138 -188 -126 188
rect -92 -188 -80 188
rect -138 -200 -80 -188
rect 80 188 138 200
rect 80 -188 92 188
rect 126 -188 138 188
rect 80 -200 138 -188
rect 298 188 356 200
rect 298 -188 310 188
rect 344 -188 356 188
rect 298 -200 356 -188
rect 516 188 574 200
rect 516 -188 528 188
rect 562 -188 574 188
rect 516 -200 574 -188
rect 734 188 792 200
rect 734 -188 746 188
rect 780 -188 792 188
rect 734 -200 792 -188
<< mvndiffc >>
rect -780 -188 -746 188
rect -562 -188 -528 188
rect -344 -188 -310 188
rect -126 -188 -92 188
rect 92 -188 126 188
rect 310 -188 344 188
rect 528 -188 562 188
rect 746 -188 780 188
<< mvpsubdiff >>
rect -926 410 926 422
rect -926 376 -818 410
rect 818 376 926 410
rect -926 364 926 376
rect -926 314 -868 364
rect -926 -314 -914 314
rect -880 -314 -868 314
rect 868 314 926 364
rect -926 -364 -868 -314
rect 868 -314 880 314
rect 914 -314 926 314
rect 868 -364 926 -314
rect -926 -376 926 -364
rect -926 -410 -818 -376
rect 818 -410 926 -376
rect -926 -422 926 -410
<< mvpsubdiffcont >>
rect -818 376 818 410
rect -914 -314 -880 314
rect 880 -314 914 314
rect -818 -410 818 -376
<< poly >>
rect -734 272 -574 288
rect -734 238 -718 272
rect -590 238 -574 272
rect -734 200 -574 238
rect -516 272 -356 288
rect -516 238 -500 272
rect -372 238 -356 272
rect -516 200 -356 238
rect -298 272 -138 288
rect -298 238 -282 272
rect -154 238 -138 272
rect -298 200 -138 238
rect -80 272 80 288
rect -80 238 -64 272
rect 64 238 80 272
rect -80 200 80 238
rect 138 272 298 288
rect 138 238 154 272
rect 282 238 298 272
rect 138 200 298 238
rect 356 272 516 288
rect 356 238 372 272
rect 500 238 516 272
rect 356 200 516 238
rect 574 272 734 288
rect 574 238 590 272
rect 718 238 734 272
rect 574 200 734 238
rect -734 -238 -574 -200
rect -734 -272 -718 -238
rect -590 -272 -574 -238
rect -734 -288 -574 -272
rect -516 -238 -356 -200
rect -516 -272 -500 -238
rect -372 -272 -356 -238
rect -516 -288 -356 -272
rect -298 -238 -138 -200
rect -298 -272 -282 -238
rect -154 -272 -138 -238
rect -298 -288 -138 -272
rect -80 -238 80 -200
rect -80 -272 -64 -238
rect 64 -272 80 -238
rect -80 -288 80 -272
rect 138 -238 298 -200
rect 138 -272 154 -238
rect 282 -272 298 -238
rect 138 -288 298 -272
rect 356 -238 516 -200
rect 356 -272 372 -238
rect 500 -272 516 -238
rect 356 -288 516 -272
rect 574 -238 734 -200
rect 574 -272 590 -238
rect 718 -272 734 -238
rect 574 -288 734 -272
<< polycont >>
rect -718 238 -590 272
rect -500 238 -372 272
rect -282 238 -154 272
rect -64 238 64 272
rect 154 238 282 272
rect 372 238 500 272
rect 590 238 718 272
rect -718 -272 -590 -238
rect -500 -272 -372 -238
rect -282 -272 -154 -238
rect -64 -272 64 -238
rect 154 -272 282 -238
rect 372 -272 500 -238
rect 590 -272 718 -238
<< locali >>
rect -914 376 -818 410
rect 818 376 914 410
rect -914 314 -880 376
rect 880 314 914 376
rect -734 238 -718 272
rect -590 238 -574 272
rect -516 238 -500 272
rect -372 238 -356 272
rect -298 238 -282 272
rect -154 238 -138 272
rect -80 238 -64 272
rect 64 238 80 272
rect 138 238 154 272
rect 282 238 298 272
rect 356 238 372 272
rect 500 238 516 272
rect 574 238 590 272
rect 718 238 734 272
rect -780 188 -746 204
rect -780 -204 -746 -188
rect -562 188 -528 204
rect -562 -204 -528 -188
rect -344 188 -310 204
rect -344 -204 -310 -188
rect -126 188 -92 204
rect -126 -204 -92 -188
rect 92 188 126 204
rect 92 -204 126 -188
rect 310 188 344 204
rect 310 -204 344 -188
rect 528 188 562 204
rect 528 -204 562 -188
rect 746 188 780 204
rect 746 -204 780 -188
rect -734 -272 -718 -238
rect -590 -272 -574 -238
rect -516 -272 -500 -238
rect -372 -272 -356 -238
rect -298 -272 -282 -238
rect -154 -272 -138 -238
rect -80 -272 -64 -238
rect 64 -272 80 -238
rect 138 -272 154 -238
rect 282 -272 298 -238
rect 356 -272 372 -238
rect 500 -272 516 -238
rect 574 -272 590 -238
rect 718 -272 734 -238
rect -914 -376 -880 -314
rect 880 -376 914 -314
rect -914 -410 -818 -376
rect 818 -410 914 -376
<< viali >>
rect -718 238 -590 272
rect -500 238 -372 272
rect -282 238 -154 272
rect -64 238 64 272
rect 154 238 282 272
rect 372 238 500 272
rect 590 238 718 272
rect -780 21 -746 171
rect -562 -171 -528 -21
rect -344 21 -310 171
rect -126 -171 -92 -21
rect 92 21 126 171
rect 310 -171 344 -21
rect 528 21 562 171
rect 746 -171 780 -21
rect -718 -272 -590 -238
rect -500 -272 -372 -238
rect -282 -272 -154 -238
rect -64 -272 64 -238
rect 154 -272 282 -238
rect 372 -272 500 -238
rect 590 -272 718 -238
<< metal1 >>
rect -730 272 -578 278
rect -730 238 -718 272
rect -590 238 -578 272
rect -730 232 -578 238
rect -512 272 -360 278
rect -512 238 -500 272
rect -372 238 -360 272
rect -512 232 -360 238
rect -294 272 -142 278
rect -294 238 -282 272
rect -154 238 -142 272
rect -294 232 -142 238
rect -76 272 76 278
rect -76 238 -64 272
rect 64 238 76 272
rect -76 232 76 238
rect 142 272 294 278
rect 142 238 154 272
rect 282 238 294 272
rect 142 232 294 238
rect 360 272 512 278
rect 360 238 372 272
rect 500 238 512 272
rect 360 232 512 238
rect 578 272 730 278
rect 578 238 590 272
rect 718 238 730 272
rect 578 232 730 238
rect -786 171 -740 183
rect -786 21 -780 171
rect -746 21 -740 171
rect -786 9 -740 21
rect -350 171 -304 183
rect -350 21 -344 171
rect -310 21 -304 171
rect -350 9 -304 21
rect 86 171 132 183
rect 86 21 92 171
rect 126 21 132 171
rect 86 9 132 21
rect 522 171 568 183
rect 522 21 528 171
rect 562 21 568 171
rect 522 9 568 21
rect -568 -21 -522 -9
rect -568 -171 -562 -21
rect -528 -171 -522 -21
rect -568 -183 -522 -171
rect -132 -21 -86 -9
rect -132 -171 -126 -21
rect -92 -171 -86 -21
rect -132 -183 -86 -171
rect 304 -21 350 -9
rect 304 -171 310 -21
rect 344 -171 350 -21
rect 304 -183 350 -171
rect 740 -21 786 -9
rect 740 -171 746 -21
rect 780 -171 786 -21
rect 740 -183 786 -171
rect -730 -238 -578 -232
rect -730 -272 -718 -238
rect -590 -272 -578 -238
rect -730 -278 -578 -272
rect -512 -238 -360 -232
rect -512 -272 -500 -238
rect -372 -272 -360 -238
rect -512 -278 -360 -272
rect -294 -238 -142 -232
rect -294 -272 -282 -238
rect -154 -272 -142 -238
rect -294 -278 -142 -272
rect -76 -238 76 -232
rect -76 -272 -64 -238
rect 64 -272 76 -238
rect -76 -278 76 -272
rect 142 -238 294 -232
rect 142 -272 154 -238
rect 282 -272 294 -238
rect 142 -278 294 -272
rect 360 -238 512 -232
rect 360 -272 372 -238
rect 500 -272 512 -238
rect 360 -278 512 -272
rect 578 -238 730 -232
rect 578 -272 590 -238
rect 718 -272 730 -238
rect 578 -278 730 -272
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -897 -393 897 393
string parameters w 2.00 l 0.80 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
