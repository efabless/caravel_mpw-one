magic
tech sky130A
magscale 1 2
timestamp 1608231460
<< viali >>
rect 2881 11169 2915 11203
rect 4721 11169 4755 11203
rect 5641 11169 5675 11203
rect 5733 11169 5767 11203
rect 5917 11169 5951 11203
rect 6377 11169 6411 11203
rect 135 11101 169 11135
rect 5089 11101 5123 11135
rect 6469 11101 6503 11135
rect 3065 10965 3099 10999
rect 4813 10965 4847 10999
rect 4721 10761 4755 10795
rect 4445 10625 4479 10659
rect 5181 10625 5215 10659
rect 6653 10625 6687 10659
rect 1685 10557 1719 10591
rect 3893 10557 3927 10591
rect 4537 10557 4571 10591
rect 6561 10557 6595 10591
rect 1961 10489 1995 10523
rect 3709 10489 3743 10523
rect 4077 10421 4111 10455
rect 6377 10217 6411 10251
rect 1777 10149 1811 10183
rect 3525 10149 3559 10183
rect 3985 10081 4019 10115
rect 5825 10081 5859 10115
rect 6193 10081 6227 10115
rect 1501 10013 1535 10047
rect 3617 10013 3651 10047
rect 5733 9877 5767 9911
rect 6009 9877 6043 9911
rect 4261 9673 4295 9707
rect 6653 9673 6687 9707
rect 3617 9537 3651 9571
rect 4445 9537 4479 9571
rect 2697 9469 2731 9503
rect 2973 9469 3007 9503
rect 3157 9469 3191 9503
rect 3525 9469 3559 9503
rect 4077 9469 4111 9503
rect 6561 9469 6595 9503
rect 2237 9401 2271 9435
rect 4721 9401 4755 9435
rect 6469 9401 6503 9435
rect 2789 9129 2823 9163
rect 5365 9129 5399 9163
rect 6377 9129 6411 9163
rect 3249 9061 3283 9095
rect 5089 9061 5123 9095
rect 1961 8993 1995 9027
rect 2513 8993 2547 9027
rect 2605 8993 2639 9027
rect 5273 8993 5307 9027
rect 6285 8993 6319 9027
rect 2973 8925 3007 8959
rect 4997 8925 5031 8959
rect 2329 8857 2363 8891
rect 2145 8789 2179 8823
rect 6653 8585 6687 8619
rect 3525 8517 3559 8551
rect 4169 8517 4203 8551
rect 1501 8449 1535 8483
rect 1225 8381 1259 8415
rect 3341 8381 3375 8415
rect 3985 8381 4019 8415
rect 4353 8381 4387 8415
rect 6469 8381 6503 8415
rect 3249 8313 3283 8347
rect 4629 8313 4663 8347
rect 6377 8313 6411 8347
rect 2329 7973 2363 8007
rect 1317 7905 1351 7939
rect 1685 7905 1719 7939
rect 2053 7905 2087 7939
rect 4169 7905 4203 7939
rect 4077 7837 4111 7871
rect 4537 7837 4571 7871
rect 5917 7837 5951 7871
rect 1501 7701 1535 7735
rect 1869 7701 1903 7735
rect 1225 7361 1259 7395
rect 1501 7361 1535 7395
rect 3893 7361 3927 7395
rect 4169 7361 4203 7395
rect 5917 7361 5951 7395
rect 3433 7293 3467 7327
rect 6377 7293 6411 7327
rect 3249 7225 3283 7259
rect 3617 7157 3651 7191
rect 6193 7157 6227 7191
rect 6561 7157 6595 7191
rect 5917 6885 5951 6919
rect 1869 6817 1903 6851
rect 2237 6817 2271 6851
rect 5089 6817 5123 6851
rect 2973 6749 3007 6783
rect 3249 6749 3283 6783
rect 4997 6749 5031 6783
rect 5825 6749 5859 6783
rect 6469 6749 6503 6783
rect 2053 6613 2087 6647
rect 2421 6613 2455 6647
rect 5273 6613 5307 6647
rect 3617 6409 3651 6443
rect 1501 6273 1535 6307
rect 4353 6273 4387 6307
rect 1225 6205 1259 6239
rect 3433 6205 3467 6239
rect 3893 6205 3927 6239
rect 6469 6205 6503 6239
rect 3249 6137 3283 6171
rect 4629 6137 4663 6171
rect 6377 6137 6411 6171
rect 4077 6069 4111 6103
rect 6653 6069 6687 6103
rect 6101 5865 6135 5899
rect 1501 5797 1535 5831
rect 5549 5729 5583 5763
rect 5917 5729 5951 5763
rect 6285 5729 6319 5763
rect 1225 5661 1259 5695
rect 3249 5661 3283 5695
rect 3341 5661 3375 5695
rect 3617 5661 3651 5695
rect 5365 5661 5399 5695
rect 5733 5525 5767 5559
rect 6377 5525 6411 5559
rect 4169 5321 4203 5355
rect 1501 5185 1535 5219
rect 4629 5185 4663 5219
rect 4997 5185 5031 5219
rect 6377 5185 6411 5219
rect 1225 5117 1259 5151
rect 3341 5117 3375 5151
rect 3985 5117 4019 5151
rect 3249 5049 3283 5083
rect 3525 4981 3559 5015
rect 1685 4777 1719 4811
rect 6009 4777 6043 4811
rect 1409 4641 1443 4675
rect 1526 4641 1560 4675
rect 1869 4641 1903 4675
rect 2237 4641 2271 4675
rect 2605 4641 2639 4675
rect 4721 4641 4755 4675
rect 2881 4573 2915 4607
rect 4629 4573 4663 4607
rect 1225 4437 1259 4471
rect 2053 4437 2087 4471
rect 2421 4437 2455 4471
rect 3525 4233 3559 4267
rect 1501 4097 1535 4131
rect 3893 4097 3927 4131
rect 6009 4097 6043 4131
rect 1225 4029 1259 4063
rect 3341 4029 3375 4063
rect 5917 4029 5951 4063
rect 6193 4029 6227 4063
rect 6285 4029 6319 4063
rect 3249 3961 3283 3995
rect 4169 3961 4203 3995
rect 6745 3961 6779 3995
rect 2881 3621 2915 3655
rect 5089 3621 5123 3655
rect 2237 3553 2271 3587
rect 2605 3553 2639 3587
rect 4721 3553 4755 3587
rect 5273 3553 5307 3587
rect 5641 3553 5675 3587
rect 6009 3553 6043 3587
rect 6469 3553 6503 3587
rect 4629 3485 4663 3519
rect 4905 3417 4939 3451
rect 5825 3417 5859 3451
rect 2421 3349 2455 3383
rect 6653 3145 6687 3179
rect 1685 3009 1719 3043
rect 1961 3009 1995 3043
rect 3709 3009 3743 3043
rect 3893 2941 3927 2975
rect 4445 2941 4479 2975
rect 4537 2941 4571 2975
rect 4905 2941 4939 2975
rect 4077 2805 4111 2839
rect 4261 2805 4295 2839
rect 4077 2601 4111 2635
rect 3709 2533 3743 2567
rect 4813 2533 4847 2567
rect 6561 2533 6595 2567
rect 1685 2465 1719 2499
rect 3893 2465 3927 2499
rect 4537 2465 4571 2499
rect 1961 2397 1995 2431
<< metal1 >>
rect 6362 12520 6368 12572
rect 6420 12560 6426 12572
rect 16574 12560 16580 12572
rect 6420 12532 16580 12560
rect 6420 12520 6426 12532
rect 16574 12520 16580 12532
rect 16632 12520 16638 12572
rect 3970 12452 3976 12504
rect 4028 12492 4034 12504
rect 16666 12492 16672 12504
rect 4028 12464 16672 12492
rect 4028 12452 4034 12464
rect 16666 12452 16672 12464
rect 16724 12452 16730 12504
rect -1630 11464 680 11472
rect -1630 11386 -1606 11464
rect -1318 11386 680 11464
rect -1630 11376 680 11386
rect 896 11450 7084 11472
rect 896 11398 3598 11450
rect 3650 11398 3662 11450
rect 3714 11398 3726 11450
rect 3778 11398 3790 11450
rect 3842 11398 7084 11450
rect 896 11376 7084 11398
rect 2869 11203 2927 11209
rect 2869 11169 2881 11203
rect 2915 11200 2927 11203
rect 3878 11200 3884 11212
rect 2915 11172 3884 11200
rect 2915 11169 2927 11172
rect 2869 11163 2927 11169
rect 3878 11160 3884 11172
rect 3936 11160 3942 11212
rect 4706 11200 4712 11212
rect 4667 11172 4712 11200
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5626 11200 5632 11212
rect 5587 11172 5632 11200
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5721 11203 5779 11209
rect 5721 11169 5733 11203
rect 5767 11169 5779 11203
rect 5902 11200 5908 11212
rect 5863 11172 5908 11200
rect 5721 11163 5779 11169
rect 123 11135 181 11141
rect 123 11101 135 11135
rect 169 11132 181 11135
rect 4982 11132 4988 11144
rect 169 11104 4988 11132
rect 169 11101 181 11104
rect 123 11095 181 11101
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5442 11132 5448 11144
rect 5123 11104 5448 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 5736 11132 5764 11163
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 6362 11200 6368 11212
rect 6323 11172 6368 11200
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 6178 11132 6184 11144
rect 5736 11104 6184 11132
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 6454 11132 6460 11144
rect 6415 11104 6460 11132
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 1762 11024 1768 11076
rect 1820 11064 1826 11076
rect 16574 11064 16580 11076
rect 1820 11036 16580 11064
rect 1820 11024 1826 11036
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 3050 10996 3056 11008
rect 3011 10968 3056 10996
rect 3050 10956 3056 10968
rect 3108 10956 3114 11008
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 4801 10999 4859 11005
rect 4801 10996 4813 10999
rect 4580 10968 4813 10996
rect 4580 10956 4586 10968
rect 4801 10965 4813 10968
rect 4847 10965 4859 10999
rect 4801 10959 4859 10965
rect -988 10918 680 10928
rect -988 10844 -948 10918
rect -658 10844 680 10918
rect -988 10832 680 10844
rect 896 10906 7084 10928
rect 896 10854 2098 10906
rect 2150 10854 2162 10906
rect 2214 10854 2226 10906
rect 2278 10854 2290 10906
rect 2342 10854 5098 10906
rect 5150 10854 5162 10906
rect 5214 10854 5226 10906
rect 5278 10854 5290 10906
rect 5342 10854 7084 10906
rect 896 10832 7084 10854
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 4709 10795 4767 10801
rect 4709 10792 4721 10795
rect 4488 10764 4721 10792
rect 4488 10752 4494 10764
rect 4709 10761 4721 10764
rect 4755 10761 4767 10795
rect 4709 10755 4767 10761
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10656 4491 10659
rect 4614 10656 4620 10668
rect 4479 10628 4620 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5169 10659 5227 10665
rect 5169 10656 5181 10659
rect 5040 10628 5181 10656
rect 5040 10616 5046 10628
rect 5169 10625 5181 10628
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 16758 10656 16764 10668
rect 6687 10628 16764 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 1486 10548 1492 10600
rect 1544 10588 1550 10600
rect 1673 10591 1731 10597
rect 1673 10588 1685 10591
rect 1544 10560 1685 10588
rect 1544 10548 1550 10560
rect 1673 10557 1685 10560
rect 1719 10557 1731 10591
rect 3878 10588 3884 10600
rect 3839 10560 3884 10588
rect 1673 10551 1731 10557
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4522 10548 4528 10600
rect 4580 10588 4586 10600
rect 6546 10588 6552 10600
rect 4580 10560 4625 10588
rect 6507 10560 6552 10588
rect 4580 10548 4586 10560
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 1946 10520 1952 10532
rect 1907 10492 1952 10520
rect 1946 10480 1952 10492
rect 2004 10480 2010 10532
rect 3697 10523 3755 10529
rect 3160 10452 3188 10506
rect 3697 10489 3709 10523
rect 3743 10520 3755 10523
rect 4338 10520 4344 10532
rect 3743 10492 4344 10520
rect 3743 10489 3755 10492
rect 3697 10483 3755 10489
rect 4338 10480 4344 10492
rect 4396 10480 4402 10532
rect 4065 10455 4123 10461
rect 4065 10452 4077 10455
rect 3160 10424 4077 10452
rect 4065 10421 4077 10424
rect 4111 10421 4123 10455
rect 4065 10415 4123 10421
rect 4706 10412 4712 10464
rect 4764 10452 4770 10464
rect 16574 10452 16580 10464
rect 4764 10424 16580 10452
rect 4764 10412 4770 10424
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 920 10362 7084 10384
rect 920 10310 3598 10362
rect 3650 10310 3662 10362
rect 3714 10310 3726 10362
rect 3778 10310 3790 10362
rect 3842 10310 7084 10362
rect 920 10288 7084 10310
rect 1946 10208 1952 10260
rect 2004 10248 2010 10260
rect 6365 10251 6423 10257
rect 2004 10220 3556 10248
rect 2004 10208 2010 10220
rect 1762 10180 1768 10192
rect 1723 10152 1768 10180
rect 1762 10140 1768 10152
rect 1820 10140 1826 10192
rect 3050 10180 3056 10192
rect 2990 10152 3056 10180
rect 3050 10140 3056 10152
rect 3108 10140 3114 10192
rect 3528 10189 3556 10220
rect 6365 10217 6377 10251
rect 6411 10217 6423 10251
rect 6365 10211 6423 10217
rect 3513 10183 3571 10189
rect 3513 10149 3525 10183
rect 3559 10149 3571 10183
rect 6380 10180 6408 10211
rect 5014 10152 6408 10180
rect 3513 10143 3571 10149
rect 3528 10112 3556 10143
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 3528 10084 3985 10112
rect 3973 10081 3985 10084
rect 4019 10081 4031 10115
rect 5810 10112 5816 10124
rect 5771 10084 5816 10112
rect 3973 10075 4031 10081
rect 5810 10072 5816 10084
rect 5868 10112 5874 10124
rect 6181 10115 6239 10121
rect 6181 10112 6193 10115
rect 5868 10084 6193 10112
rect 5868 10072 5874 10084
rect 6181 10081 6193 10084
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 1486 10044 1492 10056
rect 1447 10016 1492 10044
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10044 3663 10047
rect 4430 10044 4436 10056
rect 3651 10016 4436 10044
rect 3651 10013 3663 10016
rect 3605 10007 3663 10013
rect 4430 10004 4436 10016
rect 4488 10004 4494 10056
rect 5718 9908 5724 9920
rect 5679 9880 5724 9908
rect 5718 9868 5724 9880
rect 5776 9868 5782 9920
rect 5994 9908 6000 9920
rect 5955 9880 6000 9908
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 920 9818 7084 9840
rect 920 9766 2098 9818
rect 2150 9766 2162 9818
rect 2214 9766 2226 9818
rect 2278 9766 2290 9818
rect 2342 9766 5098 9818
rect 5150 9766 5162 9818
rect 5214 9766 5226 9818
rect 5278 9766 5290 9818
rect 5342 9766 7084 9818
rect 920 9744 7084 9766
rect 4249 9707 4307 9713
rect 4249 9704 4261 9707
rect 3068 9676 4261 9704
rect 2866 9596 2872 9648
rect 2924 9636 2930 9648
rect 3068 9636 3096 9676
rect 4249 9673 4261 9676
rect 4295 9704 4307 9707
rect 5810 9704 5816 9716
rect 4295 9676 5816 9704
rect 4295 9673 4307 9676
rect 4249 9667 4307 9673
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 6641 9707 6699 9713
rect 6641 9704 6653 9707
rect 6604 9676 6653 9704
rect 6604 9664 6610 9676
rect 6641 9673 6653 9676
rect 6687 9673 6699 9707
rect 6641 9667 6699 9673
rect 2924 9608 3096 9636
rect 3160 9608 4568 9636
rect 2924 9596 2930 9608
rect 2682 9500 2688 9512
rect 2643 9472 2688 9500
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 2958 9500 2964 9512
rect 2919 9472 2964 9500
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3160 9509 3188 9608
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9568 3663 9571
rect 3970 9568 3976 9580
rect 3651 9540 3976 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 3970 9528 3976 9540
rect 4028 9528 4034 9580
rect 4430 9568 4436 9580
rect 4391 9540 4436 9568
rect 4430 9528 4436 9540
rect 4488 9528 4494 9580
rect 4540 9568 4568 9608
rect 5718 9568 5724 9580
rect 4540 9540 5724 9568
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9500 3571 9503
rect 4062 9500 4068 9512
rect 3559 9472 3832 9500
rect 4023 9472 4068 9500
rect 3559 9469 3571 9472
rect 3513 9463 3571 9469
rect 2225 9435 2283 9441
rect 2225 9401 2237 9435
rect 2271 9432 2283 9435
rect 2498 9432 2504 9444
rect 2271 9404 2504 9432
rect 2271 9401 2283 9404
rect 2225 9395 2283 9401
rect 2498 9392 2504 9404
rect 2556 9392 2562 9444
rect 3804 9364 3832 9472
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 6546 9500 6552 9512
rect 6507 9472 6552 9500
rect 6546 9460 6552 9472
rect 6604 9460 6610 9512
rect 4154 9392 4160 9444
rect 4212 9432 4218 9444
rect 4709 9435 4767 9441
rect 4709 9432 4721 9435
rect 4212 9404 4721 9432
rect 4212 9392 4218 9404
rect 4709 9401 4721 9404
rect 4755 9401 4767 9435
rect 5994 9432 6000 9444
rect 5934 9404 6000 9432
rect 4709 9395 4767 9401
rect 5994 9392 6000 9404
rect 6052 9392 6058 9444
rect 6457 9435 6515 9441
rect 6457 9401 6469 9435
rect 6503 9432 6515 9435
rect 26234 9432 26240 9444
rect 6503 9404 26240 9432
rect 6503 9401 6515 9404
rect 6457 9395 6515 9401
rect 26234 9392 26240 9404
rect 26292 9392 26298 9444
rect 6362 9364 6368 9376
rect 3804 9336 6368 9364
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 920 9274 7084 9296
rect 920 9222 3598 9274
rect 3650 9222 3662 9274
rect 3714 9222 3726 9274
rect 3778 9222 3790 9274
rect 3842 9222 7084 9274
rect 920 9200 7084 9222
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 3142 9160 3148 9172
rect 2823 9132 3148 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 3418 9160 3424 9172
rect 3252 9132 3424 9160
rect 3252 9101 3280 9132
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 5353 9163 5411 9169
rect 5353 9160 5365 9163
rect 4120 9132 5365 9160
rect 4120 9120 4126 9132
rect 5353 9129 5365 9132
rect 5399 9129 5411 9163
rect 5353 9123 5411 9129
rect 6365 9163 6423 9169
rect 6365 9129 6377 9163
rect 6411 9160 6423 9163
rect 6454 9160 6460 9172
rect 6411 9132 6460 9160
rect 6411 9129 6423 9132
rect 6365 9123 6423 9129
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 3237 9095 3295 9101
rect 3237 9061 3249 9095
rect 3283 9061 3295 9095
rect 3237 9055 3295 9061
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 3384 9064 3726 9092
rect 3384 9052 3390 9064
rect 4706 9052 4712 9104
rect 4764 9092 4770 9104
rect 5077 9095 5135 9101
rect 5077 9092 5089 9095
rect 4764 9064 5089 9092
rect 4764 9052 4770 9064
rect 5077 9061 5089 9064
rect 5123 9061 5135 9095
rect 5077 9055 5135 9061
rect 5442 9052 5448 9104
rect 5500 9092 5506 9104
rect 16574 9092 16580 9104
rect 5500 9064 16580 9092
rect 5500 9052 5506 9064
rect 16574 9052 16580 9064
rect 16632 9052 16638 9104
rect 1762 8984 1768 9036
rect 1820 9024 1826 9036
rect 1949 9027 2007 9033
rect 1949 9024 1961 9027
rect 1820 8996 1961 9024
rect 1820 8984 1826 8996
rect 1949 8993 1961 8996
rect 1995 8993 2007 9027
rect 1949 8987 2007 8993
rect 2406 8984 2412 9036
rect 2464 9024 2470 9036
rect 2501 9027 2559 9033
rect 2501 9024 2513 9027
rect 2464 8996 2513 9024
rect 2464 8984 2470 8996
rect 2501 8993 2513 8996
rect 2547 8993 2559 9027
rect 2501 8987 2559 8993
rect 2593 9027 2651 9033
rect 2593 8993 2605 9027
rect 2639 9024 2651 9027
rect 2866 9024 2872 9036
rect 2639 8996 2872 9024
rect 2639 8993 2651 8996
rect 2593 8987 2651 8993
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 4614 8984 4620 9036
rect 4672 9024 4678 9036
rect 5261 9027 5319 9033
rect 5261 9024 5273 9027
rect 4672 8996 5273 9024
rect 4672 8984 4678 8996
rect 5261 8993 5273 8996
rect 5307 8993 5319 9027
rect 5261 8987 5319 8993
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 6273 9027 6331 9033
rect 6273 9024 6285 9027
rect 5776 8996 6285 9024
rect 5776 8984 5782 8996
rect 6273 8993 6285 8996
rect 6319 8993 6331 9027
rect 6273 8987 6331 8993
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 4430 8956 4436 8968
rect 3007 8928 4436 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 16666 8956 16672 8968
rect 5031 8928 16672 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 16666 8916 16672 8928
rect 16724 8916 16730 8968
rect 1210 8848 1216 8900
rect 1268 8888 1274 8900
rect 1486 8888 1492 8900
rect 1268 8860 1492 8888
rect 1268 8848 1274 8860
rect 1486 8848 1492 8860
rect 1544 8888 1550 8900
rect 2317 8891 2375 8897
rect 2317 8888 2329 8891
rect 1544 8860 2329 8888
rect 1544 8848 1550 8860
rect 2317 8857 2329 8860
rect 2363 8857 2375 8891
rect 2317 8851 2375 8857
rect 1946 8780 1952 8832
rect 2004 8820 2010 8832
rect 2133 8823 2191 8829
rect 2133 8820 2145 8823
rect 2004 8792 2145 8820
rect 2004 8780 2010 8792
rect 2133 8789 2145 8792
rect 2179 8789 2191 8823
rect 2133 8783 2191 8789
rect 2958 8780 2964 8832
rect 3016 8820 3022 8832
rect 5626 8820 5632 8832
rect 3016 8792 5632 8820
rect 3016 8780 3022 8792
rect 5626 8780 5632 8792
rect 5684 8780 5690 8832
rect 920 8730 7084 8752
rect 920 8678 2098 8730
rect 2150 8678 2162 8730
rect 2214 8678 2226 8730
rect 2278 8678 2290 8730
rect 2342 8678 5098 8730
rect 5150 8678 5162 8730
rect 5214 8678 5226 8730
rect 5278 8678 5290 8730
rect 5342 8678 7084 8730
rect 920 8656 7084 8678
rect 3068 8588 4292 8616
rect 1489 8483 1547 8489
rect 1489 8449 1501 8483
rect 1535 8480 1547 8483
rect 3068 8480 3096 8588
rect 3142 8508 3148 8560
rect 3200 8548 3206 8560
rect 3513 8551 3571 8557
rect 3513 8548 3525 8551
rect 3200 8520 3525 8548
rect 3200 8508 3206 8520
rect 3513 8517 3525 8520
rect 3559 8548 3571 8551
rect 3878 8548 3884 8560
rect 3559 8520 3884 8548
rect 3559 8517 3571 8520
rect 3513 8511 3571 8517
rect 3878 8508 3884 8520
rect 3936 8508 3942 8560
rect 4157 8551 4215 8557
rect 4157 8517 4169 8551
rect 4203 8517 4215 8551
rect 4264 8548 4292 8588
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 6641 8619 6699 8625
rect 6641 8616 6653 8619
rect 4856 8588 6653 8616
rect 4856 8576 4862 8588
rect 6641 8585 6653 8588
rect 6687 8585 6699 8619
rect 6641 8579 6699 8585
rect 4338 8548 4344 8560
rect 4264 8520 4344 8548
rect 4157 8511 4215 8517
rect 4172 8480 4200 8511
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 4614 8480 4620 8492
rect 1535 8452 3096 8480
rect 3344 8452 4200 8480
rect 4356 8452 4620 8480
rect 1535 8449 1547 8452
rect 1489 8443 1547 8449
rect 3344 8424 3372 8452
rect 1210 8412 1216 8424
rect 1171 8384 1216 8412
rect 1210 8372 1216 8384
rect 1268 8372 1274 8424
rect 3326 8412 3332 8424
rect 3239 8384 3332 8412
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 4062 8412 4068 8424
rect 4019 8384 4068 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4356 8421 4384 8452
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 4341 8415 4399 8421
rect 4341 8381 4353 8415
rect 4387 8381 4399 8415
rect 5828 8412 5856 8440
rect 6457 8415 6515 8421
rect 6457 8412 6469 8415
rect 5828 8384 6469 8412
rect 4341 8375 4399 8381
rect 6457 8381 6469 8384
rect 6503 8381 6515 8415
rect 6457 8375 6515 8381
rect 1946 8304 1952 8356
rect 2004 8304 2010 8356
rect 3234 8344 3240 8356
rect 3195 8316 3240 8344
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 3878 8304 3884 8356
rect 3936 8344 3942 8356
rect 4356 8344 4384 8375
rect 3936 8316 4384 8344
rect 3936 8304 3942 8316
rect 4522 8304 4528 8356
rect 4580 8344 4586 8356
rect 4617 8347 4675 8353
rect 4617 8344 4629 8347
rect 4580 8316 4629 8344
rect 4580 8304 4586 8316
rect 4617 8313 4629 8316
rect 4663 8313 4675 8347
rect 4617 8307 4675 8313
rect 4706 8304 4712 8356
rect 4764 8344 4770 8356
rect 6362 8344 6368 8356
rect 4764 8316 5106 8344
rect 6323 8316 6368 8344
rect 4764 8304 4770 8316
rect 6362 8304 6368 8316
rect 6420 8344 6426 8356
rect 26326 8344 26332 8356
rect 6420 8316 26332 8344
rect 6420 8304 6426 8316
rect 26326 8304 26332 8316
rect 26384 8304 26390 8356
rect 2498 8236 2504 8288
rect 2556 8276 2562 8288
rect 16574 8276 16580 8288
rect 2556 8248 16580 8276
rect 2556 8236 2562 8248
rect 16574 8236 16580 8248
rect 16632 8236 16638 8288
rect 920 8186 7084 8208
rect 920 8134 3598 8186
rect 3650 8134 3662 8186
rect 3714 8134 3726 8186
rect 3778 8134 3790 8186
rect 3842 8134 7084 8186
rect 920 8112 7084 8134
rect 3234 8072 3240 8084
rect 2332 8044 3240 8072
rect 2332 8013 2360 8044
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 4798 8072 4804 8084
rect 3528 8044 4804 8072
rect 2317 8007 2375 8013
rect 2317 7973 2329 8007
rect 2363 7973 2375 8007
rect 3528 7990 3556 8044
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 2317 7967 2375 7973
rect 5442 7964 5448 8016
rect 5500 7964 5506 8016
rect 1305 7939 1363 7945
rect 1305 7905 1317 7939
rect 1351 7905 1363 7939
rect 1305 7899 1363 7905
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 1719 7908 1900 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 1320 7868 1348 7899
rect 1320 7840 1808 7868
rect 1780 7744 1808 7840
rect 1872 7800 1900 7908
rect 1946 7896 1952 7948
rect 2004 7936 2010 7948
rect 2041 7939 2099 7945
rect 2041 7936 2053 7939
rect 2004 7908 2053 7936
rect 2004 7896 2010 7908
rect 2041 7905 2053 7908
rect 2087 7905 2099 7939
rect 2041 7899 2099 7905
rect 4157 7939 4215 7945
rect 4157 7905 4169 7939
rect 4203 7936 4215 7939
rect 4430 7936 4436 7948
rect 4203 7908 4436 7936
rect 4203 7905 4215 7908
rect 4157 7899 4215 7905
rect 3050 7868 3056 7880
rect 2148 7840 3056 7868
rect 2148 7800 2176 7840
rect 3050 7828 3056 7840
rect 3108 7868 3114 7880
rect 3326 7868 3332 7880
rect 3108 7840 3332 7868
rect 3108 7828 3114 7840
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 1872 7772 2176 7800
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 1857 7735 1915 7741
rect 1857 7732 1869 7735
rect 1820 7704 1869 7732
rect 1820 7692 1826 7704
rect 1857 7701 1869 7704
rect 1903 7701 1915 7735
rect 1857 7695 1915 7701
rect 1946 7692 1952 7744
rect 2004 7732 2010 7744
rect 2958 7732 2964 7744
rect 2004 7704 2964 7732
rect 2004 7692 2010 7704
rect 2958 7692 2964 7704
rect 3016 7732 3022 7744
rect 4172 7732 4200 7899
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 4396 7840 4537 7868
rect 4396 7828 4402 7840
rect 4525 7837 4537 7840
rect 4571 7837 4583 7871
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 4525 7831 4583 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 3016 7704 4200 7732
rect 3016 7692 3022 7704
rect 6270 7692 6276 7744
rect 6328 7732 6334 7744
rect 6546 7732 6552 7744
rect 6328 7704 6552 7732
rect 6328 7692 6334 7704
rect 6546 7692 6552 7704
rect 6604 7732 6610 7744
rect 16666 7732 16672 7744
rect 6604 7704 16672 7732
rect 6604 7692 6610 7704
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 920 7642 7084 7664
rect 920 7590 2098 7642
rect 2150 7590 2162 7642
rect 2214 7590 2226 7642
rect 2278 7590 2290 7642
rect 2342 7590 5098 7642
rect 5150 7590 5162 7642
rect 5214 7590 5226 7642
rect 5278 7590 5290 7642
rect 5342 7590 7084 7642
rect 920 7568 7084 7590
rect 1210 7528 1216 7540
rect 1123 7500 1216 7528
rect 1210 7488 1216 7500
rect 1268 7528 1274 7540
rect 1268 7500 2544 7528
rect 1268 7488 1274 7500
rect 1228 7401 1256 7488
rect 2516 7460 2544 7500
rect 3142 7488 3148 7540
rect 3200 7528 3206 7540
rect 3326 7528 3332 7540
rect 3200 7500 3332 7528
rect 3200 7488 3206 7500
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 2516 7432 3924 7460
rect 3896 7404 3924 7432
rect 1213 7395 1271 7401
rect 1213 7361 1225 7395
rect 1259 7361 1271 7395
rect 1213 7355 1271 7361
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7392 1547 7395
rect 3234 7392 3240 7404
rect 1535 7364 3240 7392
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 3878 7392 3884 7404
rect 3839 7364 3884 7392
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 4154 7392 4160 7404
rect 4115 7364 4160 7392
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 5905 7395 5963 7401
rect 5905 7392 5917 7395
rect 4856 7364 5917 7392
rect 4856 7352 4862 7364
rect 5905 7361 5917 7364
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 2866 7284 2872 7336
rect 2924 7324 2930 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 2924 7296 3433 7324
rect 2924 7284 2930 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 3421 7287 3479 7293
rect 6196 7296 6377 7324
rect 1486 7216 1492 7268
rect 1544 7256 1550 7268
rect 3234 7256 3240 7268
rect 1544 7228 1978 7256
rect 3195 7228 3240 7256
rect 1544 7216 1550 7228
rect 3234 7216 3240 7228
rect 3292 7216 3298 7268
rect 4614 7216 4620 7268
rect 4672 7216 4678 7268
rect 3605 7191 3663 7197
rect 3605 7157 3617 7191
rect 3651 7188 3663 7191
rect 3970 7188 3976 7200
rect 3651 7160 3976 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 6196 7197 6224 7296
rect 6365 7293 6377 7296
rect 6411 7324 6423 7327
rect 16574 7324 16580 7336
rect 6411 7296 16580 7324
rect 6411 7293 6423 7296
rect 6365 7287 6423 7293
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 5592 7160 6193 7188
rect 5592 7148 5598 7160
rect 6181 7157 6193 7160
rect 6227 7157 6239 7191
rect 6546 7188 6552 7200
rect 6507 7160 6552 7188
rect 6181 7151 6239 7157
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 920 7098 7084 7120
rect 920 7046 3598 7098
rect 3650 7046 3662 7098
rect 3714 7046 3726 7098
rect 3778 7046 3790 7098
rect 3842 7046 7084 7098
rect 920 7024 7084 7046
rect 2590 6876 2596 6928
rect 2648 6916 2654 6928
rect 2648 6888 3004 6916
rect 2648 6876 2654 6888
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 1857 6851 1915 6857
rect 1857 6848 1869 6851
rect 1820 6820 1869 6848
rect 1820 6808 1826 6820
rect 1857 6817 1869 6820
rect 1903 6848 1915 6851
rect 2225 6851 2283 6857
rect 2225 6848 2237 6851
rect 1903 6820 2237 6848
rect 1903 6817 1915 6820
rect 1857 6811 1915 6817
rect 2225 6817 2237 6820
rect 2271 6817 2283 6851
rect 2225 6811 2283 6817
rect 2976 6792 3004 6888
rect 3970 6876 3976 6928
rect 4028 6876 4034 6928
rect 5905 6919 5963 6925
rect 5905 6885 5917 6919
rect 5951 6916 5963 6919
rect 6546 6916 6552 6928
rect 5951 6888 6552 6916
rect 5951 6885 5963 6888
rect 5905 6879 5963 6885
rect 6546 6876 6552 6888
rect 6604 6876 6610 6928
rect 5077 6851 5135 6857
rect 5077 6848 5089 6851
rect 4448 6820 5089 6848
rect 2958 6780 2964 6792
rect 2871 6752 2964 6780
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 3234 6780 3240 6792
rect 3195 6752 3240 6780
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3602 6740 3608 6792
rect 3660 6780 3666 6792
rect 4448 6780 4476 6820
rect 5077 6817 5089 6820
rect 5123 6817 5135 6851
rect 5077 6811 5135 6817
rect 3660 6752 4476 6780
rect 4985 6783 5043 6789
rect 3660 6740 3666 6752
rect 4985 6749 4997 6783
rect 5031 6780 5043 6783
rect 5534 6780 5540 6792
rect 5031 6752 5540 6780
rect 5031 6749 5043 6752
rect 4985 6743 5043 6749
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 6270 6780 6276 6792
rect 5859 6752 6276 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 6454 6780 6460 6792
rect 6415 6752 6460 6780
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 5718 6712 5724 6724
rect 4264 6684 5724 6712
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2041 6647 2099 6653
rect 2041 6644 2053 6647
rect 2004 6616 2053 6644
rect 2004 6604 2010 6616
rect 2041 6613 2053 6616
rect 2087 6613 2099 6647
rect 2041 6607 2099 6613
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 2498 6644 2504 6656
rect 2455 6616 2504 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4264 6644 4292 6684
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 4028 6616 4292 6644
rect 4028 6604 4034 6616
rect 4890 6604 4896 6656
rect 4948 6644 4954 6656
rect 5261 6647 5319 6653
rect 5261 6644 5273 6647
rect 4948 6616 5273 6644
rect 4948 6604 4954 6616
rect 5261 6613 5273 6616
rect 5307 6613 5319 6647
rect 5261 6607 5319 6613
rect 920 6554 7084 6576
rect 920 6502 2098 6554
rect 2150 6502 2162 6554
rect 2214 6502 2226 6554
rect 2278 6502 2290 6554
rect 2342 6502 5098 6554
rect 5150 6502 5162 6554
rect 5214 6502 5226 6554
rect 5278 6502 5290 6554
rect 5342 6502 7084 6554
rect 920 6480 7084 6502
rect 3605 6443 3663 6449
rect 3605 6409 3617 6443
rect 3651 6440 3663 6443
rect 4706 6440 4712 6452
rect 3651 6412 4712 6440
rect 3651 6409 3663 6412
rect 3605 6403 3663 6409
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 16574 6440 16580 6452
rect 5776 6412 16580 6440
rect 5776 6400 5782 6412
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 1489 6307 1547 6313
rect 1489 6273 1501 6307
rect 1535 6304 1547 6307
rect 3234 6304 3240 6316
rect 1535 6276 3240 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 4338 6304 4344 6316
rect 4299 6276 4344 6304
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 1210 6236 1216 6248
rect 1171 6208 1216 6236
rect 1210 6196 1216 6208
rect 1268 6196 1274 6248
rect 3050 6196 3056 6248
rect 3108 6236 3114 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3108 6208 3433 6236
rect 3108 6196 3114 6208
rect 3421 6205 3433 6208
rect 3467 6236 3479 6239
rect 3602 6236 3608 6248
rect 3467 6208 3608 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 3878 6236 3884 6248
rect 3839 6208 3884 6236
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 5902 6196 5908 6248
rect 5960 6236 5966 6248
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 5960 6208 6469 6236
rect 5960 6196 5966 6208
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 2498 6128 2504 6180
rect 2556 6128 2562 6180
rect 3234 6168 3240 6180
rect 3195 6140 3240 6168
rect 3234 6128 3240 6140
rect 3292 6168 3298 6180
rect 4617 6171 4675 6177
rect 4617 6168 4629 6171
rect 3292 6140 4629 6168
rect 3292 6128 3298 6140
rect 4617 6137 4629 6140
rect 4663 6137 4675 6171
rect 6086 6168 6092 6180
rect 5842 6140 6092 6168
rect 4617 6131 4675 6137
rect 6086 6128 6092 6140
rect 6144 6128 6150 6180
rect 6365 6171 6423 6177
rect 6365 6137 6377 6171
rect 6411 6168 6423 6171
rect 16666 6168 16672 6180
rect 6411 6140 16672 6168
rect 6411 6137 6423 6140
rect 6365 6131 6423 6137
rect 16666 6128 16672 6140
rect 16724 6128 16730 6180
rect 4062 6100 4068 6112
rect 4023 6072 4068 6100
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 5442 6060 5448 6112
rect 5500 6100 5506 6112
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 5500 6072 6653 6100
rect 5500 6060 5506 6072
rect 6641 6069 6653 6072
rect 6687 6069 6699 6103
rect 6641 6063 6699 6069
rect 920 6010 7084 6032
rect 920 5958 3598 6010
rect 3650 5958 3662 6010
rect 3714 5958 3726 6010
rect 3778 5958 3790 6010
rect 3842 5958 7084 6010
rect 920 5936 7084 5958
rect 3234 5896 3240 5908
rect 1504 5868 3240 5896
rect 1504 5837 1532 5868
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 6086 5896 6092 5908
rect 6047 5868 6092 5896
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 1489 5831 1547 5837
rect 1489 5797 1501 5831
rect 1535 5797 1547 5831
rect 1489 5791 1547 5797
rect 1946 5788 1952 5840
rect 2004 5788 2010 5840
rect 4062 5788 4068 5840
rect 4120 5788 4126 5840
rect 4890 5720 4896 5772
rect 4948 5760 4954 5772
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 4948 5732 5549 5760
rect 4948 5720 4954 5732
rect 5537 5729 5549 5732
rect 5583 5760 5595 5763
rect 5902 5760 5908 5772
rect 5583 5732 5908 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 5902 5720 5908 5732
rect 5960 5720 5966 5772
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 6362 5760 6368 5772
rect 6319 5732 6368 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 6362 5720 6368 5732
rect 6420 5720 6426 5772
rect 1210 5692 1216 5704
rect 1171 5664 1216 5692
rect 1210 5652 1216 5664
rect 1268 5652 1274 5704
rect 3234 5692 3240 5704
rect 3195 5664 3240 5692
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 3329 5695 3387 5701
rect 3329 5661 3341 5695
rect 3375 5692 3387 5695
rect 3602 5692 3608 5704
rect 3375 5664 3464 5692
rect 3515 5664 3608 5692
rect 3375 5661 3387 5664
rect 3329 5655 3387 5661
rect 3436 5568 3464 5664
rect 3602 5652 3608 5664
rect 3660 5692 3666 5704
rect 3970 5692 3976 5704
rect 3660 5664 3976 5692
rect 3660 5652 3666 5664
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 5353 5695 5411 5701
rect 5353 5692 5365 5695
rect 4212 5664 5365 5692
rect 4212 5652 4218 5664
rect 5353 5661 5365 5664
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 3418 5516 3424 5568
rect 3476 5516 3482 5568
rect 5718 5556 5724 5568
rect 5679 5528 5724 5556
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 6178 5516 6184 5568
rect 6236 5556 6242 5568
rect 6365 5559 6423 5565
rect 6365 5556 6377 5559
rect 6236 5528 6377 5556
rect 6236 5516 6242 5528
rect 6365 5525 6377 5528
rect 6411 5525 6423 5559
rect 6365 5519 6423 5525
rect 920 5466 7084 5488
rect 920 5414 2098 5466
rect 2150 5414 2162 5466
rect 2214 5414 2226 5466
rect 2278 5414 2290 5466
rect 2342 5414 5098 5466
rect 5150 5414 5162 5466
rect 5214 5414 5226 5466
rect 5278 5414 5290 5466
rect 5342 5414 7084 5466
rect 920 5392 7084 5414
rect 4157 5355 4215 5361
rect 4157 5321 4169 5355
rect 4203 5352 4215 5355
rect 4614 5352 4620 5364
rect 4203 5324 4620 5352
rect 4203 5321 4215 5324
rect 4157 5315 4215 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 6270 5284 6276 5296
rect 6196 5256 6276 5284
rect 1489 5219 1547 5225
rect 1489 5185 1501 5219
rect 1535 5216 1547 5219
rect 2774 5216 2780 5228
rect 1535 5188 2780 5216
rect 1535 5185 1547 5188
rect 1489 5179 1547 5185
rect 2774 5176 2780 5188
rect 2832 5216 2838 5228
rect 3234 5216 3240 5228
rect 2832 5188 3240 5216
rect 2832 5176 2838 5188
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 4246 5176 4252 5228
rect 4304 5216 4310 5228
rect 4522 5216 4528 5228
rect 4304 5188 4528 5216
rect 4304 5176 4310 5188
rect 4522 5176 4528 5188
rect 4580 5216 4586 5228
rect 4617 5219 4675 5225
rect 4617 5216 4629 5219
rect 4580 5188 4629 5216
rect 4580 5176 4586 5188
rect 4617 5185 4629 5188
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 6196 5216 6224 5256
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 6362 5216 6368 5228
rect 5031 5188 6224 5216
rect 6323 5188 6368 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 6362 5176 6368 5188
rect 6420 5176 6426 5228
rect 1210 5148 1216 5160
rect 1171 5120 1216 5148
rect 1210 5108 1216 5120
rect 1268 5108 1274 5160
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 3329 5151 3387 5157
rect 3329 5148 3341 5151
rect 3108 5120 3341 5148
rect 3108 5108 3114 5120
rect 3329 5117 3341 5120
rect 3375 5117 3387 5151
rect 3878 5148 3884 5160
rect 3329 5111 3387 5117
rect 3528 5120 3884 5148
rect 1946 5040 1952 5092
rect 2004 5040 2010 5092
rect 3234 5080 3240 5092
rect 3195 5052 3240 5080
rect 3234 5040 3240 5052
rect 3292 5040 3298 5092
rect 2958 4972 2964 5024
rect 3016 5012 3022 5024
rect 3528 5021 3556 5120
rect 3878 5108 3884 5120
rect 3936 5148 3942 5160
rect 3973 5151 4031 5157
rect 3973 5148 3985 5151
rect 3936 5120 3985 5148
rect 3936 5108 3942 5120
rect 3973 5117 3985 5120
rect 4019 5117 4031 5151
rect 3973 5111 4031 5117
rect 5718 5040 5724 5092
rect 5776 5040 5782 5092
rect 3513 5015 3571 5021
rect 3513 5012 3525 5015
rect 3016 4984 3525 5012
rect 3016 4972 3022 4984
rect 3513 4981 3525 4984
rect 3559 4981 3571 5015
rect 3513 4975 3571 4981
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 16574 5012 16580 5024
rect 6420 4984 16580 5012
rect 6420 4972 6426 4984
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 920 4922 7084 4944
rect 920 4870 3598 4922
rect 3650 4870 3662 4922
rect 3714 4870 3726 4922
rect 3778 4870 3790 4922
rect 3842 4870 7084 4922
rect 920 4848 7084 4870
rect 1673 4811 1731 4817
rect 1673 4777 1685 4811
rect 1719 4808 1731 4811
rect 1946 4808 1952 4820
rect 1719 4780 1952 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2406 4808 2412 4820
rect 2056 4780 2412 4808
rect 2056 4740 2084 4780
rect 2406 4768 2412 4780
rect 2464 4808 2470 4820
rect 5997 4811 6055 4817
rect 5997 4808 6009 4811
rect 2464 4780 6009 4808
rect 2464 4768 2470 4780
rect 5997 4777 6009 4780
rect 6043 4777 6055 4811
rect 5997 4771 6055 4777
rect 2958 4740 2964 4752
rect 1320 4712 2084 4740
rect 2240 4712 2964 4740
rect 1320 4672 1348 4712
rect 1397 4675 1455 4681
rect 1397 4672 1409 4675
rect 1320 4644 1409 4672
rect 1397 4641 1409 4644
rect 1443 4641 1455 4675
rect 1397 4635 1455 4641
rect 1514 4675 1572 4681
rect 1514 4641 1526 4675
rect 1560 4672 1572 4675
rect 1762 4672 1768 4684
rect 1560 4644 1768 4672
rect 1560 4641 1572 4644
rect 1514 4635 1572 4641
rect 1762 4632 1768 4644
rect 1820 4632 1826 4684
rect 2240 4681 2268 4712
rect 2958 4700 2964 4712
rect 3016 4700 3022 4752
rect 3510 4700 3516 4752
rect 3568 4700 3574 4752
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 2225 4675 2283 4681
rect 2225 4672 2237 4675
rect 1903 4644 2237 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 2225 4641 2237 4644
rect 2271 4641 2283 4675
rect 2590 4672 2596 4684
rect 2551 4644 2596 4672
rect 2225 4635 2283 4641
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 4709 4675 4767 4681
rect 4709 4641 4721 4675
rect 4755 4672 4767 4675
rect 26418 4672 26424 4684
rect 4755 4644 26424 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 26418 4632 26424 4644
rect 26476 4632 26482 4684
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2700 4576 2881 4604
rect 1486 4496 1492 4548
rect 1544 4536 1550 4548
rect 2700 4536 2728 4576
rect 2869 4573 2881 4576
rect 2915 4604 2927 4607
rect 3234 4604 3240 4616
rect 2915 4576 3240 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4604 4675 4607
rect 5442 4604 5448 4616
rect 4663 4576 5448 4604
rect 4663 4573 4675 4576
rect 4617 4567 4675 4573
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 1544 4508 2728 4536
rect 1544 4496 1550 4508
rect 1210 4468 1216 4480
rect 1171 4440 1216 4468
rect 1210 4428 1216 4440
rect 1268 4428 1274 4480
rect 1946 4428 1952 4480
rect 2004 4468 2010 4480
rect 2041 4471 2099 4477
rect 2041 4468 2053 4471
rect 2004 4440 2053 4468
rect 2004 4428 2010 4440
rect 2041 4437 2053 4440
rect 2087 4437 2099 4471
rect 2041 4431 2099 4437
rect 2409 4471 2467 4477
rect 2409 4437 2421 4471
rect 2455 4468 2467 4471
rect 2866 4468 2872 4480
rect 2455 4440 2872 4468
rect 2455 4437 2467 4440
rect 2409 4431 2467 4437
rect 2866 4428 2872 4440
rect 2924 4428 2930 4480
rect 920 4378 7084 4400
rect 920 4326 2098 4378
rect 2150 4326 2162 4378
rect 2214 4326 2226 4378
rect 2278 4326 2290 4378
rect 2342 4326 5098 4378
rect 5150 4326 5162 4378
rect 5214 4326 5226 4378
rect 5278 4326 5290 4378
rect 5342 4326 7084 4378
rect 920 4304 7084 4326
rect 3510 4264 3516 4276
rect 3471 4236 3516 4264
rect 3510 4224 3516 4236
rect 3568 4224 3574 4276
rect 3970 4224 3976 4276
rect 4028 4224 4034 4276
rect 1486 4128 1492 4140
rect 1447 4100 1492 4128
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 3418 4128 3424 4140
rect 2792 4100 3424 4128
rect 1210 4060 1216 4072
rect 1171 4032 1216 4060
rect 1210 4020 1216 4032
rect 1268 4020 1274 4072
rect 1946 3952 1952 4004
rect 2004 3952 2010 4004
rect 1210 3884 1216 3936
rect 1268 3924 1274 3936
rect 2792 3924 2820 4100
rect 3418 4088 3424 4100
rect 3476 4128 3482 4140
rect 3881 4131 3939 4137
rect 3881 4128 3893 4131
rect 3476 4100 3893 4128
rect 3476 4088 3482 4100
rect 3881 4097 3893 4100
rect 3927 4097 3939 4131
rect 3988 4128 4016 4224
rect 6362 4196 6368 4208
rect 6196 4168 6368 4196
rect 5994 4128 6000 4140
rect 3988 4100 5396 4128
rect 5955 4100 6000 4128
rect 3881 4091 3939 4097
rect 3326 4060 3332 4072
rect 3287 4032 3332 4060
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 5368 4060 5396 4100
rect 5994 4088 6000 4100
rect 6052 4128 6058 4140
rect 6196 4128 6224 4168
rect 6362 4156 6368 4168
rect 6420 4156 6426 4208
rect 6638 4128 6644 4140
rect 6052 4100 6224 4128
rect 6288 4100 6644 4128
rect 6052 4088 6058 4100
rect 5905 4063 5963 4069
rect 5905 4060 5917 4063
rect 5368 4032 5917 4060
rect 5905 4029 5917 4032
rect 5951 4029 5963 4063
rect 6178 4060 6184 4072
rect 6139 4032 6184 4060
rect 5905 4023 5963 4029
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 6288 4069 6316 4100
rect 6638 4088 6644 4100
rect 6696 4128 6702 4140
rect 16666 4128 16672 4140
rect 6696 4100 16672 4128
rect 6696 4088 6702 4100
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 6273 4063 6331 4069
rect 6273 4029 6285 4063
rect 6319 4029 6331 4063
rect 6273 4023 6331 4029
rect 6362 4020 6368 4072
rect 6420 4060 6426 4072
rect 16850 4060 16856 4072
rect 6420 4032 16856 4060
rect 6420 4020 6426 4032
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 3234 3992 3240 4004
rect 3195 3964 3240 3992
rect 3234 3952 3240 3964
rect 3292 3992 3298 4004
rect 4157 3995 4215 4001
rect 4157 3992 4169 3995
rect 3292 3964 4169 3992
rect 3292 3952 3298 3964
rect 4157 3961 4169 3964
rect 4203 3961 4215 3995
rect 4157 3955 4215 3961
rect 1268 3896 2820 3924
rect 1268 3884 1274 3896
rect 2866 3884 2872 3936
rect 2924 3924 2930 3936
rect 4632 3924 4660 3978
rect 6086 3952 6092 4004
rect 6144 3992 6150 4004
rect 6733 3995 6791 4001
rect 6733 3992 6745 3995
rect 6144 3964 6745 3992
rect 6144 3952 6150 3964
rect 6733 3961 6745 3964
rect 6779 3961 6791 3995
rect 6733 3955 6791 3961
rect 2924 3896 4660 3924
rect 2924 3884 2930 3896
rect 5442 3884 5448 3936
rect 5500 3924 5506 3936
rect 16574 3924 16580 3936
rect 5500 3896 16580 3924
rect 5500 3884 5506 3896
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 920 3834 7084 3856
rect 920 3782 3598 3834
rect 3650 3782 3662 3834
rect 3714 3782 3726 3834
rect 3778 3782 3790 3834
rect 3842 3782 7084 3834
rect 920 3760 7084 3782
rect 2682 3680 2688 3732
rect 2740 3720 2746 3732
rect 5810 3720 5816 3732
rect 2740 3692 5816 3720
rect 2740 3680 2746 3692
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 2869 3655 2927 3661
rect 2869 3652 2881 3655
rect 2832 3624 2881 3652
rect 2832 3612 2838 3624
rect 2869 3621 2881 3624
rect 2915 3621 2927 3655
rect 2869 3615 2927 3621
rect 5077 3655 5135 3661
rect 5077 3621 5089 3655
rect 5123 3652 5135 3655
rect 5123 3624 6040 3652
rect 5123 3621 5135 3624
rect 5077 3615 5135 3621
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3553 2283 3587
rect 2590 3584 2596 3596
rect 2551 3556 2596 3584
rect 2225 3547 2283 3553
rect 2240 3448 2268 3547
rect 2590 3544 2596 3556
rect 2648 3544 2654 3596
rect 3970 3544 3976 3596
rect 4028 3544 4034 3596
rect 4709 3587 4767 3593
rect 4709 3584 4721 3587
rect 4540 3556 4721 3584
rect 4540 3516 4568 3556
rect 4709 3553 4721 3556
rect 4755 3584 4767 3587
rect 4890 3584 4896 3596
rect 4755 3556 4896 3584
rect 4755 3553 4767 3556
rect 4709 3547 4767 3553
rect 4890 3544 4896 3556
rect 4948 3544 4954 3596
rect 4982 3544 4988 3596
rect 5040 3584 5046 3596
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 5040 3556 5273 3584
rect 5040 3544 5046 3556
rect 5261 3553 5273 3556
rect 5307 3553 5319 3587
rect 5626 3584 5632 3596
rect 5587 3556 5632 3584
rect 5261 3547 5319 3553
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 6012 3593 6040 3624
rect 5997 3587 6055 3593
rect 5997 3553 6009 3587
rect 6043 3584 6055 3587
rect 6086 3584 6092 3596
rect 6043 3556 6092 3584
rect 6043 3553 6055 3556
rect 5997 3547 6055 3553
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3584 6515 3587
rect 6546 3584 6552 3596
rect 6503 3556 6552 3584
rect 6503 3553 6515 3556
rect 6457 3547 6515 3553
rect 6546 3544 6552 3556
rect 6604 3584 6610 3596
rect 16758 3584 16764 3596
rect 6604 3556 16764 3584
rect 6604 3544 6610 3556
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 2700 3488 4568 3516
rect 4617 3519 4675 3525
rect 2700 3448 2728 3488
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 16666 3516 16672 3528
rect 4663 3488 16672 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 2240 3420 2728 3448
rect 4893 3451 4951 3457
rect 4893 3417 4905 3451
rect 4939 3448 4951 3451
rect 5442 3448 5448 3460
rect 4939 3420 5448 3448
rect 4939 3417 4951 3420
rect 4893 3411 4951 3417
rect 5442 3408 5448 3420
rect 5500 3408 5506 3460
rect 5810 3448 5816 3460
rect 5771 3420 5816 3448
rect 5810 3408 5816 3420
rect 5868 3408 5874 3460
rect 2409 3383 2467 3389
rect 2409 3349 2421 3383
rect 2455 3380 2467 3383
rect 5534 3380 5540 3392
rect 2455 3352 5540 3380
rect 2455 3349 2467 3352
rect 2409 3343 2467 3349
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 920 3290 7084 3312
rect 920 3238 2098 3290
rect 2150 3238 2162 3290
rect 2214 3238 2226 3290
rect 2278 3238 2290 3290
rect 2342 3238 5098 3290
rect 5150 3238 5162 3290
rect 5214 3238 5226 3290
rect 5278 3238 5290 3290
rect 5342 3238 7084 3290
rect 920 3216 7084 3238
rect 2590 3176 2596 3188
rect 1688 3148 2596 3176
rect 1688 3049 1716 3148
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 4890 3176 4896 3188
rect 4488 3148 4896 3176
rect 4488 3136 4494 3148
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 6638 3176 6644 3188
rect 6599 3148 6644 3176
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3040 2007 3043
rect 3234 3040 3240 3052
rect 1995 3012 3240 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 16574 3040 16580 3052
rect 3743 3012 16580 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 3326 2932 3332 2984
rect 3384 2972 3390 2984
rect 3878 2972 3884 2984
rect 3384 2944 3884 2972
rect 3384 2932 3390 2944
rect 3878 2932 3884 2944
rect 3936 2932 3942 2984
rect 4430 2972 4436 2984
rect 4391 2944 4436 2972
rect 4430 2932 4436 2944
rect 4488 2932 4494 2984
rect 4522 2932 4528 2984
rect 4580 2972 4586 2984
rect 4890 2972 4896 2984
rect 4580 2944 4625 2972
rect 4851 2944 4896 2972
rect 4580 2932 4586 2944
rect 4890 2932 4896 2944
rect 4948 2932 4954 2984
rect 3160 2836 3188 2890
rect 5442 2864 5448 2916
rect 5500 2864 5506 2916
rect 4065 2839 4123 2845
rect 4065 2836 4077 2839
rect 3160 2808 4077 2836
rect 4065 2805 4077 2808
rect 4111 2805 4123 2839
rect 4246 2836 4252 2848
rect 4207 2808 4252 2836
rect 4065 2799 4123 2805
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 920 2746 7084 2768
rect 920 2694 3598 2746
rect 3650 2694 3662 2746
rect 3714 2694 3726 2746
rect 3778 2694 3790 2746
rect 3842 2694 7084 2746
rect 920 2672 7084 2694
rect 3970 2592 3976 2644
rect 4028 2632 4034 2644
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 4028 2604 4077 2632
rect 4028 2592 4034 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 4065 2595 4123 2601
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 16574 2632 16580 2644
rect 5040 2604 16580 2632
rect 5040 2592 5046 2604
rect 16574 2592 16580 2604
rect 16632 2592 16638 2644
rect 2958 2524 2964 2576
rect 3016 2524 3022 2576
rect 3697 2567 3755 2573
rect 3697 2533 3709 2567
rect 3743 2564 3755 2567
rect 4338 2564 4344 2576
rect 3743 2536 4344 2564
rect 3743 2533 3755 2536
rect 3697 2527 3755 2533
rect 4338 2524 4344 2536
rect 4396 2524 4402 2576
rect 4798 2564 4804 2576
rect 4759 2536 4804 2564
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 5534 2524 5540 2576
rect 5592 2524 5598 2576
rect 6546 2564 6552 2576
rect 6507 2536 6552 2564
rect 6546 2524 6552 2536
rect 6604 2524 6610 2576
rect 1210 2456 1216 2508
rect 1268 2496 1274 2508
rect 1673 2499 1731 2505
rect 1673 2496 1685 2499
rect 1268 2468 1685 2496
rect 1268 2456 1274 2468
rect 1673 2465 1685 2468
rect 1719 2465 1731 2499
rect 3878 2496 3884 2508
rect 3839 2468 3884 2496
rect 1673 2459 1731 2465
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 4522 2496 4528 2508
rect 4483 2468 4528 2496
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 4798 2428 4804 2440
rect 1995 2400 4804 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 920 2202 7084 2224
rect 920 2150 2098 2202
rect 2150 2150 2162 2202
rect 2214 2150 2226 2202
rect 2278 2150 2290 2202
rect 2342 2150 5098 2202
rect 5150 2150 5162 2202
rect 5214 2150 5226 2202
rect 5278 2150 5290 2202
rect 5342 2150 7084 2202
rect 920 2128 7084 2150
rect 4246 1300 4252 1352
rect 4304 1340 4310 1352
rect 16666 1340 16672 1352
rect 4304 1312 16672 1340
rect 4304 1300 4310 1312
rect 16666 1300 16672 1312
rect 16724 1300 16730 1352
rect 4430 1232 4436 1284
rect 4488 1272 4494 1284
rect 16758 1272 16764 1284
rect 4488 1244 16764 1272
rect 4488 1232 4494 1244
rect 16758 1232 16764 1244
rect 16816 1232 16822 1284
rect 6454 1164 6460 1216
rect 6512 1204 6518 1216
rect 16574 1204 16580 1216
rect 6512 1176 16580 1204
rect 6512 1164 6518 1176
rect 16574 1164 16580 1176
rect 16632 1164 16638 1216
<< via1 >>
rect 6368 12520 6420 12572
rect 16580 12520 16632 12572
rect 3976 12452 4028 12504
rect 16672 12452 16724 12504
rect -1606 11386 -1318 11464
rect 3598 11398 3650 11450
rect 3662 11398 3714 11450
rect 3726 11398 3778 11450
rect 3790 11398 3842 11450
rect 3884 11160 3936 11212
rect 4712 11203 4764 11212
rect 4712 11169 4721 11203
rect 4721 11169 4755 11203
rect 4755 11169 4764 11203
rect 4712 11160 4764 11169
rect 5632 11203 5684 11212
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 5908 11203 5960 11212
rect 4988 11092 5040 11144
rect 5448 11092 5500 11144
rect 5908 11169 5917 11203
rect 5917 11169 5951 11203
rect 5951 11169 5960 11203
rect 5908 11160 5960 11169
rect 6368 11203 6420 11212
rect 6368 11169 6377 11203
rect 6377 11169 6411 11203
rect 6411 11169 6420 11203
rect 6368 11160 6420 11169
rect 6184 11092 6236 11144
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 1768 11024 1820 11076
rect 16580 11024 16632 11076
rect 3056 10999 3108 11008
rect 3056 10965 3065 10999
rect 3065 10965 3099 10999
rect 3099 10965 3108 10999
rect 3056 10956 3108 10965
rect 4528 10956 4580 11008
rect -948 10844 -658 10918
rect 2098 10854 2150 10906
rect 2162 10854 2214 10906
rect 2226 10854 2278 10906
rect 2290 10854 2342 10906
rect 5098 10854 5150 10906
rect 5162 10854 5214 10906
rect 5226 10854 5278 10906
rect 5290 10854 5342 10906
rect 4436 10752 4488 10804
rect 4620 10616 4672 10668
rect 4988 10616 5040 10668
rect 16764 10616 16816 10668
rect 1492 10548 1544 10600
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 4528 10591 4580 10600
rect 4528 10557 4537 10591
rect 4537 10557 4571 10591
rect 4571 10557 4580 10591
rect 6552 10591 6604 10600
rect 4528 10548 4580 10557
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 1952 10523 2004 10532
rect 1952 10489 1961 10523
rect 1961 10489 1995 10523
rect 1995 10489 2004 10523
rect 1952 10480 2004 10489
rect 4344 10480 4396 10532
rect 4712 10412 4764 10464
rect 16580 10412 16632 10464
rect 3598 10310 3650 10362
rect 3662 10310 3714 10362
rect 3726 10310 3778 10362
rect 3790 10310 3842 10362
rect 1952 10208 2004 10260
rect 1768 10183 1820 10192
rect 1768 10149 1777 10183
rect 1777 10149 1811 10183
rect 1811 10149 1820 10183
rect 1768 10140 1820 10149
rect 3056 10140 3108 10192
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 4436 10004 4488 10056
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 6000 9911 6052 9920
rect 6000 9877 6009 9911
rect 6009 9877 6043 9911
rect 6043 9877 6052 9911
rect 6000 9868 6052 9877
rect 2098 9766 2150 9818
rect 2162 9766 2214 9818
rect 2226 9766 2278 9818
rect 2290 9766 2342 9818
rect 5098 9766 5150 9818
rect 5162 9766 5214 9818
rect 5226 9766 5278 9818
rect 5290 9766 5342 9818
rect 2872 9596 2924 9648
rect 5816 9664 5868 9716
rect 6552 9664 6604 9716
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 2964 9503 3016 9512
rect 2964 9469 2973 9503
rect 2973 9469 3007 9503
rect 3007 9469 3016 9503
rect 2964 9460 3016 9469
rect 3976 9528 4028 9580
rect 4436 9571 4488 9580
rect 4436 9537 4445 9571
rect 4445 9537 4479 9571
rect 4479 9537 4488 9571
rect 4436 9528 4488 9537
rect 5724 9528 5776 9580
rect 4068 9503 4120 9512
rect 2504 9392 2556 9444
rect 4068 9469 4077 9503
rect 4077 9469 4111 9503
rect 4111 9469 4120 9503
rect 4068 9460 4120 9469
rect 6552 9503 6604 9512
rect 6552 9469 6561 9503
rect 6561 9469 6595 9503
rect 6595 9469 6604 9503
rect 6552 9460 6604 9469
rect 4160 9392 4212 9444
rect 6000 9392 6052 9444
rect 26240 9392 26292 9444
rect 6368 9324 6420 9376
rect 3598 9222 3650 9274
rect 3662 9222 3714 9274
rect 3726 9222 3778 9274
rect 3790 9222 3842 9274
rect 3148 9120 3200 9172
rect 3424 9120 3476 9172
rect 4068 9120 4120 9172
rect 6460 9120 6512 9172
rect 3332 9052 3384 9104
rect 4712 9052 4764 9104
rect 5448 9052 5500 9104
rect 16580 9052 16632 9104
rect 1768 8984 1820 9036
rect 2412 8984 2464 9036
rect 2872 8984 2924 9036
rect 4620 8984 4672 9036
rect 5724 8984 5776 9036
rect 4436 8916 4488 8968
rect 16672 8916 16724 8968
rect 1216 8848 1268 8900
rect 1492 8848 1544 8900
rect 1952 8780 2004 8832
rect 2964 8780 3016 8832
rect 5632 8780 5684 8832
rect 2098 8678 2150 8730
rect 2162 8678 2214 8730
rect 2226 8678 2278 8730
rect 2290 8678 2342 8730
rect 5098 8678 5150 8730
rect 5162 8678 5214 8730
rect 5226 8678 5278 8730
rect 5290 8678 5342 8730
rect 3148 8508 3200 8560
rect 3884 8508 3936 8560
rect 4804 8576 4856 8628
rect 4344 8508 4396 8560
rect 1216 8415 1268 8424
rect 1216 8381 1225 8415
rect 1225 8381 1259 8415
rect 1259 8381 1268 8415
rect 1216 8372 1268 8381
rect 3332 8415 3384 8424
rect 3332 8381 3341 8415
rect 3341 8381 3375 8415
rect 3375 8381 3384 8415
rect 3332 8372 3384 8381
rect 4068 8372 4120 8424
rect 4620 8440 4672 8492
rect 5816 8440 5868 8492
rect 1952 8304 2004 8356
rect 3240 8347 3292 8356
rect 3240 8313 3249 8347
rect 3249 8313 3283 8347
rect 3283 8313 3292 8347
rect 3240 8304 3292 8313
rect 3884 8304 3936 8356
rect 4528 8304 4580 8356
rect 4712 8304 4764 8356
rect 6368 8347 6420 8356
rect 6368 8313 6377 8347
rect 6377 8313 6411 8347
rect 6411 8313 6420 8347
rect 6368 8304 6420 8313
rect 26332 8304 26384 8356
rect 2504 8236 2556 8288
rect 16580 8236 16632 8288
rect 3598 8134 3650 8186
rect 3662 8134 3714 8186
rect 3726 8134 3778 8186
rect 3790 8134 3842 8186
rect 3240 8032 3292 8084
rect 4804 8032 4856 8084
rect 5448 7964 5500 8016
rect 1952 7896 2004 7948
rect 3056 7828 3108 7880
rect 3332 7828 3384 7880
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 1768 7692 1820 7744
rect 1952 7692 2004 7744
rect 2964 7692 3016 7744
rect 4436 7896 4488 7948
rect 4344 7828 4396 7880
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 6276 7692 6328 7744
rect 6552 7692 6604 7744
rect 16672 7692 16724 7744
rect 2098 7590 2150 7642
rect 2162 7590 2214 7642
rect 2226 7590 2278 7642
rect 2290 7590 2342 7642
rect 5098 7590 5150 7642
rect 5162 7590 5214 7642
rect 5226 7590 5278 7642
rect 5290 7590 5342 7642
rect 1216 7488 1268 7540
rect 3148 7488 3200 7540
rect 3332 7488 3384 7540
rect 3240 7352 3292 7404
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 4160 7395 4212 7404
rect 4160 7361 4169 7395
rect 4169 7361 4203 7395
rect 4203 7361 4212 7395
rect 4160 7352 4212 7361
rect 4804 7352 4856 7404
rect 2872 7284 2924 7336
rect 1492 7216 1544 7268
rect 3240 7259 3292 7268
rect 3240 7225 3249 7259
rect 3249 7225 3283 7259
rect 3283 7225 3292 7259
rect 3240 7216 3292 7225
rect 4620 7216 4672 7268
rect 3976 7148 4028 7200
rect 5540 7148 5592 7200
rect 16580 7284 16632 7336
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 6552 7148 6604 7157
rect 3598 7046 3650 7098
rect 3662 7046 3714 7098
rect 3726 7046 3778 7098
rect 3790 7046 3842 7098
rect 2596 6876 2648 6928
rect 1768 6808 1820 6860
rect 3976 6876 4028 6928
rect 6552 6876 6604 6928
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 3608 6740 3660 6792
rect 5540 6740 5592 6792
rect 6276 6740 6328 6792
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 1952 6604 2004 6656
rect 2504 6604 2556 6656
rect 3976 6604 4028 6656
rect 5724 6672 5776 6724
rect 4896 6604 4948 6656
rect 2098 6502 2150 6554
rect 2162 6502 2214 6554
rect 2226 6502 2278 6554
rect 2290 6502 2342 6554
rect 5098 6502 5150 6554
rect 5162 6502 5214 6554
rect 5226 6502 5278 6554
rect 5290 6502 5342 6554
rect 4712 6400 4764 6452
rect 5724 6400 5776 6452
rect 16580 6400 16632 6452
rect 3240 6264 3292 6316
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 1216 6239 1268 6248
rect 1216 6205 1225 6239
rect 1225 6205 1259 6239
rect 1259 6205 1268 6239
rect 1216 6196 1268 6205
rect 3056 6196 3108 6248
rect 3608 6196 3660 6248
rect 3884 6239 3936 6248
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 5908 6196 5960 6248
rect 2504 6128 2556 6180
rect 3240 6171 3292 6180
rect 3240 6137 3249 6171
rect 3249 6137 3283 6171
rect 3283 6137 3292 6171
rect 3240 6128 3292 6137
rect 6092 6128 6144 6180
rect 16672 6128 16724 6180
rect 4068 6103 4120 6112
rect 4068 6069 4077 6103
rect 4077 6069 4111 6103
rect 4111 6069 4120 6103
rect 4068 6060 4120 6069
rect 5448 6060 5500 6112
rect 3598 5958 3650 6010
rect 3662 5958 3714 6010
rect 3726 5958 3778 6010
rect 3790 5958 3842 6010
rect 3240 5856 3292 5908
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 1952 5788 2004 5840
rect 4068 5788 4120 5840
rect 4896 5720 4948 5772
rect 5908 5763 5960 5772
rect 5908 5729 5917 5763
rect 5917 5729 5951 5763
rect 5951 5729 5960 5763
rect 5908 5720 5960 5729
rect 6368 5720 6420 5772
rect 1216 5695 1268 5704
rect 1216 5661 1225 5695
rect 1225 5661 1259 5695
rect 1259 5661 1268 5695
rect 1216 5652 1268 5661
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 3608 5695 3660 5704
rect 3608 5661 3617 5695
rect 3617 5661 3651 5695
rect 3651 5661 3660 5695
rect 3608 5652 3660 5661
rect 3976 5652 4028 5704
rect 4160 5652 4212 5704
rect 3424 5516 3476 5568
rect 5724 5559 5776 5568
rect 5724 5525 5733 5559
rect 5733 5525 5767 5559
rect 5767 5525 5776 5559
rect 5724 5516 5776 5525
rect 6184 5516 6236 5568
rect 2098 5414 2150 5466
rect 2162 5414 2214 5466
rect 2226 5414 2278 5466
rect 2290 5414 2342 5466
rect 5098 5414 5150 5466
rect 5162 5414 5214 5466
rect 5226 5414 5278 5466
rect 5290 5414 5342 5466
rect 4620 5312 4672 5364
rect 2780 5176 2832 5228
rect 3240 5176 3292 5228
rect 4252 5176 4304 5228
rect 4528 5176 4580 5228
rect 6276 5244 6328 5296
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 1216 5151 1268 5160
rect 1216 5117 1225 5151
rect 1225 5117 1259 5151
rect 1259 5117 1268 5151
rect 1216 5108 1268 5117
rect 3056 5108 3108 5160
rect 1952 5040 2004 5092
rect 3240 5083 3292 5092
rect 3240 5049 3249 5083
rect 3249 5049 3283 5083
rect 3283 5049 3292 5083
rect 3240 5040 3292 5049
rect 2964 4972 3016 5024
rect 3884 5108 3936 5160
rect 5724 5040 5776 5092
rect 6368 4972 6420 5024
rect 16580 4972 16632 5024
rect 3598 4870 3650 4922
rect 3662 4870 3714 4922
rect 3726 4870 3778 4922
rect 3790 4870 3842 4922
rect 1952 4768 2004 4820
rect 2412 4768 2464 4820
rect 1768 4632 1820 4684
rect 2964 4700 3016 4752
rect 3516 4700 3568 4752
rect 2596 4675 2648 4684
rect 2596 4641 2605 4675
rect 2605 4641 2639 4675
rect 2639 4641 2648 4675
rect 2596 4632 2648 4641
rect 26424 4632 26476 4684
rect 1492 4496 1544 4548
rect 3240 4564 3292 4616
rect 5448 4564 5500 4616
rect 1216 4471 1268 4480
rect 1216 4437 1225 4471
rect 1225 4437 1259 4471
rect 1259 4437 1268 4471
rect 1216 4428 1268 4437
rect 1952 4428 2004 4480
rect 2872 4428 2924 4480
rect 2098 4326 2150 4378
rect 2162 4326 2214 4378
rect 2226 4326 2278 4378
rect 2290 4326 2342 4378
rect 5098 4326 5150 4378
rect 5162 4326 5214 4378
rect 5226 4326 5278 4378
rect 5290 4326 5342 4378
rect 3516 4267 3568 4276
rect 3516 4233 3525 4267
rect 3525 4233 3559 4267
rect 3559 4233 3568 4267
rect 3516 4224 3568 4233
rect 3976 4224 4028 4276
rect 1492 4131 1544 4140
rect 1492 4097 1501 4131
rect 1501 4097 1535 4131
rect 1535 4097 1544 4131
rect 1492 4088 1544 4097
rect 1216 4063 1268 4072
rect 1216 4029 1225 4063
rect 1225 4029 1259 4063
rect 1259 4029 1268 4063
rect 1216 4020 1268 4029
rect 1952 3952 2004 4004
rect 1216 3884 1268 3936
rect 3424 4088 3476 4140
rect 6000 4131 6052 4140
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6368 4156 6420 4208
rect 6000 4088 6052 4097
rect 6184 4063 6236 4072
rect 6184 4029 6193 4063
rect 6193 4029 6227 4063
rect 6227 4029 6236 4063
rect 6184 4020 6236 4029
rect 6644 4088 6696 4140
rect 16672 4088 16724 4140
rect 6368 4020 6420 4072
rect 16856 4020 16908 4072
rect 3240 3995 3292 4004
rect 3240 3961 3249 3995
rect 3249 3961 3283 3995
rect 3283 3961 3292 3995
rect 3240 3952 3292 3961
rect 2872 3884 2924 3936
rect 6092 3952 6144 4004
rect 5448 3884 5500 3936
rect 16580 3884 16632 3936
rect 3598 3782 3650 3834
rect 3662 3782 3714 3834
rect 3726 3782 3778 3834
rect 3790 3782 3842 3834
rect 2688 3680 2740 3732
rect 5816 3680 5868 3732
rect 2780 3612 2832 3664
rect 2596 3587 2648 3596
rect 2596 3553 2605 3587
rect 2605 3553 2639 3587
rect 2639 3553 2648 3587
rect 2596 3544 2648 3553
rect 3976 3544 4028 3596
rect 4896 3544 4948 3596
rect 4988 3544 5040 3596
rect 5632 3587 5684 3596
rect 5632 3553 5641 3587
rect 5641 3553 5675 3587
rect 5675 3553 5684 3587
rect 5632 3544 5684 3553
rect 6092 3544 6144 3596
rect 6552 3544 6604 3596
rect 16764 3544 16816 3596
rect 16672 3476 16724 3528
rect 5448 3408 5500 3460
rect 5816 3451 5868 3460
rect 5816 3417 5825 3451
rect 5825 3417 5859 3451
rect 5859 3417 5868 3451
rect 5816 3408 5868 3417
rect 5540 3340 5592 3392
rect 2098 3238 2150 3290
rect 2162 3238 2214 3290
rect 2226 3238 2278 3290
rect 2290 3238 2342 3290
rect 5098 3238 5150 3290
rect 5162 3238 5214 3290
rect 5226 3238 5278 3290
rect 5290 3238 5342 3290
rect 2596 3136 2648 3188
rect 4436 3136 4488 3188
rect 4896 3136 4948 3188
rect 6644 3179 6696 3188
rect 6644 3145 6653 3179
rect 6653 3145 6687 3179
rect 6687 3145 6696 3179
rect 6644 3136 6696 3145
rect 3240 3000 3292 3052
rect 16580 3000 16632 3052
rect 3332 2932 3384 2984
rect 3884 2975 3936 2984
rect 3884 2941 3893 2975
rect 3893 2941 3927 2975
rect 3927 2941 3936 2975
rect 3884 2932 3936 2941
rect 4436 2975 4488 2984
rect 4436 2941 4445 2975
rect 4445 2941 4479 2975
rect 4479 2941 4488 2975
rect 4436 2932 4488 2941
rect 4528 2975 4580 2984
rect 4528 2941 4537 2975
rect 4537 2941 4571 2975
rect 4571 2941 4580 2975
rect 4896 2975 4948 2984
rect 4528 2932 4580 2941
rect 4896 2941 4905 2975
rect 4905 2941 4939 2975
rect 4939 2941 4948 2975
rect 4896 2932 4948 2941
rect 5448 2864 5500 2916
rect 4252 2839 4304 2848
rect 4252 2805 4261 2839
rect 4261 2805 4295 2839
rect 4295 2805 4304 2839
rect 4252 2796 4304 2805
rect 3598 2694 3650 2746
rect 3662 2694 3714 2746
rect 3726 2694 3778 2746
rect 3790 2694 3842 2746
rect 3976 2592 4028 2644
rect 4988 2592 5040 2644
rect 16580 2592 16632 2644
rect 2964 2524 3016 2576
rect 4344 2524 4396 2576
rect 4804 2567 4856 2576
rect 4804 2533 4813 2567
rect 4813 2533 4847 2567
rect 4847 2533 4856 2567
rect 4804 2524 4856 2533
rect 5540 2524 5592 2576
rect 6552 2567 6604 2576
rect 6552 2533 6561 2567
rect 6561 2533 6595 2567
rect 6595 2533 6604 2567
rect 6552 2524 6604 2533
rect 1216 2456 1268 2508
rect 3884 2499 3936 2508
rect 3884 2465 3893 2499
rect 3893 2465 3927 2499
rect 3927 2465 3936 2499
rect 3884 2456 3936 2465
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 4528 2456 4580 2465
rect 4804 2388 4856 2440
rect 2098 2150 2150 2202
rect 2162 2150 2214 2202
rect 2226 2150 2278 2202
rect 2290 2150 2342 2202
rect 5098 2150 5150 2202
rect 5162 2150 5214 2202
rect 5226 2150 5278 2202
rect 5290 2150 5342 2202
rect 4252 1300 4304 1352
rect 16672 1300 16724 1352
rect 4436 1232 4488 1284
rect 16764 1232 16816 1284
rect 6460 1164 6512 1216
rect 16580 1164 16632 1216
<< metal2 >>
rect 16670 13696 16726 13705
rect 16670 13631 16726 13640
rect 16578 13152 16634 13161
rect 16578 13087 16634 13096
rect 16592 12578 16620 13087
rect 6368 12572 6420 12578
rect 6368 12514 6420 12520
rect 16580 12572 16632 12578
rect 16580 12514 16632 12520
rect 3976 12504 4028 12510
rect 3976 12446 4028 12452
rect -1620 11464 -1300 11472
rect -1620 11386 -1606 11464
rect -1318 11386 -1300 11464
rect -1620 11376 -1300 11386
rect 3572 11452 3868 11472
rect 3628 11450 3652 11452
rect 3708 11450 3732 11452
rect 3788 11450 3812 11452
rect 3650 11398 3652 11450
rect 3714 11398 3726 11450
rect 3788 11398 3790 11450
rect 3628 11396 3652 11398
rect 3708 11396 3732 11398
rect 3788 11396 3812 11398
rect 3572 11376 3868 11396
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 1768 11076 1820 11082
rect 1768 11018 1820 11024
rect -960 10918 -640 10928
rect -960 10844 -948 10918
rect -658 10844 -640 10918
rect -960 10832 -640 10844
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1504 10062 1532 10542
rect 1780 10198 1808 11018
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 2072 10908 2368 10928
rect 2128 10906 2152 10908
rect 2208 10906 2232 10908
rect 2288 10906 2312 10908
rect 2150 10854 2152 10906
rect 2214 10854 2226 10906
rect 2288 10854 2290 10906
rect 2128 10852 2152 10854
rect 2208 10852 2232 10854
rect 2288 10852 2312 10854
rect 2072 10832 2368 10852
rect 1952 10532 2004 10538
rect 1952 10474 2004 10480
rect 1964 10266 1992 10474
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 3068 10198 3096 10950
rect 3896 10606 3924 11154
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3572 10364 3868 10384
rect 3628 10362 3652 10364
rect 3708 10362 3732 10364
rect 3788 10362 3812 10364
rect 3650 10310 3652 10362
rect 3714 10310 3726 10362
rect 3788 10310 3790 10362
rect 3628 10308 3652 10310
rect 3708 10308 3732 10310
rect 3788 10308 3812 10310
rect 3572 10288 3868 10308
rect 1768 10192 1820 10198
rect 1768 10134 1820 10140
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1504 8906 1532 9998
rect 2072 9820 2368 9840
rect 2128 9818 2152 9820
rect 2208 9818 2232 9820
rect 2288 9818 2312 9820
rect 2150 9766 2152 9818
rect 2214 9766 2226 9818
rect 2288 9766 2290 9818
rect 2128 9764 2152 9766
rect 2208 9764 2232 9766
rect 2288 9764 2312 9766
rect 2072 9744 2368 9764
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 1216 8900 1268 8906
rect 1216 8842 1268 8848
rect 1492 8900 1544 8906
rect 1492 8842 1544 8848
rect 1228 8430 1256 8842
rect 1216 8424 1268 8430
rect 1216 8366 1268 8372
rect 1228 7546 1256 8366
rect 1780 7750 1808 8978
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1964 8362 1992 8774
rect 2072 8732 2368 8752
rect 2128 8730 2152 8732
rect 2208 8730 2232 8732
rect 2288 8730 2312 8732
rect 2150 8678 2152 8730
rect 2214 8678 2226 8730
rect 2288 8678 2290 8730
rect 2128 8676 2152 8678
rect 2208 8676 2232 8678
rect 2288 8676 2312 8678
rect 2072 8656 2368 8676
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1964 7750 1992 7890
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1216 7540 1268 7546
rect 1216 7482 1268 7488
rect 1504 7274 1532 7686
rect 1492 7268 1544 7274
rect 1492 7210 1544 7216
rect 1780 6866 1808 7686
rect 2072 7644 2368 7664
rect 2128 7642 2152 7644
rect 2208 7642 2232 7644
rect 2288 7642 2312 7644
rect 2150 7590 2152 7642
rect 2214 7590 2226 7642
rect 2288 7590 2290 7642
rect 2128 7588 2152 7590
rect 2208 7588 2232 7590
rect 2288 7588 2312 7590
rect 2072 7568 2368 7588
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1216 6248 1268 6254
rect 1216 6190 1268 6196
rect 1228 5710 1256 6190
rect 1216 5704 1268 5710
rect 1216 5646 1268 5652
rect 1228 5166 1256 5646
rect 1216 5160 1268 5166
rect 1216 5102 1268 5108
rect 1228 4486 1256 5102
rect 1780 4690 1808 6802
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1964 5846 1992 6598
rect 2072 6556 2368 6576
rect 2128 6554 2152 6556
rect 2208 6554 2232 6556
rect 2288 6554 2312 6556
rect 2150 6502 2152 6554
rect 2214 6502 2226 6554
rect 2288 6502 2290 6554
rect 2128 6500 2152 6502
rect 2208 6500 2232 6502
rect 2288 6500 2312 6502
rect 2072 6480 2368 6500
rect 1952 5840 2004 5846
rect 1952 5782 2004 5788
rect 2072 5468 2368 5488
rect 2128 5466 2152 5468
rect 2208 5466 2232 5468
rect 2288 5466 2312 5468
rect 2150 5414 2152 5466
rect 2214 5414 2226 5466
rect 2288 5414 2290 5466
rect 2128 5412 2152 5414
rect 2208 5412 2232 5414
rect 2288 5412 2312 5414
rect 2072 5392 2368 5412
rect 1952 5092 2004 5098
rect 1952 5034 2004 5040
rect 1964 4826 1992 5034
rect 2424 4826 2452 8978
rect 2516 8294 2544 9386
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2596 6928 2648 6934
rect 2596 6870 2648 6876
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 6186 2544 6598
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2608 4690 2636 6870
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 1492 4548 1544 4554
rect 1492 4490 1544 4496
rect 1216 4480 1268 4486
rect 1216 4422 1268 4428
rect 1228 4078 1256 4422
rect 1504 4146 1532 4490
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1216 4072 1268 4078
rect 1216 4014 1268 4020
rect 1228 3942 1256 4014
rect 1964 4010 1992 4422
rect 2072 4380 2368 4400
rect 2128 4378 2152 4380
rect 2208 4378 2232 4380
rect 2288 4378 2312 4380
rect 2150 4326 2152 4378
rect 2214 4326 2226 4378
rect 2288 4326 2290 4378
rect 2128 4324 2152 4326
rect 2208 4324 2232 4326
rect 2288 4324 2312 4326
rect 2072 4304 2368 4324
rect 1952 4004 2004 4010
rect 1952 3946 2004 3952
rect 1216 3936 1268 3942
rect 1216 3878 1268 3884
rect 1228 2514 1256 3878
rect 2608 3602 2636 4626
rect 2700 3738 2728 9454
rect 2884 9042 2912 9590
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2884 7342 2912 8978
rect 2976 8838 3004 9454
rect 3572 9276 3868 9296
rect 3628 9274 3652 9276
rect 3708 9274 3732 9276
rect 3788 9274 3812 9276
rect 3650 9222 3652 9274
rect 3714 9222 3726 9274
rect 3788 9222 3790 9274
rect 3628 9220 3652 9222
rect 3708 9220 3732 9222
rect 3788 9220 3812 9222
rect 3572 9200 3868 9220
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3160 9058 3188 9114
rect 3332 9104 3384 9110
rect 3160 9052 3332 9058
rect 3160 9046 3384 9052
rect 3160 9030 3372 9046
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2976 6798 3004 7686
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 3068 6254 3096 7822
rect 3160 7546 3188 8502
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3252 8090 3280 8298
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3252 7410 3280 8026
rect 3344 7886 3372 8366
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3252 6798 3280 7210
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3252 6322 3280 6734
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2792 3670 2820 5170
rect 3068 5166 3096 6190
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3252 5914 3280 6122
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3252 5234 3280 5646
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3240 5092 3292 5098
rect 3240 5034 3292 5040
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2976 4758 3004 4966
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2884 3942 2912 4422
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2072 3292 2368 3312
rect 2128 3290 2152 3292
rect 2208 3290 2232 3292
rect 2288 3290 2312 3292
rect 2150 3238 2152 3290
rect 2214 3238 2226 3290
rect 2288 3238 2290 3290
rect 2128 3236 2152 3238
rect 2208 3236 2232 3238
rect 2288 3236 2312 3238
rect 2072 3216 2368 3236
rect 2608 3194 2636 3538
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2976 2582 3004 4694
rect 3252 4622 3280 5034
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3344 4078 3372 7482
rect 3436 5794 3464 9114
rect 3896 8566 3924 10542
rect 3988 9586 4016 12446
rect 6380 11218 6408 12514
rect 16684 12510 16712 13631
rect 16762 12608 16818 12617
rect 16762 12543 16818 12552
rect 16672 12504 16724 12510
rect 16672 12446 16724 12452
rect 16578 11520 16634 11529
rect 16578 11455 16634 11464
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4080 9178 4108 9454
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 4080 8430 4108 9114
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 3572 8188 3868 8208
rect 3628 8186 3652 8188
rect 3708 8186 3732 8188
rect 3788 8186 3812 8188
rect 3650 8134 3652 8186
rect 3714 8134 3726 8186
rect 3788 8134 3790 8186
rect 3628 8132 3652 8134
rect 3708 8132 3732 8134
rect 3788 8132 3812 8134
rect 3572 8112 3868 8132
rect 3896 7410 3924 8298
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3572 7100 3868 7120
rect 3628 7098 3652 7100
rect 3708 7098 3732 7100
rect 3788 7098 3812 7100
rect 3650 7046 3652 7098
rect 3714 7046 3726 7098
rect 3788 7046 3790 7098
rect 3628 7044 3652 7046
rect 3708 7044 3732 7046
rect 3788 7044 3812 7046
rect 3572 7024 3868 7044
rect 3988 6934 4016 7142
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3608 6792 3660 6798
rect 4080 6746 4108 7822
rect 4172 7410 4200 9386
rect 4356 8566 4384 10474
rect 4448 10062 4476 10746
rect 4540 10606 4568 10950
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4448 9586 4476 9998
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4448 8974 4476 9522
rect 4632 9042 4660 10610
rect 4724 10470 4752 11154
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5000 10674 5028 11086
rect 5072 10908 5368 10928
rect 5128 10906 5152 10908
rect 5208 10906 5232 10908
rect 5288 10906 5312 10908
rect 5150 10854 5152 10906
rect 5214 10854 5226 10906
rect 5288 10854 5290 10906
rect 5128 10852 5152 10854
rect 5208 10852 5232 10854
rect 5288 10852 5312 10854
rect 5072 10832 5368 10852
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4724 9110 4752 10406
rect 5072 9820 5368 9840
rect 5128 9818 5152 9820
rect 5208 9818 5232 9820
rect 5288 9818 5312 9820
rect 5150 9766 5152 9818
rect 5214 9766 5226 9818
rect 5288 9766 5290 9818
rect 5128 9764 5152 9766
rect 5208 9764 5232 9766
rect 5288 9764 5312 9766
rect 5072 9744 5368 9764
rect 5460 9110 5488 11086
rect 5644 10010 5672 11154
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5644 9982 5764 10010
rect 5736 9926 5764 9982
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5736 9586 5764 9862
rect 5828 9722 5856 10066
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5736 9042 5764 9522
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4356 7886 4384 8502
rect 4448 7954 4476 8910
rect 4632 8498 4660 8978
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5072 8732 5368 8752
rect 5128 8730 5152 8732
rect 5208 8730 5232 8732
rect 5288 8730 5312 8732
rect 5150 8678 5152 8730
rect 5214 8678 5226 8730
rect 5288 8678 5290 8730
rect 5128 8676 5152 8678
rect 5208 8676 5232 8678
rect 5288 8676 5312 8678
rect 5072 8656 5368 8676
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 3608 6734 3660 6740
rect 3620 6254 3648 6734
rect 3988 6718 4108 6746
rect 3988 6662 4016 6718
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3572 6012 3868 6032
rect 3628 6010 3652 6012
rect 3708 6010 3732 6012
rect 3788 6010 3812 6012
rect 3650 5958 3652 6010
rect 3714 5958 3726 6010
rect 3788 5958 3790 6010
rect 3628 5956 3652 5958
rect 3708 5956 3732 5958
rect 3788 5956 3812 5958
rect 3572 5936 3868 5956
rect 3436 5766 3648 5794
rect 3620 5710 3648 5766
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3436 4146 3464 5510
rect 3896 5166 3924 6190
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5846 4108 6054
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4172 5710 4200 7346
rect 4448 6338 4476 7890
rect 4264 6316 4476 6338
rect 4264 6310 4344 6316
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3572 4924 3868 4944
rect 3628 4922 3652 4924
rect 3708 4922 3732 4924
rect 3788 4922 3812 4924
rect 3650 4870 3652 4922
rect 3714 4870 3726 4922
rect 3788 4870 3790 4922
rect 3628 4868 3652 4870
rect 3708 4868 3732 4870
rect 3788 4868 3812 4870
rect 3572 4848 3868 4868
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 3528 4282 3556 4694
rect 3988 4282 4016 5646
rect 4264 5234 4292 6310
rect 4396 6310 4476 6316
rect 4344 6258 4396 6264
rect 4540 5386 4568 8298
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4448 5358 4568 5386
rect 4632 5370 4660 7210
rect 4724 6458 4752 8298
rect 4816 8090 4844 8570
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5072 7644 5368 7664
rect 5128 7642 5152 7644
rect 5208 7642 5232 7644
rect 5288 7642 5312 7644
rect 5150 7590 5152 7642
rect 5214 7590 5226 7642
rect 5288 7590 5290 7642
rect 5128 7588 5152 7590
rect 5208 7588 5232 7590
rect 5288 7588 5312 7590
rect 5072 7568 5368 7588
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4620 5364 4672 5370
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3252 3058 3280 3946
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3344 2990 3372 4014
rect 3572 3836 3868 3856
rect 3628 3834 3652 3836
rect 3708 3834 3732 3836
rect 3788 3834 3812 3836
rect 3650 3782 3652 3834
rect 3714 3782 3726 3834
rect 3788 3782 3790 3834
rect 3628 3780 3652 3782
rect 3708 3780 3732 3782
rect 3788 3780 3812 3782
rect 3572 3760 3868 3780
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3572 2748 3868 2768
rect 3628 2746 3652 2748
rect 3708 2746 3732 2748
rect 3788 2746 3812 2748
rect 3650 2694 3652 2746
rect 3714 2694 3726 2746
rect 3788 2694 3790 2746
rect 3628 2692 3652 2694
rect 3708 2692 3732 2694
rect 3788 2692 3812 2694
rect 3572 2672 3868 2692
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 3896 2514 3924 2926
rect 3988 2650 4016 3538
rect 4448 3194 4476 5358
rect 4620 5306 4672 5312
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4448 3074 4476 3130
rect 4356 3046 4476 3074
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 1216 2508 1268 2514
rect 1216 2450 1268 2456
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 2072 2204 2368 2224
rect 2128 2202 2152 2204
rect 2208 2202 2232 2204
rect 2288 2202 2312 2204
rect 2150 2150 2152 2202
rect 2214 2150 2226 2202
rect 2288 2150 2290 2202
rect 2128 2148 2152 2150
rect 2208 2148 2232 2150
rect 2288 2148 2312 2150
rect 2072 2128 2368 2148
rect 4264 1358 4292 2790
rect 4356 2582 4384 3046
rect 4540 2990 4568 5170
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 4252 1352 4304 1358
rect 4252 1294 4304 1300
rect 4448 1290 4476 2926
rect 4540 2514 4568 2926
rect 4816 2582 4844 7346
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 5778 4936 6598
rect 5072 6556 5368 6576
rect 5128 6554 5152 6556
rect 5208 6554 5232 6556
rect 5288 6554 5312 6556
rect 5150 6502 5152 6554
rect 5214 6502 5226 6554
rect 5288 6502 5290 6554
rect 5128 6500 5152 6502
rect 5208 6500 5232 6502
rect 5288 6500 5312 6502
rect 5072 6480 5368 6500
rect 5460 6118 5488 7958
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 6798 5580 7142
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4908 3602 4936 5714
rect 5072 5468 5368 5488
rect 5128 5466 5152 5468
rect 5208 5466 5232 5468
rect 5288 5466 5312 5468
rect 5150 5414 5152 5466
rect 5214 5414 5226 5466
rect 5288 5414 5290 5466
rect 5128 5412 5152 5414
rect 5208 5412 5232 5414
rect 5288 5412 5312 5414
rect 5072 5392 5368 5412
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5072 4380 5368 4400
rect 5128 4378 5152 4380
rect 5208 4378 5232 4380
rect 5288 4378 5312 4380
rect 5150 4326 5152 4378
rect 5214 4326 5226 4378
rect 5288 4326 5290 4378
rect 5128 4324 5152 4326
rect 5208 4324 5232 4326
rect 5288 4324 5312 4326
rect 5072 4304 5368 4324
rect 5460 3942 5488 4558
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5644 3602 5672 8774
rect 5828 8498 5856 9658
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5920 7886 5948 11154
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6012 9450 6040 9862
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 6196 9058 6224 11086
rect 6368 9376 6420 9382
rect 6472 9330 6500 11086
rect 16592 11082 16620 11455
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16776 10674 16804 12543
rect 26330 12064 26386 12073
rect 26330 11999 26386 12008
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6564 9722 6592 10542
rect 16580 10464 16632 10470
rect 16578 10432 16580 10441
rect 16632 10432 16634 10441
rect 16578 10367 16634 10376
rect 26238 9888 26294 9897
rect 26238 9823 26294 9832
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6420 9324 6500 9330
rect 6368 9318 6500 9324
rect 6380 9302 6500 9318
rect 6472 9178 6500 9302
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6012 9030 6224 9058
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5736 6458 5764 6666
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5920 5778 5948 6190
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5736 5098 5764 5510
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 6012 4146 6040 9030
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 6798 6316 7686
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 6104 5914 6132 6122
rect 6380 6066 6408 8298
rect 6564 7750 6592 9454
rect 26252 9450 26280 9823
rect 26240 9444 26292 9450
rect 26240 9386 26292 9392
rect 16670 9344 16726 9353
rect 16670 9279 16726 9288
rect 16580 9104 16632 9110
rect 16580 9046 16632 9052
rect 16592 8809 16620 9046
rect 16684 8974 16712 9279
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16578 8800 16634 8809
rect 16578 8735 16634 8744
rect 26344 8362 26372 11999
rect 26422 10976 26478 10985
rect 26422 10911 26478 10920
rect 26332 8356 26384 8362
rect 26332 8298 26384 8304
rect 16580 8288 16632 8294
rect 16578 8256 16580 8265
rect 16632 8256 16634 8265
rect 16578 8191 16634 8200
rect 6552 7744 6604 7750
rect 16672 7744 16724 7750
rect 6552 7686 6604 7692
rect 16578 7712 16634 7721
rect 16672 7686 16724 7692
rect 16578 7647 16634 7656
rect 16592 7342 16620 7647
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 6552 7200 6604 7206
rect 16684 7177 16712 7686
rect 6552 7142 6604 7148
rect 16670 7168 16726 7177
rect 6564 6934 6592 7142
rect 16670 7103 16726 7112
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6288 6038 6408 6066
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6196 4078 6224 5510
rect 6288 5302 6316 6038
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6380 5234 6408 5714
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6380 5030 6408 5170
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6380 4078 6408 4150
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4908 2990 4936 3130
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 5000 2650 5028 3538
rect 5828 3466 5856 3674
rect 6104 3602 6132 3946
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5072 3292 5368 3312
rect 5128 3290 5152 3292
rect 5208 3290 5232 3292
rect 5288 3290 5312 3292
rect 5150 3238 5152 3290
rect 5214 3238 5226 3290
rect 5288 3238 5290 3290
rect 5128 3236 5152 3238
rect 5208 3236 5232 3238
rect 5288 3236 5312 3238
rect 5072 3216 5368 3236
rect 5460 2922 5488 3402
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5552 2582 5580 3334
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4816 2446 4844 2518
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 5072 2204 5368 2224
rect 5128 2202 5152 2204
rect 5208 2202 5232 2204
rect 5288 2202 5312 2204
rect 5150 2150 5152 2202
rect 5214 2150 5226 2202
rect 5288 2150 5290 2202
rect 5128 2148 5152 2150
rect 5208 2148 5232 2150
rect 5288 2148 5312 2150
rect 5072 2128 5368 2148
rect 4436 1284 4488 1290
rect 4436 1226 4488 1232
rect 6472 1222 6500 6734
rect 16670 6624 16726 6633
rect 16670 6559 16726 6568
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16592 6089 16620 6394
rect 16684 6186 16712 6559
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16578 6080 16634 6089
rect 16578 6015 16634 6024
rect 16578 5536 16634 5545
rect 16578 5471 16634 5480
rect 16592 5030 16620 5471
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16670 4992 16726 5001
rect 16670 4927 16726 4936
rect 16684 4146 16712 4927
rect 26436 4690 26464 10911
rect 26424 4684 26476 4690
rect 26424 4626 26476 4632
rect 16762 4448 16818 4457
rect 16762 4383 16818 4392
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6564 2582 6592 3538
rect 6656 3194 6684 4082
rect 16580 3936 16632 3942
rect 16578 3904 16580 3913
rect 16632 3904 16634 3913
rect 16578 3839 16634 3848
rect 16776 3602 16804 4383
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16578 3360 16634 3369
rect 16578 3295 16634 3304
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 16592 3058 16620 3295
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16684 2825 16712 3470
rect 16670 2816 16726 2825
rect 16670 2751 16726 2760
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 16592 2281 16620 2586
rect 16578 2272 16634 2281
rect 16578 2207 16634 2216
rect 16868 1737 16896 4014
rect 16854 1728 16910 1737
rect 16854 1663 16910 1672
rect 16672 1352 16724 1358
rect 16672 1294 16724 1300
rect 6460 1216 6512 1222
rect 16580 1216 16632 1222
rect 6460 1158 6512 1164
rect 16578 1184 16580 1193
rect 16632 1184 16634 1193
rect 16578 1119 16634 1128
rect 16684 649 16712 1294
rect 16764 1284 16816 1290
rect 16764 1226 16816 1232
rect 16670 640 16726 649
rect 16670 575 16726 584
rect 16776 241 16804 1226
rect 16762 232 16818 241
rect 16762 167 16818 176
<< via2 >>
rect 16670 13640 16726 13696
rect 16578 13096 16634 13152
rect -1606 11386 -1318 11464
rect 3572 11450 3628 11452
rect 3652 11450 3708 11452
rect 3732 11450 3788 11452
rect 3812 11450 3868 11452
rect 3572 11398 3598 11450
rect 3598 11398 3628 11450
rect 3652 11398 3662 11450
rect 3662 11398 3708 11450
rect 3732 11398 3778 11450
rect 3778 11398 3788 11450
rect 3812 11398 3842 11450
rect 3842 11398 3868 11450
rect 3572 11396 3628 11398
rect 3652 11396 3708 11398
rect 3732 11396 3788 11398
rect 3812 11396 3868 11398
rect -948 10844 -658 10918
rect 2072 10906 2128 10908
rect 2152 10906 2208 10908
rect 2232 10906 2288 10908
rect 2312 10906 2368 10908
rect 2072 10854 2098 10906
rect 2098 10854 2128 10906
rect 2152 10854 2162 10906
rect 2162 10854 2208 10906
rect 2232 10854 2278 10906
rect 2278 10854 2288 10906
rect 2312 10854 2342 10906
rect 2342 10854 2368 10906
rect 2072 10852 2128 10854
rect 2152 10852 2208 10854
rect 2232 10852 2288 10854
rect 2312 10852 2368 10854
rect 3572 10362 3628 10364
rect 3652 10362 3708 10364
rect 3732 10362 3788 10364
rect 3812 10362 3868 10364
rect 3572 10310 3598 10362
rect 3598 10310 3628 10362
rect 3652 10310 3662 10362
rect 3662 10310 3708 10362
rect 3732 10310 3778 10362
rect 3778 10310 3788 10362
rect 3812 10310 3842 10362
rect 3842 10310 3868 10362
rect 3572 10308 3628 10310
rect 3652 10308 3708 10310
rect 3732 10308 3788 10310
rect 3812 10308 3868 10310
rect 2072 9818 2128 9820
rect 2152 9818 2208 9820
rect 2232 9818 2288 9820
rect 2312 9818 2368 9820
rect 2072 9766 2098 9818
rect 2098 9766 2128 9818
rect 2152 9766 2162 9818
rect 2162 9766 2208 9818
rect 2232 9766 2278 9818
rect 2278 9766 2288 9818
rect 2312 9766 2342 9818
rect 2342 9766 2368 9818
rect 2072 9764 2128 9766
rect 2152 9764 2208 9766
rect 2232 9764 2288 9766
rect 2312 9764 2368 9766
rect 2072 8730 2128 8732
rect 2152 8730 2208 8732
rect 2232 8730 2288 8732
rect 2312 8730 2368 8732
rect 2072 8678 2098 8730
rect 2098 8678 2128 8730
rect 2152 8678 2162 8730
rect 2162 8678 2208 8730
rect 2232 8678 2278 8730
rect 2278 8678 2288 8730
rect 2312 8678 2342 8730
rect 2342 8678 2368 8730
rect 2072 8676 2128 8678
rect 2152 8676 2208 8678
rect 2232 8676 2288 8678
rect 2312 8676 2368 8678
rect 2072 7642 2128 7644
rect 2152 7642 2208 7644
rect 2232 7642 2288 7644
rect 2312 7642 2368 7644
rect 2072 7590 2098 7642
rect 2098 7590 2128 7642
rect 2152 7590 2162 7642
rect 2162 7590 2208 7642
rect 2232 7590 2278 7642
rect 2278 7590 2288 7642
rect 2312 7590 2342 7642
rect 2342 7590 2368 7642
rect 2072 7588 2128 7590
rect 2152 7588 2208 7590
rect 2232 7588 2288 7590
rect 2312 7588 2368 7590
rect 2072 6554 2128 6556
rect 2152 6554 2208 6556
rect 2232 6554 2288 6556
rect 2312 6554 2368 6556
rect 2072 6502 2098 6554
rect 2098 6502 2128 6554
rect 2152 6502 2162 6554
rect 2162 6502 2208 6554
rect 2232 6502 2278 6554
rect 2278 6502 2288 6554
rect 2312 6502 2342 6554
rect 2342 6502 2368 6554
rect 2072 6500 2128 6502
rect 2152 6500 2208 6502
rect 2232 6500 2288 6502
rect 2312 6500 2368 6502
rect 2072 5466 2128 5468
rect 2152 5466 2208 5468
rect 2232 5466 2288 5468
rect 2312 5466 2368 5468
rect 2072 5414 2098 5466
rect 2098 5414 2128 5466
rect 2152 5414 2162 5466
rect 2162 5414 2208 5466
rect 2232 5414 2278 5466
rect 2278 5414 2288 5466
rect 2312 5414 2342 5466
rect 2342 5414 2368 5466
rect 2072 5412 2128 5414
rect 2152 5412 2208 5414
rect 2232 5412 2288 5414
rect 2312 5412 2368 5414
rect 2072 4378 2128 4380
rect 2152 4378 2208 4380
rect 2232 4378 2288 4380
rect 2312 4378 2368 4380
rect 2072 4326 2098 4378
rect 2098 4326 2128 4378
rect 2152 4326 2162 4378
rect 2162 4326 2208 4378
rect 2232 4326 2278 4378
rect 2278 4326 2288 4378
rect 2312 4326 2342 4378
rect 2342 4326 2368 4378
rect 2072 4324 2128 4326
rect 2152 4324 2208 4326
rect 2232 4324 2288 4326
rect 2312 4324 2368 4326
rect 3572 9274 3628 9276
rect 3652 9274 3708 9276
rect 3732 9274 3788 9276
rect 3812 9274 3868 9276
rect 3572 9222 3598 9274
rect 3598 9222 3628 9274
rect 3652 9222 3662 9274
rect 3662 9222 3708 9274
rect 3732 9222 3778 9274
rect 3778 9222 3788 9274
rect 3812 9222 3842 9274
rect 3842 9222 3868 9274
rect 3572 9220 3628 9222
rect 3652 9220 3708 9222
rect 3732 9220 3788 9222
rect 3812 9220 3868 9222
rect 2072 3290 2128 3292
rect 2152 3290 2208 3292
rect 2232 3290 2288 3292
rect 2312 3290 2368 3292
rect 2072 3238 2098 3290
rect 2098 3238 2128 3290
rect 2152 3238 2162 3290
rect 2162 3238 2208 3290
rect 2232 3238 2278 3290
rect 2278 3238 2288 3290
rect 2312 3238 2342 3290
rect 2342 3238 2368 3290
rect 2072 3236 2128 3238
rect 2152 3236 2208 3238
rect 2232 3236 2288 3238
rect 2312 3236 2368 3238
rect 16762 12552 16818 12608
rect 16578 11464 16634 11520
rect 3572 8186 3628 8188
rect 3652 8186 3708 8188
rect 3732 8186 3788 8188
rect 3812 8186 3868 8188
rect 3572 8134 3598 8186
rect 3598 8134 3628 8186
rect 3652 8134 3662 8186
rect 3662 8134 3708 8186
rect 3732 8134 3778 8186
rect 3778 8134 3788 8186
rect 3812 8134 3842 8186
rect 3842 8134 3868 8186
rect 3572 8132 3628 8134
rect 3652 8132 3708 8134
rect 3732 8132 3788 8134
rect 3812 8132 3868 8134
rect 3572 7098 3628 7100
rect 3652 7098 3708 7100
rect 3732 7098 3788 7100
rect 3812 7098 3868 7100
rect 3572 7046 3598 7098
rect 3598 7046 3628 7098
rect 3652 7046 3662 7098
rect 3662 7046 3708 7098
rect 3732 7046 3778 7098
rect 3778 7046 3788 7098
rect 3812 7046 3842 7098
rect 3842 7046 3868 7098
rect 3572 7044 3628 7046
rect 3652 7044 3708 7046
rect 3732 7044 3788 7046
rect 3812 7044 3868 7046
rect 5072 10906 5128 10908
rect 5152 10906 5208 10908
rect 5232 10906 5288 10908
rect 5312 10906 5368 10908
rect 5072 10854 5098 10906
rect 5098 10854 5128 10906
rect 5152 10854 5162 10906
rect 5162 10854 5208 10906
rect 5232 10854 5278 10906
rect 5278 10854 5288 10906
rect 5312 10854 5342 10906
rect 5342 10854 5368 10906
rect 5072 10852 5128 10854
rect 5152 10852 5208 10854
rect 5232 10852 5288 10854
rect 5312 10852 5368 10854
rect 5072 9818 5128 9820
rect 5152 9818 5208 9820
rect 5232 9818 5288 9820
rect 5312 9818 5368 9820
rect 5072 9766 5098 9818
rect 5098 9766 5128 9818
rect 5152 9766 5162 9818
rect 5162 9766 5208 9818
rect 5232 9766 5278 9818
rect 5278 9766 5288 9818
rect 5312 9766 5342 9818
rect 5342 9766 5368 9818
rect 5072 9764 5128 9766
rect 5152 9764 5208 9766
rect 5232 9764 5288 9766
rect 5312 9764 5368 9766
rect 5072 8730 5128 8732
rect 5152 8730 5208 8732
rect 5232 8730 5288 8732
rect 5312 8730 5368 8732
rect 5072 8678 5098 8730
rect 5098 8678 5128 8730
rect 5152 8678 5162 8730
rect 5162 8678 5208 8730
rect 5232 8678 5278 8730
rect 5278 8678 5288 8730
rect 5312 8678 5342 8730
rect 5342 8678 5368 8730
rect 5072 8676 5128 8678
rect 5152 8676 5208 8678
rect 5232 8676 5288 8678
rect 5312 8676 5368 8678
rect 3572 6010 3628 6012
rect 3652 6010 3708 6012
rect 3732 6010 3788 6012
rect 3812 6010 3868 6012
rect 3572 5958 3598 6010
rect 3598 5958 3628 6010
rect 3652 5958 3662 6010
rect 3662 5958 3708 6010
rect 3732 5958 3778 6010
rect 3778 5958 3788 6010
rect 3812 5958 3842 6010
rect 3842 5958 3868 6010
rect 3572 5956 3628 5958
rect 3652 5956 3708 5958
rect 3732 5956 3788 5958
rect 3812 5956 3868 5958
rect 3572 4922 3628 4924
rect 3652 4922 3708 4924
rect 3732 4922 3788 4924
rect 3812 4922 3868 4924
rect 3572 4870 3598 4922
rect 3598 4870 3628 4922
rect 3652 4870 3662 4922
rect 3662 4870 3708 4922
rect 3732 4870 3778 4922
rect 3778 4870 3788 4922
rect 3812 4870 3842 4922
rect 3842 4870 3868 4922
rect 3572 4868 3628 4870
rect 3652 4868 3708 4870
rect 3732 4868 3788 4870
rect 3812 4868 3868 4870
rect 5072 7642 5128 7644
rect 5152 7642 5208 7644
rect 5232 7642 5288 7644
rect 5312 7642 5368 7644
rect 5072 7590 5098 7642
rect 5098 7590 5128 7642
rect 5152 7590 5162 7642
rect 5162 7590 5208 7642
rect 5232 7590 5278 7642
rect 5278 7590 5288 7642
rect 5312 7590 5342 7642
rect 5342 7590 5368 7642
rect 5072 7588 5128 7590
rect 5152 7588 5208 7590
rect 5232 7588 5288 7590
rect 5312 7588 5368 7590
rect 3572 3834 3628 3836
rect 3652 3834 3708 3836
rect 3732 3834 3788 3836
rect 3812 3834 3868 3836
rect 3572 3782 3598 3834
rect 3598 3782 3628 3834
rect 3652 3782 3662 3834
rect 3662 3782 3708 3834
rect 3732 3782 3778 3834
rect 3778 3782 3788 3834
rect 3812 3782 3842 3834
rect 3842 3782 3868 3834
rect 3572 3780 3628 3782
rect 3652 3780 3708 3782
rect 3732 3780 3788 3782
rect 3812 3780 3868 3782
rect 3572 2746 3628 2748
rect 3652 2746 3708 2748
rect 3732 2746 3788 2748
rect 3812 2746 3868 2748
rect 3572 2694 3598 2746
rect 3598 2694 3628 2746
rect 3652 2694 3662 2746
rect 3662 2694 3708 2746
rect 3732 2694 3778 2746
rect 3778 2694 3788 2746
rect 3812 2694 3842 2746
rect 3842 2694 3868 2746
rect 3572 2692 3628 2694
rect 3652 2692 3708 2694
rect 3732 2692 3788 2694
rect 3812 2692 3868 2694
rect 2072 2202 2128 2204
rect 2152 2202 2208 2204
rect 2232 2202 2288 2204
rect 2312 2202 2368 2204
rect 2072 2150 2098 2202
rect 2098 2150 2128 2202
rect 2152 2150 2162 2202
rect 2162 2150 2208 2202
rect 2232 2150 2278 2202
rect 2278 2150 2288 2202
rect 2312 2150 2342 2202
rect 2342 2150 2368 2202
rect 2072 2148 2128 2150
rect 2152 2148 2208 2150
rect 2232 2148 2288 2150
rect 2312 2148 2368 2150
rect 5072 6554 5128 6556
rect 5152 6554 5208 6556
rect 5232 6554 5288 6556
rect 5312 6554 5368 6556
rect 5072 6502 5098 6554
rect 5098 6502 5128 6554
rect 5152 6502 5162 6554
rect 5162 6502 5208 6554
rect 5232 6502 5278 6554
rect 5278 6502 5288 6554
rect 5312 6502 5342 6554
rect 5342 6502 5368 6554
rect 5072 6500 5128 6502
rect 5152 6500 5208 6502
rect 5232 6500 5288 6502
rect 5312 6500 5368 6502
rect 5072 5466 5128 5468
rect 5152 5466 5208 5468
rect 5232 5466 5288 5468
rect 5312 5466 5368 5468
rect 5072 5414 5098 5466
rect 5098 5414 5128 5466
rect 5152 5414 5162 5466
rect 5162 5414 5208 5466
rect 5232 5414 5278 5466
rect 5278 5414 5288 5466
rect 5312 5414 5342 5466
rect 5342 5414 5368 5466
rect 5072 5412 5128 5414
rect 5152 5412 5208 5414
rect 5232 5412 5288 5414
rect 5312 5412 5368 5414
rect 5072 4378 5128 4380
rect 5152 4378 5208 4380
rect 5232 4378 5288 4380
rect 5312 4378 5368 4380
rect 5072 4326 5098 4378
rect 5098 4326 5128 4378
rect 5152 4326 5162 4378
rect 5162 4326 5208 4378
rect 5232 4326 5278 4378
rect 5278 4326 5288 4378
rect 5312 4326 5342 4378
rect 5342 4326 5368 4378
rect 5072 4324 5128 4326
rect 5152 4324 5208 4326
rect 5232 4324 5288 4326
rect 5312 4324 5368 4326
rect 26330 12008 26386 12064
rect 16578 10412 16580 10432
rect 16580 10412 16632 10432
rect 16632 10412 16634 10432
rect 16578 10376 16634 10412
rect 26238 9832 26294 9888
rect 16670 9288 16726 9344
rect 16578 8744 16634 8800
rect 26422 10920 26478 10976
rect 16578 8236 16580 8256
rect 16580 8236 16632 8256
rect 16632 8236 16634 8256
rect 16578 8200 16634 8236
rect 16578 7656 16634 7712
rect 16670 7112 16726 7168
rect 5072 3290 5128 3292
rect 5152 3290 5208 3292
rect 5232 3290 5288 3292
rect 5312 3290 5368 3292
rect 5072 3238 5098 3290
rect 5098 3238 5128 3290
rect 5152 3238 5162 3290
rect 5162 3238 5208 3290
rect 5232 3238 5278 3290
rect 5278 3238 5288 3290
rect 5312 3238 5342 3290
rect 5342 3238 5368 3290
rect 5072 3236 5128 3238
rect 5152 3236 5208 3238
rect 5232 3236 5288 3238
rect 5312 3236 5368 3238
rect 5072 2202 5128 2204
rect 5152 2202 5208 2204
rect 5232 2202 5288 2204
rect 5312 2202 5368 2204
rect 5072 2150 5098 2202
rect 5098 2150 5128 2202
rect 5152 2150 5162 2202
rect 5162 2150 5208 2202
rect 5232 2150 5278 2202
rect 5278 2150 5288 2202
rect 5312 2150 5342 2202
rect 5342 2150 5368 2202
rect 5072 2148 5128 2150
rect 5152 2148 5208 2150
rect 5232 2148 5288 2150
rect 5312 2148 5368 2150
rect 16670 6568 16726 6624
rect 16578 6024 16634 6080
rect 16578 5480 16634 5536
rect 16670 4936 16726 4992
rect 16762 4392 16818 4448
rect 16578 3884 16580 3904
rect 16580 3884 16632 3904
rect 16632 3884 16634 3904
rect 16578 3848 16634 3884
rect 16578 3304 16634 3360
rect 16670 2760 16726 2816
rect 16578 2216 16634 2272
rect 16854 1672 16910 1728
rect 16578 1164 16580 1184
rect 16580 1164 16632 1184
rect 16632 1164 16634 1184
rect 16578 1128 16634 1164
rect 16670 584 16726 640
rect 16762 176 16818 232
<< metal3 >>
rect 14000 13696 34000 13728
rect 14000 13640 16670 13696
rect 16726 13640 34000 13696
rect 14000 13608 34000 13640
rect 14000 13152 34000 13184
rect 14000 13096 16578 13152
rect 16634 13096 34000 13152
rect 14000 13064 34000 13096
rect 14000 12608 34000 12640
rect 14000 12552 16762 12608
rect 16818 12552 34000 12608
rect 14000 12520 34000 12552
rect 14000 12064 34000 12096
rect 14000 12008 26330 12064
rect 26386 12008 34000 12064
rect 14000 11976 34000 12008
rect 14000 11520 34000 11552
rect -1620 11464 -1300 11472
rect -1620 11386 -1606 11464
rect -1318 11386 -1300 11464
rect 14000 11464 16578 11520
rect 16634 11464 34000 11520
rect 3560 11456 3880 11457
rect 3560 11392 3568 11456
rect 3632 11392 3648 11456
rect 3712 11392 3728 11456
rect 3792 11392 3808 11456
rect 3872 11392 3880 11456
rect 14000 11432 34000 11464
rect 3560 11391 3880 11392
rect -1620 11376 -1300 11386
rect 14000 10976 34000 11008
rect -960 10918 -640 10928
rect -960 10844 -948 10918
rect -658 10844 -640 10918
rect 14000 10920 26422 10976
rect 26478 10920 34000 10976
rect 2060 10912 2380 10913
rect 2060 10848 2068 10912
rect 2132 10848 2148 10912
rect 2212 10848 2228 10912
rect 2292 10848 2308 10912
rect 2372 10848 2380 10912
rect 2060 10847 2380 10848
rect 5060 10912 5380 10913
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 14000 10888 34000 10920
rect 5060 10847 5380 10848
rect -960 10832 -640 10844
rect 14000 10432 34000 10464
rect 14000 10376 16578 10432
rect 16634 10376 34000 10432
rect 3560 10368 3880 10369
rect 3560 10304 3568 10368
rect 3632 10304 3648 10368
rect 3712 10304 3728 10368
rect 3792 10304 3808 10368
rect 3872 10304 3880 10368
rect 14000 10344 34000 10376
rect 3560 10303 3880 10304
rect 14000 9888 34000 9920
rect 14000 9832 26238 9888
rect 26294 9832 34000 9888
rect 2060 9824 2380 9825
rect 2060 9760 2068 9824
rect 2132 9760 2148 9824
rect 2212 9760 2228 9824
rect 2292 9760 2308 9824
rect 2372 9760 2380 9824
rect 2060 9759 2380 9760
rect 5060 9824 5380 9825
rect 5060 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5380 9824
rect 14000 9800 34000 9832
rect 5060 9759 5380 9760
rect 14000 9344 34000 9376
rect 14000 9288 16670 9344
rect 16726 9288 34000 9344
rect 3560 9280 3880 9281
rect 3560 9216 3568 9280
rect 3632 9216 3648 9280
rect 3712 9216 3728 9280
rect 3792 9216 3808 9280
rect 3872 9216 3880 9280
rect 14000 9256 34000 9288
rect 3560 9215 3880 9216
rect 14000 8800 34000 8832
rect 14000 8744 16578 8800
rect 16634 8744 34000 8800
rect 2060 8736 2380 8737
rect 2060 8672 2068 8736
rect 2132 8672 2148 8736
rect 2212 8672 2228 8736
rect 2292 8672 2308 8736
rect 2372 8672 2380 8736
rect 2060 8671 2380 8672
rect 5060 8736 5380 8737
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 14000 8712 34000 8744
rect 5060 8671 5380 8672
rect 14000 8256 34000 8288
rect 14000 8200 16578 8256
rect 16634 8200 34000 8256
rect 3560 8192 3880 8193
rect 3560 8128 3568 8192
rect 3632 8128 3648 8192
rect 3712 8128 3728 8192
rect 3792 8128 3808 8192
rect 3872 8128 3880 8192
rect 14000 8168 34000 8200
rect 3560 8127 3880 8128
rect 14000 7712 34000 7744
rect 14000 7656 16578 7712
rect 16634 7656 34000 7712
rect 2060 7648 2380 7649
rect 2060 7584 2068 7648
rect 2132 7584 2148 7648
rect 2212 7584 2228 7648
rect 2292 7584 2308 7648
rect 2372 7584 2380 7648
rect 2060 7583 2380 7584
rect 5060 7648 5380 7649
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 14000 7624 34000 7656
rect 5060 7583 5380 7584
rect 14000 7168 34000 7200
rect 14000 7112 16670 7168
rect 16726 7112 34000 7168
rect 3560 7104 3880 7105
rect 3560 7040 3568 7104
rect 3632 7040 3648 7104
rect 3712 7040 3728 7104
rect 3792 7040 3808 7104
rect 3872 7040 3880 7104
rect 14000 7080 34000 7112
rect 3560 7039 3880 7040
rect 14000 6624 34000 6656
rect 14000 6568 16670 6624
rect 16726 6568 34000 6624
rect 2060 6560 2380 6561
rect 2060 6496 2068 6560
rect 2132 6496 2148 6560
rect 2212 6496 2228 6560
rect 2292 6496 2308 6560
rect 2372 6496 2380 6560
rect 2060 6495 2380 6496
rect 5060 6560 5380 6561
rect 5060 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5380 6560
rect 14000 6536 34000 6568
rect 5060 6495 5380 6496
rect 14000 6080 34000 6112
rect 14000 6024 16578 6080
rect 16634 6024 34000 6080
rect 3560 6016 3880 6017
rect 3560 5952 3568 6016
rect 3632 5952 3648 6016
rect 3712 5952 3728 6016
rect 3792 5952 3808 6016
rect 3872 5952 3880 6016
rect 14000 5992 34000 6024
rect 3560 5951 3880 5952
rect 14000 5536 34000 5568
rect 14000 5480 16578 5536
rect 16634 5480 34000 5536
rect 2060 5472 2380 5473
rect 2060 5408 2068 5472
rect 2132 5408 2148 5472
rect 2212 5408 2228 5472
rect 2292 5408 2308 5472
rect 2372 5408 2380 5472
rect 2060 5407 2380 5408
rect 5060 5472 5380 5473
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 14000 5448 34000 5480
rect 5060 5407 5380 5408
rect 14000 4992 34000 5024
rect 14000 4936 16670 4992
rect 16726 4936 34000 4992
rect 3560 4928 3880 4929
rect 3560 4864 3568 4928
rect 3632 4864 3648 4928
rect 3712 4864 3728 4928
rect 3792 4864 3808 4928
rect 3872 4864 3880 4928
rect 14000 4904 34000 4936
rect 3560 4863 3880 4864
rect 14000 4448 34000 4480
rect 14000 4392 16762 4448
rect 16818 4392 34000 4448
rect 2060 4384 2380 4385
rect 2060 4320 2068 4384
rect 2132 4320 2148 4384
rect 2212 4320 2228 4384
rect 2292 4320 2308 4384
rect 2372 4320 2380 4384
rect 2060 4319 2380 4320
rect 5060 4384 5380 4385
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 14000 4360 34000 4392
rect 5060 4319 5380 4320
rect 14000 3904 34000 3936
rect 14000 3848 16578 3904
rect 16634 3848 34000 3904
rect 3560 3840 3880 3841
rect 3560 3776 3568 3840
rect 3632 3776 3648 3840
rect 3712 3776 3728 3840
rect 3792 3776 3808 3840
rect 3872 3776 3880 3840
rect 14000 3816 34000 3848
rect 3560 3775 3880 3776
rect 14000 3360 34000 3392
rect 14000 3304 16578 3360
rect 16634 3304 34000 3360
rect 2060 3296 2380 3297
rect 2060 3232 2068 3296
rect 2132 3232 2148 3296
rect 2212 3232 2228 3296
rect 2292 3232 2308 3296
rect 2372 3232 2380 3296
rect 2060 3231 2380 3232
rect 5060 3296 5380 3297
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 14000 3272 34000 3304
rect 5060 3231 5380 3232
rect 14000 2816 34000 2848
rect 14000 2760 16670 2816
rect 16726 2760 34000 2816
rect 3560 2752 3880 2753
rect 3560 2688 3568 2752
rect 3632 2688 3648 2752
rect 3712 2688 3728 2752
rect 3792 2688 3808 2752
rect 3872 2688 3880 2752
rect 14000 2728 34000 2760
rect 3560 2687 3880 2688
rect 14000 2272 34000 2304
rect 14000 2216 16578 2272
rect 16634 2216 34000 2272
rect 2060 2208 2380 2209
rect 2060 2144 2068 2208
rect 2132 2144 2148 2208
rect 2212 2144 2228 2208
rect 2292 2144 2308 2208
rect 2372 2144 2380 2208
rect 2060 2143 2380 2144
rect 5060 2208 5380 2209
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 14000 2184 34000 2216
rect 5060 2143 5380 2144
rect 14000 1728 34000 1760
rect 14000 1672 16854 1728
rect 16910 1672 34000 1728
rect 14000 1640 34000 1672
rect 14000 1184 34000 1216
rect 14000 1128 16578 1184
rect 16634 1128 34000 1184
rect 14000 1096 34000 1128
rect 14000 640 34000 672
rect 14000 584 16670 640
rect 16726 584 34000 640
rect 14000 552 34000 584
rect 14000 232 34000 264
rect 14000 176 16762 232
rect 16818 176 34000 232
rect 14000 144 34000 176
<< via3 >>
rect -1606 11386 -1318 11464
rect 3568 11452 3632 11456
rect 3568 11396 3572 11452
rect 3572 11396 3628 11452
rect 3628 11396 3632 11452
rect 3568 11392 3632 11396
rect 3648 11452 3712 11456
rect 3648 11396 3652 11452
rect 3652 11396 3708 11452
rect 3708 11396 3712 11452
rect 3648 11392 3712 11396
rect 3728 11452 3792 11456
rect 3728 11396 3732 11452
rect 3732 11396 3788 11452
rect 3788 11396 3792 11452
rect 3728 11392 3792 11396
rect 3808 11452 3872 11456
rect 3808 11396 3812 11452
rect 3812 11396 3868 11452
rect 3868 11396 3872 11452
rect 3808 11392 3872 11396
rect -948 10844 -658 10918
rect 2068 10908 2132 10912
rect 2068 10852 2072 10908
rect 2072 10852 2128 10908
rect 2128 10852 2132 10908
rect 2068 10848 2132 10852
rect 2148 10908 2212 10912
rect 2148 10852 2152 10908
rect 2152 10852 2208 10908
rect 2208 10852 2212 10908
rect 2148 10848 2212 10852
rect 2228 10908 2292 10912
rect 2228 10852 2232 10908
rect 2232 10852 2288 10908
rect 2288 10852 2292 10908
rect 2228 10848 2292 10852
rect 2308 10908 2372 10912
rect 2308 10852 2312 10908
rect 2312 10852 2368 10908
rect 2368 10852 2372 10908
rect 2308 10848 2372 10852
rect 5068 10908 5132 10912
rect 5068 10852 5072 10908
rect 5072 10852 5128 10908
rect 5128 10852 5132 10908
rect 5068 10848 5132 10852
rect 5148 10908 5212 10912
rect 5148 10852 5152 10908
rect 5152 10852 5208 10908
rect 5208 10852 5212 10908
rect 5148 10848 5212 10852
rect 5228 10908 5292 10912
rect 5228 10852 5232 10908
rect 5232 10852 5288 10908
rect 5288 10852 5292 10908
rect 5228 10848 5292 10852
rect 5308 10908 5372 10912
rect 5308 10852 5312 10908
rect 5312 10852 5368 10908
rect 5368 10852 5372 10908
rect 5308 10848 5372 10852
rect 3568 10364 3632 10368
rect 3568 10308 3572 10364
rect 3572 10308 3628 10364
rect 3628 10308 3632 10364
rect 3568 10304 3632 10308
rect 3648 10364 3712 10368
rect 3648 10308 3652 10364
rect 3652 10308 3708 10364
rect 3708 10308 3712 10364
rect 3648 10304 3712 10308
rect 3728 10364 3792 10368
rect 3728 10308 3732 10364
rect 3732 10308 3788 10364
rect 3788 10308 3792 10364
rect 3728 10304 3792 10308
rect 3808 10364 3872 10368
rect 3808 10308 3812 10364
rect 3812 10308 3868 10364
rect 3868 10308 3872 10364
rect 3808 10304 3872 10308
rect 2068 9820 2132 9824
rect 2068 9764 2072 9820
rect 2072 9764 2128 9820
rect 2128 9764 2132 9820
rect 2068 9760 2132 9764
rect 2148 9820 2212 9824
rect 2148 9764 2152 9820
rect 2152 9764 2208 9820
rect 2208 9764 2212 9820
rect 2148 9760 2212 9764
rect 2228 9820 2292 9824
rect 2228 9764 2232 9820
rect 2232 9764 2288 9820
rect 2288 9764 2292 9820
rect 2228 9760 2292 9764
rect 2308 9820 2372 9824
rect 2308 9764 2312 9820
rect 2312 9764 2368 9820
rect 2368 9764 2372 9820
rect 2308 9760 2372 9764
rect 5068 9820 5132 9824
rect 5068 9764 5072 9820
rect 5072 9764 5128 9820
rect 5128 9764 5132 9820
rect 5068 9760 5132 9764
rect 5148 9820 5212 9824
rect 5148 9764 5152 9820
rect 5152 9764 5208 9820
rect 5208 9764 5212 9820
rect 5148 9760 5212 9764
rect 5228 9820 5292 9824
rect 5228 9764 5232 9820
rect 5232 9764 5288 9820
rect 5288 9764 5292 9820
rect 5228 9760 5292 9764
rect 5308 9820 5372 9824
rect 5308 9764 5312 9820
rect 5312 9764 5368 9820
rect 5368 9764 5372 9820
rect 5308 9760 5372 9764
rect 3568 9276 3632 9280
rect 3568 9220 3572 9276
rect 3572 9220 3628 9276
rect 3628 9220 3632 9276
rect 3568 9216 3632 9220
rect 3648 9276 3712 9280
rect 3648 9220 3652 9276
rect 3652 9220 3708 9276
rect 3708 9220 3712 9276
rect 3648 9216 3712 9220
rect 3728 9276 3792 9280
rect 3728 9220 3732 9276
rect 3732 9220 3788 9276
rect 3788 9220 3792 9276
rect 3728 9216 3792 9220
rect 3808 9276 3872 9280
rect 3808 9220 3812 9276
rect 3812 9220 3868 9276
rect 3868 9220 3872 9276
rect 3808 9216 3872 9220
rect 2068 8732 2132 8736
rect 2068 8676 2072 8732
rect 2072 8676 2128 8732
rect 2128 8676 2132 8732
rect 2068 8672 2132 8676
rect 2148 8732 2212 8736
rect 2148 8676 2152 8732
rect 2152 8676 2208 8732
rect 2208 8676 2212 8732
rect 2148 8672 2212 8676
rect 2228 8732 2292 8736
rect 2228 8676 2232 8732
rect 2232 8676 2288 8732
rect 2288 8676 2292 8732
rect 2228 8672 2292 8676
rect 2308 8732 2372 8736
rect 2308 8676 2312 8732
rect 2312 8676 2368 8732
rect 2368 8676 2372 8732
rect 2308 8672 2372 8676
rect 5068 8732 5132 8736
rect 5068 8676 5072 8732
rect 5072 8676 5128 8732
rect 5128 8676 5132 8732
rect 5068 8672 5132 8676
rect 5148 8732 5212 8736
rect 5148 8676 5152 8732
rect 5152 8676 5208 8732
rect 5208 8676 5212 8732
rect 5148 8672 5212 8676
rect 5228 8732 5292 8736
rect 5228 8676 5232 8732
rect 5232 8676 5288 8732
rect 5288 8676 5292 8732
rect 5228 8672 5292 8676
rect 5308 8732 5372 8736
rect 5308 8676 5312 8732
rect 5312 8676 5368 8732
rect 5368 8676 5372 8732
rect 5308 8672 5372 8676
rect 3568 8188 3632 8192
rect 3568 8132 3572 8188
rect 3572 8132 3628 8188
rect 3628 8132 3632 8188
rect 3568 8128 3632 8132
rect 3648 8188 3712 8192
rect 3648 8132 3652 8188
rect 3652 8132 3708 8188
rect 3708 8132 3712 8188
rect 3648 8128 3712 8132
rect 3728 8188 3792 8192
rect 3728 8132 3732 8188
rect 3732 8132 3788 8188
rect 3788 8132 3792 8188
rect 3728 8128 3792 8132
rect 3808 8188 3872 8192
rect 3808 8132 3812 8188
rect 3812 8132 3868 8188
rect 3868 8132 3872 8188
rect 3808 8128 3872 8132
rect 2068 7644 2132 7648
rect 2068 7588 2072 7644
rect 2072 7588 2128 7644
rect 2128 7588 2132 7644
rect 2068 7584 2132 7588
rect 2148 7644 2212 7648
rect 2148 7588 2152 7644
rect 2152 7588 2208 7644
rect 2208 7588 2212 7644
rect 2148 7584 2212 7588
rect 2228 7644 2292 7648
rect 2228 7588 2232 7644
rect 2232 7588 2288 7644
rect 2288 7588 2292 7644
rect 2228 7584 2292 7588
rect 2308 7644 2372 7648
rect 2308 7588 2312 7644
rect 2312 7588 2368 7644
rect 2368 7588 2372 7644
rect 2308 7584 2372 7588
rect 5068 7644 5132 7648
rect 5068 7588 5072 7644
rect 5072 7588 5128 7644
rect 5128 7588 5132 7644
rect 5068 7584 5132 7588
rect 5148 7644 5212 7648
rect 5148 7588 5152 7644
rect 5152 7588 5208 7644
rect 5208 7588 5212 7644
rect 5148 7584 5212 7588
rect 5228 7644 5292 7648
rect 5228 7588 5232 7644
rect 5232 7588 5288 7644
rect 5288 7588 5292 7644
rect 5228 7584 5292 7588
rect 5308 7644 5372 7648
rect 5308 7588 5312 7644
rect 5312 7588 5368 7644
rect 5368 7588 5372 7644
rect 5308 7584 5372 7588
rect 3568 7100 3632 7104
rect 3568 7044 3572 7100
rect 3572 7044 3628 7100
rect 3628 7044 3632 7100
rect 3568 7040 3632 7044
rect 3648 7100 3712 7104
rect 3648 7044 3652 7100
rect 3652 7044 3708 7100
rect 3708 7044 3712 7100
rect 3648 7040 3712 7044
rect 3728 7100 3792 7104
rect 3728 7044 3732 7100
rect 3732 7044 3788 7100
rect 3788 7044 3792 7100
rect 3728 7040 3792 7044
rect 3808 7100 3872 7104
rect 3808 7044 3812 7100
rect 3812 7044 3868 7100
rect 3868 7044 3872 7100
rect 3808 7040 3872 7044
rect 2068 6556 2132 6560
rect 2068 6500 2072 6556
rect 2072 6500 2128 6556
rect 2128 6500 2132 6556
rect 2068 6496 2132 6500
rect 2148 6556 2212 6560
rect 2148 6500 2152 6556
rect 2152 6500 2208 6556
rect 2208 6500 2212 6556
rect 2148 6496 2212 6500
rect 2228 6556 2292 6560
rect 2228 6500 2232 6556
rect 2232 6500 2288 6556
rect 2288 6500 2292 6556
rect 2228 6496 2292 6500
rect 2308 6556 2372 6560
rect 2308 6500 2312 6556
rect 2312 6500 2368 6556
rect 2368 6500 2372 6556
rect 2308 6496 2372 6500
rect 5068 6556 5132 6560
rect 5068 6500 5072 6556
rect 5072 6500 5128 6556
rect 5128 6500 5132 6556
rect 5068 6496 5132 6500
rect 5148 6556 5212 6560
rect 5148 6500 5152 6556
rect 5152 6500 5208 6556
rect 5208 6500 5212 6556
rect 5148 6496 5212 6500
rect 5228 6556 5292 6560
rect 5228 6500 5232 6556
rect 5232 6500 5288 6556
rect 5288 6500 5292 6556
rect 5228 6496 5292 6500
rect 5308 6556 5372 6560
rect 5308 6500 5312 6556
rect 5312 6500 5368 6556
rect 5368 6500 5372 6556
rect 5308 6496 5372 6500
rect 3568 6012 3632 6016
rect 3568 5956 3572 6012
rect 3572 5956 3628 6012
rect 3628 5956 3632 6012
rect 3568 5952 3632 5956
rect 3648 6012 3712 6016
rect 3648 5956 3652 6012
rect 3652 5956 3708 6012
rect 3708 5956 3712 6012
rect 3648 5952 3712 5956
rect 3728 6012 3792 6016
rect 3728 5956 3732 6012
rect 3732 5956 3788 6012
rect 3788 5956 3792 6012
rect 3728 5952 3792 5956
rect 3808 6012 3872 6016
rect 3808 5956 3812 6012
rect 3812 5956 3868 6012
rect 3868 5956 3872 6012
rect 3808 5952 3872 5956
rect 2068 5468 2132 5472
rect 2068 5412 2072 5468
rect 2072 5412 2128 5468
rect 2128 5412 2132 5468
rect 2068 5408 2132 5412
rect 2148 5468 2212 5472
rect 2148 5412 2152 5468
rect 2152 5412 2208 5468
rect 2208 5412 2212 5468
rect 2148 5408 2212 5412
rect 2228 5468 2292 5472
rect 2228 5412 2232 5468
rect 2232 5412 2288 5468
rect 2288 5412 2292 5468
rect 2228 5408 2292 5412
rect 2308 5468 2372 5472
rect 2308 5412 2312 5468
rect 2312 5412 2368 5468
rect 2368 5412 2372 5468
rect 2308 5408 2372 5412
rect 5068 5468 5132 5472
rect 5068 5412 5072 5468
rect 5072 5412 5128 5468
rect 5128 5412 5132 5468
rect 5068 5408 5132 5412
rect 5148 5468 5212 5472
rect 5148 5412 5152 5468
rect 5152 5412 5208 5468
rect 5208 5412 5212 5468
rect 5148 5408 5212 5412
rect 5228 5468 5292 5472
rect 5228 5412 5232 5468
rect 5232 5412 5288 5468
rect 5288 5412 5292 5468
rect 5228 5408 5292 5412
rect 5308 5468 5372 5472
rect 5308 5412 5312 5468
rect 5312 5412 5368 5468
rect 5368 5412 5372 5468
rect 5308 5408 5372 5412
rect 3568 4924 3632 4928
rect 3568 4868 3572 4924
rect 3572 4868 3628 4924
rect 3628 4868 3632 4924
rect 3568 4864 3632 4868
rect 3648 4924 3712 4928
rect 3648 4868 3652 4924
rect 3652 4868 3708 4924
rect 3708 4868 3712 4924
rect 3648 4864 3712 4868
rect 3728 4924 3792 4928
rect 3728 4868 3732 4924
rect 3732 4868 3788 4924
rect 3788 4868 3792 4924
rect 3728 4864 3792 4868
rect 3808 4924 3872 4928
rect 3808 4868 3812 4924
rect 3812 4868 3868 4924
rect 3868 4868 3872 4924
rect 3808 4864 3872 4868
rect 2068 4380 2132 4384
rect 2068 4324 2072 4380
rect 2072 4324 2128 4380
rect 2128 4324 2132 4380
rect 2068 4320 2132 4324
rect 2148 4380 2212 4384
rect 2148 4324 2152 4380
rect 2152 4324 2208 4380
rect 2208 4324 2212 4380
rect 2148 4320 2212 4324
rect 2228 4380 2292 4384
rect 2228 4324 2232 4380
rect 2232 4324 2288 4380
rect 2288 4324 2292 4380
rect 2228 4320 2292 4324
rect 2308 4380 2372 4384
rect 2308 4324 2312 4380
rect 2312 4324 2368 4380
rect 2368 4324 2372 4380
rect 2308 4320 2372 4324
rect 5068 4380 5132 4384
rect 5068 4324 5072 4380
rect 5072 4324 5128 4380
rect 5128 4324 5132 4380
rect 5068 4320 5132 4324
rect 5148 4380 5212 4384
rect 5148 4324 5152 4380
rect 5152 4324 5208 4380
rect 5208 4324 5212 4380
rect 5148 4320 5212 4324
rect 5228 4380 5292 4384
rect 5228 4324 5232 4380
rect 5232 4324 5288 4380
rect 5288 4324 5292 4380
rect 5228 4320 5292 4324
rect 5308 4380 5372 4384
rect 5308 4324 5312 4380
rect 5312 4324 5368 4380
rect 5368 4324 5372 4380
rect 5308 4320 5372 4324
rect 3568 3836 3632 3840
rect 3568 3780 3572 3836
rect 3572 3780 3628 3836
rect 3628 3780 3632 3836
rect 3568 3776 3632 3780
rect 3648 3836 3712 3840
rect 3648 3780 3652 3836
rect 3652 3780 3708 3836
rect 3708 3780 3712 3836
rect 3648 3776 3712 3780
rect 3728 3836 3792 3840
rect 3728 3780 3732 3836
rect 3732 3780 3788 3836
rect 3788 3780 3792 3836
rect 3728 3776 3792 3780
rect 3808 3836 3872 3840
rect 3808 3780 3812 3836
rect 3812 3780 3868 3836
rect 3868 3780 3872 3836
rect 3808 3776 3872 3780
rect 2068 3292 2132 3296
rect 2068 3236 2072 3292
rect 2072 3236 2128 3292
rect 2128 3236 2132 3292
rect 2068 3232 2132 3236
rect 2148 3292 2212 3296
rect 2148 3236 2152 3292
rect 2152 3236 2208 3292
rect 2208 3236 2212 3292
rect 2148 3232 2212 3236
rect 2228 3292 2292 3296
rect 2228 3236 2232 3292
rect 2232 3236 2288 3292
rect 2288 3236 2292 3292
rect 2228 3232 2292 3236
rect 2308 3292 2372 3296
rect 2308 3236 2312 3292
rect 2312 3236 2368 3292
rect 2368 3236 2372 3292
rect 2308 3232 2372 3236
rect 5068 3292 5132 3296
rect 5068 3236 5072 3292
rect 5072 3236 5128 3292
rect 5128 3236 5132 3292
rect 5068 3232 5132 3236
rect 5148 3292 5212 3296
rect 5148 3236 5152 3292
rect 5152 3236 5208 3292
rect 5208 3236 5212 3292
rect 5148 3232 5212 3236
rect 5228 3292 5292 3296
rect 5228 3236 5232 3292
rect 5232 3236 5288 3292
rect 5288 3236 5292 3292
rect 5228 3232 5292 3236
rect 5308 3292 5372 3296
rect 5308 3236 5312 3292
rect 5312 3236 5368 3292
rect 5368 3236 5372 3292
rect 5308 3232 5372 3236
rect 3568 2748 3632 2752
rect 3568 2692 3572 2748
rect 3572 2692 3628 2748
rect 3628 2692 3632 2748
rect 3568 2688 3632 2692
rect 3648 2748 3712 2752
rect 3648 2692 3652 2748
rect 3652 2692 3708 2748
rect 3708 2692 3712 2748
rect 3648 2688 3712 2692
rect 3728 2748 3792 2752
rect 3728 2692 3732 2748
rect 3732 2692 3788 2748
rect 3788 2692 3792 2748
rect 3728 2688 3792 2692
rect 3808 2748 3872 2752
rect 3808 2692 3812 2748
rect 3812 2692 3868 2748
rect 3868 2692 3872 2748
rect 3808 2688 3872 2692
rect 2068 2204 2132 2208
rect 2068 2148 2072 2204
rect 2072 2148 2128 2204
rect 2128 2148 2132 2204
rect 2068 2144 2132 2148
rect 2148 2204 2212 2208
rect 2148 2148 2152 2204
rect 2152 2148 2208 2204
rect 2208 2148 2212 2204
rect 2148 2144 2212 2148
rect 2228 2204 2292 2208
rect 2228 2148 2232 2204
rect 2232 2148 2288 2204
rect 2288 2148 2292 2204
rect 2228 2144 2292 2148
rect 2308 2204 2372 2208
rect 2308 2148 2312 2204
rect 2312 2148 2368 2204
rect 2368 2148 2372 2204
rect 2308 2144 2372 2148
rect 5068 2204 5132 2208
rect 5068 2148 5072 2204
rect 5072 2148 5128 2204
rect 5128 2148 5132 2204
rect 5068 2144 5132 2148
rect 5148 2204 5212 2208
rect 5148 2148 5152 2204
rect 5152 2148 5208 2204
rect 5208 2148 5212 2204
rect 5148 2144 5212 2148
rect 5228 2204 5292 2208
rect 5228 2148 5232 2204
rect 5232 2148 5288 2204
rect 5288 2148 5292 2204
rect 5228 2144 5292 2148
rect 5308 2204 5372 2208
rect 5308 2148 5312 2204
rect 5312 2148 5368 2204
rect 5368 2148 5372 2204
rect 5308 2144 5372 2148
<< metal4 >>
rect -1620 13922 -1300 13964
rect -1620 13686 -1578 13922
rect -1342 13686 -1300 13922
rect -1620 11464 -1300 13686
rect -1620 11386 -1606 11464
rect -1318 11386 -1300 11464
rect -1620 9694 -1300 11386
rect -1620 9458 -1578 9694
rect -1342 9458 -1300 9694
rect -1620 6494 -1300 9458
rect -1620 6258 -1578 6494
rect -1342 6258 -1300 6494
rect -1620 -86 -1300 6258
rect -960 13262 -640 13304
rect -960 13026 -918 13262
rect -682 13026 -640 13262
rect -960 10918 -640 13026
rect 2960 13262 3280 13964
rect 2960 13026 3002 13262
rect 3238 13026 3280 13262
rect -960 10844 -948 10918
rect -658 10844 -640 10918
rect -960 8094 -640 10844
rect -960 7858 -918 8094
rect -682 7858 -640 8094
rect -960 4894 -640 7858
rect -960 4658 -918 4894
rect -682 4658 -640 4894
rect -960 574 -640 4658
rect -300 12602 20 12644
rect -300 12366 -258 12602
rect -22 12366 20 12602
rect -300 8794 20 12366
rect -300 8558 -258 8794
rect -22 8558 20 8794
rect -300 5594 20 8558
rect -300 5358 -258 5594
rect -22 5358 20 5594
rect -300 1234 20 5358
rect 360 11942 680 11984
rect 360 11706 402 11942
rect 638 11706 680 11942
rect 360 10394 680 11706
rect 360 10158 402 10394
rect 638 10158 680 10394
rect 360 7194 680 10158
rect 360 6958 402 7194
rect 638 6958 680 7194
rect 360 3994 680 6958
rect 360 3758 402 3994
rect 638 3758 680 3994
rect 360 1894 680 3758
rect 360 1658 402 1894
rect 638 1658 680 1894
rect 360 1616 680 1658
rect 2060 11942 2380 12644
rect 2060 11706 2102 11942
rect 2338 11706 2380 11942
rect 2060 10912 2380 11706
rect 2060 10848 2068 10912
rect 2132 10848 2148 10912
rect 2212 10848 2228 10912
rect 2292 10848 2308 10912
rect 2372 10848 2380 10912
rect 2060 10394 2380 10848
rect 2060 10158 2102 10394
rect 2338 10158 2380 10394
rect 2060 9824 2380 10158
rect 2060 9760 2068 9824
rect 2132 9760 2148 9824
rect 2212 9760 2228 9824
rect 2292 9760 2308 9824
rect 2372 9760 2380 9824
rect 2060 8736 2380 9760
rect 2060 8672 2068 8736
rect 2132 8672 2148 8736
rect 2212 8672 2228 8736
rect 2292 8672 2308 8736
rect 2372 8672 2380 8736
rect 2060 7648 2380 8672
rect 2060 7584 2068 7648
rect 2132 7584 2148 7648
rect 2212 7584 2228 7648
rect 2292 7584 2308 7648
rect 2372 7584 2380 7648
rect 2060 7194 2380 7584
rect 2060 6958 2102 7194
rect 2338 6958 2380 7194
rect 2060 6560 2380 6958
rect 2060 6496 2068 6560
rect 2132 6496 2148 6560
rect 2212 6496 2228 6560
rect 2292 6496 2308 6560
rect 2372 6496 2380 6560
rect 2060 5472 2380 6496
rect 2060 5408 2068 5472
rect 2132 5408 2148 5472
rect 2212 5408 2228 5472
rect 2292 5408 2308 5472
rect 2372 5408 2380 5472
rect 2060 4384 2380 5408
rect 2060 4320 2068 4384
rect 2132 4320 2148 4384
rect 2212 4320 2228 4384
rect 2292 4320 2308 4384
rect 2372 4320 2380 4384
rect 2060 3994 2380 4320
rect 2060 3758 2102 3994
rect 2338 3758 2380 3994
rect 2060 3296 2380 3758
rect 2060 3232 2068 3296
rect 2132 3232 2148 3296
rect 2212 3232 2228 3296
rect 2292 3232 2308 3296
rect 2372 3232 2380 3296
rect 2060 2208 2380 3232
rect 2060 2144 2068 2208
rect 2132 2144 2148 2208
rect 2212 2144 2228 2208
rect 2292 2144 2308 2208
rect 2372 2144 2380 2208
rect 2060 1894 2380 2144
rect 2060 1658 2102 1894
rect 2338 1658 2380 1894
rect -300 998 -258 1234
rect -22 998 20 1234
rect -300 956 20 998
rect 2060 956 2380 1658
rect 2960 8094 3280 13026
rect 4460 13922 4780 13964
rect 4460 13686 4502 13922
rect 4738 13686 4780 13922
rect 2960 7858 3002 8094
rect 3238 7858 3280 8094
rect 2960 4894 3280 7858
rect 2960 4658 3002 4894
rect 3238 4658 3280 4894
rect -960 338 -918 574
rect -682 338 -640 574
rect -960 296 -640 338
rect 2960 574 3280 4658
rect 3560 12602 3880 12644
rect 3560 12366 3602 12602
rect 3838 12366 3880 12602
rect 3560 11456 3880 12366
rect 3560 11392 3568 11456
rect 3632 11392 3648 11456
rect 3712 11392 3728 11456
rect 3792 11392 3808 11456
rect 3872 11392 3880 11456
rect 3560 10368 3880 11392
rect 3560 10304 3568 10368
rect 3632 10304 3648 10368
rect 3712 10304 3728 10368
rect 3792 10304 3808 10368
rect 3872 10304 3880 10368
rect 3560 9280 3880 10304
rect 3560 9216 3568 9280
rect 3632 9216 3648 9280
rect 3712 9216 3728 9280
rect 3792 9216 3808 9280
rect 3872 9216 3880 9280
rect 3560 8794 3880 9216
rect 3560 8558 3602 8794
rect 3838 8558 3880 8794
rect 3560 8192 3880 8558
rect 3560 8128 3568 8192
rect 3632 8128 3648 8192
rect 3712 8128 3728 8192
rect 3792 8128 3808 8192
rect 3872 8128 3880 8192
rect 3560 7104 3880 8128
rect 3560 7040 3568 7104
rect 3632 7040 3648 7104
rect 3712 7040 3728 7104
rect 3792 7040 3808 7104
rect 3872 7040 3880 7104
rect 3560 6016 3880 7040
rect 3560 5952 3568 6016
rect 3632 5952 3648 6016
rect 3712 5952 3728 6016
rect 3792 5952 3808 6016
rect 3872 5952 3880 6016
rect 3560 5594 3880 5952
rect 3560 5358 3602 5594
rect 3838 5358 3880 5594
rect 3560 4928 3880 5358
rect 3560 4864 3568 4928
rect 3632 4864 3648 4928
rect 3712 4864 3728 4928
rect 3792 4864 3808 4928
rect 3872 4864 3880 4928
rect 3560 3840 3880 4864
rect 3560 3776 3568 3840
rect 3632 3776 3648 3840
rect 3712 3776 3728 3840
rect 3792 3776 3808 3840
rect 3872 3776 3880 3840
rect 3560 2752 3880 3776
rect 3560 2688 3568 2752
rect 3632 2688 3648 2752
rect 3712 2688 3728 2752
rect 3792 2688 3808 2752
rect 3872 2688 3880 2752
rect 3560 1234 3880 2688
rect 3560 998 3602 1234
rect 3838 998 3880 1234
rect 3560 956 3880 998
rect 4460 9694 4780 13686
rect 5960 13262 6280 13964
rect 9304 13922 9624 13964
rect 9304 13686 9346 13922
rect 9582 13686 9624 13922
rect 5960 13026 6002 13262
rect 6238 13026 6280 13262
rect 4460 9458 4502 9694
rect 4738 9458 4780 9694
rect 4460 6494 4780 9458
rect 4460 6258 4502 6494
rect 4738 6258 4780 6494
rect 2960 338 3002 574
rect 3238 338 3280 574
rect -1620 -322 -1578 -86
rect -1342 -322 -1300 -86
rect -1620 -364 -1300 -322
rect 2960 -364 3280 338
rect 4460 -86 4780 6258
rect 5060 11942 5380 12644
rect 5060 11706 5102 11942
rect 5338 11706 5380 11942
rect 5060 10912 5380 11706
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 10394 5380 10848
rect 5060 10158 5102 10394
rect 5338 10158 5380 10394
rect 5060 9824 5380 10158
rect 5060 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5380 9824
rect 5060 8736 5380 9760
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 7648 5380 8672
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 7194 5380 7584
rect 5060 6958 5102 7194
rect 5338 6958 5380 7194
rect 5060 6560 5380 6958
rect 5060 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5380 6560
rect 5060 5472 5380 6496
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 4384 5380 5408
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 3994 5380 4320
rect 5060 3758 5102 3994
rect 5338 3758 5380 3994
rect 5060 3296 5380 3758
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 5060 2208 5380 3232
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 1894 5380 2144
rect 5060 1658 5102 1894
rect 5338 1658 5380 1894
rect 5060 956 5380 1658
rect 5960 8094 6280 13026
rect 8644 13262 8964 13304
rect 8644 13026 8686 13262
rect 8922 13026 8964 13262
rect 7984 12602 8304 12644
rect 7984 12366 8026 12602
rect 8262 12366 8304 12602
rect 5960 7858 6002 8094
rect 6238 7858 6280 8094
rect 5960 4894 6280 7858
rect 5960 4658 6002 4894
rect 6238 4658 6280 4894
rect 4460 -322 4502 -86
rect 4738 -322 4780 -86
rect 4460 -364 4780 -322
rect 5960 574 6280 4658
rect 7324 11942 7644 11984
rect 7324 11706 7366 11942
rect 7602 11706 7644 11942
rect 7324 10394 7644 11706
rect 7324 10158 7366 10394
rect 7602 10158 7644 10394
rect 7324 7194 7644 10158
rect 7324 6958 7366 7194
rect 7602 6958 7644 7194
rect 7324 3994 7644 6958
rect 7324 3758 7366 3994
rect 7602 3758 7644 3994
rect 7324 1894 7644 3758
rect 7324 1658 7366 1894
rect 7602 1658 7644 1894
rect 7324 1616 7644 1658
rect 7984 8794 8304 12366
rect 7984 8558 8026 8794
rect 8262 8558 8304 8794
rect 7984 5594 8304 8558
rect 7984 5358 8026 5594
rect 8262 5358 8304 5594
rect 7984 1234 8304 5358
rect 7984 998 8026 1234
rect 8262 998 8304 1234
rect 7984 956 8304 998
rect 8644 8094 8964 13026
rect 8644 7858 8686 8094
rect 8922 7858 8964 8094
rect 8644 4894 8964 7858
rect 8644 4658 8686 4894
rect 8922 4658 8964 4894
rect 5960 338 6002 574
rect 6238 338 6280 574
rect 5960 -364 6280 338
rect 8644 574 8964 4658
rect 8644 338 8686 574
rect 8922 338 8964 574
rect 8644 296 8964 338
rect 9304 9694 9624 13686
rect 9304 9458 9346 9694
rect 9582 9458 9624 9694
rect 9304 6494 9624 9458
rect 9304 6258 9346 6494
rect 9582 6258 9624 6494
rect 9304 -86 9624 6258
rect 9304 -322 9346 -86
rect 9582 -322 9624 -86
rect 9304 -364 9624 -322
<< via4 >>
rect -1578 13686 -1342 13922
rect -1578 9458 -1342 9694
rect -1578 6258 -1342 6494
rect -918 13026 -682 13262
rect 3002 13026 3238 13262
rect -918 7858 -682 8094
rect -918 4658 -682 4894
rect -258 12366 -22 12602
rect -258 8558 -22 8794
rect -258 5358 -22 5594
rect 402 11706 638 11942
rect 402 10158 638 10394
rect 402 6958 638 7194
rect 402 3758 638 3994
rect 402 1658 638 1894
rect 2102 11706 2338 11942
rect 2102 10158 2338 10394
rect 2102 6958 2338 7194
rect 2102 3758 2338 3994
rect 2102 1658 2338 1894
rect -258 998 -22 1234
rect 4502 13686 4738 13922
rect 3002 7858 3238 8094
rect 3002 4658 3238 4894
rect -918 338 -682 574
rect 3602 12366 3838 12602
rect 3602 8558 3838 8794
rect 3602 5358 3838 5594
rect 3602 998 3838 1234
rect 9346 13686 9582 13922
rect 6002 13026 6238 13262
rect 4502 9458 4738 9694
rect 4502 6258 4738 6494
rect 3002 338 3238 574
rect -1578 -322 -1342 -86
rect 5102 11706 5338 11942
rect 5102 10158 5338 10394
rect 5102 6958 5338 7194
rect 5102 3758 5338 3994
rect 5102 1658 5338 1894
rect 8686 13026 8922 13262
rect 8026 12366 8262 12602
rect 6002 7858 6238 8094
rect 6002 4658 6238 4894
rect 4502 -322 4738 -86
rect 7366 11706 7602 11942
rect 7366 10158 7602 10394
rect 7366 6958 7602 7194
rect 7366 3758 7602 3994
rect 7366 1658 7602 1894
rect 8026 8558 8262 8794
rect 8026 5358 8262 5594
rect 8026 998 8262 1234
rect 8686 7858 8922 8094
rect 8686 4658 8922 4894
rect 6002 338 6238 574
rect 8686 338 8922 574
rect 9346 9458 9582 9694
rect 9346 6258 9582 6494
rect 9346 -322 9582 -86
<< metal5 >>
rect -1620 13922 9624 13964
rect -1620 13686 -1578 13922
rect -1342 13686 4502 13922
rect 4738 13686 9346 13922
rect 9582 13686 9624 13922
rect -1620 13644 9624 13686
rect -960 13262 8964 13304
rect -960 13026 -918 13262
rect -682 13026 3002 13262
rect 3238 13026 6002 13262
rect 6238 13026 8686 13262
rect 8922 13026 8964 13262
rect -960 12984 8964 13026
rect -300 12602 8304 12644
rect -300 12366 -258 12602
rect -22 12366 3602 12602
rect 3838 12366 8026 12602
rect 8262 12366 8304 12602
rect -300 12324 8304 12366
rect 360 11942 7644 11984
rect 360 11706 402 11942
rect 638 11706 2102 11942
rect 2338 11706 5102 11942
rect 5338 11706 7366 11942
rect 7602 11706 7644 11942
rect 360 11664 7644 11706
rect -300 10394 8304 10436
rect -300 10158 402 10394
rect 638 10158 2102 10394
rect 2338 10158 5102 10394
rect 5338 10158 7366 10394
rect 7602 10158 8304 10394
rect -300 10116 8304 10158
rect -1620 9694 9624 9736
rect -1620 9458 -1578 9694
rect -1342 9458 4502 9694
rect 4738 9458 9346 9694
rect 9582 9458 9624 9694
rect -1620 9416 9624 9458
rect -300 8794 8304 8836
rect -300 8558 -258 8794
rect -22 8558 3602 8794
rect 3838 8558 8026 8794
rect 8262 8558 8304 8794
rect -300 8516 8304 8558
rect -1620 8094 9624 8136
rect -1620 7858 -918 8094
rect -682 7858 3002 8094
rect 3238 7858 6002 8094
rect 6238 7858 8686 8094
rect 8922 7858 9624 8094
rect -1620 7816 9624 7858
rect -300 7194 8304 7236
rect -300 6958 402 7194
rect 638 6958 2102 7194
rect 2338 6958 5102 7194
rect 5338 6958 7366 7194
rect 7602 6958 8304 7194
rect -300 6916 8304 6958
rect -1620 6494 9624 6536
rect -1620 6258 -1578 6494
rect -1342 6258 4502 6494
rect 4738 6258 9346 6494
rect 9582 6258 9624 6494
rect -1620 6216 9624 6258
rect -300 5594 8304 5636
rect -300 5358 -258 5594
rect -22 5358 3602 5594
rect 3838 5358 8026 5594
rect 8262 5358 8304 5594
rect -300 5316 8304 5358
rect -1620 4894 9624 4936
rect -1620 4658 -918 4894
rect -682 4658 3002 4894
rect 3238 4658 6002 4894
rect 6238 4658 8686 4894
rect 8922 4658 9624 4894
rect -1620 4616 9624 4658
rect -300 3994 8304 4036
rect -300 3758 402 3994
rect 638 3758 2102 3994
rect 2338 3758 5102 3994
rect 5338 3758 7366 3994
rect 7602 3758 8304 3994
rect -300 3716 8304 3758
rect 360 1894 7644 1936
rect 360 1658 402 1894
rect 638 1658 2102 1894
rect 2338 1658 5102 1894
rect 5338 1658 7366 1894
rect 7602 1658 7644 1894
rect 360 1616 7644 1658
rect -300 1234 8304 1276
rect -300 998 -258 1234
rect -22 998 3602 1234
rect 3838 998 8026 1234
rect 8262 998 8304 1234
rect -300 956 8304 998
rect -960 574 8964 616
rect -960 338 -918 574
rect -682 338 3002 574
rect 3238 338 6002 574
rect 6238 338 8686 574
rect 8922 338 8964 574
rect -960 296 8964 338
rect -1620 -86 9624 -44
rect -1620 -322 -1578 -86
rect -1342 -322 4502 -86
rect 4738 -322 9346 -86
rect 9582 -322 9624 -86
rect -1620 -364 9624 -322
use sky130_fd_sc_hd__dfrtp_4  _096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 1656 0 1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _108_
timestamp 1608231460
transform 1 0 1656 0 -1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 920 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608231460
transform 1 0 920 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 1196 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 1564 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1608231460
transform 1 0 1196 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1608231460
transform 1 0 1564 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _056_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1608231460
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _091_
timestamp 1608231460
transform 1 0 4508 0 -1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_4  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 4508 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 4232 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1608231460
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36
timestamp 1608231460
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608231460
transform -1 0 7084 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608231460
transform -1 0 7084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1608231460
transform 1 0 6624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1608231460
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_63
timestamp 1608231460
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1608231460
transform 1 0 2208 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _094_
timestamp 1608231460
transform 1 0 2576 0 -1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608231460
transform 1 0 920 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 1196 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_11
timestamp 1608231460
transform 1 0 1932 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1608231460
transform 1 0 4692 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 5060 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 5704 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608231460
transform -1 0 7084 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1608231460
transform 1 0 6532 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _104_
timestamp 1608231460
transform 1 0 1196 0 1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608231460
transform 1 0 920 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1608231460
transform 1 0 3312 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _105_
timestamp 1608231460
transform 1 0 3864 0 1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1608231460
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_30
timestamp 1608231460
transform 1 0 3680 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 5980 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608231460
transform -1 0 7084 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _045_
timestamp 1608231460
transform 1 0 2208 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _046_
timestamp 1608231460
transform 1 0 1840 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _048_
timestamp 1608231460
transform 1 0 1472 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _095_
timestamp 1608231460
transform 1 0 2576 0 -1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608231460
transform 1 0 920 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 1196 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 4692 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608231460
transform -1 0 7084 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1608231460
transform 1 0 6532 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_62
timestamp 1608231460
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _103_
timestamp 1608231460
transform 1 0 1196 0 1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608231460
transform 1 0 920 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _042_
timestamp 1608231460
transform 1 0 3312 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _043_
timestamp 1608231460
transform 1 0 3956 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_4  _093_
timestamp 1608231460
transform 1 0 4600 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1608231460
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_30
timestamp 1608231460
transform 1 0 3680 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_32
timestamp 1608231460
transform 1 0 3864 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_37
timestamp 1608231460
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608231460
transform -1 0 7084 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _101_
timestamp 1608231460
transform 1 0 1196 0 1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _102_
timestamp 1608231460
transform 1 0 1196 0 -1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608231460
transform 1 0 920 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608231460
transform 1 0 920 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _044_
timestamp 1608231460
transform 1 0 3864 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608231460
transform 1 0 3404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _089_
timestamp 1608231460
transform 1 0 4324 0 1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _106_
timestamp 1608231460
transform 1 0 3312 0 -1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1608231460
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_49
timestamp 1608231460
transform 1 0 5428 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_26
timestamp 1608231460
transform 1 0 3312 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_36
timestamp 1608231460
transform 1 0 4232 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1608231460
transform 1 0 5520 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1608231460
transform 1 0 6440 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1608231460
transform 1 0 5888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 6256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608231460
transform -1 0 7084 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608231460
transform -1 0 7084 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1608231460
transform 1 0 6532 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_62
timestamp 1608231460
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _049_
timestamp 1608231460
transform 1 0 1840 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _050_
timestamp 1608231460
transform 1 0 2208 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _088_
timestamp 1608231460
transform 1 0 2944 0 -1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608231460
transform 1 0 920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 1196 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1608231460
transform 1 0 1748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_18
timestamp 1608231460
transform 1 0 2576 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1608231460
transform 1 0 5060 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_49
timestamp 1608231460
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _083_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 5704 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608231460
transform -1 0 7084 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1608231460
transform 1 0 6532 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_62
timestamp 1608231460
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _100_
timestamp 1608231460
transform 1 0 1196 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608231460
transform 1 0 920 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1608231460
transform 1 0 3404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _107_
timestamp 1608231460
transform 1 0 3864 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1608231460
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_26
timestamp 1608231460
transform 1 0 3312 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608231460
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608231460
transform -1 0 7084 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_55
timestamp 1608231460
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_63
timestamp 1608231460
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _047_
timestamp 1608231460
transform 1 0 1656 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _051_
timestamp 1608231460
transform 1 0 1288 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _085_
timestamp 1608231460
transform 1 0 2024 0 -1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608231460
transform 1 0 920 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1608231460
transform 1 0 1196 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _090_
timestamp 1608231460
transform 1 0 4140 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608231460
transform -1 0 7084 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1608231460
transform 1 0 6532 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1608231460
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_62
timestamp 1608231460
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _099_
timestamp 1608231460
transform 1 0 1196 0 1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608231460
transform 1 0 920 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _041_
timestamp 1608231460
transform 1 0 3956 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _053_
timestamp 1608231460
transform 1 0 3312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _109_
timestamp 1608231460
transform 1 0 4324 0 1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1608231460
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_30
timestamp 1608231460
transform 1 0 3680 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_32
timestamp 1608231460
transform 1 0 3864 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608231460
transform 1 0 6440 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608231460
transform -1 0 7084 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _052_
timestamp 1608231460
transform 1 0 1932 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608231460
transform 1 0 2576 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _086_
timestamp 1608231460
transform 1 0 2944 0 -1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608231460
transform 1 0 920 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_serial_clock
timestamp 1608231460
transform 1 0 2300 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1608231460
transform 1 0 1196 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _040_
timestamp 1608231460
transform 1 0 5060 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _072_
timestamp 1608231460
transform 1 0 6256 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608231460
transform -1 0 7084 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1608231460
transform 1 0 6532 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_52
timestamp 1608231460
transform 1 0 5704 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_62
timestamp 1608231460
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 2208 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_4  _097_
timestamp 1608231460
transform 1 0 1472 0 -1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608231460
transform 1 0 920 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608231460
transform 1 0 920 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1608231460
transform 1 0 1196 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_11
timestamp 1608231460
transform 1 0 1932 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1608231460
transform 1 0 1196 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1608231460
transform 1 0 4048 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_4  _084_
timestamp 1608231460
transform 1 0 3588 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_4  _087_
timestamp 1608231460
transform 1 0 4416 0 1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1608231460
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_32
timestamp 1608231460
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1608231460
transform 1 0 5796 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608231460
transform 1 0 6164 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _079_
timestamp 1608231460
transform 1 0 6532 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608231460
transform -1 0 7084 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608231460
transform -1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1608231460
transform 1 0 6532 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_62
timestamp 1608231460
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _098_
timestamp 1608231460
transform 1 0 1656 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608231460
transform 1 0 920 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1608231460
transform 1 0 1196 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1608231460
transform 1 0 1564 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _054_
timestamp 1608231460
transform 1 0 3864 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 4416 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 5152 0 1 10336
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1608231460
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1608231460
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_45
timestamp 1608231460
transform 1 0 5060 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608231460
transform -1 0 7084 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608231460
transform 1 0 1196 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _055_
timestamp 1608231460
transform 1 0 2852 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608231460
transform 1 0 1472 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_18
timestamp 1608231460
transform 1 0 2576 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_4  _073_
timestamp 1608231460
transform 1 0 5060 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _080_
timestamp 1608231460
transform 1 0 4692 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1608231460
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_25
timestamp 1608231460
transform 1 0 3220 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_32
timestamp 1608231460
transform 1 0 3864 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_40
timestamp 1608231460
transform 1 0 4600 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_44
timestamp 1608231460
transform 1 0 4968 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608231460
transform -1 0 7084 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1608231460
transform 1 0 6624 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_63
timestamp 1608231460
transform 1 0 6716 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1608231460
transform -1 0 460 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  gpio_logic_high
timestamp 1608231460
transform 1 0 92 0 -1 11424
box -38 -48 314 592
<< labels >>
rlabel metal3 s 14000 1096 34000 1216 6 mgmt_gpio_in
port 0 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 1 nsew signal input
rlabel metal3 s 14000 2184 34000 2304 6 mgmt_gpio_out
port 2 nsew signal input
rlabel metal3 s 14000 552 34000 672 6 one
port 3 nsew signal tristate
rlabel metal3 s 14000 2728 34000 2848 6 pad_gpio_ana_en
port 4 nsew signal tristate
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_pol
port 5 nsew signal tristate
rlabel metal3 s 14000 3816 34000 3936 6 pad_gpio_ana_sel
port 6 nsew signal tristate
rlabel metal3 s 14000 4360 34000 4480 6 pad_gpio_dm[0]
port 7 nsew signal tristate
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_dm[1]
port 8 nsew signal tristate
rlabel metal3 s 14000 5448 34000 5568 6 pad_gpio_dm[2]
port 9 nsew signal tristate
rlabel metal3 s 14000 5992 34000 6112 6 pad_gpio_holdover
port 10 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_ib_mode_sel
port 11 nsew signal tristate
rlabel metal3 s 14000 7080 34000 7200 6 pad_gpio_in
port 12 nsew signal input
rlabel metal3 s 14000 7624 34000 7744 6 pad_gpio_inenb
port 13 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 pad_gpio_out
port 14 nsew signal tristate
rlabel metal3 s 14000 8712 34000 8832 6 pad_gpio_outenb
port 15 nsew signal tristate
rlabel metal3 s 14000 9256 34000 9376 6 pad_gpio_slow_sel
port 16 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 pad_gpio_vtrip_sel
port 17 nsew signal tristate
rlabel metal3 s 14000 10344 34000 10464 6 resetn
port 18 nsew signal input
rlabel metal3 s 14000 10888 34000 11008 6 serial_clock
port 19 nsew signal input
rlabel metal3 s 14000 11432 34000 11552 6 serial_data_in
port 20 nsew signal input
rlabel metal3 s 14000 11976 34000 12096 6 serial_data_out
port 21 nsew signal tristate
rlabel metal3 s 14000 12520 34000 12640 6 user_gpio_in
port 22 nsew signal tristate
rlabel metal3 s 14000 13064 34000 13184 6 user_gpio_oeb
port 23 nsew signal input
rlabel metal3 s 14000 13608 34000 13728 6 user_gpio_out
port 24 nsew signal input
rlabel metal3 s 14000 144 34000 264 6 zero
port 25 nsew signal tristate
rlabel metal4 s 5060 956 5380 12644 6 vccd
port 26 nsew power bidirectional
rlabel metal4 s 2060 956 2380 12644 6 vccd
port 27 nsew power bidirectional
rlabel metal4 s 7324 1616 7644 11984 6 vccd
port 28 nsew power bidirectional
rlabel metal4 s 360 1616 680 11984 6 vccd
port 29 nsew power bidirectional
rlabel metal5 s 360 11664 7644 11984 6 vccd
port 30 nsew power bidirectional
rlabel metal5 s -300 10116 8304 10436 6 vccd
port 31 nsew power bidirectional
rlabel metal5 s -300 6916 8304 7236 6 vccd
port 32 nsew power bidirectional
rlabel metal5 s -300 3716 8304 4036 6 vccd
port 33 nsew power bidirectional
rlabel metal5 s 360 1616 7644 1936 6 vccd
port 34 nsew power bidirectional
rlabel metal4 s 7984 956 8304 12644 6 vssd
port 35 nsew ground bidirectional
rlabel metal4 s 3560 956 3880 12644 6 vssd
port 36 nsew ground bidirectional
rlabel metal4 s -300 956 20 12644 4 vssd
port 37 nsew ground bidirectional
rlabel metal5 s -300 12324 8304 12644 6 vssd
port 38 nsew ground bidirectional
rlabel metal5 s -300 8516 8304 8836 6 vssd
port 39 nsew ground bidirectional
rlabel metal5 s -300 5316 8304 5636 6 vssd
port 40 nsew ground bidirectional
rlabel metal5 s -300 956 8304 1276 6 vssd
port 41 nsew ground bidirectional
rlabel metal4 s 5960 -364 6280 13964 6 vccd1
port 42 nsew power bidirectional
rlabel metal4 s 2960 -364 3280 13964 6 vccd1
port 43 nsew power bidirectional
rlabel metal4 s 8644 296 8964 13304 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s -960 296 -640 13304 4 vccd1
port 45 nsew power bidirectional
rlabel metal5 s -960 12984 8964 13304 6 vccd1
port 46 nsew power bidirectional
rlabel metal5 s -1620 7816 9624 8136 6 vccd1
port 47 nsew power bidirectional
rlabel metal5 s -1620 4616 9624 4936 6 vccd1
port 48 nsew power bidirectional
rlabel metal5 s -960 296 8964 616 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 9304 -364 9624 13964 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 4460 -364 4780 13964 6 vssd1
port 51 nsew ground bidirectional
rlabel metal4 s -1620 -364 -1300 13964 4 vssd1
port 52 nsew ground bidirectional
rlabel metal5 s -1620 13644 9624 13964 6 vssd1
port 53 nsew ground bidirectional
rlabel metal5 s -1620 9416 9624 9736 6 vssd1
port 54 nsew ground bidirectional
rlabel metal5 s -1620 6216 9624 6536 6 vssd1
port 55 nsew ground bidirectional
rlabel metal5 s -1620 -364 9624 -44 8 vssd1
port 56 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 34000 14000
<< end >>
