VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1426.380000 2924.800000 1427.580000 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490000 3520.400000 2231.050000 3524.800000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730000 3520.400000 1906.290000 3524.800000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430000 3520.400000 1581.990000 3524.800000 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130000 3520.400000 1257.690000 3524.800000 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370000 3520.400000 932.930000 3524.800000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070000 3520.400000 608.630000 3524.800000 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770000 3520.400000 284.330000 3524.800000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3486.100000 -0.400000 3487.300000 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3224.980000 -0.400000 3226.180000 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2964.540000 -0.400000 2965.740000 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1692.260000 2924.800000 1693.460000 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2703.420000 -0.400000 2704.620000 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2442.980000 -0.400000 2444.180000 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2182.540000 -0.400000 2183.740000 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1921.420000 -0.400000 1922.620000 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1660.980000 -0.400000 1662.180000 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1399.860000 -0.400000 1401.060000 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1139.420000 -0.400000 1140.620000 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 878.980000 -0.400000 880.180000 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 617.860000 -0.400000 619.060000 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1958.140000 2924.800000 1959.340000 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2223.340000 2924.800000 2224.540000 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2489.220000 2924.800000 2490.420000 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2755.100000 2924.800000 2756.300000 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3020.300000 2924.800000 3021.500000 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3286.180000 2924.800000 3287.380000 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090000 3520.400000 2879.650000 3524.800000 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790000 3520.400000 2555.350000 3524.800000 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 32.380000 2924.800000 33.580000 ;
    END
  END io_in[0]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 98.340000 2924.800000 99.540000 ;
    END
  END io_out[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2289.980000 2924.800000 2291.180000 ;
    END
  END io_in[10]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2356.620000 2924.800000 2357.820000 ;
    END
  END io_out[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2555.860000 2924.800000 2557.060000 ;
    END
  END io_in[11]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2621.820000 2924.800000 2623.020000 ;
    END
  END io_out[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2821.060000 2924.800000 2822.260000 ;
    END
  END io_in[12]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2887.700000 2924.800000 2888.900000 ;
    END
  END io_out[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3086.940000 2924.800000 3088.140000 ;
    END
  END io_in[13]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3153.580000 2924.800000 3154.780000 ;
    END
  END io_out[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3352.820000 2924.800000 3354.020000 ;
    END
  END io_in[14]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3418.780000 2924.800000 3419.980000 ;
    END
  END io_out[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130000 3520.400000 2798.690000 3524.800000 ;
    END
  END io_in[15]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170000 3520.400000 2717.730000 3524.800000 ;
    END
  END io_out[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830000 3520.400000 2474.390000 3524.800000 ;
    END
  END io_in[16]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410000 3520.400000 2392.970000 3524.800000 ;
    END
  END io_out[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070000 3520.400000 2149.630000 3524.800000 ;
    END
  END io_in[17]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110000 3520.400000 2068.670000 3524.800000 ;
    END
  END io_out[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770000 3520.400000 1825.330000 3524.800000 ;
    END
  END io_in[18]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810000 3520.400000 1744.370000 3524.800000 ;
    END
  END io_out[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470000 3520.400000 1501.030000 3524.800000 ;
    END
  END io_in[19]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050000 3520.400000 1419.610000 3524.800000 ;
    END
  END io_out[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 230.940000 2924.800000 232.140000 ;
    END
  END io_in[1]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 297.580000 2924.800000 298.780000 ;
    END
  END io_out[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710000 3520.400000 1176.270000 3524.800000 ;
    END
  END io_in[20]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750000 3520.400000 1095.310000 3524.800000 ;
    END
  END io_out[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410000 3520.400000 851.970000 3524.800000 ;
    END
  END io_in[21]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450000 3520.400000 771.010000 3524.800000 ;
    END
  END io_out[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110000 3520.400000 527.670000 3524.800000 ;
    END
  END io_in[22]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690000 3520.400000 446.250000 3524.800000 ;
    END
  END io_out[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350000 3520.400000 202.910000 3524.800000 ;
    END
  END io_in[23]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390000 3520.400000 121.950000 3524.800000 ;
    END
  END io_out[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3420.820000 -0.400000 3422.020000 ;
    END
  END io_in[24]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3355.540000 -0.400000 3356.740000 ;
    END
  END io_out[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3159.700000 -0.400000 3160.900000 ;
    END
  END io_in[25]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3095.100000 -0.400000 3096.300000 ;
    END
  END io_out[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2899.260000 -0.400000 2900.460000 ;
    END
  END io_in[26]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2833.980000 -0.400000 2835.180000 ;
    END
  END io_out[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2638.820000 -0.400000 2640.020000 ;
    END
  END io_in[27]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2573.540000 -0.400000 2574.740000 ;
    END
  END io_out[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2377.700000 -0.400000 2378.900000 ;
    END
  END io_in[28]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2312.420000 -0.400000 2313.620000 ;
    END
  END io_out[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2117.260000 -0.400000 2118.460000 ;
    END
  END io_in[29]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2051.980000 -0.400000 2053.180000 ;
    END
  END io_out[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 430.180000 2924.800000 431.380000 ;
    END
  END io_in[2]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 496.820000 2924.800000 498.020000 ;
    END
  END io_out[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1856.140000 -0.400000 1857.340000 ;
    END
  END io_in[30]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1791.540000 -0.400000 1792.740000 ;
    END
  END io_out[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1595.700000 -0.400000 1596.900000 ;
    END
  END io_in[31]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1530.420000 -0.400000 1531.620000 ;
    END
  END io_out[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1335.260000 -0.400000 1336.460000 ;
    END
  END io_in[32]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1269.980000 -0.400000 1271.180000 ;
    END
  END io_out[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1074.140000 -0.400000 1075.340000 ;
    END
  END io_in[33]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1008.860000 -0.400000 1010.060000 ;
    END
  END io_out[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 813.700000 -0.400000 814.900000 ;
    END
  END io_in[34]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 748.420000 -0.400000 749.620000 ;
    END
  END io_out[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 552.580000 -0.400000 553.780000 ;
    END
  END io_in[35]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 487.300000 -0.400000 488.500000 ;
    END
  END io_out[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 357.420000 -0.400000 358.620000 ;
    END
  END io_in[36]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 292.140000 -0.400000 293.340000 ;
    END
  END io_out[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 161.580000 -0.400000 162.780000 ;
    END
  END io_in[37]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 96.300000 -0.400000 97.500000 ;
    END
  END io_out[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 629.420000 2924.800000 630.620000 ;
    END
  END io_in[3]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 696.060000 2924.800000 697.260000 ;
    END
  END io_out[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 828.660000 2924.800000 829.860000 ;
    END
  END io_in[4]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 895.300000 2924.800000 896.500000 ;
    END
  END io_out[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1027.900000 2924.800000 1029.100000 ;
    END
  END io_in[5]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1094.540000 2924.800000 1095.740000 ;
    END
  END io_out[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1227.140000 2924.800000 1228.340000 ;
    END
  END io_in[6]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1293.780000 2924.800000 1294.980000 ;
    END
  END io_out[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1493.020000 2924.800000 1494.220000 ;
    END
  END io_in[7]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1559.660000 2924.800000 1560.860000 ;
    END
  END io_out[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1758.900000 2924.800000 1760.100000 ;
    END
  END io_in[8]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1824.860000 2924.800000 1826.060000 ;
    END
  END io_out[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2024.100000 2924.800000 2025.300000 ;
    END
  END io_in[9]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2090.740000 2924.800000 2091.940000 ;
    END
  END io_out[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 164.980000 2924.800000 166.180000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2422.580000 2924.800000 2423.780000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2688.460000 2924.800000 2689.660000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2954.340000 2924.800000 2955.540000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3219.540000 2924.800000 3220.740000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3485.420000 2924.800000 3486.620000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750000 3520.400000 2636.310000 3524.800000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450000 3520.400000 2312.010000 3524.800000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150000 3520.400000 1987.710000 3524.800000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390000 3520.400000 1662.950000 3524.800000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090000 3520.400000 1338.650000 3524.800000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 364.220000 2924.800000 365.420000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790000 3520.400000 1014.350000 3524.800000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030000 3520.400000 689.590000 3524.800000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730000 3520.400000 365.290000 3524.800000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430000 3520.400000 40.990000 3524.800000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3290.260000 -0.400000 3291.460000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3029.820000 -0.400000 3031.020000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2768.700000 -0.400000 2769.900000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2508.260000 -0.400000 2509.460000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2247.140000 -0.400000 2248.340000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1986.700000 -0.400000 1987.900000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 563.460000 2924.800000 564.660000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1726.260000 -0.400000 1727.460000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1465.140000 -0.400000 1466.340000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1204.700000 -0.400000 1205.900000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 943.580000 -0.400000 944.780000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 683.140000 -0.400000 684.340000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 422.700000 -0.400000 423.900000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 226.860000 -0.400000 228.060000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800000 31.700000 -0.400000 32.900000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 762.700000 2924.800000 763.900000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 961.940000 2924.800000 963.140000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1161.180000 2924.800000 1162.380000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1360.420000 2924.800000 1361.620000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1625.620000 2924.800000 1626.820000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1891.500000 2924.800000 1892.700000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2157.380000 2924.800000 2158.580000 ;
    END
  END io_oeb[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230000 -4.800000 629.790000 -0.400000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530000 -4.800000 2403.090000 -0.400000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010000 -4.800000 2420.570000 -0.400000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950000 -4.800000 2438.510000 -0.400000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430000 -4.800000 2455.990000 -0.400000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370000 -4.800000 2473.930000 -0.400000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850000 -4.800000 2491.410000 -0.400000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790000 -4.800000 2509.350000 -0.400000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730000 -4.800000 2527.290000 -0.400000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210000 -4.800000 2544.770000 -0.400000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150000 -4.800000 2562.710000 -0.400000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330000 -4.800000 806.890000 -0.400000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630000 -4.800000 2580.190000 -0.400000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570000 -4.800000 2598.130000 -0.400000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050000 -4.800000 2615.610000 -0.400000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990000 -4.800000 2633.550000 -0.400000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470000 -4.800000 2651.030000 -0.400000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410000 -4.800000 2668.970000 -0.400000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890000 -4.800000 2686.450000 -0.400000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830000 -4.800000 2704.390000 -0.400000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770000 -4.800000 2722.330000 -0.400000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250000 -4.800000 2739.810000 -0.400000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270000 -4.800000 824.830000 -0.400000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190000 -4.800000 2757.750000 -0.400000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670000 -4.800000 2775.230000 -0.400000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610000 -4.800000 2793.170000 -0.400000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090000 -4.800000 2810.650000 -0.400000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030000 -4.800000 2828.590000 -0.400000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510000 -4.800000 2846.070000 -0.400000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450000 -4.800000 2864.010000 -0.400000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390000 -4.800000 2881.950000 -0.400000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750000 -4.800000 842.310000 -0.400000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690000 -4.800000 860.250000 -0.400000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170000 -4.800000 877.730000 -0.400000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110000 -4.800000 895.670000 -0.400000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590000 -4.800000 913.150000 -0.400000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530000 -4.800000 931.090000 -0.400000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470000 -4.800000 949.030000 -0.400000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950000 -4.800000 966.510000 -0.400000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710000 -4.800000 647.270000 -0.400000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890000 -4.800000 984.450000 -0.400000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370000 -4.800000 1001.930000 -0.400000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310000 -4.800000 1019.870000 -0.400000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790000 -4.800000 1037.350000 -0.400000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730000 -4.800000 1055.290000 -0.400000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210000 -4.800000 1072.770000 -0.400000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150000 -4.800000 1090.710000 -0.400000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630000 -4.800000 1108.190000 -0.400000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570000 -4.800000 1126.130000 -0.400000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510000 -4.800000 1144.070000 -0.400000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650000 -4.800000 665.210000 -0.400000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990000 -4.800000 1161.550000 -0.400000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930000 -4.800000 1179.490000 -0.400000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410000 -4.800000 1196.970000 -0.400000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350000 -4.800000 1214.910000 -0.400000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830000 -4.800000 1232.390000 -0.400000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770000 -4.800000 1250.330000 -0.400000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250000 -4.800000 1267.810000 -0.400000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190000 -4.800000 1285.750000 -0.400000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130000 -4.800000 1303.690000 -0.400000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610000 -4.800000 1321.170000 -0.400000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130000 -4.800000 682.690000 -0.400000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550000 -4.800000 1339.110000 -0.400000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030000 -4.800000 1356.590000 -0.400000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970000 -4.800000 1374.530000 -0.400000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450000 -4.800000 1392.010000 -0.400000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390000 -4.800000 1409.950000 -0.400000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870000 -4.800000 1427.430000 -0.400000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810000 -4.800000 1445.370000 -0.400000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750000 -4.800000 1463.310000 -0.400000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230000 -4.800000 1480.790000 -0.400000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170000 -4.800000 1498.730000 -0.400000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070000 -4.800000 700.630000 -0.400000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650000 -4.800000 1516.210000 -0.400000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590000 -4.800000 1534.150000 -0.400000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070000 -4.800000 1551.630000 -0.400000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010000 -4.800000 1569.570000 -0.400000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490000 -4.800000 1587.050000 -0.400000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430000 -4.800000 1604.990000 -0.400000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910000 -4.800000 1622.470000 -0.400000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850000 -4.800000 1640.410000 -0.400000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790000 -4.800000 1658.350000 -0.400000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270000 -4.800000 1675.830000 -0.400000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550000 -4.800000 718.110000 -0.400000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210000 -4.800000 1693.770000 -0.400000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690000 -4.800000 1711.250000 -0.400000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630000 -4.800000 1729.190000 -0.400000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110000 -4.800000 1746.670000 -0.400000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050000 -4.800000 1764.610000 -0.400000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530000 -4.800000 1782.090000 -0.400000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470000 -4.800000 1800.030000 -0.400000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410000 -4.800000 1817.970000 -0.400000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890000 -4.800000 1835.450000 -0.400000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830000 -4.800000 1853.390000 -0.400000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490000 -4.800000 736.050000 -0.400000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310000 -4.800000 1870.870000 -0.400000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250000 -4.800000 1888.810000 -0.400000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730000 -4.800000 1906.290000 -0.400000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670000 -4.800000 1924.230000 -0.400000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150000 -4.800000 1941.710000 -0.400000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090000 -4.800000 1959.650000 -0.400000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570000 -4.800000 1977.130000 -0.400000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510000 -4.800000 1995.070000 -0.400000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450000 -4.800000 2013.010000 -0.400000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930000 -4.800000 2030.490000 -0.400000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970000 -4.800000 753.530000 -0.400000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870000 -4.800000 2048.430000 -0.400000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350000 -4.800000 2065.910000 -0.400000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290000 -4.800000 2083.850000 -0.400000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770000 -4.800000 2101.330000 -0.400000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710000 -4.800000 2119.270000 -0.400000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190000 -4.800000 2136.750000 -0.400000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130000 -4.800000 2154.690000 -0.400000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070000 -4.800000 2172.630000 -0.400000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550000 -4.800000 2190.110000 -0.400000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490000 -4.800000 2208.050000 -0.400000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910000 -4.800000 771.470000 -0.400000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970000 -4.800000 2225.530000 -0.400000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910000 -4.800000 2243.470000 -0.400000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390000 -4.800000 2260.950000 -0.400000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330000 -4.800000 2278.890000 -0.400000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810000 -4.800000 2296.370000 -0.400000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750000 -4.800000 2314.310000 -0.400000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230000 -4.800000 2331.790000 -0.400000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170000 -4.800000 2349.730000 -0.400000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110000 -4.800000 2367.670000 -0.400000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590000 -4.800000 2385.150000 -0.400000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850000 -4.800000 789.410000 -0.400000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750000 -4.800000 635.310000 -0.400000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510000 -4.800000 2409.070000 -0.400000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990000 -4.800000 2426.550000 -0.400000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930000 -4.800000 2444.490000 -0.400000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410000 -4.800000 2461.970000 -0.400000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350000 -4.800000 2479.910000 -0.400000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830000 -4.800000 2497.390000 -0.400000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770000 -4.800000 2515.330000 -0.400000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250000 -4.800000 2532.810000 -0.400000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190000 -4.800000 2550.750000 -0.400000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670000 -4.800000 2568.230000 -0.400000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310000 -4.800000 812.870000 -0.400000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610000 -4.800000 2586.170000 -0.400000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550000 -4.800000 2604.110000 -0.400000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030000 -4.800000 2621.590000 -0.400000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970000 -4.800000 2639.530000 -0.400000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450000 -4.800000 2657.010000 -0.400000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390000 -4.800000 2674.950000 -0.400000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870000 -4.800000 2692.430000 -0.400000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810000 -4.800000 2710.370000 -0.400000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290000 -4.800000 2727.850000 -0.400000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230000 -4.800000 2745.790000 -0.400000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250000 -4.800000 830.810000 -0.400000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170000 -4.800000 2763.730000 -0.400000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650000 -4.800000 2781.210000 -0.400000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590000 -4.800000 2799.150000 -0.400000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070000 -4.800000 2816.630000 -0.400000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010000 -4.800000 2834.570000 -0.400000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490000 -4.800000 2852.050000 -0.400000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430000 -4.800000 2869.990000 -0.400000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910000 -4.800000 2887.470000 -0.400000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730000 -4.800000 848.290000 -0.400000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670000 -4.800000 866.230000 -0.400000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150000 -4.800000 883.710000 -0.400000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090000 -4.800000 901.650000 -0.400000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570000 -4.800000 919.130000 -0.400000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510000 -4.800000 937.070000 -0.400000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990000 -4.800000 954.550000 -0.400000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930000 -4.800000 972.490000 -0.400000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690000 -4.800000 653.250000 -0.400000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410000 -4.800000 989.970000 -0.400000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350000 -4.800000 1007.910000 -0.400000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290000 -4.800000 1025.850000 -0.400000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770000 -4.800000 1043.330000 -0.400000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710000 -4.800000 1061.270000 -0.400000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190000 -4.800000 1078.750000 -0.400000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130000 -4.800000 1096.690000 -0.400000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610000 -4.800000 1114.170000 -0.400000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550000 -4.800000 1132.110000 -0.400000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030000 -4.800000 1149.590000 -0.400000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630000 -4.800000 671.190000 -0.400000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970000 -4.800000 1167.530000 -0.400000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910000 -4.800000 1185.470000 -0.400000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390000 -4.800000 1202.950000 -0.400000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330000 -4.800000 1220.890000 -0.400000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810000 -4.800000 1238.370000 -0.400000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750000 -4.800000 1256.310000 -0.400000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230000 -4.800000 1273.790000 -0.400000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170000 -4.800000 1291.730000 -0.400000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650000 -4.800000 1309.210000 -0.400000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590000 -4.800000 1327.150000 -0.400000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110000 -4.800000 688.670000 -0.400000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070000 -4.800000 1344.630000 -0.400000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010000 -4.800000 1362.570000 -0.400000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950000 -4.800000 1380.510000 -0.400000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430000 -4.800000 1397.990000 -0.400000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370000 -4.800000 1415.930000 -0.400000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850000 -4.800000 1433.410000 -0.400000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790000 -4.800000 1451.350000 -0.400000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270000 -4.800000 1468.830000 -0.400000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210000 -4.800000 1486.770000 -0.400000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690000 -4.800000 1504.250000 -0.400000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050000 -4.800000 706.610000 -0.400000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630000 -4.800000 1522.190000 -0.400000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570000 -4.800000 1540.130000 -0.400000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050000 -4.800000 1557.610000 -0.400000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990000 -4.800000 1575.550000 -0.400000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470000 -4.800000 1593.030000 -0.400000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410000 -4.800000 1610.970000 -0.400000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890000 -4.800000 1628.450000 -0.400000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830000 -4.800000 1646.390000 -0.400000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310000 -4.800000 1663.870000 -0.400000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250000 -4.800000 1681.810000 -0.400000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530000 -4.800000 724.090000 -0.400000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190000 -4.800000 1699.750000 -0.400000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670000 -4.800000 1717.230000 -0.400000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610000 -4.800000 1735.170000 -0.400000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090000 -4.800000 1752.650000 -0.400000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030000 -4.800000 1770.590000 -0.400000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510000 -4.800000 1788.070000 -0.400000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450000 -4.800000 1806.010000 -0.400000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930000 -4.800000 1823.490000 -0.400000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870000 -4.800000 1841.430000 -0.400000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350000 -4.800000 1858.910000 -0.400000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470000 -4.800000 742.030000 -0.400000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290000 -4.800000 1876.850000 -0.400000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230000 -4.800000 1894.790000 -0.400000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710000 -4.800000 1912.270000 -0.400000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650000 -4.800000 1930.210000 -0.400000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130000 -4.800000 1947.690000 -0.400000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070000 -4.800000 1965.630000 -0.400000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550000 -4.800000 1983.110000 -0.400000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490000 -4.800000 2001.050000 -0.400000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970000 -4.800000 2018.530000 -0.400000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910000 -4.800000 2036.470000 -0.400000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950000 -4.800000 759.510000 -0.400000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850000 -4.800000 2054.410000 -0.400000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330000 -4.800000 2071.890000 -0.400000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270000 -4.800000 2089.830000 -0.400000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750000 -4.800000 2107.310000 -0.400000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690000 -4.800000 2125.250000 -0.400000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170000 -4.800000 2142.730000 -0.400000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110000 -4.800000 2160.670000 -0.400000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590000 -4.800000 2178.150000 -0.400000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530000 -4.800000 2196.090000 -0.400000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010000 -4.800000 2213.570000 -0.400000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890000 -4.800000 777.450000 -0.400000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950000 -4.800000 2231.510000 -0.400000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890000 -4.800000 2249.450000 -0.400000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370000 -4.800000 2266.930000 -0.400000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310000 -4.800000 2284.870000 -0.400000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790000 -4.800000 2302.350000 -0.400000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730000 -4.800000 2320.290000 -0.400000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210000 -4.800000 2337.770000 -0.400000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150000 -4.800000 2355.710000 -0.400000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630000 -4.800000 2373.190000 -0.400000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570000 -4.800000 2391.130000 -0.400000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370000 -4.800000 794.930000 -0.400000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730000 -4.800000 641.290000 -0.400000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030000 -4.800000 2414.590000 -0.400000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970000 -4.800000 2432.530000 -0.400000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450000 -4.800000 2450.010000 -0.400000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390000 -4.800000 2467.950000 -0.400000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330000 -4.800000 2485.890000 -0.400000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810000 -4.800000 2503.370000 -0.400000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750000 -4.800000 2521.310000 -0.400000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230000 -4.800000 2538.790000 -0.400000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170000 -4.800000 2556.730000 -0.400000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650000 -4.800000 2574.210000 -0.400000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290000 -4.800000 818.850000 -0.400000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590000 -4.800000 2592.150000 -0.400000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070000 -4.800000 2609.630000 -0.400000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010000 -4.800000 2627.570000 -0.400000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950000 -4.800000 2645.510000 -0.400000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430000 -4.800000 2662.990000 -0.400000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370000 -4.800000 2680.930000 -0.400000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850000 -4.800000 2698.410000 -0.400000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790000 -4.800000 2716.350000 -0.400000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270000 -4.800000 2733.830000 -0.400000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210000 -4.800000 2751.770000 -0.400000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770000 -4.800000 836.330000 -0.400000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690000 -4.800000 2769.250000 -0.400000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630000 -4.800000 2787.190000 -0.400000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110000 -4.800000 2804.670000 -0.400000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050000 -4.800000 2822.610000 -0.400000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990000 -4.800000 2840.550000 -0.400000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470000 -4.800000 2858.030000 -0.400000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410000 -4.800000 2875.970000 -0.400000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890000 -4.800000 2893.450000 -0.400000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710000 -4.800000 854.270000 -0.400000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190000 -4.800000 871.750000 -0.400000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130000 -4.800000 889.690000 -0.400000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070000 -4.800000 907.630000 -0.400000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550000 -4.800000 925.110000 -0.400000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490000 -4.800000 943.050000 -0.400000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970000 -4.800000 960.530000 -0.400000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910000 -4.800000 978.470000 -0.400000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670000 -4.800000 659.230000 -0.400000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390000 -4.800000 995.950000 -0.400000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330000 -4.800000 1013.890000 -0.400000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810000 -4.800000 1031.370000 -0.400000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750000 -4.800000 1049.310000 -0.400000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690000 -4.800000 1067.250000 -0.400000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170000 -4.800000 1084.730000 -0.400000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110000 -4.800000 1102.670000 -0.400000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590000 -4.800000 1120.150000 -0.400000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530000 -4.800000 1138.090000 -0.400000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010000 -4.800000 1155.570000 -0.400000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150000 -4.800000 676.710000 -0.400000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950000 -4.800000 1173.510000 -0.400000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430000 -4.800000 1190.990000 -0.400000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370000 -4.800000 1208.930000 -0.400000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850000 -4.800000 1226.410000 -0.400000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790000 -4.800000 1244.350000 -0.400000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730000 -4.800000 1262.290000 -0.400000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210000 -4.800000 1279.770000 -0.400000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150000 -4.800000 1297.710000 -0.400000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630000 -4.800000 1315.190000 -0.400000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570000 -4.800000 1333.130000 -0.400000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090000 -4.800000 694.650000 -0.400000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050000 -4.800000 1350.610000 -0.400000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990000 -4.800000 1368.550000 -0.400000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470000 -4.800000 1386.030000 -0.400000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410000 -4.800000 1403.970000 -0.400000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350000 -4.800000 1421.910000 -0.400000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830000 -4.800000 1439.390000 -0.400000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770000 -4.800000 1457.330000 -0.400000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250000 -4.800000 1474.810000 -0.400000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190000 -4.800000 1492.750000 -0.400000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670000 -4.800000 1510.230000 -0.400000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030000 -4.800000 712.590000 -0.400000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610000 -4.800000 1528.170000 -0.400000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090000 -4.800000 1545.650000 -0.400000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030000 -4.800000 1563.590000 -0.400000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970000 -4.800000 1581.530000 -0.400000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450000 -4.800000 1599.010000 -0.400000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390000 -4.800000 1616.950000 -0.400000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870000 -4.800000 1634.430000 -0.400000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810000 -4.800000 1652.370000 -0.400000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290000 -4.800000 1669.850000 -0.400000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230000 -4.800000 1687.790000 -0.400000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510000 -4.800000 730.070000 -0.400000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710000 -4.800000 1705.270000 -0.400000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650000 -4.800000 1723.210000 -0.400000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130000 -4.800000 1740.690000 -0.400000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070000 -4.800000 1758.630000 -0.400000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010000 -4.800000 1776.570000 -0.400000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490000 -4.800000 1794.050000 -0.400000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430000 -4.800000 1811.990000 -0.400000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910000 -4.800000 1829.470000 -0.400000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850000 -4.800000 1847.410000 -0.400000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330000 -4.800000 1864.890000 -0.400000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450000 -4.800000 748.010000 -0.400000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270000 -4.800000 1882.830000 -0.400000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750000 -4.800000 1900.310000 -0.400000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690000 -4.800000 1918.250000 -0.400000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630000 -4.800000 1936.190000 -0.400000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110000 -4.800000 1953.670000 -0.400000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050000 -4.800000 1971.610000 -0.400000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530000 -4.800000 1989.090000 -0.400000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470000 -4.800000 2007.030000 -0.400000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950000 -4.800000 2024.510000 -0.400000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890000 -4.800000 2042.450000 -0.400000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930000 -4.800000 765.490000 -0.400000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370000 -4.800000 2059.930000 -0.400000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310000 -4.800000 2077.870000 -0.400000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790000 -4.800000 2095.350000 -0.400000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730000 -4.800000 2113.290000 -0.400000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670000 -4.800000 2131.230000 -0.400000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150000 -4.800000 2148.710000 -0.400000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090000 -4.800000 2166.650000 -0.400000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570000 -4.800000 2184.130000 -0.400000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510000 -4.800000 2202.070000 -0.400000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990000 -4.800000 2219.550000 -0.400000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870000 -4.800000 783.430000 -0.400000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930000 -4.800000 2237.490000 -0.400000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410000 -4.800000 2254.970000 -0.400000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350000 -4.800000 2272.910000 -0.400000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290000 -4.800000 2290.850000 -0.400000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770000 -4.800000 2308.330000 -0.400000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710000 -4.800000 2326.270000 -0.400000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190000 -4.800000 2343.750000 -0.400000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130000 -4.800000 2361.690000 -0.400000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610000 -4.800000 2379.170000 -0.400000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550000 -4.800000 2397.110000 -0.400000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350000 -4.800000 800.910000 -0.400000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870000 -4.800000 2899.430000 -0.400000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850000 -4.800000 2905.410000 -0.400000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830000 -4.800000 2911.390000 -0.400000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810000 -4.800000 2917.370000 -0.400000 ;
    END
  END user_irq[2]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710000 -4.800000 3.270000 -0.400000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230000 -4.800000 8.790000 -0.400000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210000 -4.800000 14.770000 -0.400000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130000 -4.800000 38.690000 -0.400000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150000 -4.800000 239.710000 -0.400000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630000 -4.800000 257.190000 -0.400000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570000 -4.800000 275.130000 -0.400000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050000 -4.800000 292.610000 -0.400000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990000 -4.800000 310.550000 -0.400000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470000 -4.800000 328.030000 -0.400000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410000 -4.800000 345.970000 -0.400000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890000 -4.800000 363.450000 -0.400000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830000 -4.800000 381.390000 -0.400000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310000 -4.800000 398.870000 -0.400000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590000 -4.800000 62.150000 -0.400000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250000 -4.800000 416.810000 -0.400000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190000 -4.800000 434.750000 -0.400000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670000 -4.800000 452.230000 -0.400000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610000 -4.800000 470.170000 -0.400000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090000 -4.800000 487.650000 -0.400000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030000 -4.800000 505.590000 -0.400000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510000 -4.800000 523.070000 -0.400000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450000 -4.800000 541.010000 -0.400000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930000 -4.800000 558.490000 -0.400000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870000 -4.800000 576.430000 -0.400000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050000 -4.800000 85.610000 -0.400000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810000 -4.800000 594.370000 -0.400000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290000 -4.800000 611.850000 -0.400000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970000 -4.800000 109.530000 -0.400000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430000 -4.800000 132.990000 -0.400000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370000 -4.800000 150.930000 -0.400000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850000 -4.800000 168.410000 -0.400000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790000 -4.800000 186.350000 -0.400000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270000 -4.800000 203.830000 -0.400000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210000 -4.800000 221.770000 -0.400000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190000 -4.800000 20.750000 -0.400000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650000 -4.800000 44.210000 -0.400000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670000 -4.800000 245.230000 -0.400000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610000 -4.800000 263.170000 -0.400000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090000 -4.800000 280.650000 -0.400000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030000 -4.800000 298.590000 -0.400000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970000 -4.800000 316.530000 -0.400000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450000 -4.800000 334.010000 -0.400000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390000 -4.800000 351.950000 -0.400000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870000 -4.800000 369.430000 -0.400000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810000 -4.800000 387.370000 -0.400000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290000 -4.800000 404.850000 -0.400000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570000 -4.800000 68.130000 -0.400000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230000 -4.800000 422.790000 -0.400000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710000 -4.800000 440.270000 -0.400000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650000 -4.800000 458.210000 -0.400000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590000 -4.800000 476.150000 -0.400000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070000 -4.800000 493.630000 -0.400000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010000 -4.800000 511.570000 -0.400000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490000 -4.800000 529.050000 -0.400000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430000 -4.800000 546.990000 -0.400000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910000 -4.800000 564.470000 -0.400000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850000 -4.800000 582.410000 -0.400000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030000 -4.800000 91.590000 -0.400000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330000 -4.800000 599.890000 -0.400000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270000 -4.800000 617.830000 -0.400000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950000 -4.800000 115.510000 -0.400000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410000 -4.800000 138.970000 -0.400000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350000 -4.800000 156.910000 -0.400000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830000 -4.800000 174.390000 -0.400000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770000 -4.800000 192.330000 -0.400000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250000 -4.800000 209.810000 -0.400000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190000 -4.800000 227.750000 -0.400000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630000 -4.800000 50.190000 -0.400000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650000 -4.800000 251.210000 -0.400000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590000 -4.800000 269.150000 -0.400000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070000 -4.800000 286.630000 -0.400000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010000 -4.800000 304.570000 -0.400000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490000 -4.800000 322.050000 -0.400000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430000 -4.800000 339.990000 -0.400000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370000 -4.800000 357.930000 -0.400000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850000 -4.800000 375.410000 -0.400000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790000 -4.800000 393.350000 -0.400000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270000 -4.800000 410.830000 -0.400000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550000 -4.800000 74.110000 -0.400000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210000 -4.800000 428.770000 -0.400000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690000 -4.800000 446.250000 -0.400000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630000 -4.800000 464.190000 -0.400000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110000 -4.800000 481.670000 -0.400000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050000 -4.800000 499.610000 -0.400000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530000 -4.800000 517.090000 -0.400000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470000 -4.800000 535.030000 -0.400000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410000 -4.800000 552.970000 -0.400000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890000 -4.800000 570.450000 -0.400000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830000 -4.800000 588.390000 -0.400000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010000 -4.800000 97.570000 -0.400000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310000 -4.800000 605.870000 -0.400000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250000 -4.800000 623.810000 -0.400000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930000 -4.800000 121.490000 -0.400000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390000 -4.800000 144.950000 -0.400000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870000 -4.800000 162.430000 -0.400000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810000 -4.800000 180.370000 -0.400000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750000 -4.800000 198.310000 -0.400000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230000 -4.800000 215.790000 -0.400000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170000 -4.800000 233.730000 -0.400000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610000 -4.800000 56.170000 -0.400000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530000 -4.800000 80.090000 -0.400000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990000 -4.800000 103.550000 -0.400000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450000 -4.800000 127.010000 -0.400000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170000 -4.800000 26.730000 -0.400000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150000 -4.800000 32.710000 -0.400000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2889.020000 -9.320000 2892.020000 -0.400000 ;
        RECT 2889.020000 3520.400000 2892.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2709.020000 -9.320000 2712.020000 -0.400000 ;
        RECT 2709.020000 3520.400000 2712.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2529.020000 -9.320000 2532.020000 -0.400000 ;
        RECT 2529.020000 3520.400000 2532.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2349.020000 -9.320000 2352.020000 -0.400000 ;
        RECT 2349.020000 3520.400000 2352.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2169.020000 -9.320000 2172.020000 -0.400000 ;
        RECT 2169.020000 3520.400000 2172.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1989.020000 -9.320000 1992.020000 -0.400000 ;
        RECT 1989.020000 3520.400000 1992.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1809.020000 -9.320000 1812.020000 -0.400000 ;
        RECT 1809.020000 3520.400000 1812.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1629.020000 -9.320000 1632.020000 -0.400000 ;
        RECT 1629.020000 3520.400000 1632.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1449.020000 -9.320000 1452.020000 -0.400000 ;
        RECT 1449.020000 3520.400000 1452.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1269.020000 -9.320000 1272.020000 -0.400000 ;
        RECT 1269.020000 3520.400000 1272.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1089.020000 -9.320000 1092.020000 -0.400000 ;
        RECT 1089.020000 3520.400000 1092.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 909.020000 -9.320000 912.020000 -0.400000 ;
        RECT 909.020000 3520.400000 912.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 729.020000 -9.320000 732.020000 -0.400000 ;
        RECT 729.020000 3520.400000 732.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 549.020000 -9.320000 552.020000 -0.400000 ;
        RECT 549.020000 3520.400000 552.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 369.020000 -9.320000 372.020000 -0.400000 ;
        RECT 369.020000 3520.400000 372.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 189.020000 -9.320000 192.020000 -0.400000 ;
        RECT 189.020000 3520.400000 192.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.020000 -9.320000 12.020000 -0.400000 ;
        RECT 9.020000 3520.400000 12.020000 3529.000000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2926.600000 -4.620000 2929.600000 3524.300000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980000 -4.620000 -6.980000 3524.300000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -9.980000 3521.300000 2929.600000 3524.300000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 3434.140000 -0.400000 3437.140000 ;
        RECT 2920.400000 3434.140000 2934.300000 3437.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 3254.140000 -0.400000 3257.140000 ;
        RECT 2920.400000 3254.140000 2934.300000 3257.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 3074.140000 -0.400000 3077.140000 ;
        RECT 2920.400000 3074.140000 2934.300000 3077.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 2894.140000 -0.400000 2897.140000 ;
        RECT 2920.400000 2894.140000 2934.300000 2897.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 2714.140000 -0.400000 2717.140000 ;
        RECT 2920.400000 2714.140000 2934.300000 2717.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 2534.140000 -0.400000 2537.140000 ;
        RECT 2920.400000 2534.140000 2934.300000 2537.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 2354.140000 -0.400000 2357.140000 ;
        RECT 2920.400000 2354.140000 2934.300000 2357.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 2174.140000 -0.400000 2177.140000 ;
        RECT 2920.400000 2174.140000 2934.300000 2177.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1994.140000 -0.400000 1997.140000 ;
        RECT 2920.400000 1994.140000 2934.300000 1997.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1814.140000 -0.400000 1817.140000 ;
        RECT 2920.400000 1814.140000 2934.300000 1817.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1634.140000 -0.400000 1637.140000 ;
        RECT 2920.400000 1634.140000 2934.300000 1637.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1454.140000 -0.400000 1457.140000 ;
        RECT 2920.400000 1454.140000 2934.300000 1457.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1274.140000 -0.400000 1277.140000 ;
        RECT 2920.400000 1274.140000 2934.300000 1277.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1094.140000 -0.400000 1097.140000 ;
        RECT 2920.400000 1094.140000 2934.300000 1097.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 914.140000 -0.400000 917.140000 ;
        RECT 2920.400000 914.140000 2934.300000 917.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 734.140000 -0.400000 737.140000 ;
        RECT 2920.400000 734.140000 2934.300000 737.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 554.140000 -0.400000 557.140000 ;
        RECT 2920.400000 554.140000 2934.300000 557.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 374.140000 -0.400000 377.140000 ;
        RECT 2920.400000 374.140000 2934.300000 377.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 194.140000 -0.400000 197.140000 ;
        RECT 2920.400000 194.140000 2934.300000 197.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680000 14.140000 -0.400000 17.140000 ;
        RECT 2920.400000 14.140000 2934.300000 17.140000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -9.980000 -4.620000 2929.600000 -1.620000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2931.300000 -9.320000 2934.300000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2799.020000 -9.320000 2802.020000 -0.400000 ;
        RECT 2799.020000 3520.400000 2802.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2619.020000 -9.320000 2622.020000 -0.400000 ;
        RECT 2619.020000 3520.400000 2622.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2439.020000 -9.320000 2442.020000 -0.400000 ;
        RECT 2439.020000 3520.400000 2442.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2259.020000 -9.320000 2262.020000 -0.400000 ;
        RECT 2259.020000 3520.400000 2262.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2079.020000 -9.320000 2082.020000 -0.400000 ;
        RECT 2079.020000 3520.400000 2082.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1899.020000 -9.320000 1902.020000 -0.400000 ;
        RECT 1899.020000 3520.400000 1902.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1719.020000 -9.320000 1722.020000 -0.400000 ;
        RECT 1719.020000 3520.400000 1722.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1539.020000 -9.320000 1542.020000 -0.400000 ;
        RECT 1539.020000 3520.400000 1542.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1359.020000 -9.320000 1362.020000 -0.400000 ;
        RECT 1359.020000 3520.400000 1362.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1179.020000 -9.320000 1182.020000 -0.400000 ;
        RECT 1179.020000 3520.400000 1182.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 999.020000 -9.320000 1002.020000 -0.400000 ;
        RECT 999.020000 3520.400000 1002.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 819.020000 -9.320000 822.020000 -0.400000 ;
        RECT 819.020000 3520.400000 822.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 639.020000 -9.320000 642.020000 -0.400000 ;
        RECT 639.020000 3520.400000 642.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 459.020000 -9.320000 462.020000 -0.400000 ;
        RECT 459.020000 3520.400000 462.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 279.020000 -9.320000 282.020000 -0.400000 ;
        RECT 279.020000 3520.400000 282.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 99.020000 -9.320000 102.020000 -0.400000 ;
        RECT 99.020000 3520.400000 102.020000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.680000 -9.320000 -11.680000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 3526.000000 2934.300000 3529.000000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 3344.140000 -0.400000 3347.140000 ;
        RECT 2920.400000 3344.140000 2934.300000 3347.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 3164.140000 -0.400000 3167.140000 ;
        RECT 2920.400000 3164.140000 2934.300000 3167.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 2984.140000 -0.400000 2987.140000 ;
        RECT 2920.400000 2984.140000 2934.300000 2987.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 2804.140000 -0.400000 2807.140000 ;
        RECT 2920.400000 2804.140000 2934.300000 2807.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 2624.140000 -0.400000 2627.140000 ;
        RECT 2920.400000 2624.140000 2934.300000 2627.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 2444.140000 -0.400000 2447.140000 ;
        RECT 2920.400000 2444.140000 2934.300000 2447.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 2264.140000 -0.400000 2267.140000 ;
        RECT 2920.400000 2264.140000 2934.300000 2267.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 2084.140000 -0.400000 2087.140000 ;
        RECT 2920.400000 2084.140000 2934.300000 2087.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1904.140000 -0.400000 1907.140000 ;
        RECT 2920.400000 1904.140000 2934.300000 1907.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1724.140000 -0.400000 1727.140000 ;
        RECT 2920.400000 1724.140000 2934.300000 1727.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1544.140000 -0.400000 1547.140000 ;
        RECT 2920.400000 1544.140000 2934.300000 1547.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1364.140000 -0.400000 1367.140000 ;
        RECT 2920.400000 1364.140000 2934.300000 1367.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1184.140000 -0.400000 1187.140000 ;
        RECT 2920.400000 1184.140000 2934.300000 1187.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 1004.140000 -0.400000 1007.140000 ;
        RECT 2920.400000 1004.140000 2934.300000 1007.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 824.140000 -0.400000 827.140000 ;
        RECT 2920.400000 824.140000 2934.300000 827.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 644.140000 -0.400000 647.140000 ;
        RECT 2920.400000 644.140000 2934.300000 647.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 464.140000 -0.400000 467.140000 ;
        RECT 2920.400000 464.140000 2934.300000 467.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 284.140000 -0.400000 287.140000 ;
        RECT 2920.400000 284.140000 2934.300000 287.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 104.140000 -0.400000 107.140000 ;
        RECT 2920.400000 104.140000 2934.300000 107.140000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680000 -9.320000 2934.300000 -6.320000 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2907.020000 -18.720000 2910.020000 -0.400000 ;
        RECT 2907.020000 3520.400000 2910.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2727.020000 -18.720000 2730.020000 -0.400000 ;
        RECT 2727.020000 3520.400000 2730.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2547.020000 -18.720000 2550.020000 -0.400000 ;
        RECT 2547.020000 3520.400000 2550.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2367.020000 -18.720000 2370.020000 -0.400000 ;
        RECT 2367.020000 3520.400000 2370.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2187.020000 -18.720000 2190.020000 -0.400000 ;
        RECT 2187.020000 3520.400000 2190.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2007.020000 -18.720000 2010.020000 -0.400000 ;
        RECT 2007.020000 3520.400000 2010.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1827.020000 -18.720000 1830.020000 -0.400000 ;
        RECT 1827.020000 3520.400000 1830.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1647.020000 -18.720000 1650.020000 -0.400000 ;
        RECT 1647.020000 3520.400000 1650.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1467.020000 -18.720000 1470.020000 -0.400000 ;
        RECT 1467.020000 3520.400000 1470.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1287.020000 -18.720000 1290.020000 -0.400000 ;
        RECT 1287.020000 3520.400000 1290.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1107.020000 -18.720000 1110.020000 -0.400000 ;
        RECT 1107.020000 3520.400000 1110.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 927.020000 -18.720000 930.020000 -0.400000 ;
        RECT 927.020000 3520.400000 930.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 747.020000 -18.720000 750.020000 -0.400000 ;
        RECT 747.020000 3520.400000 750.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 567.020000 -18.720000 570.020000 -0.400000 ;
        RECT 567.020000 3520.400000 570.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 387.020000 -18.720000 390.020000 -0.400000 ;
        RECT 387.020000 3520.400000 390.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 207.020000 -18.720000 210.020000 -0.400000 ;
        RECT 207.020000 3520.400000 210.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.020000 -18.720000 30.020000 -0.400000 ;
        RECT 27.020000 3520.400000 30.020000 3538.400000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2936.000000 -14.020000 2939.000000 3533.700000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.380000 -14.020000 -16.380000 3533.700000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.380000 3530.700000 2939.000000 3533.700000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 3452.380000 -0.400000 3455.380000 ;
        RECT 2920.400000 3452.380000 2943.700000 3455.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 3272.380000 -0.400000 3275.380000 ;
        RECT 2920.400000 3272.380000 2943.700000 3275.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 3092.380000 -0.400000 3095.380000 ;
        RECT 2920.400000 3092.380000 2943.700000 3095.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 2912.380000 -0.400000 2915.380000 ;
        RECT 2920.400000 2912.380000 2943.700000 2915.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 2732.380000 -0.400000 2735.380000 ;
        RECT 2920.400000 2732.380000 2943.700000 2735.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 2552.380000 -0.400000 2555.380000 ;
        RECT 2920.400000 2552.380000 2943.700000 2555.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 2372.380000 -0.400000 2375.380000 ;
        RECT 2920.400000 2372.380000 2943.700000 2375.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 2192.380000 -0.400000 2195.380000 ;
        RECT 2920.400000 2192.380000 2943.700000 2195.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 2012.380000 -0.400000 2015.380000 ;
        RECT 2920.400000 2012.380000 2943.700000 2015.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 1832.380000 -0.400000 1835.380000 ;
        RECT 2920.400000 1832.380000 2943.700000 1835.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 1652.380000 -0.400000 1655.380000 ;
        RECT 2920.400000 1652.380000 2943.700000 1655.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 1472.380000 -0.400000 1475.380000 ;
        RECT 2920.400000 1472.380000 2943.700000 1475.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 1292.380000 -0.400000 1295.380000 ;
        RECT 2920.400000 1292.380000 2943.700000 1295.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 1112.380000 -0.400000 1115.380000 ;
        RECT 2920.400000 1112.380000 2943.700000 1115.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 932.380000 -0.400000 935.380000 ;
        RECT 2920.400000 932.380000 2943.700000 935.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 752.380000 -0.400000 755.380000 ;
        RECT 2920.400000 752.380000 2943.700000 755.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 572.380000 -0.400000 575.380000 ;
        RECT 2920.400000 572.380000 2943.700000 575.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 392.380000 -0.400000 395.380000 ;
        RECT 2920.400000 392.380000 2943.700000 395.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 212.380000 -0.400000 215.380000 ;
        RECT 2920.400000 212.380000 2943.700000 215.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080000 32.380000 -0.400000 35.380000 ;
        RECT 2920.400000 32.380000 2943.700000 35.380000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.380000 -14.020000 2939.000000 -11.020000 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2940.700000 -18.720000 2943.700000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2817.020000 -18.720000 2820.020000 -0.400000 ;
        RECT 2817.020000 3520.400000 2820.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2637.020000 -18.720000 2640.020000 -0.400000 ;
        RECT 2637.020000 3520.400000 2640.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2457.020000 -18.720000 2460.020000 -0.400000 ;
        RECT 2457.020000 3520.400000 2460.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2277.020000 -18.720000 2280.020000 -0.400000 ;
        RECT 2277.020000 3520.400000 2280.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.020000 -18.720000 2100.020000 -0.400000 ;
        RECT 2097.020000 3520.400000 2100.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1917.020000 -18.720000 1920.020000 -0.400000 ;
        RECT 1917.020000 3520.400000 1920.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1737.020000 -18.720000 1740.020000 -0.400000 ;
        RECT 1737.020000 3520.400000 1740.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1557.020000 -18.720000 1560.020000 -0.400000 ;
        RECT 1557.020000 3520.400000 1560.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1377.020000 -18.720000 1380.020000 -0.400000 ;
        RECT 1377.020000 3520.400000 1380.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1197.020000 -18.720000 1200.020000 -0.400000 ;
        RECT 1197.020000 3520.400000 1200.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1017.020000 -18.720000 1020.020000 -0.400000 ;
        RECT 1017.020000 3520.400000 1020.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 837.020000 -18.720000 840.020000 -0.400000 ;
        RECT 837.020000 3520.400000 840.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 657.020000 -18.720000 660.020000 -0.400000 ;
        RECT 657.020000 3520.400000 660.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 477.020000 -18.720000 480.020000 -0.400000 ;
        RECT 477.020000 3520.400000 480.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 297.020000 -18.720000 300.020000 -0.400000 ;
        RECT 297.020000 3520.400000 300.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 117.020000 -18.720000 120.020000 -0.400000 ;
        RECT 117.020000 3520.400000 120.020000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.080000 -18.720000 -21.080000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 3535.400000 2943.700000 3538.400000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 3362.380000 -0.400000 3365.380000 ;
        RECT 2920.400000 3362.380000 2943.700000 3365.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 3182.380000 -0.400000 3185.380000 ;
        RECT 2920.400000 3182.380000 2943.700000 3185.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 3002.380000 -0.400000 3005.380000 ;
        RECT 2920.400000 3002.380000 2943.700000 3005.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 2822.380000 -0.400000 2825.380000 ;
        RECT 2920.400000 2822.380000 2943.700000 2825.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 2642.380000 -0.400000 2645.380000 ;
        RECT 2920.400000 2642.380000 2943.700000 2645.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 2462.380000 -0.400000 2465.380000 ;
        RECT 2920.400000 2462.380000 2943.700000 2465.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 2282.380000 -0.400000 2285.380000 ;
        RECT 2920.400000 2282.380000 2943.700000 2285.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 2102.380000 -0.400000 2105.380000 ;
        RECT 2920.400000 2102.380000 2943.700000 2105.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 1922.380000 -0.400000 1925.380000 ;
        RECT 2920.400000 1922.380000 2943.700000 1925.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 1742.380000 -0.400000 1745.380000 ;
        RECT 2920.400000 1742.380000 2943.700000 1745.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 1562.380000 -0.400000 1565.380000 ;
        RECT 2920.400000 1562.380000 2943.700000 1565.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 1382.380000 -0.400000 1385.380000 ;
        RECT 2920.400000 1382.380000 2943.700000 1385.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 1202.380000 -0.400000 1205.380000 ;
        RECT 2920.400000 1202.380000 2943.700000 1205.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 1022.380000 -0.400000 1025.380000 ;
        RECT 2920.400000 1022.380000 2943.700000 1025.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 842.380000 -0.400000 845.380000 ;
        RECT 2920.400000 842.380000 2943.700000 845.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 662.380000 -0.400000 665.380000 ;
        RECT 2920.400000 662.380000 2943.700000 665.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 482.380000 -0.400000 485.380000 ;
        RECT 2920.400000 482.380000 2943.700000 485.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 302.380000 -0.400000 305.380000 ;
        RECT 2920.400000 302.380000 2943.700000 305.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 122.380000 -0.400000 125.380000 ;
        RECT 2920.400000 122.380000 2943.700000 125.380000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080000 -18.720000 2943.700000 -15.720000 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2745.020000 -28.120000 2748.020000 -0.400000 ;
        RECT 2745.020000 3520.400000 2748.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2565.020000 -28.120000 2568.020000 -0.400000 ;
        RECT 2565.020000 3520.400000 2568.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2385.020000 -28.120000 2388.020000 -0.400000 ;
        RECT 2385.020000 3520.400000 2388.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2205.020000 -28.120000 2208.020000 -0.400000 ;
        RECT 2205.020000 3520.400000 2208.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2025.020000 -28.120000 2028.020000 -0.400000 ;
        RECT 2025.020000 3520.400000 2028.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1845.020000 -28.120000 1848.020000 -0.400000 ;
        RECT 1845.020000 3520.400000 1848.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1665.020000 -28.120000 1668.020000 -0.400000 ;
        RECT 1665.020000 3520.400000 1668.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1485.020000 -28.120000 1488.020000 -0.400000 ;
        RECT 1485.020000 3520.400000 1488.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1305.020000 -28.120000 1308.020000 -0.400000 ;
        RECT 1305.020000 3520.400000 1308.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1125.020000 -28.120000 1128.020000 -0.400000 ;
        RECT 1125.020000 3520.400000 1128.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 945.020000 -28.120000 948.020000 -0.400000 ;
        RECT 945.020000 3520.400000 948.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 765.020000 -28.120000 768.020000 -0.400000 ;
        RECT 765.020000 3520.400000 768.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 585.020000 -28.120000 588.020000 -0.400000 ;
        RECT 585.020000 3520.400000 588.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 405.020000 -28.120000 408.020000 -0.400000 ;
        RECT 405.020000 3520.400000 408.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 225.020000 -28.120000 228.020000 -0.400000 ;
        RECT 225.020000 3520.400000 228.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 45.020000 -28.120000 48.020000 -0.400000 ;
        RECT 45.020000 3520.400000 48.020000 3547.800000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2945.400000 -23.420000 2948.400000 3543.100000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -28.780000 -23.420000 -25.780000 3543.100000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -28.780000 3540.100000 2948.400000 3543.100000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 3470.380000 -0.400000 3473.380000 ;
        RECT 2920.400000 3470.380000 2953.100000 3473.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 3290.380000 -0.400000 3293.380000 ;
        RECT 2920.400000 3290.380000 2953.100000 3293.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 3110.380000 -0.400000 3113.380000 ;
        RECT 2920.400000 3110.380000 2953.100000 3113.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 2930.380000 -0.400000 2933.380000 ;
        RECT 2920.400000 2930.380000 2953.100000 2933.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 2750.380000 -0.400000 2753.380000 ;
        RECT 2920.400000 2750.380000 2953.100000 2753.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 2570.380000 -0.400000 2573.380000 ;
        RECT 2920.400000 2570.380000 2953.100000 2573.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 2390.380000 -0.400000 2393.380000 ;
        RECT 2920.400000 2390.380000 2953.100000 2393.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 2210.380000 -0.400000 2213.380000 ;
        RECT 2920.400000 2210.380000 2953.100000 2213.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 2030.380000 -0.400000 2033.380000 ;
        RECT 2920.400000 2030.380000 2953.100000 2033.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 1850.380000 -0.400000 1853.380000 ;
        RECT 2920.400000 1850.380000 2953.100000 1853.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 1670.380000 -0.400000 1673.380000 ;
        RECT 2920.400000 1670.380000 2953.100000 1673.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 1490.380000 -0.400000 1493.380000 ;
        RECT 2920.400000 1490.380000 2953.100000 1493.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 1310.380000 -0.400000 1313.380000 ;
        RECT 2920.400000 1310.380000 2953.100000 1313.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 1130.380000 -0.400000 1133.380000 ;
        RECT 2920.400000 1130.380000 2953.100000 1133.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 950.380000 -0.400000 953.380000 ;
        RECT 2920.400000 950.380000 2953.100000 953.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 770.380000 -0.400000 773.380000 ;
        RECT 2920.400000 770.380000 2953.100000 773.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 590.380000 -0.400000 593.380000 ;
        RECT 2920.400000 590.380000 2953.100000 593.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 410.380000 -0.400000 413.380000 ;
        RECT 2920.400000 410.380000 2953.100000 413.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 230.380000 -0.400000 233.380000 ;
        RECT 2920.400000 230.380000 2953.100000 233.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480000 50.380000 -0.400000 53.380000 ;
        RECT 2920.400000 50.380000 2953.100000 53.380000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -28.780000 -23.420000 2948.400000 -20.420000 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2950.100000 -28.120000 2953.100000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2835.020000 -28.120000 2838.020000 -0.400000 ;
        RECT 2835.020000 3520.400000 2838.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2655.020000 -28.120000 2658.020000 -0.400000 ;
        RECT 2655.020000 3520.400000 2658.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2475.020000 -28.120000 2478.020000 -0.400000 ;
        RECT 2475.020000 3520.400000 2478.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2295.020000 -28.120000 2298.020000 -0.400000 ;
        RECT 2295.020000 3520.400000 2298.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2115.020000 -28.120000 2118.020000 -0.400000 ;
        RECT 2115.020000 3520.400000 2118.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1935.020000 -28.120000 1938.020000 -0.400000 ;
        RECT 1935.020000 3520.400000 1938.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1755.020000 -28.120000 1758.020000 -0.400000 ;
        RECT 1755.020000 3520.400000 1758.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1575.020000 -28.120000 1578.020000 -0.400000 ;
        RECT 1575.020000 3520.400000 1578.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1395.020000 -28.120000 1398.020000 -0.400000 ;
        RECT 1395.020000 3520.400000 1398.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1215.020000 -28.120000 1218.020000 -0.400000 ;
        RECT 1215.020000 3520.400000 1218.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1035.020000 -28.120000 1038.020000 -0.400000 ;
        RECT 1035.020000 3520.400000 1038.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 855.020000 -28.120000 858.020000 -0.400000 ;
        RECT 855.020000 3520.400000 858.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 675.020000 -28.120000 678.020000 -0.400000 ;
        RECT 675.020000 3520.400000 678.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 495.020000 -28.120000 498.020000 -0.400000 ;
        RECT 495.020000 3520.400000 498.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 315.020000 -28.120000 318.020000 -0.400000 ;
        RECT 315.020000 3520.400000 318.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 135.020000 -28.120000 138.020000 -0.400000 ;
        RECT 135.020000 3520.400000 138.020000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -33.480000 -28.120000 -30.480000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 3544.800000 2953.100000 3547.800000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 3380.380000 -0.400000 3383.380000 ;
        RECT 2920.400000 3380.380000 2953.100000 3383.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 3200.380000 -0.400000 3203.380000 ;
        RECT 2920.400000 3200.380000 2953.100000 3203.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 3020.380000 -0.400000 3023.380000 ;
        RECT 2920.400000 3020.380000 2953.100000 3023.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 2840.380000 -0.400000 2843.380000 ;
        RECT 2920.400000 2840.380000 2953.100000 2843.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 2660.380000 -0.400000 2663.380000 ;
        RECT 2920.400000 2660.380000 2953.100000 2663.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 2480.380000 -0.400000 2483.380000 ;
        RECT 2920.400000 2480.380000 2953.100000 2483.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 2300.380000 -0.400000 2303.380000 ;
        RECT 2920.400000 2300.380000 2953.100000 2303.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 2120.380000 -0.400000 2123.380000 ;
        RECT 2920.400000 2120.380000 2953.100000 2123.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 1940.380000 -0.400000 1943.380000 ;
        RECT 2920.400000 1940.380000 2953.100000 1943.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 1760.380000 -0.400000 1763.380000 ;
        RECT 2920.400000 1760.380000 2953.100000 1763.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 1580.380000 -0.400000 1583.380000 ;
        RECT 2920.400000 1580.380000 2953.100000 1583.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 1400.380000 -0.400000 1403.380000 ;
        RECT 2920.400000 1400.380000 2953.100000 1403.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 1220.380000 -0.400000 1223.380000 ;
        RECT 2920.400000 1220.380000 2953.100000 1223.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 1040.380000 -0.400000 1043.380000 ;
        RECT 2920.400000 1040.380000 2953.100000 1043.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 860.380000 -0.400000 863.380000 ;
        RECT 2920.400000 860.380000 2953.100000 863.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 680.380000 -0.400000 683.380000 ;
        RECT 2920.400000 680.380000 2953.100000 683.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 500.380000 -0.400000 503.380000 ;
        RECT 2920.400000 500.380000 2953.100000 503.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 320.380000 -0.400000 323.380000 ;
        RECT 2920.400000 320.380000 2953.100000 323.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 140.380000 -0.400000 143.380000 ;
        RECT 2920.400000 140.380000 2953.100000 143.380000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480000 -28.120000 2953.100000 -25.120000 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2763.020000 -37.520000 2766.020000 -0.400000 ;
        RECT 2763.020000 3520.400000 2766.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2583.020000 -37.520000 2586.020000 -0.400000 ;
        RECT 2583.020000 3520.400000 2586.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2403.020000 -37.520000 2406.020000 -0.400000 ;
        RECT 2403.020000 3520.400000 2406.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2223.020000 -37.520000 2226.020000 -0.400000 ;
        RECT 2223.020000 3520.400000 2226.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2043.020000 -37.520000 2046.020000 -0.400000 ;
        RECT 2043.020000 3520.400000 2046.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1863.020000 -37.520000 1866.020000 -0.400000 ;
        RECT 1863.020000 3520.400000 1866.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1683.020000 -37.520000 1686.020000 -0.400000 ;
        RECT 1683.020000 3520.400000 1686.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1503.020000 -37.520000 1506.020000 -0.400000 ;
        RECT 1503.020000 3520.400000 1506.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1323.020000 -37.520000 1326.020000 -0.400000 ;
        RECT 1323.020000 3520.400000 1326.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1143.020000 -37.520000 1146.020000 -0.400000 ;
        RECT 1143.020000 3520.400000 1146.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 963.020000 -37.520000 966.020000 -0.400000 ;
        RECT 963.020000 3520.400000 966.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 783.020000 -37.520000 786.020000 -0.400000 ;
        RECT 783.020000 3520.400000 786.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 603.020000 -37.520000 606.020000 -0.400000 ;
        RECT 603.020000 3520.400000 606.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 423.020000 -37.520000 426.020000 -0.400000 ;
        RECT 423.020000 3520.400000 426.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 243.020000 -37.520000 246.020000 -0.400000 ;
        RECT 243.020000 3520.400000 246.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 63.020000 -37.520000 66.020000 -0.400000 ;
        RECT 63.020000 3520.400000 66.020000 3557.200000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2954.800000 -32.820000 2957.800000 3552.500000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180000 -32.820000 -35.180000 3552.500000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.180000 3549.500000 2957.800000 3552.500000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 3488.380000 -0.400000 3491.380000 ;
        RECT 2920.400000 3488.380000 2962.500000 3491.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 3308.380000 -0.400000 3311.380000 ;
        RECT 2920.400000 3308.380000 2962.500000 3311.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 3128.380000 -0.400000 3131.380000 ;
        RECT 2920.400000 3128.380000 2962.500000 3131.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 2948.380000 -0.400000 2951.380000 ;
        RECT 2920.400000 2948.380000 2962.500000 2951.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 2768.380000 -0.400000 2771.380000 ;
        RECT 2920.400000 2768.380000 2962.500000 2771.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 2588.380000 -0.400000 2591.380000 ;
        RECT 2920.400000 2588.380000 2962.500000 2591.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 2408.380000 -0.400000 2411.380000 ;
        RECT 2920.400000 2408.380000 2962.500000 2411.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 2228.380000 -0.400000 2231.380000 ;
        RECT 2920.400000 2228.380000 2962.500000 2231.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 2048.380000 -0.400000 2051.380000 ;
        RECT 2920.400000 2048.380000 2962.500000 2051.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 1868.380000 -0.400000 1871.380000 ;
        RECT 2920.400000 1868.380000 2962.500000 1871.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 1688.380000 -0.400000 1691.380000 ;
        RECT 2920.400000 1688.380000 2962.500000 1691.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 1508.380000 -0.400000 1511.380000 ;
        RECT 2920.400000 1508.380000 2962.500000 1511.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 1328.380000 -0.400000 1331.380000 ;
        RECT 2920.400000 1328.380000 2962.500000 1331.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 1148.380000 -0.400000 1151.380000 ;
        RECT 2920.400000 1148.380000 2962.500000 1151.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 968.380000 -0.400000 971.380000 ;
        RECT 2920.400000 968.380000 2962.500000 971.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 788.380000 -0.400000 791.380000 ;
        RECT 2920.400000 788.380000 2962.500000 791.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 608.380000 -0.400000 611.380000 ;
        RECT 2920.400000 608.380000 2962.500000 611.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 428.380000 -0.400000 431.380000 ;
        RECT 2920.400000 428.380000 2962.500000 431.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 248.380000 -0.400000 251.380000 ;
        RECT 2920.400000 248.380000 2962.500000 251.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880000 68.380000 -0.400000 71.380000 ;
        RECT 2920.400000 68.380000 2962.500000 71.380000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.180000 -32.820000 2957.800000 -29.820000 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2959.500000 -37.520000 2962.500000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2853.020000 -37.520000 2856.020000 -0.400000 ;
        RECT 2853.020000 3520.400000 2856.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2673.020000 -37.520000 2676.020000 -0.400000 ;
        RECT 2673.020000 3520.400000 2676.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2493.020000 -37.520000 2496.020000 -0.400000 ;
        RECT 2493.020000 3520.400000 2496.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2313.020000 -37.520000 2316.020000 -0.400000 ;
        RECT 2313.020000 3520.400000 2316.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2133.020000 -37.520000 2136.020000 -0.400000 ;
        RECT 2133.020000 3520.400000 2136.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1953.020000 -37.520000 1956.020000 -0.400000 ;
        RECT 1953.020000 3520.400000 1956.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1773.020000 -37.520000 1776.020000 -0.400000 ;
        RECT 1773.020000 3520.400000 1776.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1593.020000 -37.520000 1596.020000 -0.400000 ;
        RECT 1593.020000 3520.400000 1596.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1413.020000 -37.520000 1416.020000 -0.400000 ;
        RECT 1413.020000 3520.400000 1416.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1233.020000 -37.520000 1236.020000 -0.400000 ;
        RECT 1233.020000 3520.400000 1236.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1053.020000 -37.520000 1056.020000 -0.400000 ;
        RECT 1053.020000 3520.400000 1056.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 873.020000 -37.520000 876.020000 -0.400000 ;
        RECT 873.020000 3520.400000 876.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 693.020000 -37.520000 696.020000 -0.400000 ;
        RECT 693.020000 3520.400000 696.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 513.020000 -37.520000 516.020000 -0.400000 ;
        RECT 513.020000 3520.400000 516.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 333.020000 -37.520000 336.020000 -0.400000 ;
        RECT 333.020000 3520.400000 336.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 153.020000 -37.520000 156.020000 -0.400000 ;
        RECT 153.020000 3520.400000 156.020000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.880000 -37.520000 -39.880000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 3554.200000 2962.500000 3557.200000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 3398.380000 -0.400000 3401.380000 ;
        RECT 2920.400000 3398.380000 2962.500000 3401.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 3218.380000 -0.400000 3221.380000 ;
        RECT 2920.400000 3218.380000 2962.500000 3221.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 3038.380000 -0.400000 3041.380000 ;
        RECT 2920.400000 3038.380000 2962.500000 3041.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 2858.380000 -0.400000 2861.380000 ;
        RECT 2920.400000 2858.380000 2962.500000 2861.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 2678.380000 -0.400000 2681.380000 ;
        RECT 2920.400000 2678.380000 2962.500000 2681.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 2498.380000 -0.400000 2501.380000 ;
        RECT 2920.400000 2498.380000 2962.500000 2501.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 2318.380000 -0.400000 2321.380000 ;
        RECT 2920.400000 2318.380000 2962.500000 2321.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 2138.380000 -0.400000 2141.380000 ;
        RECT 2920.400000 2138.380000 2962.500000 2141.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 1958.380000 -0.400000 1961.380000 ;
        RECT 2920.400000 1958.380000 2962.500000 1961.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 1778.380000 -0.400000 1781.380000 ;
        RECT 2920.400000 1778.380000 2962.500000 1781.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 1598.380000 -0.400000 1601.380000 ;
        RECT 2920.400000 1598.380000 2962.500000 1601.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 1418.380000 -0.400000 1421.380000 ;
        RECT 2920.400000 1418.380000 2962.500000 1421.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 1238.380000 -0.400000 1241.380000 ;
        RECT 2920.400000 1238.380000 2962.500000 1241.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 1058.380000 -0.400000 1061.380000 ;
        RECT 2920.400000 1058.380000 2962.500000 1061.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 878.380000 -0.400000 881.380000 ;
        RECT 2920.400000 878.380000 2962.500000 881.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 698.380000 -0.400000 701.380000 ;
        RECT 2920.400000 698.380000 2962.500000 701.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 518.380000 -0.400000 521.380000 ;
        RECT 2920.400000 518.380000 2962.500000 521.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 338.380000 -0.400000 341.380000 ;
        RECT 2920.400000 338.380000 2962.500000 341.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 158.380000 -0.400000 161.380000 ;
        RECT 2920.400000 158.380000 2962.500000 161.380000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880000 -37.520000 2962.500000 -34.520000 ;
    END
  END vssa2
  OBS
      LAYER met5 ;
       RECT 0.000 0.000 2920.000 3520.000 ;
       RECT -42.880 -37.530 2962.500 3557.210 ;
        RECT -42.880000 3557.200000 -39.880000 3557.210000 ;
        RECT 153.020000 3557.200000 156.020000 3557.210000 ;
        RECT 333.020000 3557.200000 336.020000 3557.210000 ;
        RECT 513.020000 3557.200000 516.020000 3557.210000 ;
        RECT 693.020000 3557.200000 696.020000 3557.210000 ;
        RECT 873.020000 3557.200000 876.020000 3557.210000 ;
        RECT 1053.020000 3557.200000 1056.020000 3557.210000 ;
        RECT 1233.020000 3557.200000 1236.020000 3557.210000 ;
        RECT 1413.020000 3557.200000 1416.020000 3557.210000 ;
        RECT 1593.020000 3557.200000 1596.020000 3557.210000 ;
        RECT 1773.020000 3557.200000 1776.020000 3557.210000 ;
        RECT 1953.020000 3557.200000 1956.020000 3557.210000 ;
        RECT 2133.020000 3557.200000 2136.020000 3557.210000 ;
        RECT 2313.020000 3557.200000 2316.020000 3557.210000 ;
        RECT 2493.020000 3557.200000 2496.020000 3557.210000 ;
        RECT 2673.020000 3557.200000 2676.020000 3557.210000 ;
        RECT 2853.020000 3557.200000 2856.020000 3557.210000 ;
        RECT 2959.500000 3557.200000 2962.500000 3557.210000 ;
        RECT -42.880000 3554.190000 -39.880000 3554.200000 ;
        RECT 153.020000 3554.190000 156.020000 3554.200000 ;
        RECT 333.020000 3554.190000 336.020000 3554.200000 ;
        RECT 513.020000 3554.190000 516.020000 3554.200000 ;
        RECT 693.020000 3554.190000 696.020000 3554.200000 ;
        RECT 873.020000 3554.190000 876.020000 3554.200000 ;
        RECT 1053.020000 3554.190000 1056.020000 3554.200000 ;
        RECT 1233.020000 3554.190000 1236.020000 3554.200000 ;
        RECT 1413.020000 3554.190000 1416.020000 3554.200000 ;
        RECT 1593.020000 3554.190000 1596.020000 3554.200000 ;
        RECT 1773.020000 3554.190000 1776.020000 3554.200000 ;
        RECT 1953.020000 3554.190000 1956.020000 3554.200000 ;
        RECT 2133.020000 3554.190000 2136.020000 3554.200000 ;
        RECT 2313.020000 3554.190000 2316.020000 3554.200000 ;
        RECT 2493.020000 3554.190000 2496.020000 3554.200000 ;
        RECT 2673.020000 3554.190000 2676.020000 3554.200000 ;
        RECT 2853.020000 3554.190000 2856.020000 3554.200000 ;
        RECT 2959.500000 3554.190000 2962.500000 3554.200000 ;
        RECT -38.180000 3552.500000 -35.180000 3552.510000 ;
        RECT 63.020000 3552.500000 66.020000 3552.510000 ;
        RECT 243.020000 3552.500000 246.020000 3552.510000 ;
        RECT 423.020000 3552.500000 426.020000 3552.510000 ;
        RECT 603.020000 3552.500000 606.020000 3552.510000 ;
        RECT 783.020000 3552.500000 786.020000 3552.510000 ;
        RECT 963.020000 3552.500000 966.020000 3552.510000 ;
        RECT 1143.020000 3552.500000 1146.020000 3552.510000 ;
        RECT 1323.020000 3552.500000 1326.020000 3552.510000 ;
        RECT 1503.020000 3552.500000 1506.020000 3552.510000 ;
        RECT 1683.020000 3552.500000 1686.020000 3552.510000 ;
        RECT 1863.020000 3552.500000 1866.020000 3552.510000 ;
        RECT 2043.020000 3552.500000 2046.020000 3552.510000 ;
        RECT 2223.020000 3552.500000 2226.020000 3552.510000 ;
        RECT 2403.020000 3552.500000 2406.020000 3552.510000 ;
        RECT 2583.020000 3552.500000 2586.020000 3552.510000 ;
        RECT 2763.020000 3552.500000 2766.020000 3552.510000 ;
        RECT 2954.800000 3552.500000 2957.800000 3552.510000 ;
        RECT -38.180000 3549.490000 -35.180000 3549.500000 ;
        RECT 63.020000 3549.490000 66.020000 3549.500000 ;
        RECT 243.020000 3549.490000 246.020000 3549.500000 ;
        RECT 423.020000 3549.490000 426.020000 3549.500000 ;
        RECT 603.020000 3549.490000 606.020000 3549.500000 ;
        RECT 783.020000 3549.490000 786.020000 3549.500000 ;
        RECT 963.020000 3549.490000 966.020000 3549.500000 ;
        RECT 1143.020000 3549.490000 1146.020000 3549.500000 ;
        RECT 1323.020000 3549.490000 1326.020000 3549.500000 ;
        RECT 1503.020000 3549.490000 1506.020000 3549.500000 ;
        RECT 1683.020000 3549.490000 1686.020000 3549.500000 ;
        RECT 1863.020000 3549.490000 1866.020000 3549.500000 ;
        RECT 2043.020000 3549.490000 2046.020000 3549.500000 ;
        RECT 2223.020000 3549.490000 2226.020000 3549.500000 ;
        RECT 2403.020000 3549.490000 2406.020000 3549.500000 ;
        RECT 2583.020000 3549.490000 2586.020000 3549.500000 ;
        RECT 2763.020000 3549.490000 2766.020000 3549.500000 ;
        RECT 2954.800000 3549.490000 2957.800000 3549.500000 ;
        RECT -33.480000 3547.800000 -30.480000 3547.810000 ;
        RECT 135.020000 3547.800000 138.020000 3547.810000 ;
        RECT 315.020000 3547.800000 318.020000 3547.810000 ;
        RECT 495.020000 3547.800000 498.020000 3547.810000 ;
        RECT 675.020000 3547.800000 678.020000 3547.810000 ;
        RECT 855.020000 3547.800000 858.020000 3547.810000 ;
        RECT 1035.020000 3547.800000 1038.020000 3547.810000 ;
        RECT 1215.020000 3547.800000 1218.020000 3547.810000 ;
        RECT 1395.020000 3547.800000 1398.020000 3547.810000 ;
        RECT 1575.020000 3547.800000 1578.020000 3547.810000 ;
        RECT 1755.020000 3547.800000 1758.020000 3547.810000 ;
        RECT 1935.020000 3547.800000 1938.020000 3547.810000 ;
        RECT 2115.020000 3547.800000 2118.020000 3547.810000 ;
        RECT 2295.020000 3547.800000 2298.020000 3547.810000 ;
        RECT 2475.020000 3547.800000 2478.020000 3547.810000 ;
        RECT 2655.020000 3547.800000 2658.020000 3547.810000 ;
        RECT 2835.020000 3547.800000 2838.020000 3547.810000 ;
        RECT 2950.100000 3547.800000 2953.100000 3547.810000 ;
        RECT -33.480000 3544.790000 -30.480000 3544.800000 ;
        RECT 135.020000 3544.790000 138.020000 3544.800000 ;
        RECT 315.020000 3544.790000 318.020000 3544.800000 ;
        RECT 495.020000 3544.790000 498.020000 3544.800000 ;
        RECT 675.020000 3544.790000 678.020000 3544.800000 ;
        RECT 855.020000 3544.790000 858.020000 3544.800000 ;
        RECT 1035.020000 3544.790000 1038.020000 3544.800000 ;
        RECT 1215.020000 3544.790000 1218.020000 3544.800000 ;
        RECT 1395.020000 3544.790000 1398.020000 3544.800000 ;
        RECT 1575.020000 3544.790000 1578.020000 3544.800000 ;
        RECT 1755.020000 3544.790000 1758.020000 3544.800000 ;
        RECT 1935.020000 3544.790000 1938.020000 3544.800000 ;
        RECT 2115.020000 3544.790000 2118.020000 3544.800000 ;
        RECT 2295.020000 3544.790000 2298.020000 3544.800000 ;
        RECT 2475.020000 3544.790000 2478.020000 3544.800000 ;
        RECT 2655.020000 3544.790000 2658.020000 3544.800000 ;
        RECT 2835.020000 3544.790000 2838.020000 3544.800000 ;
        RECT 2950.100000 3544.790000 2953.100000 3544.800000 ;
        RECT -28.780000 3543.100000 -25.780000 3543.110000 ;
        RECT 45.020000 3543.100000 48.020000 3543.110000 ;
        RECT 225.020000 3543.100000 228.020000 3543.110000 ;
        RECT 405.020000 3543.100000 408.020000 3543.110000 ;
        RECT 585.020000 3543.100000 588.020000 3543.110000 ;
        RECT 765.020000 3543.100000 768.020000 3543.110000 ;
        RECT 945.020000 3543.100000 948.020000 3543.110000 ;
        RECT 1125.020000 3543.100000 1128.020000 3543.110000 ;
        RECT 1305.020000 3543.100000 1308.020000 3543.110000 ;
        RECT 1485.020000 3543.100000 1488.020000 3543.110000 ;
        RECT 1665.020000 3543.100000 1668.020000 3543.110000 ;
        RECT 1845.020000 3543.100000 1848.020000 3543.110000 ;
        RECT 2025.020000 3543.100000 2028.020000 3543.110000 ;
        RECT 2205.020000 3543.100000 2208.020000 3543.110000 ;
        RECT 2385.020000 3543.100000 2388.020000 3543.110000 ;
        RECT 2565.020000 3543.100000 2568.020000 3543.110000 ;
        RECT 2745.020000 3543.100000 2748.020000 3543.110000 ;
        RECT 2945.400000 3543.100000 2948.400000 3543.110000 ;
        RECT -28.780000 3540.090000 -25.780000 3540.100000 ;
        RECT 45.020000 3540.090000 48.020000 3540.100000 ;
        RECT 225.020000 3540.090000 228.020000 3540.100000 ;
        RECT 405.020000 3540.090000 408.020000 3540.100000 ;
        RECT 585.020000 3540.090000 588.020000 3540.100000 ;
        RECT 765.020000 3540.090000 768.020000 3540.100000 ;
        RECT 945.020000 3540.090000 948.020000 3540.100000 ;
        RECT 1125.020000 3540.090000 1128.020000 3540.100000 ;
        RECT 1305.020000 3540.090000 1308.020000 3540.100000 ;
        RECT 1485.020000 3540.090000 1488.020000 3540.100000 ;
        RECT 1665.020000 3540.090000 1668.020000 3540.100000 ;
        RECT 1845.020000 3540.090000 1848.020000 3540.100000 ;
        RECT 2025.020000 3540.090000 2028.020000 3540.100000 ;
        RECT 2205.020000 3540.090000 2208.020000 3540.100000 ;
        RECT 2385.020000 3540.090000 2388.020000 3540.100000 ;
        RECT 2565.020000 3540.090000 2568.020000 3540.100000 ;
        RECT 2745.020000 3540.090000 2748.020000 3540.100000 ;
        RECT 2945.400000 3540.090000 2948.400000 3540.100000 ;
        RECT -24.080000 3538.400000 -21.080000 3538.410000 ;
        RECT 117.020000 3538.400000 120.020000 3538.410000 ;
        RECT 297.020000 3538.400000 300.020000 3538.410000 ;
        RECT 477.020000 3538.400000 480.020000 3538.410000 ;
        RECT 657.020000 3538.400000 660.020000 3538.410000 ;
        RECT 837.020000 3538.400000 840.020000 3538.410000 ;
        RECT 1017.020000 3538.400000 1020.020000 3538.410000 ;
        RECT 1197.020000 3538.400000 1200.020000 3538.410000 ;
        RECT 1377.020000 3538.400000 1380.020000 3538.410000 ;
        RECT 1557.020000 3538.400000 1560.020000 3538.410000 ;
        RECT 1737.020000 3538.400000 1740.020000 3538.410000 ;
        RECT 1917.020000 3538.400000 1920.020000 3538.410000 ;
        RECT 2097.020000 3538.400000 2100.020000 3538.410000 ;
        RECT 2277.020000 3538.400000 2280.020000 3538.410000 ;
        RECT 2457.020000 3538.400000 2460.020000 3538.410000 ;
        RECT 2637.020000 3538.400000 2640.020000 3538.410000 ;
        RECT 2817.020000 3538.400000 2820.020000 3538.410000 ;
        RECT 2940.700000 3538.400000 2943.700000 3538.410000 ;
        RECT -24.080000 3535.390000 -21.080000 3535.400000 ;
        RECT 117.020000 3535.390000 120.020000 3535.400000 ;
        RECT 297.020000 3535.390000 300.020000 3535.400000 ;
        RECT 477.020000 3535.390000 480.020000 3535.400000 ;
        RECT 657.020000 3535.390000 660.020000 3535.400000 ;
        RECT 837.020000 3535.390000 840.020000 3535.400000 ;
        RECT 1017.020000 3535.390000 1020.020000 3535.400000 ;
        RECT 1197.020000 3535.390000 1200.020000 3535.400000 ;
        RECT 1377.020000 3535.390000 1380.020000 3535.400000 ;
        RECT 1557.020000 3535.390000 1560.020000 3535.400000 ;
        RECT 1737.020000 3535.390000 1740.020000 3535.400000 ;
        RECT 1917.020000 3535.390000 1920.020000 3535.400000 ;
        RECT 2097.020000 3535.390000 2100.020000 3535.400000 ;
        RECT 2277.020000 3535.390000 2280.020000 3535.400000 ;
        RECT 2457.020000 3535.390000 2460.020000 3535.400000 ;
        RECT 2637.020000 3535.390000 2640.020000 3535.400000 ;
        RECT 2817.020000 3535.390000 2820.020000 3535.400000 ;
        RECT 2940.700000 3535.390000 2943.700000 3535.400000 ;
        RECT -19.380000 3533.700000 -16.380000 3533.710000 ;
        RECT 27.020000 3533.700000 30.020000 3533.710000 ;
        RECT 207.020000 3533.700000 210.020000 3533.710000 ;
        RECT 387.020000 3533.700000 390.020000 3533.710000 ;
        RECT 567.020000 3533.700000 570.020000 3533.710000 ;
        RECT 747.020000 3533.700000 750.020000 3533.710000 ;
        RECT 927.020000 3533.700000 930.020000 3533.710000 ;
        RECT 1107.020000 3533.700000 1110.020000 3533.710000 ;
        RECT 1287.020000 3533.700000 1290.020000 3533.710000 ;
        RECT 1467.020000 3533.700000 1470.020000 3533.710000 ;
        RECT 1647.020000 3533.700000 1650.020000 3533.710000 ;
        RECT 1827.020000 3533.700000 1830.020000 3533.710000 ;
        RECT 2007.020000 3533.700000 2010.020000 3533.710000 ;
        RECT 2187.020000 3533.700000 2190.020000 3533.710000 ;
        RECT 2367.020000 3533.700000 2370.020000 3533.710000 ;
        RECT 2547.020000 3533.700000 2550.020000 3533.710000 ;
        RECT 2727.020000 3533.700000 2730.020000 3533.710000 ;
        RECT 2907.020000 3533.700000 2910.020000 3533.710000 ;
        RECT 2936.000000 3533.700000 2939.000000 3533.710000 ;
        RECT -19.380000 3530.690000 -16.380000 3530.700000 ;
        RECT 27.020000 3530.690000 30.020000 3530.700000 ;
        RECT 207.020000 3530.690000 210.020000 3530.700000 ;
        RECT 387.020000 3530.690000 390.020000 3530.700000 ;
        RECT 567.020000 3530.690000 570.020000 3530.700000 ;
        RECT 747.020000 3530.690000 750.020000 3530.700000 ;
        RECT 927.020000 3530.690000 930.020000 3530.700000 ;
        RECT 1107.020000 3530.690000 1110.020000 3530.700000 ;
        RECT 1287.020000 3530.690000 1290.020000 3530.700000 ;
        RECT 1467.020000 3530.690000 1470.020000 3530.700000 ;
        RECT 1647.020000 3530.690000 1650.020000 3530.700000 ;
        RECT 1827.020000 3530.690000 1830.020000 3530.700000 ;
        RECT 2007.020000 3530.690000 2010.020000 3530.700000 ;
        RECT 2187.020000 3530.690000 2190.020000 3530.700000 ;
        RECT 2367.020000 3530.690000 2370.020000 3530.700000 ;
        RECT 2547.020000 3530.690000 2550.020000 3530.700000 ;
        RECT 2727.020000 3530.690000 2730.020000 3530.700000 ;
        RECT 2907.020000 3530.690000 2910.020000 3530.700000 ;
        RECT 2936.000000 3530.690000 2939.000000 3530.700000 ;
        RECT -14.680000 3529.000000 -11.680000 3529.010000 ;
        RECT 99.020000 3529.000000 102.020000 3529.010000 ;
        RECT 279.020000 3529.000000 282.020000 3529.010000 ;
        RECT 459.020000 3529.000000 462.020000 3529.010000 ;
        RECT 639.020000 3529.000000 642.020000 3529.010000 ;
        RECT 819.020000 3529.000000 822.020000 3529.010000 ;
        RECT 999.020000 3529.000000 1002.020000 3529.010000 ;
        RECT 1179.020000 3529.000000 1182.020000 3529.010000 ;
        RECT 1359.020000 3529.000000 1362.020000 3529.010000 ;
        RECT 1539.020000 3529.000000 1542.020000 3529.010000 ;
        RECT 1719.020000 3529.000000 1722.020000 3529.010000 ;
        RECT 1899.020000 3529.000000 1902.020000 3529.010000 ;
        RECT 2079.020000 3529.000000 2082.020000 3529.010000 ;
        RECT 2259.020000 3529.000000 2262.020000 3529.010000 ;
        RECT 2439.020000 3529.000000 2442.020000 3529.010000 ;
        RECT 2619.020000 3529.000000 2622.020000 3529.010000 ;
        RECT 2799.020000 3529.000000 2802.020000 3529.010000 ;
        RECT 2931.300000 3529.000000 2934.300000 3529.010000 ;
        RECT -14.680000 3525.990000 -11.680000 3526.000000 ;
        RECT 99.020000 3525.990000 102.020000 3526.000000 ;
        RECT 279.020000 3525.990000 282.020000 3526.000000 ;
        RECT 459.020000 3525.990000 462.020000 3526.000000 ;
        RECT 639.020000 3525.990000 642.020000 3526.000000 ;
        RECT 819.020000 3525.990000 822.020000 3526.000000 ;
        RECT 999.020000 3525.990000 1002.020000 3526.000000 ;
        RECT 1179.020000 3525.990000 1182.020000 3526.000000 ;
        RECT 1359.020000 3525.990000 1362.020000 3526.000000 ;
        RECT 1539.020000 3525.990000 1542.020000 3526.000000 ;
        RECT 1719.020000 3525.990000 1722.020000 3526.000000 ;
        RECT 1899.020000 3525.990000 1902.020000 3526.000000 ;
        RECT 2079.020000 3525.990000 2082.020000 3526.000000 ;
        RECT 2259.020000 3525.990000 2262.020000 3526.000000 ;
        RECT 2439.020000 3525.990000 2442.020000 3526.000000 ;
        RECT 2619.020000 3525.990000 2622.020000 3526.000000 ;
        RECT 2799.020000 3525.990000 2802.020000 3526.000000 ;
        RECT 2931.300000 3525.990000 2934.300000 3526.000000 ;
        RECT -9.980000 3524.300000 -6.980000 3524.310000 ;
        RECT 9.020000 3524.300000 12.020000 3524.310000 ;
        RECT 189.020000 3524.300000 192.020000 3524.310000 ;
        RECT 369.020000 3524.300000 372.020000 3524.310000 ;
        RECT 549.020000 3524.300000 552.020000 3524.310000 ;
        RECT 729.020000 3524.300000 732.020000 3524.310000 ;
        RECT 909.020000 3524.300000 912.020000 3524.310000 ;
        RECT 1089.020000 3524.300000 1092.020000 3524.310000 ;
        RECT 1269.020000 3524.300000 1272.020000 3524.310000 ;
        RECT 1449.020000 3524.300000 1452.020000 3524.310000 ;
        RECT 1629.020000 3524.300000 1632.020000 3524.310000 ;
        RECT 1809.020000 3524.300000 1812.020000 3524.310000 ;
        RECT 1989.020000 3524.300000 1992.020000 3524.310000 ;
        RECT 2169.020000 3524.300000 2172.020000 3524.310000 ;
        RECT 2349.020000 3524.300000 2352.020000 3524.310000 ;
        RECT 2529.020000 3524.300000 2532.020000 3524.310000 ;
        RECT 2709.020000 3524.300000 2712.020000 3524.310000 ;
        RECT 2889.020000 3524.300000 2892.020000 3524.310000 ;
        RECT 2926.600000 3524.300000 2929.600000 3524.310000 ;
        RECT -9.980000 3521.290000 -6.980000 3521.300000 ;
        RECT 9.020000 3521.290000 12.020000 3521.300000 ;
        RECT 189.020000 3521.290000 192.020000 3521.300000 ;
        RECT 369.020000 3521.290000 372.020000 3521.300000 ;
        RECT 549.020000 3521.290000 552.020000 3521.300000 ;
        RECT 729.020000 3521.290000 732.020000 3521.300000 ;
        RECT 909.020000 3521.290000 912.020000 3521.300000 ;
        RECT 1089.020000 3521.290000 1092.020000 3521.300000 ;
        RECT 1269.020000 3521.290000 1272.020000 3521.300000 ;
        RECT 1449.020000 3521.290000 1452.020000 3521.300000 ;
        RECT 1629.020000 3521.290000 1632.020000 3521.300000 ;
        RECT 1809.020000 3521.290000 1812.020000 3521.300000 ;
        RECT 1989.020000 3521.290000 1992.020000 3521.300000 ;
        RECT 2169.020000 3521.290000 2172.020000 3521.300000 ;
        RECT 2349.020000 3521.290000 2352.020000 3521.300000 ;
        RECT 2529.020000 3521.290000 2532.020000 3521.300000 ;
        RECT 2709.020000 3521.290000 2712.020000 3521.300000 ;
        RECT 2889.020000 3521.290000 2892.020000 3521.300000 ;
        RECT 2926.600000 3521.290000 2929.600000 3521.300000 ;
        RECT -38.180000 3491.380000 -35.180000 3491.390000 ;
        RECT 2954.800000 3491.380000 2957.800000 3491.390000 ;
        RECT -38.180000 3488.370000 -35.180000 3488.380000 ;
        RECT 2954.800000 3488.370000 2957.800000 3488.380000 ;
        RECT -28.780000 3473.380000 -25.780000 3473.390000 ;
        RECT 2945.400000 3473.380000 2948.400000 3473.390000 ;
        RECT -28.780000 3470.370000 -25.780000 3470.380000 ;
        RECT 2945.400000 3470.370000 2948.400000 3470.380000 ;
        RECT -19.380000 3455.380000 -16.380000 3455.390000 ;
        RECT 2936.000000 3455.380000 2939.000000 3455.390000 ;
        RECT -19.380000 3452.370000 -16.380000 3452.380000 ;
        RECT 2936.000000 3452.370000 2939.000000 3452.380000 ;
        RECT -9.980000 3437.140000 -6.980000 3437.150000 ;
        RECT 2926.600000 3437.140000 2929.600000 3437.150000 ;
        RECT -9.980000 3434.130000 -6.980000 3434.140000 ;
        RECT 2926.600000 3434.130000 2929.600000 3434.140000 ;
        RECT -42.880000 3401.380000 -39.880000 3401.390000 ;
        RECT 2959.500000 3401.380000 2962.500000 3401.390000 ;
        RECT -42.880000 3398.370000 -39.880000 3398.380000 ;
        RECT 2959.500000 3398.370000 2962.500000 3398.380000 ;
        RECT -33.480000 3383.380000 -30.480000 3383.390000 ;
        RECT 2950.100000 3383.380000 2953.100000 3383.390000 ;
        RECT -33.480000 3380.370000 -30.480000 3380.380000 ;
        RECT 2950.100000 3380.370000 2953.100000 3380.380000 ;
        RECT -24.080000 3365.380000 -21.080000 3365.390000 ;
        RECT 2940.700000 3365.380000 2943.700000 3365.390000 ;
        RECT -24.080000 3362.370000 -21.080000 3362.380000 ;
        RECT 2940.700000 3362.370000 2943.700000 3362.380000 ;
        RECT -14.680000 3347.140000 -11.680000 3347.150000 ;
        RECT 2931.300000 3347.140000 2934.300000 3347.150000 ;
        RECT -14.680000 3344.130000 -11.680000 3344.140000 ;
        RECT 2931.300000 3344.130000 2934.300000 3344.140000 ;
        RECT -38.180000 3311.380000 -35.180000 3311.390000 ;
        RECT 2954.800000 3311.380000 2957.800000 3311.390000 ;
        RECT -38.180000 3308.370000 -35.180000 3308.380000 ;
        RECT 2954.800000 3308.370000 2957.800000 3308.380000 ;
        RECT -28.780000 3293.380000 -25.780000 3293.390000 ;
        RECT 2945.400000 3293.380000 2948.400000 3293.390000 ;
        RECT -28.780000 3290.370000 -25.780000 3290.380000 ;
        RECT 2945.400000 3290.370000 2948.400000 3290.380000 ;
        RECT -19.380000 3275.380000 -16.380000 3275.390000 ;
        RECT 2936.000000 3275.380000 2939.000000 3275.390000 ;
        RECT -19.380000 3272.370000 -16.380000 3272.380000 ;
        RECT 2936.000000 3272.370000 2939.000000 3272.380000 ;
        RECT -9.980000 3257.140000 -6.980000 3257.150000 ;
        RECT 2926.600000 3257.140000 2929.600000 3257.150000 ;
        RECT -9.980000 3254.130000 -6.980000 3254.140000 ;
        RECT 2926.600000 3254.130000 2929.600000 3254.140000 ;
        RECT -42.880000 3221.380000 -39.880000 3221.390000 ;
        RECT 2959.500000 3221.380000 2962.500000 3221.390000 ;
        RECT -42.880000 3218.370000 -39.880000 3218.380000 ;
        RECT 2959.500000 3218.370000 2962.500000 3218.380000 ;
        RECT -33.480000 3203.380000 -30.480000 3203.390000 ;
        RECT 2950.100000 3203.380000 2953.100000 3203.390000 ;
        RECT -33.480000 3200.370000 -30.480000 3200.380000 ;
        RECT 2950.100000 3200.370000 2953.100000 3200.380000 ;
        RECT -24.080000 3185.380000 -21.080000 3185.390000 ;
        RECT 2940.700000 3185.380000 2943.700000 3185.390000 ;
        RECT -24.080000 3182.370000 -21.080000 3182.380000 ;
        RECT 2940.700000 3182.370000 2943.700000 3182.380000 ;
        RECT -14.680000 3167.140000 -11.680000 3167.150000 ;
        RECT 2931.300000 3167.140000 2934.300000 3167.150000 ;
        RECT -14.680000 3164.130000 -11.680000 3164.140000 ;
        RECT 2931.300000 3164.130000 2934.300000 3164.140000 ;
        RECT -38.180000 3131.380000 -35.180000 3131.390000 ;
        RECT 2954.800000 3131.380000 2957.800000 3131.390000 ;
        RECT -38.180000 3128.370000 -35.180000 3128.380000 ;
        RECT 2954.800000 3128.370000 2957.800000 3128.380000 ;
        RECT -28.780000 3113.380000 -25.780000 3113.390000 ;
        RECT 2945.400000 3113.380000 2948.400000 3113.390000 ;
        RECT -28.780000 3110.370000 -25.780000 3110.380000 ;
        RECT 2945.400000 3110.370000 2948.400000 3110.380000 ;
        RECT -19.380000 3095.380000 -16.380000 3095.390000 ;
        RECT 2936.000000 3095.380000 2939.000000 3095.390000 ;
        RECT -19.380000 3092.370000 -16.380000 3092.380000 ;
        RECT 2936.000000 3092.370000 2939.000000 3092.380000 ;
        RECT -9.980000 3077.140000 -6.980000 3077.150000 ;
        RECT 2926.600000 3077.140000 2929.600000 3077.150000 ;
        RECT -9.980000 3074.130000 -6.980000 3074.140000 ;
        RECT 2926.600000 3074.130000 2929.600000 3074.140000 ;
        RECT -42.880000 3041.380000 -39.880000 3041.390000 ;
        RECT 2959.500000 3041.380000 2962.500000 3041.390000 ;
        RECT -42.880000 3038.370000 -39.880000 3038.380000 ;
        RECT 2959.500000 3038.370000 2962.500000 3038.380000 ;
        RECT -33.480000 3023.380000 -30.480000 3023.390000 ;
        RECT 2950.100000 3023.380000 2953.100000 3023.390000 ;
        RECT -33.480000 3020.370000 -30.480000 3020.380000 ;
        RECT 2950.100000 3020.370000 2953.100000 3020.380000 ;
        RECT -24.080000 3005.380000 -21.080000 3005.390000 ;
        RECT 2940.700000 3005.380000 2943.700000 3005.390000 ;
        RECT -24.080000 3002.370000 -21.080000 3002.380000 ;
        RECT 2940.700000 3002.370000 2943.700000 3002.380000 ;
        RECT -14.680000 2987.140000 -11.680000 2987.150000 ;
        RECT 2931.300000 2987.140000 2934.300000 2987.150000 ;
        RECT -14.680000 2984.130000 -11.680000 2984.140000 ;
        RECT 2931.300000 2984.130000 2934.300000 2984.140000 ;
        RECT -38.180000 2951.380000 -35.180000 2951.390000 ;
        RECT 2954.800000 2951.380000 2957.800000 2951.390000 ;
        RECT -38.180000 2948.370000 -35.180000 2948.380000 ;
        RECT 2954.800000 2948.370000 2957.800000 2948.380000 ;
        RECT -28.780000 2933.380000 -25.780000 2933.390000 ;
        RECT 2945.400000 2933.380000 2948.400000 2933.390000 ;
        RECT -28.780000 2930.370000 -25.780000 2930.380000 ;
        RECT 2945.400000 2930.370000 2948.400000 2930.380000 ;
        RECT -19.380000 2915.380000 -16.380000 2915.390000 ;
        RECT 2936.000000 2915.380000 2939.000000 2915.390000 ;
        RECT -19.380000 2912.370000 -16.380000 2912.380000 ;
        RECT 2936.000000 2912.370000 2939.000000 2912.380000 ;
        RECT -9.980000 2897.140000 -6.980000 2897.150000 ;
        RECT 2926.600000 2897.140000 2929.600000 2897.150000 ;
        RECT -9.980000 2894.130000 -6.980000 2894.140000 ;
        RECT 2926.600000 2894.130000 2929.600000 2894.140000 ;
        RECT -42.880000 2861.380000 -39.880000 2861.390000 ;
        RECT 2959.500000 2861.380000 2962.500000 2861.390000 ;
        RECT -42.880000 2858.370000 -39.880000 2858.380000 ;
        RECT 2959.500000 2858.370000 2962.500000 2858.380000 ;
        RECT -33.480000 2843.380000 -30.480000 2843.390000 ;
        RECT 2950.100000 2843.380000 2953.100000 2843.390000 ;
        RECT -33.480000 2840.370000 -30.480000 2840.380000 ;
        RECT 2950.100000 2840.370000 2953.100000 2840.380000 ;
        RECT -24.080000 2825.380000 -21.080000 2825.390000 ;
        RECT 2940.700000 2825.380000 2943.700000 2825.390000 ;
        RECT -24.080000 2822.370000 -21.080000 2822.380000 ;
        RECT 2940.700000 2822.370000 2943.700000 2822.380000 ;
        RECT -14.680000 2807.140000 -11.680000 2807.150000 ;
        RECT 2931.300000 2807.140000 2934.300000 2807.150000 ;
        RECT -14.680000 2804.130000 -11.680000 2804.140000 ;
        RECT 2931.300000 2804.130000 2934.300000 2804.140000 ;
        RECT -38.180000 2771.380000 -35.180000 2771.390000 ;
        RECT 2954.800000 2771.380000 2957.800000 2771.390000 ;
        RECT -38.180000 2768.370000 -35.180000 2768.380000 ;
        RECT 2954.800000 2768.370000 2957.800000 2768.380000 ;
        RECT -28.780000 2753.380000 -25.780000 2753.390000 ;
        RECT 2945.400000 2753.380000 2948.400000 2753.390000 ;
        RECT -28.780000 2750.370000 -25.780000 2750.380000 ;
        RECT 2945.400000 2750.370000 2948.400000 2750.380000 ;
        RECT -19.380000 2735.380000 -16.380000 2735.390000 ;
        RECT 2936.000000 2735.380000 2939.000000 2735.390000 ;
        RECT -19.380000 2732.370000 -16.380000 2732.380000 ;
        RECT 2936.000000 2732.370000 2939.000000 2732.380000 ;
        RECT -9.980000 2717.140000 -6.980000 2717.150000 ;
        RECT 2926.600000 2717.140000 2929.600000 2717.150000 ;
        RECT -9.980000 2714.130000 -6.980000 2714.140000 ;
        RECT 2926.600000 2714.130000 2929.600000 2714.140000 ;
        RECT -42.880000 2681.380000 -39.880000 2681.390000 ;
        RECT 2959.500000 2681.380000 2962.500000 2681.390000 ;
        RECT -42.880000 2678.370000 -39.880000 2678.380000 ;
        RECT 2959.500000 2678.370000 2962.500000 2678.380000 ;
        RECT -33.480000 2663.380000 -30.480000 2663.390000 ;
        RECT 2950.100000 2663.380000 2953.100000 2663.390000 ;
        RECT -33.480000 2660.370000 -30.480000 2660.380000 ;
        RECT 2950.100000 2660.370000 2953.100000 2660.380000 ;
        RECT -24.080000 2645.380000 -21.080000 2645.390000 ;
        RECT 2940.700000 2645.380000 2943.700000 2645.390000 ;
        RECT -24.080000 2642.370000 -21.080000 2642.380000 ;
        RECT 2940.700000 2642.370000 2943.700000 2642.380000 ;
        RECT -14.680000 2627.140000 -11.680000 2627.150000 ;
        RECT 2931.300000 2627.140000 2934.300000 2627.150000 ;
        RECT -14.680000 2624.130000 -11.680000 2624.140000 ;
        RECT 2931.300000 2624.130000 2934.300000 2624.140000 ;
        RECT -38.180000 2591.380000 -35.180000 2591.390000 ;
        RECT 2954.800000 2591.380000 2957.800000 2591.390000 ;
        RECT -38.180000 2588.370000 -35.180000 2588.380000 ;
        RECT 2954.800000 2588.370000 2957.800000 2588.380000 ;
        RECT -28.780000 2573.380000 -25.780000 2573.390000 ;
        RECT 2945.400000 2573.380000 2948.400000 2573.390000 ;
        RECT -28.780000 2570.370000 -25.780000 2570.380000 ;
        RECT 2945.400000 2570.370000 2948.400000 2570.380000 ;
        RECT -19.380000 2555.380000 -16.380000 2555.390000 ;
        RECT 2936.000000 2555.380000 2939.000000 2555.390000 ;
        RECT -19.380000 2552.370000 -16.380000 2552.380000 ;
        RECT 2936.000000 2552.370000 2939.000000 2552.380000 ;
        RECT -9.980000 2537.140000 -6.980000 2537.150000 ;
        RECT 2926.600000 2537.140000 2929.600000 2537.150000 ;
        RECT -9.980000 2534.130000 -6.980000 2534.140000 ;
        RECT 2926.600000 2534.130000 2929.600000 2534.140000 ;
        RECT -42.880000 2501.380000 -39.880000 2501.390000 ;
        RECT 2959.500000 2501.380000 2962.500000 2501.390000 ;
        RECT -42.880000 2498.370000 -39.880000 2498.380000 ;
        RECT 2959.500000 2498.370000 2962.500000 2498.380000 ;
        RECT -33.480000 2483.380000 -30.480000 2483.390000 ;
        RECT 2950.100000 2483.380000 2953.100000 2483.390000 ;
        RECT -33.480000 2480.370000 -30.480000 2480.380000 ;
        RECT 2950.100000 2480.370000 2953.100000 2480.380000 ;
        RECT -24.080000 2465.380000 -21.080000 2465.390000 ;
        RECT 2940.700000 2465.380000 2943.700000 2465.390000 ;
        RECT -24.080000 2462.370000 -21.080000 2462.380000 ;
        RECT 2940.700000 2462.370000 2943.700000 2462.380000 ;
        RECT -14.680000 2447.140000 -11.680000 2447.150000 ;
        RECT 2931.300000 2447.140000 2934.300000 2447.150000 ;
        RECT -14.680000 2444.130000 -11.680000 2444.140000 ;
        RECT 2931.300000 2444.130000 2934.300000 2444.140000 ;
        RECT -38.180000 2411.380000 -35.180000 2411.390000 ;
        RECT 2954.800000 2411.380000 2957.800000 2411.390000 ;
        RECT -38.180000 2408.370000 -35.180000 2408.380000 ;
        RECT 2954.800000 2408.370000 2957.800000 2408.380000 ;
        RECT -28.780000 2393.380000 -25.780000 2393.390000 ;
        RECT 2945.400000 2393.380000 2948.400000 2393.390000 ;
        RECT -28.780000 2390.370000 -25.780000 2390.380000 ;
        RECT 2945.400000 2390.370000 2948.400000 2390.380000 ;
        RECT -19.380000 2375.380000 -16.380000 2375.390000 ;
        RECT 2936.000000 2375.380000 2939.000000 2375.390000 ;
        RECT -19.380000 2372.370000 -16.380000 2372.380000 ;
        RECT 2936.000000 2372.370000 2939.000000 2372.380000 ;
        RECT -9.980000 2357.140000 -6.980000 2357.150000 ;
        RECT 2926.600000 2357.140000 2929.600000 2357.150000 ;
        RECT -9.980000 2354.130000 -6.980000 2354.140000 ;
        RECT 2926.600000 2354.130000 2929.600000 2354.140000 ;
        RECT -42.880000 2321.380000 -39.880000 2321.390000 ;
        RECT 2959.500000 2321.380000 2962.500000 2321.390000 ;
        RECT -42.880000 2318.370000 -39.880000 2318.380000 ;
        RECT 2959.500000 2318.370000 2962.500000 2318.380000 ;
        RECT -33.480000 2303.380000 -30.480000 2303.390000 ;
        RECT 2950.100000 2303.380000 2953.100000 2303.390000 ;
        RECT -33.480000 2300.370000 -30.480000 2300.380000 ;
        RECT 2950.100000 2300.370000 2953.100000 2300.380000 ;
        RECT -24.080000 2285.380000 -21.080000 2285.390000 ;
        RECT 2940.700000 2285.380000 2943.700000 2285.390000 ;
        RECT -24.080000 2282.370000 -21.080000 2282.380000 ;
        RECT 2940.700000 2282.370000 2943.700000 2282.380000 ;
        RECT -14.680000 2267.140000 -11.680000 2267.150000 ;
        RECT 2931.300000 2267.140000 2934.300000 2267.150000 ;
        RECT -14.680000 2264.130000 -11.680000 2264.140000 ;
        RECT 2931.300000 2264.130000 2934.300000 2264.140000 ;
        RECT -38.180000 2231.380000 -35.180000 2231.390000 ;
        RECT 2954.800000 2231.380000 2957.800000 2231.390000 ;
        RECT -38.180000 2228.370000 -35.180000 2228.380000 ;
        RECT 2954.800000 2228.370000 2957.800000 2228.380000 ;
        RECT -28.780000 2213.380000 -25.780000 2213.390000 ;
        RECT 2945.400000 2213.380000 2948.400000 2213.390000 ;
        RECT -28.780000 2210.370000 -25.780000 2210.380000 ;
        RECT 2945.400000 2210.370000 2948.400000 2210.380000 ;
        RECT -19.380000 2195.380000 -16.380000 2195.390000 ;
        RECT 2936.000000 2195.380000 2939.000000 2195.390000 ;
        RECT -19.380000 2192.370000 -16.380000 2192.380000 ;
        RECT 2936.000000 2192.370000 2939.000000 2192.380000 ;
        RECT -9.980000 2177.140000 -6.980000 2177.150000 ;
        RECT 2926.600000 2177.140000 2929.600000 2177.150000 ;
        RECT -9.980000 2174.130000 -6.980000 2174.140000 ;
        RECT 2926.600000 2174.130000 2929.600000 2174.140000 ;
        RECT -42.880000 2141.380000 -39.880000 2141.390000 ;
        RECT 2959.500000 2141.380000 2962.500000 2141.390000 ;
        RECT -42.880000 2138.370000 -39.880000 2138.380000 ;
        RECT 2959.500000 2138.370000 2962.500000 2138.380000 ;
        RECT -33.480000 2123.380000 -30.480000 2123.390000 ;
        RECT 2950.100000 2123.380000 2953.100000 2123.390000 ;
        RECT -33.480000 2120.370000 -30.480000 2120.380000 ;
        RECT 2950.100000 2120.370000 2953.100000 2120.380000 ;
        RECT -24.080000 2105.380000 -21.080000 2105.390000 ;
        RECT 2940.700000 2105.380000 2943.700000 2105.390000 ;
        RECT -24.080000 2102.370000 -21.080000 2102.380000 ;
        RECT 2940.700000 2102.370000 2943.700000 2102.380000 ;
        RECT -14.680000 2087.140000 -11.680000 2087.150000 ;
        RECT 2931.300000 2087.140000 2934.300000 2087.150000 ;
        RECT -14.680000 2084.130000 -11.680000 2084.140000 ;
        RECT 2931.300000 2084.130000 2934.300000 2084.140000 ;
        RECT -38.180000 2051.380000 -35.180000 2051.390000 ;
        RECT 2954.800000 2051.380000 2957.800000 2051.390000 ;
        RECT -38.180000 2048.370000 -35.180000 2048.380000 ;
        RECT 2954.800000 2048.370000 2957.800000 2048.380000 ;
        RECT -28.780000 2033.380000 -25.780000 2033.390000 ;
        RECT 2945.400000 2033.380000 2948.400000 2033.390000 ;
        RECT -28.780000 2030.370000 -25.780000 2030.380000 ;
        RECT 2945.400000 2030.370000 2948.400000 2030.380000 ;
        RECT -19.380000 2015.380000 -16.380000 2015.390000 ;
        RECT 2936.000000 2015.380000 2939.000000 2015.390000 ;
        RECT -19.380000 2012.370000 -16.380000 2012.380000 ;
        RECT 2936.000000 2012.370000 2939.000000 2012.380000 ;
        RECT -9.980000 1997.140000 -6.980000 1997.150000 ;
        RECT 2926.600000 1997.140000 2929.600000 1997.150000 ;
        RECT -9.980000 1994.130000 -6.980000 1994.140000 ;
        RECT 2926.600000 1994.130000 2929.600000 1994.140000 ;
        RECT -42.880000 1961.380000 -39.880000 1961.390000 ;
        RECT 2959.500000 1961.380000 2962.500000 1961.390000 ;
        RECT -42.880000 1958.370000 -39.880000 1958.380000 ;
        RECT 2959.500000 1958.370000 2962.500000 1958.380000 ;
        RECT -33.480000 1943.380000 -30.480000 1943.390000 ;
        RECT 2950.100000 1943.380000 2953.100000 1943.390000 ;
        RECT -33.480000 1940.370000 -30.480000 1940.380000 ;
        RECT 2950.100000 1940.370000 2953.100000 1940.380000 ;
        RECT -24.080000 1925.380000 -21.080000 1925.390000 ;
        RECT 2940.700000 1925.380000 2943.700000 1925.390000 ;
        RECT -24.080000 1922.370000 -21.080000 1922.380000 ;
        RECT 2940.700000 1922.370000 2943.700000 1922.380000 ;
        RECT -14.680000 1907.140000 -11.680000 1907.150000 ;
        RECT 2931.300000 1907.140000 2934.300000 1907.150000 ;
        RECT -14.680000 1904.130000 -11.680000 1904.140000 ;
        RECT 2931.300000 1904.130000 2934.300000 1904.140000 ;
        RECT -38.180000 1871.380000 -35.180000 1871.390000 ;
        RECT 2954.800000 1871.380000 2957.800000 1871.390000 ;
        RECT -38.180000 1868.370000 -35.180000 1868.380000 ;
        RECT 2954.800000 1868.370000 2957.800000 1868.380000 ;
        RECT -28.780000 1853.380000 -25.780000 1853.390000 ;
        RECT 2945.400000 1853.380000 2948.400000 1853.390000 ;
        RECT -28.780000 1850.370000 -25.780000 1850.380000 ;
        RECT 2945.400000 1850.370000 2948.400000 1850.380000 ;
        RECT -19.380000 1835.380000 -16.380000 1835.390000 ;
        RECT 2936.000000 1835.380000 2939.000000 1835.390000 ;
        RECT -19.380000 1832.370000 -16.380000 1832.380000 ;
        RECT 2936.000000 1832.370000 2939.000000 1832.380000 ;
        RECT -9.980000 1817.140000 -6.980000 1817.150000 ;
        RECT 2926.600000 1817.140000 2929.600000 1817.150000 ;
        RECT -9.980000 1814.130000 -6.980000 1814.140000 ;
        RECT 2926.600000 1814.130000 2929.600000 1814.140000 ;
        RECT -42.880000 1781.380000 -39.880000 1781.390000 ;
        RECT 2959.500000 1781.380000 2962.500000 1781.390000 ;
        RECT -42.880000 1778.370000 -39.880000 1778.380000 ;
        RECT 2959.500000 1778.370000 2962.500000 1778.380000 ;
        RECT -33.480000 1763.380000 -30.480000 1763.390000 ;
        RECT 2950.100000 1763.380000 2953.100000 1763.390000 ;
        RECT -33.480000 1760.370000 -30.480000 1760.380000 ;
        RECT 2950.100000 1760.370000 2953.100000 1760.380000 ;
        RECT -24.080000 1745.380000 -21.080000 1745.390000 ;
        RECT 2940.700000 1745.380000 2943.700000 1745.390000 ;
        RECT -24.080000 1742.370000 -21.080000 1742.380000 ;
        RECT 2940.700000 1742.370000 2943.700000 1742.380000 ;
        RECT -14.680000 1727.140000 -11.680000 1727.150000 ;
        RECT 2931.300000 1727.140000 2934.300000 1727.150000 ;
        RECT -14.680000 1724.130000 -11.680000 1724.140000 ;
        RECT 2931.300000 1724.130000 2934.300000 1724.140000 ;
        RECT -38.180000 1691.380000 -35.180000 1691.390000 ;
        RECT 2954.800000 1691.380000 2957.800000 1691.390000 ;
        RECT -38.180000 1688.370000 -35.180000 1688.380000 ;
        RECT 2954.800000 1688.370000 2957.800000 1688.380000 ;
        RECT -28.780000 1673.380000 -25.780000 1673.390000 ;
        RECT 2945.400000 1673.380000 2948.400000 1673.390000 ;
        RECT -28.780000 1670.370000 -25.780000 1670.380000 ;
        RECT 2945.400000 1670.370000 2948.400000 1670.380000 ;
        RECT -19.380000 1655.380000 -16.380000 1655.390000 ;
        RECT 2936.000000 1655.380000 2939.000000 1655.390000 ;
        RECT -19.380000 1652.370000 -16.380000 1652.380000 ;
        RECT 2936.000000 1652.370000 2939.000000 1652.380000 ;
        RECT -9.980000 1637.140000 -6.980000 1637.150000 ;
        RECT 2926.600000 1637.140000 2929.600000 1637.150000 ;
        RECT -9.980000 1634.130000 -6.980000 1634.140000 ;
        RECT 2926.600000 1634.130000 2929.600000 1634.140000 ;
        RECT -42.880000 1601.380000 -39.880000 1601.390000 ;
        RECT 2959.500000 1601.380000 2962.500000 1601.390000 ;
        RECT -42.880000 1598.370000 -39.880000 1598.380000 ;
        RECT 2959.500000 1598.370000 2962.500000 1598.380000 ;
        RECT -33.480000 1583.380000 -30.480000 1583.390000 ;
        RECT 2950.100000 1583.380000 2953.100000 1583.390000 ;
        RECT -33.480000 1580.370000 -30.480000 1580.380000 ;
        RECT 2950.100000 1580.370000 2953.100000 1580.380000 ;
        RECT -24.080000 1565.380000 -21.080000 1565.390000 ;
        RECT 2940.700000 1565.380000 2943.700000 1565.390000 ;
        RECT -24.080000 1562.370000 -21.080000 1562.380000 ;
        RECT 2940.700000 1562.370000 2943.700000 1562.380000 ;
        RECT -14.680000 1547.140000 -11.680000 1547.150000 ;
        RECT 2931.300000 1547.140000 2934.300000 1547.150000 ;
        RECT -14.680000 1544.130000 -11.680000 1544.140000 ;
        RECT 2931.300000 1544.130000 2934.300000 1544.140000 ;
        RECT -38.180000 1511.380000 -35.180000 1511.390000 ;
        RECT 2954.800000 1511.380000 2957.800000 1511.390000 ;
        RECT -38.180000 1508.370000 -35.180000 1508.380000 ;
        RECT 2954.800000 1508.370000 2957.800000 1508.380000 ;
        RECT -28.780000 1493.380000 -25.780000 1493.390000 ;
        RECT 2945.400000 1493.380000 2948.400000 1493.390000 ;
        RECT -28.780000 1490.370000 -25.780000 1490.380000 ;
        RECT 2945.400000 1490.370000 2948.400000 1490.380000 ;
        RECT -19.380000 1475.380000 -16.380000 1475.390000 ;
        RECT 2936.000000 1475.380000 2939.000000 1475.390000 ;
        RECT -19.380000 1472.370000 -16.380000 1472.380000 ;
        RECT 2936.000000 1472.370000 2939.000000 1472.380000 ;
        RECT -9.980000 1457.140000 -6.980000 1457.150000 ;
        RECT 2926.600000 1457.140000 2929.600000 1457.150000 ;
        RECT -9.980000 1454.130000 -6.980000 1454.140000 ;
        RECT 2926.600000 1454.130000 2929.600000 1454.140000 ;
        RECT -42.880000 1421.380000 -39.880000 1421.390000 ;
        RECT 2959.500000 1421.380000 2962.500000 1421.390000 ;
        RECT -42.880000 1418.370000 -39.880000 1418.380000 ;
        RECT 2959.500000 1418.370000 2962.500000 1418.380000 ;
        RECT -33.480000 1403.380000 -30.480000 1403.390000 ;
        RECT 2950.100000 1403.380000 2953.100000 1403.390000 ;
        RECT -33.480000 1400.370000 -30.480000 1400.380000 ;
        RECT 2950.100000 1400.370000 2953.100000 1400.380000 ;
        RECT -24.080000 1385.380000 -21.080000 1385.390000 ;
        RECT 2940.700000 1385.380000 2943.700000 1385.390000 ;
        RECT -24.080000 1382.370000 -21.080000 1382.380000 ;
        RECT 2940.700000 1382.370000 2943.700000 1382.380000 ;
        RECT -14.680000 1367.140000 -11.680000 1367.150000 ;
        RECT 2931.300000 1367.140000 2934.300000 1367.150000 ;
        RECT -14.680000 1364.130000 -11.680000 1364.140000 ;
        RECT 2931.300000 1364.130000 2934.300000 1364.140000 ;
        RECT -38.180000 1331.380000 -35.180000 1331.390000 ;
        RECT 2954.800000 1331.380000 2957.800000 1331.390000 ;
        RECT -38.180000 1328.370000 -35.180000 1328.380000 ;
        RECT 2954.800000 1328.370000 2957.800000 1328.380000 ;
        RECT -28.780000 1313.380000 -25.780000 1313.390000 ;
        RECT 2945.400000 1313.380000 2948.400000 1313.390000 ;
        RECT -28.780000 1310.370000 -25.780000 1310.380000 ;
        RECT 2945.400000 1310.370000 2948.400000 1310.380000 ;
        RECT -19.380000 1295.380000 -16.380000 1295.390000 ;
        RECT 2936.000000 1295.380000 2939.000000 1295.390000 ;
        RECT -19.380000 1292.370000 -16.380000 1292.380000 ;
        RECT 2936.000000 1292.370000 2939.000000 1292.380000 ;
        RECT -9.980000 1277.140000 -6.980000 1277.150000 ;
        RECT 2926.600000 1277.140000 2929.600000 1277.150000 ;
        RECT -9.980000 1274.130000 -6.980000 1274.140000 ;
        RECT 2926.600000 1274.130000 2929.600000 1274.140000 ;
        RECT -42.880000 1241.380000 -39.880000 1241.390000 ;
        RECT 2959.500000 1241.380000 2962.500000 1241.390000 ;
        RECT -42.880000 1238.370000 -39.880000 1238.380000 ;
        RECT 2959.500000 1238.370000 2962.500000 1238.380000 ;
        RECT -33.480000 1223.380000 -30.480000 1223.390000 ;
        RECT 2950.100000 1223.380000 2953.100000 1223.390000 ;
        RECT -33.480000 1220.370000 -30.480000 1220.380000 ;
        RECT 2950.100000 1220.370000 2953.100000 1220.380000 ;
        RECT -24.080000 1205.380000 -21.080000 1205.390000 ;
        RECT 2940.700000 1205.380000 2943.700000 1205.390000 ;
        RECT -24.080000 1202.370000 -21.080000 1202.380000 ;
        RECT 2940.700000 1202.370000 2943.700000 1202.380000 ;
        RECT -14.680000 1187.140000 -11.680000 1187.150000 ;
        RECT 2931.300000 1187.140000 2934.300000 1187.150000 ;
        RECT -14.680000 1184.130000 -11.680000 1184.140000 ;
        RECT 2931.300000 1184.130000 2934.300000 1184.140000 ;
        RECT -38.180000 1151.380000 -35.180000 1151.390000 ;
        RECT 2954.800000 1151.380000 2957.800000 1151.390000 ;
        RECT -38.180000 1148.370000 -35.180000 1148.380000 ;
        RECT 2954.800000 1148.370000 2957.800000 1148.380000 ;
        RECT -28.780000 1133.380000 -25.780000 1133.390000 ;
        RECT 2945.400000 1133.380000 2948.400000 1133.390000 ;
        RECT -28.780000 1130.370000 -25.780000 1130.380000 ;
        RECT 2945.400000 1130.370000 2948.400000 1130.380000 ;
        RECT -19.380000 1115.380000 -16.380000 1115.390000 ;
        RECT 2936.000000 1115.380000 2939.000000 1115.390000 ;
        RECT -19.380000 1112.370000 -16.380000 1112.380000 ;
        RECT 2936.000000 1112.370000 2939.000000 1112.380000 ;
        RECT -9.980000 1097.140000 -6.980000 1097.150000 ;
        RECT 2926.600000 1097.140000 2929.600000 1097.150000 ;
        RECT -9.980000 1094.130000 -6.980000 1094.140000 ;
        RECT 2926.600000 1094.130000 2929.600000 1094.140000 ;
        RECT -42.880000 1061.380000 -39.880000 1061.390000 ;
        RECT 2959.500000 1061.380000 2962.500000 1061.390000 ;
        RECT -42.880000 1058.370000 -39.880000 1058.380000 ;
        RECT 2959.500000 1058.370000 2962.500000 1058.380000 ;
        RECT -33.480000 1043.380000 -30.480000 1043.390000 ;
        RECT 2950.100000 1043.380000 2953.100000 1043.390000 ;
        RECT -33.480000 1040.370000 -30.480000 1040.380000 ;
        RECT 2950.100000 1040.370000 2953.100000 1040.380000 ;
        RECT -24.080000 1025.380000 -21.080000 1025.390000 ;
        RECT 2940.700000 1025.380000 2943.700000 1025.390000 ;
        RECT -24.080000 1022.370000 -21.080000 1022.380000 ;
        RECT 2940.700000 1022.370000 2943.700000 1022.380000 ;
        RECT -14.680000 1007.140000 -11.680000 1007.150000 ;
        RECT 2931.300000 1007.140000 2934.300000 1007.150000 ;
        RECT -14.680000 1004.130000 -11.680000 1004.140000 ;
        RECT 2931.300000 1004.130000 2934.300000 1004.140000 ;
        RECT -38.180000 971.380000 -35.180000 971.390000 ;
        RECT 2954.800000 971.380000 2957.800000 971.390000 ;
        RECT -38.180000 968.370000 -35.180000 968.380000 ;
        RECT 2954.800000 968.370000 2957.800000 968.380000 ;
        RECT -28.780000 953.380000 -25.780000 953.390000 ;
        RECT 2945.400000 953.380000 2948.400000 953.390000 ;
        RECT -28.780000 950.370000 -25.780000 950.380000 ;
        RECT 2945.400000 950.370000 2948.400000 950.380000 ;
        RECT -19.380000 935.380000 -16.380000 935.390000 ;
        RECT 2936.000000 935.380000 2939.000000 935.390000 ;
        RECT -19.380000 932.370000 -16.380000 932.380000 ;
        RECT 2936.000000 932.370000 2939.000000 932.380000 ;
        RECT -9.980000 917.140000 -6.980000 917.150000 ;
        RECT 2926.600000 917.140000 2929.600000 917.150000 ;
        RECT -9.980000 914.130000 -6.980000 914.140000 ;
        RECT 2926.600000 914.130000 2929.600000 914.140000 ;
        RECT -42.880000 881.380000 -39.880000 881.390000 ;
        RECT 2959.500000 881.380000 2962.500000 881.390000 ;
        RECT -42.880000 878.370000 -39.880000 878.380000 ;
        RECT 2959.500000 878.370000 2962.500000 878.380000 ;
        RECT -33.480000 863.380000 -30.480000 863.390000 ;
        RECT 2950.100000 863.380000 2953.100000 863.390000 ;
        RECT -33.480000 860.370000 -30.480000 860.380000 ;
        RECT 2950.100000 860.370000 2953.100000 860.380000 ;
        RECT -24.080000 845.380000 -21.080000 845.390000 ;
        RECT 2940.700000 845.380000 2943.700000 845.390000 ;
        RECT -24.080000 842.370000 -21.080000 842.380000 ;
        RECT 2940.700000 842.370000 2943.700000 842.380000 ;
        RECT -14.680000 827.140000 -11.680000 827.150000 ;
        RECT 2931.300000 827.140000 2934.300000 827.150000 ;
        RECT -14.680000 824.130000 -11.680000 824.140000 ;
        RECT 2931.300000 824.130000 2934.300000 824.140000 ;
        RECT -38.180000 791.380000 -35.180000 791.390000 ;
        RECT 2954.800000 791.380000 2957.800000 791.390000 ;
        RECT -38.180000 788.370000 -35.180000 788.380000 ;
        RECT 2954.800000 788.370000 2957.800000 788.380000 ;
        RECT -28.780000 773.380000 -25.780000 773.390000 ;
        RECT 2945.400000 773.380000 2948.400000 773.390000 ;
        RECT -28.780000 770.370000 -25.780000 770.380000 ;
        RECT 2945.400000 770.370000 2948.400000 770.380000 ;
        RECT -19.380000 755.380000 -16.380000 755.390000 ;
        RECT 2936.000000 755.380000 2939.000000 755.390000 ;
        RECT -19.380000 752.370000 -16.380000 752.380000 ;
        RECT 2936.000000 752.370000 2939.000000 752.380000 ;
        RECT -9.980000 737.140000 -6.980000 737.150000 ;
        RECT 2926.600000 737.140000 2929.600000 737.150000 ;
        RECT -9.980000 734.130000 -6.980000 734.140000 ;
        RECT 2926.600000 734.130000 2929.600000 734.140000 ;
        RECT -42.880000 701.380000 -39.880000 701.390000 ;
        RECT 2959.500000 701.380000 2962.500000 701.390000 ;
        RECT -42.880000 698.370000 -39.880000 698.380000 ;
        RECT 2959.500000 698.370000 2962.500000 698.380000 ;
        RECT -33.480000 683.380000 -30.480000 683.390000 ;
        RECT 2950.100000 683.380000 2953.100000 683.390000 ;
        RECT -33.480000 680.370000 -30.480000 680.380000 ;
        RECT 2950.100000 680.370000 2953.100000 680.380000 ;
        RECT -24.080000 665.380000 -21.080000 665.390000 ;
        RECT 2940.700000 665.380000 2943.700000 665.390000 ;
        RECT -24.080000 662.370000 -21.080000 662.380000 ;
        RECT 2940.700000 662.370000 2943.700000 662.380000 ;
        RECT -14.680000 647.140000 -11.680000 647.150000 ;
        RECT 2931.300000 647.140000 2934.300000 647.150000 ;
        RECT -14.680000 644.130000 -11.680000 644.140000 ;
        RECT 2931.300000 644.130000 2934.300000 644.140000 ;
        RECT -38.180000 611.380000 -35.180000 611.390000 ;
        RECT 2954.800000 611.380000 2957.800000 611.390000 ;
        RECT -38.180000 608.370000 -35.180000 608.380000 ;
        RECT 2954.800000 608.370000 2957.800000 608.380000 ;
        RECT -28.780000 593.380000 -25.780000 593.390000 ;
        RECT 2945.400000 593.380000 2948.400000 593.390000 ;
        RECT -28.780000 590.370000 -25.780000 590.380000 ;
        RECT 2945.400000 590.370000 2948.400000 590.380000 ;
        RECT -19.380000 575.380000 -16.380000 575.390000 ;
        RECT 2936.000000 575.380000 2939.000000 575.390000 ;
        RECT -19.380000 572.370000 -16.380000 572.380000 ;
        RECT 2936.000000 572.370000 2939.000000 572.380000 ;
        RECT -9.980000 557.140000 -6.980000 557.150000 ;
        RECT 2926.600000 557.140000 2929.600000 557.150000 ;
        RECT -9.980000 554.130000 -6.980000 554.140000 ;
        RECT 2926.600000 554.130000 2929.600000 554.140000 ;
        RECT -42.880000 521.380000 -39.880000 521.390000 ;
        RECT 2959.500000 521.380000 2962.500000 521.390000 ;
        RECT -42.880000 518.370000 -39.880000 518.380000 ;
        RECT 2959.500000 518.370000 2962.500000 518.380000 ;
        RECT -33.480000 503.380000 -30.480000 503.390000 ;
        RECT 2950.100000 503.380000 2953.100000 503.390000 ;
        RECT -33.480000 500.370000 -30.480000 500.380000 ;
        RECT 2950.100000 500.370000 2953.100000 500.380000 ;
        RECT -24.080000 485.380000 -21.080000 485.390000 ;
        RECT 2940.700000 485.380000 2943.700000 485.390000 ;
        RECT -24.080000 482.370000 -21.080000 482.380000 ;
        RECT 2940.700000 482.370000 2943.700000 482.380000 ;
        RECT -14.680000 467.140000 -11.680000 467.150000 ;
        RECT 2931.300000 467.140000 2934.300000 467.150000 ;
        RECT -14.680000 464.130000 -11.680000 464.140000 ;
        RECT 2931.300000 464.130000 2934.300000 464.140000 ;
        RECT -38.180000 431.380000 -35.180000 431.390000 ;
        RECT 2954.800000 431.380000 2957.800000 431.390000 ;
        RECT -38.180000 428.370000 -35.180000 428.380000 ;
        RECT 2954.800000 428.370000 2957.800000 428.380000 ;
        RECT -28.780000 413.380000 -25.780000 413.390000 ;
        RECT 2945.400000 413.380000 2948.400000 413.390000 ;
        RECT -28.780000 410.370000 -25.780000 410.380000 ;
        RECT 2945.400000 410.370000 2948.400000 410.380000 ;
        RECT -19.380000 395.380000 -16.380000 395.390000 ;
        RECT 2936.000000 395.380000 2939.000000 395.390000 ;
        RECT -19.380000 392.370000 -16.380000 392.380000 ;
        RECT 2936.000000 392.370000 2939.000000 392.380000 ;
        RECT -9.980000 377.140000 -6.980000 377.150000 ;
        RECT 2926.600000 377.140000 2929.600000 377.150000 ;
        RECT -9.980000 374.130000 -6.980000 374.140000 ;
        RECT 2926.600000 374.130000 2929.600000 374.140000 ;
        RECT -42.880000 341.380000 -39.880000 341.390000 ;
        RECT 2959.500000 341.380000 2962.500000 341.390000 ;
        RECT -42.880000 338.370000 -39.880000 338.380000 ;
        RECT 2959.500000 338.370000 2962.500000 338.380000 ;
        RECT -33.480000 323.380000 -30.480000 323.390000 ;
        RECT 2950.100000 323.380000 2953.100000 323.390000 ;
        RECT -33.480000 320.370000 -30.480000 320.380000 ;
        RECT 2950.100000 320.370000 2953.100000 320.380000 ;
        RECT -24.080000 305.380000 -21.080000 305.390000 ;
        RECT 2940.700000 305.380000 2943.700000 305.390000 ;
        RECT -24.080000 302.370000 -21.080000 302.380000 ;
        RECT 2940.700000 302.370000 2943.700000 302.380000 ;
        RECT -14.680000 287.140000 -11.680000 287.150000 ;
        RECT 2931.300000 287.140000 2934.300000 287.150000 ;
        RECT -14.680000 284.130000 -11.680000 284.140000 ;
        RECT 2931.300000 284.130000 2934.300000 284.140000 ;
        RECT -38.180000 251.380000 -35.180000 251.390000 ;
        RECT 2954.800000 251.380000 2957.800000 251.390000 ;
        RECT -38.180000 248.370000 -35.180000 248.380000 ;
        RECT 2954.800000 248.370000 2957.800000 248.380000 ;
        RECT -28.780000 233.380000 -25.780000 233.390000 ;
        RECT 2945.400000 233.380000 2948.400000 233.390000 ;
        RECT -28.780000 230.370000 -25.780000 230.380000 ;
        RECT 2945.400000 230.370000 2948.400000 230.380000 ;
        RECT -19.380000 215.380000 -16.380000 215.390000 ;
        RECT 2936.000000 215.380000 2939.000000 215.390000 ;
        RECT -19.380000 212.370000 -16.380000 212.380000 ;
        RECT 2936.000000 212.370000 2939.000000 212.380000 ;
        RECT -9.980000 197.140000 -6.980000 197.150000 ;
        RECT 2926.600000 197.140000 2929.600000 197.150000 ;
        RECT -9.980000 194.130000 -6.980000 194.140000 ;
        RECT 2926.600000 194.130000 2929.600000 194.140000 ;
        RECT -42.880000 161.380000 -39.880000 161.390000 ;
        RECT 2959.500000 161.380000 2962.500000 161.390000 ;
        RECT -42.880000 158.370000 -39.880000 158.380000 ;
        RECT 2959.500000 158.370000 2962.500000 158.380000 ;
        RECT -33.480000 143.380000 -30.480000 143.390000 ;
        RECT 2950.100000 143.380000 2953.100000 143.390000 ;
        RECT -33.480000 140.370000 -30.480000 140.380000 ;
        RECT 2950.100000 140.370000 2953.100000 140.380000 ;
        RECT -24.080000 125.380000 -21.080000 125.390000 ;
        RECT 2940.700000 125.380000 2943.700000 125.390000 ;
        RECT -24.080000 122.370000 -21.080000 122.380000 ;
        RECT 2940.700000 122.370000 2943.700000 122.380000 ;
        RECT -14.680000 107.140000 -11.680000 107.150000 ;
        RECT 2931.300000 107.140000 2934.300000 107.150000 ;
        RECT -14.680000 104.130000 -11.680000 104.140000 ;
        RECT 2931.300000 104.130000 2934.300000 104.140000 ;
        RECT -38.180000 71.380000 -35.180000 71.390000 ;
        RECT 2954.800000 71.380000 2957.800000 71.390000 ;
        RECT -38.180000 68.370000 -35.180000 68.380000 ;
        RECT 2954.800000 68.370000 2957.800000 68.380000 ;
        RECT -28.780000 53.380000 -25.780000 53.390000 ;
        RECT 2945.400000 53.380000 2948.400000 53.390000 ;
        RECT -28.780000 50.370000 -25.780000 50.380000 ;
        RECT 2945.400000 50.370000 2948.400000 50.380000 ;
        RECT -19.380000 35.380000 -16.380000 35.390000 ;
        RECT 2936.000000 35.380000 2939.000000 35.390000 ;
        RECT -19.380000 32.370000 -16.380000 32.380000 ;
        RECT 2936.000000 32.370000 2939.000000 32.380000 ;
        RECT -9.980000 17.140000 -6.980000 17.150000 ;
        RECT 2926.600000 17.140000 2929.600000 17.150000 ;
        RECT -9.980000 14.130000 -6.980000 14.140000 ;
        RECT 2926.600000 14.130000 2929.600000 14.140000 ;
        RECT -9.980000 -1.620000 -6.980000 -1.610000 ;
        RECT 9.020000 -1.620000 12.020000 -1.610000 ;
        RECT 189.020000 -1.620000 192.020000 -1.610000 ;
        RECT 369.020000 -1.620000 372.020000 -1.610000 ;
        RECT 549.020000 -1.620000 552.020000 -1.610000 ;
        RECT 729.020000 -1.620000 732.020000 -1.610000 ;
        RECT 909.020000 -1.620000 912.020000 -1.610000 ;
        RECT 1089.020000 -1.620000 1092.020000 -1.610000 ;
        RECT 1269.020000 -1.620000 1272.020000 -1.610000 ;
        RECT 1449.020000 -1.620000 1452.020000 -1.610000 ;
        RECT 1629.020000 -1.620000 1632.020000 -1.610000 ;
        RECT 1809.020000 -1.620000 1812.020000 -1.610000 ;
        RECT 1989.020000 -1.620000 1992.020000 -1.610000 ;
        RECT 2169.020000 -1.620000 2172.020000 -1.610000 ;
        RECT 2349.020000 -1.620000 2352.020000 -1.610000 ;
        RECT 2529.020000 -1.620000 2532.020000 -1.610000 ;
        RECT 2709.020000 -1.620000 2712.020000 -1.610000 ;
        RECT 2889.020000 -1.620000 2892.020000 -1.610000 ;
        RECT 2926.600000 -1.620000 2929.600000 -1.610000 ;
        RECT -9.980000 -4.630000 -6.980000 -4.620000 ;
        RECT 9.020000 -4.630000 12.020000 -4.620000 ;
        RECT 189.020000 -4.630000 192.020000 -4.620000 ;
        RECT 369.020000 -4.630000 372.020000 -4.620000 ;
        RECT 549.020000 -4.630000 552.020000 -4.620000 ;
        RECT 729.020000 -4.630000 732.020000 -4.620000 ;
        RECT 909.020000 -4.630000 912.020000 -4.620000 ;
        RECT 1089.020000 -4.630000 1092.020000 -4.620000 ;
        RECT 1269.020000 -4.630000 1272.020000 -4.620000 ;
        RECT 1449.020000 -4.630000 1452.020000 -4.620000 ;
        RECT 1629.020000 -4.630000 1632.020000 -4.620000 ;
        RECT 1809.020000 -4.630000 1812.020000 -4.620000 ;
        RECT 1989.020000 -4.630000 1992.020000 -4.620000 ;
        RECT 2169.020000 -4.630000 2172.020000 -4.620000 ;
        RECT 2349.020000 -4.630000 2352.020000 -4.620000 ;
        RECT 2529.020000 -4.630000 2532.020000 -4.620000 ;
        RECT 2709.020000 -4.630000 2712.020000 -4.620000 ;
        RECT 2889.020000 -4.630000 2892.020000 -4.620000 ;
        RECT 2926.600000 -4.630000 2929.600000 -4.620000 ;
        RECT -14.680000 -6.320000 -11.680000 -6.310000 ;
        RECT 99.020000 -6.320000 102.020000 -6.310000 ;
        RECT 279.020000 -6.320000 282.020000 -6.310000 ;
        RECT 459.020000 -6.320000 462.020000 -6.310000 ;
        RECT 639.020000 -6.320000 642.020000 -6.310000 ;
        RECT 819.020000 -6.320000 822.020000 -6.310000 ;
        RECT 999.020000 -6.320000 1002.020000 -6.310000 ;
        RECT 1179.020000 -6.320000 1182.020000 -6.310000 ;
        RECT 1359.020000 -6.320000 1362.020000 -6.310000 ;
        RECT 1539.020000 -6.320000 1542.020000 -6.310000 ;
        RECT 1719.020000 -6.320000 1722.020000 -6.310000 ;
        RECT 1899.020000 -6.320000 1902.020000 -6.310000 ;
        RECT 2079.020000 -6.320000 2082.020000 -6.310000 ;
        RECT 2259.020000 -6.320000 2262.020000 -6.310000 ;
        RECT 2439.020000 -6.320000 2442.020000 -6.310000 ;
        RECT 2619.020000 -6.320000 2622.020000 -6.310000 ;
        RECT 2799.020000 -6.320000 2802.020000 -6.310000 ;
        RECT 2931.300000 -6.320000 2934.300000 -6.310000 ;
        RECT -14.680000 -9.330000 -11.680000 -9.320000 ;
        RECT 99.020000 -9.330000 102.020000 -9.320000 ;
        RECT 279.020000 -9.330000 282.020000 -9.320000 ;
        RECT 459.020000 -9.330000 462.020000 -9.320000 ;
        RECT 639.020000 -9.330000 642.020000 -9.320000 ;
        RECT 819.020000 -9.330000 822.020000 -9.320000 ;
        RECT 999.020000 -9.330000 1002.020000 -9.320000 ;
        RECT 1179.020000 -9.330000 1182.020000 -9.320000 ;
        RECT 1359.020000 -9.330000 1362.020000 -9.320000 ;
        RECT 1539.020000 -9.330000 1542.020000 -9.320000 ;
        RECT 1719.020000 -9.330000 1722.020000 -9.320000 ;
        RECT 1899.020000 -9.330000 1902.020000 -9.320000 ;
        RECT 2079.020000 -9.330000 2082.020000 -9.320000 ;
        RECT 2259.020000 -9.330000 2262.020000 -9.320000 ;
        RECT 2439.020000 -9.330000 2442.020000 -9.320000 ;
        RECT 2619.020000 -9.330000 2622.020000 -9.320000 ;
        RECT 2799.020000 -9.330000 2802.020000 -9.320000 ;
        RECT 2931.300000 -9.330000 2934.300000 -9.320000 ;
        RECT -19.380000 -11.020000 -16.380000 -11.010000 ;
        RECT 27.020000 -11.020000 30.020000 -11.010000 ;
        RECT 207.020000 -11.020000 210.020000 -11.010000 ;
        RECT 387.020000 -11.020000 390.020000 -11.010000 ;
        RECT 567.020000 -11.020000 570.020000 -11.010000 ;
        RECT 747.020000 -11.020000 750.020000 -11.010000 ;
        RECT 927.020000 -11.020000 930.020000 -11.010000 ;
        RECT 1107.020000 -11.020000 1110.020000 -11.010000 ;
        RECT 1287.020000 -11.020000 1290.020000 -11.010000 ;
        RECT 1467.020000 -11.020000 1470.020000 -11.010000 ;
        RECT 1647.020000 -11.020000 1650.020000 -11.010000 ;
        RECT 1827.020000 -11.020000 1830.020000 -11.010000 ;
        RECT 2007.020000 -11.020000 2010.020000 -11.010000 ;
        RECT 2187.020000 -11.020000 2190.020000 -11.010000 ;
        RECT 2367.020000 -11.020000 2370.020000 -11.010000 ;
        RECT 2547.020000 -11.020000 2550.020000 -11.010000 ;
        RECT 2727.020000 -11.020000 2730.020000 -11.010000 ;
        RECT 2907.020000 -11.020000 2910.020000 -11.010000 ;
        RECT 2936.000000 -11.020000 2939.000000 -11.010000 ;
        RECT -19.380000 -14.030000 -16.380000 -14.020000 ;
        RECT 27.020000 -14.030000 30.020000 -14.020000 ;
        RECT 207.020000 -14.030000 210.020000 -14.020000 ;
        RECT 387.020000 -14.030000 390.020000 -14.020000 ;
        RECT 567.020000 -14.030000 570.020000 -14.020000 ;
        RECT 747.020000 -14.030000 750.020000 -14.020000 ;
        RECT 927.020000 -14.030000 930.020000 -14.020000 ;
        RECT 1107.020000 -14.030000 1110.020000 -14.020000 ;
        RECT 1287.020000 -14.030000 1290.020000 -14.020000 ;
        RECT 1467.020000 -14.030000 1470.020000 -14.020000 ;
        RECT 1647.020000 -14.030000 1650.020000 -14.020000 ;
        RECT 1827.020000 -14.030000 1830.020000 -14.020000 ;
        RECT 2007.020000 -14.030000 2010.020000 -14.020000 ;
        RECT 2187.020000 -14.030000 2190.020000 -14.020000 ;
        RECT 2367.020000 -14.030000 2370.020000 -14.020000 ;
        RECT 2547.020000 -14.030000 2550.020000 -14.020000 ;
        RECT 2727.020000 -14.030000 2730.020000 -14.020000 ;
        RECT 2907.020000 -14.030000 2910.020000 -14.020000 ;
        RECT 2936.000000 -14.030000 2939.000000 -14.020000 ;
        RECT -24.080000 -15.720000 -21.080000 -15.710000 ;
        RECT 117.020000 -15.720000 120.020000 -15.710000 ;
        RECT 297.020000 -15.720000 300.020000 -15.710000 ;
        RECT 477.020000 -15.720000 480.020000 -15.710000 ;
        RECT 657.020000 -15.720000 660.020000 -15.710000 ;
        RECT 837.020000 -15.720000 840.020000 -15.710000 ;
        RECT 1017.020000 -15.720000 1020.020000 -15.710000 ;
        RECT 1197.020000 -15.720000 1200.020000 -15.710000 ;
        RECT 1377.020000 -15.720000 1380.020000 -15.710000 ;
        RECT 1557.020000 -15.720000 1560.020000 -15.710000 ;
        RECT 1737.020000 -15.720000 1740.020000 -15.710000 ;
        RECT 1917.020000 -15.720000 1920.020000 -15.710000 ;
        RECT 2097.020000 -15.720000 2100.020000 -15.710000 ;
        RECT 2277.020000 -15.720000 2280.020000 -15.710000 ;
        RECT 2457.020000 -15.720000 2460.020000 -15.710000 ;
        RECT 2637.020000 -15.720000 2640.020000 -15.710000 ;
        RECT 2817.020000 -15.720000 2820.020000 -15.710000 ;
        RECT 2940.700000 -15.720000 2943.700000 -15.710000 ;
        RECT -24.080000 -18.730000 -21.080000 -18.720000 ;
        RECT 117.020000 -18.730000 120.020000 -18.720000 ;
        RECT 297.020000 -18.730000 300.020000 -18.720000 ;
        RECT 477.020000 -18.730000 480.020000 -18.720000 ;
        RECT 657.020000 -18.730000 660.020000 -18.720000 ;
        RECT 837.020000 -18.730000 840.020000 -18.720000 ;
        RECT 1017.020000 -18.730000 1020.020000 -18.720000 ;
        RECT 1197.020000 -18.730000 1200.020000 -18.720000 ;
        RECT 1377.020000 -18.730000 1380.020000 -18.720000 ;
        RECT 1557.020000 -18.730000 1560.020000 -18.720000 ;
        RECT 1737.020000 -18.730000 1740.020000 -18.720000 ;
        RECT 1917.020000 -18.730000 1920.020000 -18.720000 ;
        RECT 2097.020000 -18.730000 2100.020000 -18.720000 ;
        RECT 2277.020000 -18.730000 2280.020000 -18.720000 ;
        RECT 2457.020000 -18.730000 2460.020000 -18.720000 ;
        RECT 2637.020000 -18.730000 2640.020000 -18.720000 ;
        RECT 2817.020000 -18.730000 2820.020000 -18.720000 ;
        RECT 2940.700000 -18.730000 2943.700000 -18.720000 ;
        RECT -28.780000 -20.420000 -25.780000 -20.410000 ;
        RECT 45.020000 -20.420000 48.020000 -20.410000 ;
        RECT 225.020000 -20.420000 228.020000 -20.410000 ;
        RECT 405.020000 -20.420000 408.020000 -20.410000 ;
        RECT 585.020000 -20.420000 588.020000 -20.410000 ;
        RECT 765.020000 -20.420000 768.020000 -20.410000 ;
        RECT 945.020000 -20.420000 948.020000 -20.410000 ;
        RECT 1125.020000 -20.420000 1128.020000 -20.410000 ;
        RECT 1305.020000 -20.420000 1308.020000 -20.410000 ;
        RECT 1485.020000 -20.420000 1488.020000 -20.410000 ;
        RECT 1665.020000 -20.420000 1668.020000 -20.410000 ;
        RECT 1845.020000 -20.420000 1848.020000 -20.410000 ;
        RECT 2025.020000 -20.420000 2028.020000 -20.410000 ;
        RECT 2205.020000 -20.420000 2208.020000 -20.410000 ;
        RECT 2385.020000 -20.420000 2388.020000 -20.410000 ;
        RECT 2565.020000 -20.420000 2568.020000 -20.410000 ;
        RECT 2745.020000 -20.420000 2748.020000 -20.410000 ;
        RECT 2945.400000 -20.420000 2948.400000 -20.410000 ;
        RECT -28.780000 -23.430000 -25.780000 -23.420000 ;
        RECT 45.020000 -23.430000 48.020000 -23.420000 ;
        RECT 225.020000 -23.430000 228.020000 -23.420000 ;
        RECT 405.020000 -23.430000 408.020000 -23.420000 ;
        RECT 585.020000 -23.430000 588.020000 -23.420000 ;
        RECT 765.020000 -23.430000 768.020000 -23.420000 ;
        RECT 945.020000 -23.430000 948.020000 -23.420000 ;
        RECT 1125.020000 -23.430000 1128.020000 -23.420000 ;
        RECT 1305.020000 -23.430000 1308.020000 -23.420000 ;
        RECT 1485.020000 -23.430000 1488.020000 -23.420000 ;
        RECT 1665.020000 -23.430000 1668.020000 -23.420000 ;
        RECT 1845.020000 -23.430000 1848.020000 -23.420000 ;
        RECT 2025.020000 -23.430000 2028.020000 -23.420000 ;
        RECT 2205.020000 -23.430000 2208.020000 -23.420000 ;
        RECT 2385.020000 -23.430000 2388.020000 -23.420000 ;
        RECT 2565.020000 -23.430000 2568.020000 -23.420000 ;
        RECT 2745.020000 -23.430000 2748.020000 -23.420000 ;
        RECT 2945.400000 -23.430000 2948.400000 -23.420000 ;
        RECT -33.480000 -25.120000 -30.480000 -25.110000 ;
        RECT 135.020000 -25.120000 138.020000 -25.110000 ;
        RECT 315.020000 -25.120000 318.020000 -25.110000 ;
        RECT 495.020000 -25.120000 498.020000 -25.110000 ;
        RECT 675.020000 -25.120000 678.020000 -25.110000 ;
        RECT 855.020000 -25.120000 858.020000 -25.110000 ;
        RECT 1035.020000 -25.120000 1038.020000 -25.110000 ;
        RECT 1215.020000 -25.120000 1218.020000 -25.110000 ;
        RECT 1395.020000 -25.120000 1398.020000 -25.110000 ;
        RECT 1575.020000 -25.120000 1578.020000 -25.110000 ;
        RECT 1755.020000 -25.120000 1758.020000 -25.110000 ;
        RECT 1935.020000 -25.120000 1938.020000 -25.110000 ;
        RECT 2115.020000 -25.120000 2118.020000 -25.110000 ;
        RECT 2295.020000 -25.120000 2298.020000 -25.110000 ;
        RECT 2475.020000 -25.120000 2478.020000 -25.110000 ;
        RECT 2655.020000 -25.120000 2658.020000 -25.110000 ;
        RECT 2835.020000 -25.120000 2838.020000 -25.110000 ;
        RECT 2950.100000 -25.120000 2953.100000 -25.110000 ;
        RECT -33.480000 -28.130000 -30.480000 -28.120000 ;
        RECT 135.020000 -28.130000 138.020000 -28.120000 ;
        RECT 315.020000 -28.130000 318.020000 -28.120000 ;
        RECT 495.020000 -28.130000 498.020000 -28.120000 ;
        RECT 675.020000 -28.130000 678.020000 -28.120000 ;
        RECT 855.020000 -28.130000 858.020000 -28.120000 ;
        RECT 1035.020000 -28.130000 1038.020000 -28.120000 ;
        RECT 1215.020000 -28.130000 1218.020000 -28.120000 ;
        RECT 1395.020000 -28.130000 1398.020000 -28.120000 ;
        RECT 1575.020000 -28.130000 1578.020000 -28.120000 ;
        RECT 1755.020000 -28.130000 1758.020000 -28.120000 ;
        RECT 1935.020000 -28.130000 1938.020000 -28.120000 ;
        RECT 2115.020000 -28.130000 2118.020000 -28.120000 ;
        RECT 2295.020000 -28.130000 2298.020000 -28.120000 ;
        RECT 2475.020000 -28.130000 2478.020000 -28.120000 ;
        RECT 2655.020000 -28.130000 2658.020000 -28.120000 ;
        RECT 2835.020000 -28.130000 2838.020000 -28.120000 ;
        RECT 2950.100000 -28.130000 2953.100000 -28.120000 ;
        RECT -38.180000 -29.820000 -35.180000 -29.810000 ;
        RECT 63.020000 -29.820000 66.020000 -29.810000 ;
        RECT 243.020000 -29.820000 246.020000 -29.810000 ;
        RECT 423.020000 -29.820000 426.020000 -29.810000 ;
        RECT 603.020000 -29.820000 606.020000 -29.810000 ;
        RECT 783.020000 -29.820000 786.020000 -29.810000 ;
        RECT 963.020000 -29.820000 966.020000 -29.810000 ;
        RECT 1143.020000 -29.820000 1146.020000 -29.810000 ;
        RECT 1323.020000 -29.820000 1326.020000 -29.810000 ;
        RECT 1503.020000 -29.820000 1506.020000 -29.810000 ;
        RECT 1683.020000 -29.820000 1686.020000 -29.810000 ;
        RECT 1863.020000 -29.820000 1866.020000 -29.810000 ;
        RECT 2043.020000 -29.820000 2046.020000 -29.810000 ;
        RECT 2223.020000 -29.820000 2226.020000 -29.810000 ;
        RECT 2403.020000 -29.820000 2406.020000 -29.810000 ;
        RECT 2583.020000 -29.820000 2586.020000 -29.810000 ;
        RECT 2763.020000 -29.820000 2766.020000 -29.810000 ;
        RECT 2954.800000 -29.820000 2957.800000 -29.810000 ;
        RECT -38.180000 -32.830000 -35.180000 -32.820000 ;
        RECT 63.020000 -32.830000 66.020000 -32.820000 ;
        RECT 243.020000 -32.830000 246.020000 -32.820000 ;
        RECT 423.020000 -32.830000 426.020000 -32.820000 ;
        RECT 603.020000 -32.830000 606.020000 -32.820000 ;
        RECT 783.020000 -32.830000 786.020000 -32.820000 ;
        RECT 963.020000 -32.830000 966.020000 -32.820000 ;
        RECT 1143.020000 -32.830000 1146.020000 -32.820000 ;
        RECT 1323.020000 -32.830000 1326.020000 -32.820000 ;
        RECT 1503.020000 -32.830000 1506.020000 -32.820000 ;
        RECT 1683.020000 -32.830000 1686.020000 -32.820000 ;
        RECT 1863.020000 -32.830000 1866.020000 -32.820000 ;
        RECT 2043.020000 -32.830000 2046.020000 -32.820000 ;
        RECT 2223.020000 -32.830000 2226.020000 -32.820000 ;
        RECT 2403.020000 -32.830000 2406.020000 -32.820000 ;
        RECT 2583.020000 -32.830000 2586.020000 -32.820000 ;
        RECT 2763.020000 -32.830000 2766.020000 -32.820000 ;
        RECT 2954.800000 -32.830000 2957.800000 -32.820000 ;
        RECT -42.880000 -34.520000 -39.880000 -34.510000 ;
        RECT 153.020000 -34.520000 156.020000 -34.510000 ;
        RECT 333.020000 -34.520000 336.020000 -34.510000 ;
        RECT 513.020000 -34.520000 516.020000 -34.510000 ;
        RECT 693.020000 -34.520000 696.020000 -34.510000 ;
        RECT 873.020000 -34.520000 876.020000 -34.510000 ;
        RECT 1053.020000 -34.520000 1056.020000 -34.510000 ;
        RECT 1233.020000 -34.520000 1236.020000 -34.510000 ;
        RECT 1413.020000 -34.520000 1416.020000 -34.510000 ;
        RECT 1593.020000 -34.520000 1596.020000 -34.510000 ;
        RECT 1773.020000 -34.520000 1776.020000 -34.510000 ;
        RECT 1953.020000 -34.520000 1956.020000 -34.510000 ;
        RECT 2133.020000 -34.520000 2136.020000 -34.510000 ;
        RECT 2313.020000 -34.520000 2316.020000 -34.510000 ;
        RECT 2493.020000 -34.520000 2496.020000 -34.510000 ;
        RECT 2673.020000 -34.520000 2676.020000 -34.510000 ;
        RECT 2853.020000 -34.520000 2856.020000 -34.510000 ;
        RECT 2959.500000 -34.520000 2962.500000 -34.510000 ;
        RECT -42.880000 -37.530000 -39.880000 -37.520000 ;
        RECT 153.020000 -37.530000 156.020000 -37.520000 ;
        RECT 333.020000 -37.530000 336.020000 -37.520000 ;
        RECT 513.020000 -37.530000 516.020000 -37.520000 ;
        RECT 693.020000 -37.530000 696.020000 -37.520000 ;
        RECT 873.020000 -37.530000 876.020000 -37.520000 ;
        RECT 1053.020000 -37.530000 1056.020000 -37.520000 ;
        RECT 1233.020000 -37.530000 1236.020000 -37.520000 ;
        RECT 1413.020000 -37.530000 1416.020000 -37.520000 ;
        RECT 1593.020000 -37.530000 1596.020000 -37.520000 ;
        RECT 1773.020000 -37.530000 1776.020000 -37.520000 ;
        RECT 1953.020000 -37.530000 1956.020000 -37.520000 ;
        RECT 2133.020000 -37.530000 2136.020000 -37.520000 ;
        RECT 2313.020000 -37.530000 2316.020000 -37.520000 ;
        RECT 2493.020000 -37.530000 2496.020000 -37.520000 ;
        RECT 2673.020000 -37.530000 2676.020000 -37.520000 ;
        RECT 2853.020000 -37.530000 2856.020000 -37.520000 ;
        RECT 2959.500000 -37.530000 2962.500000 -37.520000 ;
     LAYER met4 ;
       RECT 0.000 0.000 2920.000 3520.000 ;
       RECT -42.880 -37.530 2962.500 3557.210 ;
     LAYER li1 ;
       RECT 0.000 0.000 2920.000 3520.000 ;
     LAYER met1 ;
       RECT 0.000 0.000 2920.000 3520.000 ;
     LAYER met2 ;
       RECT 0.000 0.000 2920.000 3520.000 ;
     LAYER met3 ;
       RECT 0.000 0.000 2920.000 3520.000 ;
  END
END user_project_wrapper
END LIBRARY
