magic
tech sky130A
magscale 1 2
timestamp 1625092191
<< nwell >>
rect 232772 997737 244593 998041
rect 284372 997737 296193 998041
rect 335772 997737 347593 998041
rect 577972 997737 589793 998041
rect 677737 953407 678041 965228
rect 39559 872172 39863 883993
rect 678733 877778 679465 878483
rect 688918 878257 693847 878543
rect 695297 878424 696080 878483
rect 681431 865434 682216 877484
rect 688918 873697 689204 878257
rect 689636 877638 690068 878257
rect 689636 876308 689804 877638
rect 689754 875693 689804 876308
rect 693561 873437 693847 878257
rect 694716 877841 696080 878424
rect 694716 877494 695964 877841
rect 694932 877205 695964 877494
rect 694932 876716 695256 877205
rect 694932 876701 695148 876716
rect 684453 866745 684811 868617
rect 684082 865434 684811 866745
rect 681431 862310 682669 865434
rect 683557 862310 684811 865434
rect 692119 865870 692253 869012
rect 687724 862575 688010 864333
rect 690639 862575 690809 864333
rect 692119 862575 692355 865870
rect 687724 862552 692355 862575
rect 694233 862552 694469 869012
rect 696449 865870 696633 869012
rect 696347 862552 696633 865870
rect 687724 862266 696633 862552
rect 703733 869192 705676 878483
rect 703733 862312 705677 869192
rect 706576 877123 713395 878483
rect 706576 862674 706938 877123
rect 711303 876897 713395 877123
rect 711303 865006 711695 876897
rect 712309 865006 713395 876897
rect 711303 862674 713395 865006
rect 706576 862313 713395 862674
rect 706576 862312 711646 862313
rect 39559 829972 39863 841793
rect 677737 819207 678041 831028
rect 5954 800487 11024 800488
rect 4205 800126 11024 800487
rect 4205 797794 6297 800126
rect 4205 785903 5291 797794
rect 5905 785903 6297 797794
rect 4205 785677 6297 785903
rect 10662 785677 11024 800126
rect 4205 784317 11024 785677
rect 11923 793608 13867 800488
rect 11924 784317 13867 793608
rect 20967 800248 29876 800534
rect 20967 796930 21253 800248
rect 20967 793788 21151 796930
rect 23131 793788 23367 800248
rect 25245 800225 29876 800248
rect 25245 796930 25481 800225
rect 26791 798467 26961 800225
rect 29590 798467 29876 800225
rect 25347 793788 25481 796930
rect 32789 797366 34043 800490
rect 34931 797366 36169 800490
rect 32789 796055 33518 797366
rect 32789 794183 33147 796055
rect 22452 786084 22668 786099
rect 22344 785595 22668 786084
rect 21636 785306 22668 785595
rect 21636 784959 22884 785306
rect 21520 784376 22884 784959
rect 23753 784543 24039 789363
rect 27796 786492 27846 787107
rect 27796 785162 27964 786492
rect 27532 784543 27964 785162
rect 28396 784543 28682 789103
rect 35384 785316 36169 797366
rect 678733 788578 679465 789283
rect 688918 789057 693847 789343
rect 695297 789224 696080 789283
rect 21520 784317 22303 784376
rect 23753 784257 28682 784543
rect 38135 784317 38867 785022
rect 681431 776234 682216 788284
rect 688918 784497 689204 789057
rect 689636 788438 690068 789057
rect 689636 787108 689804 788438
rect 689754 786493 689804 787108
rect 693561 784237 693847 789057
rect 694716 788641 696080 789224
rect 694716 788294 695964 788641
rect 694932 788005 695964 788294
rect 694932 787516 695256 788005
rect 694932 787501 695148 787516
rect 684453 777545 684811 779417
rect 684082 776234 684811 777545
rect 681431 773110 682669 776234
rect 683557 773110 684811 776234
rect 692119 776670 692253 779812
rect 687724 773375 688010 775133
rect 690639 773375 690809 775133
rect 692119 773375 692355 776670
rect 687724 773352 692355 773375
rect 694233 773352 694469 779812
rect 696449 776670 696633 779812
rect 696347 773352 696633 776670
rect 687724 773066 696633 773352
rect 703733 779992 705676 789283
rect 703733 773112 705677 779992
rect 706576 787923 713395 789283
rect 706576 773474 706938 787923
rect 711303 787697 713395 787923
rect 711303 775806 711695 787697
rect 712309 775806 713395 787697
rect 711303 773474 713395 775806
rect 706576 773113 713395 773474
rect 706576 773112 711646 773113
rect 5954 757287 11024 757288
rect 4205 756926 11024 757287
rect 4205 754594 6297 756926
rect 4205 742703 5291 754594
rect 5905 742703 6297 754594
rect 4205 742477 6297 742703
rect 10662 742477 11024 756926
rect 4205 741117 11024 742477
rect 11923 750408 13867 757288
rect 11924 741117 13867 750408
rect 20967 757048 29876 757334
rect 20967 753730 21253 757048
rect 20967 750588 21151 753730
rect 23131 750588 23367 757048
rect 25245 757025 29876 757048
rect 25245 753730 25481 757025
rect 26791 755267 26961 757025
rect 29590 755267 29876 757025
rect 25347 750588 25481 753730
rect 32789 754166 34043 757290
rect 34931 754166 36169 757290
rect 32789 752855 33518 754166
rect 32789 750983 33147 752855
rect 22452 742884 22668 742899
rect 22344 742395 22668 742884
rect 21636 742106 22668 742395
rect 21636 741759 22884 742106
rect 21520 741176 22884 741759
rect 23753 741343 24039 746163
rect 27796 743292 27846 743907
rect 27796 741962 27964 743292
rect 27532 741343 27964 741962
rect 28396 741343 28682 745903
rect 35384 742116 36169 754166
rect 678733 743578 679465 744283
rect 688918 744057 693847 744343
rect 695297 744224 696080 744283
rect 21520 741117 22303 741176
rect 23753 741057 28682 741343
rect 38135 741117 38867 741822
rect 681431 731234 682216 743284
rect 688918 739497 689204 744057
rect 689636 743438 690068 744057
rect 689636 742108 689804 743438
rect 689754 741493 689804 742108
rect 693561 739237 693847 744057
rect 694716 743641 696080 744224
rect 694716 743294 695964 743641
rect 694932 743005 695964 743294
rect 694932 742516 695256 743005
rect 694932 742501 695148 742516
rect 684453 732545 684811 734417
rect 684082 731234 684811 732545
rect 681431 728110 682669 731234
rect 683557 728110 684811 731234
rect 692119 731670 692253 734812
rect 687724 728375 688010 730133
rect 690639 728375 690809 730133
rect 692119 728375 692355 731670
rect 687724 728352 692355 728375
rect 694233 728352 694469 734812
rect 696449 731670 696633 734812
rect 696347 728352 696633 731670
rect 687724 728066 696633 728352
rect 703733 734992 705676 744283
rect 703733 728112 705677 734992
rect 706576 742923 713395 744283
rect 706576 728474 706938 742923
rect 711303 742697 713395 742923
rect 711303 730806 711695 742697
rect 712309 730806 713395 742697
rect 711303 728474 713395 730806
rect 706576 728113 713395 728474
rect 706576 728112 711646 728113
rect 5954 714087 11024 714088
rect 4205 713726 11024 714087
rect 4205 711394 6297 713726
rect 4205 699503 5291 711394
rect 5905 699503 6297 711394
rect 4205 699277 6297 699503
rect 10662 699277 11024 713726
rect 4205 697917 11024 699277
rect 11923 707208 13867 714088
rect 11924 697917 13867 707208
rect 20967 713848 29876 714134
rect 20967 710530 21253 713848
rect 20967 707388 21151 710530
rect 23131 707388 23367 713848
rect 25245 713825 29876 713848
rect 25245 710530 25481 713825
rect 26791 712067 26961 713825
rect 29590 712067 29876 713825
rect 25347 707388 25481 710530
rect 32789 710966 34043 714090
rect 34931 710966 36169 714090
rect 32789 709655 33518 710966
rect 32789 707783 33147 709655
rect 22452 699684 22668 699699
rect 22344 699195 22668 699684
rect 21636 698906 22668 699195
rect 21636 698559 22884 698906
rect 21520 697976 22884 698559
rect 23753 698143 24039 702963
rect 27796 700092 27846 700707
rect 27796 698762 27964 700092
rect 27532 698143 27964 698762
rect 28396 698143 28682 702703
rect 35384 698916 36169 710966
rect 21520 697917 22303 697976
rect 23753 697857 28682 698143
rect 38135 697917 38867 698622
rect 678733 698578 679465 699283
rect 688918 699057 693847 699343
rect 695297 699224 696080 699283
rect 681431 686234 682216 698284
rect 688918 694497 689204 699057
rect 689636 698438 690068 699057
rect 689636 697108 689804 698438
rect 689754 696493 689804 697108
rect 693561 694237 693847 699057
rect 694716 698641 696080 699224
rect 694716 698294 695964 698641
rect 694932 698005 695964 698294
rect 694932 697516 695256 698005
rect 694932 697501 695148 697516
rect 684453 687545 684811 689417
rect 684082 686234 684811 687545
rect 681431 683110 682669 686234
rect 683557 683110 684811 686234
rect 692119 686670 692253 689812
rect 687724 683375 688010 685133
rect 690639 683375 690809 685133
rect 692119 683375 692355 686670
rect 687724 683352 692355 683375
rect 694233 683352 694469 689812
rect 696449 686670 696633 689812
rect 696347 683352 696633 686670
rect 687724 683066 696633 683352
rect 703733 689992 705676 699283
rect 703733 683112 705677 689992
rect 706576 697923 713395 699283
rect 706576 683474 706938 697923
rect 711303 697697 713395 697923
rect 711303 685806 711695 697697
rect 712309 685806 713395 697697
rect 711303 683474 713395 685806
rect 706576 683113 713395 683474
rect 706576 683112 711646 683113
rect 5954 670887 11024 670888
rect 4205 670526 11024 670887
rect 4205 668194 6297 670526
rect 4205 656303 5291 668194
rect 5905 656303 6297 668194
rect 4205 656077 6297 656303
rect 10662 656077 11024 670526
rect 4205 654717 11024 656077
rect 11923 664008 13867 670888
rect 11924 654717 13867 664008
rect 20967 670648 29876 670934
rect 20967 667330 21253 670648
rect 20967 664188 21151 667330
rect 23131 664188 23367 670648
rect 25245 670625 29876 670648
rect 25245 667330 25481 670625
rect 26791 668867 26961 670625
rect 29590 668867 29876 670625
rect 25347 664188 25481 667330
rect 32789 667766 34043 670890
rect 34931 667766 36169 670890
rect 32789 666455 33518 667766
rect 32789 664583 33147 666455
rect 22452 656484 22668 656499
rect 22344 655995 22668 656484
rect 21636 655706 22668 655995
rect 21636 655359 22884 655706
rect 21520 654776 22884 655359
rect 23753 654943 24039 659763
rect 27796 656892 27846 657507
rect 27796 655562 27964 656892
rect 27532 654943 27964 655562
rect 28396 654943 28682 659503
rect 35384 655716 36169 667766
rect 21520 654717 22303 654776
rect 23753 654657 28682 654943
rect 38135 654717 38867 655422
rect 678733 653378 679465 654083
rect 688918 653857 693847 654143
rect 695297 654024 696080 654083
rect 681431 641034 682216 653084
rect 688918 649297 689204 653857
rect 689636 653238 690068 653857
rect 689636 651908 689804 653238
rect 689754 651293 689804 651908
rect 693561 649037 693847 653857
rect 694716 653441 696080 654024
rect 694716 653094 695964 653441
rect 694932 652805 695964 653094
rect 694932 652316 695256 652805
rect 694932 652301 695148 652316
rect 684453 642345 684811 644217
rect 684082 641034 684811 642345
rect 681431 637910 682669 641034
rect 683557 637910 684811 641034
rect 692119 641470 692253 644612
rect 687724 638175 688010 639933
rect 690639 638175 690809 639933
rect 692119 638175 692355 641470
rect 687724 638152 692355 638175
rect 694233 638152 694469 644612
rect 696449 641470 696633 644612
rect 696347 638152 696633 641470
rect 687724 637866 696633 638152
rect 703733 644792 705676 654083
rect 703733 637912 705677 644792
rect 706576 652723 713395 654083
rect 706576 638274 706938 652723
rect 711303 652497 713395 652723
rect 711303 640606 711695 652497
rect 712309 640606 713395 652497
rect 711303 638274 713395 640606
rect 706576 637913 713395 638274
rect 706576 637912 711646 637913
rect 5954 627687 11024 627688
rect 4205 627326 11024 627687
rect 4205 624994 6297 627326
rect 4205 613103 5291 624994
rect 5905 613103 6297 624994
rect 4205 612877 6297 613103
rect 10662 612877 11024 627326
rect 4205 611517 11024 612877
rect 11923 620808 13867 627688
rect 11924 611517 13867 620808
rect 20967 627448 29876 627734
rect 20967 624130 21253 627448
rect 20967 620988 21151 624130
rect 23131 620988 23367 627448
rect 25245 627425 29876 627448
rect 25245 624130 25481 627425
rect 26791 625667 26961 627425
rect 29590 625667 29876 627425
rect 25347 620988 25481 624130
rect 32789 624566 34043 627690
rect 34931 624566 36169 627690
rect 32789 623255 33518 624566
rect 32789 621383 33147 623255
rect 22452 613284 22668 613299
rect 22344 612795 22668 613284
rect 21636 612506 22668 612795
rect 21636 612159 22884 612506
rect 21520 611576 22884 612159
rect 23753 611743 24039 616563
rect 27796 613692 27846 614307
rect 27796 612362 27964 613692
rect 27532 611743 27964 612362
rect 28396 611743 28682 616303
rect 35384 612516 36169 624566
rect 21520 611517 22303 611576
rect 23753 611457 28682 611743
rect 38135 611517 38867 612222
rect 678733 608378 679465 609083
rect 688918 608857 693847 609143
rect 695297 609024 696080 609083
rect 681431 596034 682216 608084
rect 688918 604297 689204 608857
rect 689636 608238 690068 608857
rect 689636 606908 689804 608238
rect 689754 606293 689804 606908
rect 693561 604037 693847 608857
rect 694716 608441 696080 609024
rect 694716 608094 695964 608441
rect 694932 607805 695964 608094
rect 694932 607316 695256 607805
rect 694932 607301 695148 607316
rect 684453 597345 684811 599217
rect 684082 596034 684811 597345
rect 681431 592910 682669 596034
rect 683557 592910 684811 596034
rect 692119 596470 692253 599612
rect 687724 593175 688010 594933
rect 690639 593175 690809 594933
rect 692119 593175 692355 596470
rect 687724 593152 692355 593175
rect 694233 593152 694469 599612
rect 696449 596470 696633 599612
rect 696347 593152 696633 596470
rect 687724 592866 696633 593152
rect 703733 599792 705676 609083
rect 703733 592912 705677 599792
rect 706576 607723 713395 609083
rect 706576 593274 706938 607723
rect 711303 607497 713395 607723
rect 711303 595606 711695 607497
rect 712309 595606 713395 607497
rect 711303 593274 713395 595606
rect 706576 592913 713395 593274
rect 706576 592912 711646 592913
rect 5954 584487 11024 584488
rect 4205 584126 11024 584487
rect 4205 581794 6297 584126
rect 4205 569903 5291 581794
rect 5905 569903 6297 581794
rect 4205 569677 6297 569903
rect 10662 569677 11024 584126
rect 4205 568317 11024 569677
rect 11923 577608 13867 584488
rect 11924 568317 13867 577608
rect 20967 584248 29876 584534
rect 20967 580930 21253 584248
rect 20967 577788 21151 580930
rect 23131 577788 23367 584248
rect 25245 584225 29876 584248
rect 25245 580930 25481 584225
rect 26791 582467 26961 584225
rect 29590 582467 29876 584225
rect 25347 577788 25481 580930
rect 32789 581366 34043 584490
rect 34931 581366 36169 584490
rect 32789 580055 33518 581366
rect 32789 578183 33147 580055
rect 22452 570084 22668 570099
rect 22344 569595 22668 570084
rect 21636 569306 22668 569595
rect 21636 568959 22884 569306
rect 21520 568376 22884 568959
rect 23753 568543 24039 573363
rect 27796 570492 27846 571107
rect 27796 569162 27964 570492
rect 27532 568543 27964 569162
rect 28396 568543 28682 573103
rect 35384 569316 36169 581366
rect 21520 568317 22303 568376
rect 23753 568257 28682 568543
rect 38135 568317 38867 569022
rect 678733 563178 679465 563883
rect 688918 563657 693847 563943
rect 695297 563824 696080 563883
rect 681431 550834 682216 562884
rect 688918 559097 689204 563657
rect 689636 563038 690068 563657
rect 689636 561708 689804 563038
rect 689754 561093 689804 561708
rect 693561 558837 693847 563657
rect 694716 563241 696080 563824
rect 694716 562894 695964 563241
rect 694932 562605 695964 562894
rect 694932 562116 695256 562605
rect 694932 562101 695148 562116
rect 684453 552145 684811 554017
rect 684082 550834 684811 552145
rect 681431 547710 682669 550834
rect 683557 547710 684811 550834
rect 692119 551270 692253 554412
rect 687724 547975 688010 549733
rect 690639 547975 690809 549733
rect 692119 547975 692355 551270
rect 687724 547952 692355 547975
rect 694233 547952 694469 554412
rect 696449 551270 696633 554412
rect 696347 547952 696633 551270
rect 687724 547666 696633 547952
rect 703733 554592 705676 563883
rect 703733 547712 705677 554592
rect 706576 562523 713395 563883
rect 706576 548074 706938 562523
rect 711303 562297 713395 562523
rect 711303 550406 711695 562297
rect 712309 550406 713395 562297
rect 711303 548074 713395 550406
rect 706576 547713 713395 548074
rect 706576 547712 711646 547713
rect 5954 541287 11024 541288
rect 4205 540926 11024 541287
rect 4205 538594 6297 540926
rect 4205 526703 5291 538594
rect 5905 526703 6297 538594
rect 4205 526477 6297 526703
rect 10662 526477 11024 540926
rect 4205 525117 11024 526477
rect 11923 534408 13867 541288
rect 11924 525117 13867 534408
rect 20967 541048 29876 541334
rect 20967 537730 21253 541048
rect 20967 534588 21151 537730
rect 23131 534588 23367 541048
rect 25245 541025 29876 541048
rect 25245 537730 25481 541025
rect 26791 539267 26961 541025
rect 29590 539267 29876 541025
rect 25347 534588 25481 537730
rect 32789 538166 34043 541290
rect 34931 538166 36169 541290
rect 32789 536855 33518 538166
rect 32789 534983 33147 536855
rect 22452 526884 22668 526899
rect 22344 526395 22668 526884
rect 21636 526106 22668 526395
rect 21636 525759 22884 526106
rect 21520 525176 22884 525759
rect 23753 525343 24039 530163
rect 27796 527292 27846 527907
rect 27796 525962 27964 527292
rect 27532 525343 27964 525962
rect 28396 525343 28682 529903
rect 35384 526116 36169 538166
rect 21520 525117 22303 525176
rect 23753 525057 28682 525343
rect 38135 525117 38867 525822
rect 677737 504607 678041 516428
rect 39559 485372 39863 497193
rect 677737 416407 678041 428228
rect 5954 413687 11024 413688
rect 4205 413326 11024 413687
rect 4205 410994 6297 413326
rect 4205 399103 5291 410994
rect 5905 399103 6297 410994
rect 4205 398877 6297 399103
rect 10662 398877 11024 413326
rect 4205 397517 11024 398877
rect 11923 406808 13867 413688
rect 11924 397517 13867 406808
rect 20967 413448 29876 413734
rect 20967 410130 21253 413448
rect 20967 406988 21151 410130
rect 23131 406988 23367 413448
rect 25245 413425 29876 413448
rect 25245 410130 25481 413425
rect 26791 411667 26961 413425
rect 29590 411667 29876 413425
rect 25347 406988 25481 410130
rect 32789 410566 34043 413690
rect 34931 410566 36169 413690
rect 32789 409255 33518 410566
rect 32789 407383 33147 409255
rect 22452 399284 22668 399299
rect 22344 398795 22668 399284
rect 21636 398506 22668 398795
rect 21636 398159 22884 398506
rect 21520 397576 22884 398159
rect 23753 397743 24039 402563
rect 27796 399692 27846 400307
rect 27796 398362 27964 399692
rect 27532 397743 27964 398362
rect 28396 397743 28682 402303
rect 35384 398516 36169 410566
rect 21520 397517 22303 397576
rect 23753 397457 28682 397743
rect 38135 397517 38867 398222
rect 678733 385978 679465 386683
rect 688918 386457 693847 386743
rect 695297 386624 696080 386683
rect 681431 373634 682216 385684
rect 688918 381897 689204 386457
rect 689636 385838 690068 386457
rect 689636 384508 689804 385838
rect 689754 383893 689804 384508
rect 693561 381637 693847 386457
rect 694716 386041 696080 386624
rect 694716 385694 695964 386041
rect 694932 385405 695964 385694
rect 694932 384916 695256 385405
rect 694932 384901 695148 384916
rect 684453 374945 684811 376817
rect 684082 373634 684811 374945
rect 5954 370487 11024 370488
rect 4205 370126 11024 370487
rect 4205 367794 6297 370126
rect 4205 355903 5291 367794
rect 5905 355903 6297 367794
rect 4205 355677 6297 355903
rect 10662 355677 11024 370126
rect 4205 354317 11024 355677
rect 11923 363608 13867 370488
rect 11924 354317 13867 363608
rect 20967 370248 29876 370534
rect 681431 370510 682669 373634
rect 683557 370510 684811 373634
rect 692119 374070 692253 377212
rect 687724 370775 688010 372533
rect 690639 370775 690809 372533
rect 692119 370775 692355 374070
rect 687724 370752 692355 370775
rect 694233 370752 694469 377212
rect 696449 374070 696633 377212
rect 696347 370752 696633 374070
rect 20967 366930 21253 370248
rect 20967 363788 21151 366930
rect 23131 363788 23367 370248
rect 25245 370225 29876 370248
rect 25245 366930 25481 370225
rect 26791 368467 26961 370225
rect 29590 368467 29876 370225
rect 25347 363788 25481 366930
rect 32789 367366 34043 370490
rect 34931 367366 36169 370490
rect 687724 370466 696633 370752
rect 703733 377392 705676 386683
rect 703733 370512 705677 377392
rect 706576 385323 713395 386683
rect 706576 370874 706938 385323
rect 711303 385097 713395 385323
rect 711303 373206 711695 385097
rect 712309 373206 713395 385097
rect 711303 370874 713395 373206
rect 706576 370513 713395 370874
rect 706576 370512 711646 370513
rect 32789 366055 33518 367366
rect 32789 364183 33147 366055
rect 22452 356084 22668 356099
rect 22344 355595 22668 356084
rect 21636 355306 22668 355595
rect 21636 354959 22884 355306
rect 21520 354376 22884 354959
rect 23753 354543 24039 359363
rect 27796 356492 27846 357107
rect 27796 355162 27964 356492
rect 27532 354543 27964 355162
rect 28396 354543 28682 359103
rect 35384 355316 36169 367366
rect 21520 354317 22303 354376
rect 23753 354257 28682 354543
rect 38135 354317 38867 355022
rect 678733 340778 679465 341483
rect 688918 341257 693847 341543
rect 695297 341424 696080 341483
rect 681431 328434 682216 340484
rect 688918 336697 689204 341257
rect 689636 340638 690068 341257
rect 689636 339308 689804 340638
rect 689754 338693 689804 339308
rect 693561 336437 693847 341257
rect 694716 340841 696080 341424
rect 694716 340494 695964 340841
rect 694932 340205 695964 340494
rect 694932 339716 695256 340205
rect 694932 339701 695148 339716
rect 684453 329745 684811 331617
rect 684082 328434 684811 329745
rect 5954 327287 11024 327288
rect 4205 326926 11024 327287
rect 4205 324594 6297 326926
rect 4205 312703 5291 324594
rect 5905 312703 6297 324594
rect 4205 312477 6297 312703
rect 10662 312477 11024 326926
rect 4205 311117 11024 312477
rect 11923 320408 13867 327288
rect 11924 311117 13867 320408
rect 20967 327048 29876 327334
rect 20967 323730 21253 327048
rect 20967 320588 21151 323730
rect 23131 320588 23367 327048
rect 25245 327025 29876 327048
rect 25245 323730 25481 327025
rect 26791 325267 26961 327025
rect 29590 325267 29876 327025
rect 25347 320588 25481 323730
rect 32789 324166 34043 327290
rect 34931 324166 36169 327290
rect 681431 325310 682669 328434
rect 683557 325310 684811 328434
rect 692119 328870 692253 332012
rect 687724 325575 688010 327333
rect 690639 325575 690809 327333
rect 692119 325575 692355 328870
rect 687724 325552 692355 325575
rect 694233 325552 694469 332012
rect 696449 328870 696633 332012
rect 696347 325552 696633 328870
rect 687724 325266 696633 325552
rect 703733 332192 705676 341483
rect 703733 325312 705677 332192
rect 706576 340123 713395 341483
rect 706576 325674 706938 340123
rect 711303 339897 713395 340123
rect 711303 328006 711695 339897
rect 712309 328006 713395 339897
rect 711303 325674 713395 328006
rect 706576 325313 713395 325674
rect 706576 325312 711646 325313
rect 32789 322855 33518 324166
rect 32789 320983 33147 322855
rect 22452 312884 22668 312899
rect 22344 312395 22668 312884
rect 21636 312106 22668 312395
rect 21636 311759 22884 312106
rect 21520 311176 22884 311759
rect 23753 311343 24039 316163
rect 27796 313292 27846 313907
rect 27796 311962 27964 313292
rect 27532 311343 27964 311962
rect 28396 311343 28682 315903
rect 35384 312116 36169 324166
rect 21520 311117 22303 311176
rect 23753 311057 28682 311343
rect 38135 311117 38867 311822
rect 678733 295778 679465 296483
rect 688918 296257 693847 296543
rect 695297 296424 696080 296483
rect 5954 284087 11024 284088
rect 4205 283726 11024 284087
rect 4205 281394 6297 283726
rect 4205 269503 5291 281394
rect 5905 269503 6297 281394
rect 4205 269277 6297 269503
rect 10662 269277 11024 283726
rect 4205 267917 11024 269277
rect 11923 277208 13867 284088
rect 11924 267917 13867 277208
rect 20967 283848 29876 284134
rect 20967 280530 21253 283848
rect 20967 277388 21151 280530
rect 23131 277388 23367 283848
rect 25245 283825 29876 283848
rect 25245 280530 25481 283825
rect 26791 282067 26961 283825
rect 29590 282067 29876 283825
rect 25347 277388 25481 280530
rect 32789 280966 34043 284090
rect 34931 280966 36169 284090
rect 32789 279655 33518 280966
rect 32789 277783 33147 279655
rect 22452 269684 22668 269699
rect 22344 269195 22668 269684
rect 21636 268906 22668 269195
rect 21636 268559 22884 268906
rect 21520 267976 22884 268559
rect 23753 268143 24039 272963
rect 27796 270092 27846 270707
rect 27796 268762 27964 270092
rect 27532 268143 27964 268762
rect 28396 268143 28682 272703
rect 35384 268916 36169 280966
rect 681431 283434 682216 295484
rect 688918 291697 689204 296257
rect 689636 295638 690068 296257
rect 689636 294308 689804 295638
rect 689754 293693 689804 294308
rect 693561 291437 693847 296257
rect 694716 295841 696080 296424
rect 694716 295494 695964 295841
rect 694932 295205 695964 295494
rect 694932 294716 695256 295205
rect 694932 294701 695148 294716
rect 684453 284745 684811 286617
rect 684082 283434 684811 284745
rect 681431 280310 682669 283434
rect 683557 280310 684811 283434
rect 692119 283870 692253 287012
rect 687724 280575 688010 282333
rect 690639 280575 690809 282333
rect 692119 280575 692355 283870
rect 687724 280552 692355 280575
rect 694233 280552 694469 287012
rect 696449 283870 696633 287012
rect 696347 280552 696633 283870
rect 687724 280266 696633 280552
rect 703733 287192 705676 296483
rect 703733 280312 705677 287192
rect 706576 295123 713395 296483
rect 706576 280674 706938 295123
rect 711303 294897 713395 295123
rect 711303 283006 711695 294897
rect 712309 283006 713395 294897
rect 711303 280674 713395 283006
rect 706576 280313 713395 280674
rect 706576 280312 711646 280313
rect 21520 267917 22303 267976
rect 23753 267857 28682 268143
rect 38135 267917 38867 268622
rect 678733 250778 679465 251483
rect 688918 251257 693847 251543
rect 695297 251424 696080 251483
rect 5954 240887 11024 240888
rect 4205 240526 11024 240887
rect 4205 238194 6297 240526
rect 4205 226303 5291 238194
rect 5905 226303 6297 238194
rect 4205 226077 6297 226303
rect 10662 226077 11024 240526
rect 4205 224717 11024 226077
rect 11923 234008 13867 240888
rect 11924 224717 13867 234008
rect 20967 240648 29876 240934
rect 20967 237330 21253 240648
rect 20967 234188 21151 237330
rect 23131 234188 23367 240648
rect 25245 240625 29876 240648
rect 25245 237330 25481 240625
rect 26791 238867 26961 240625
rect 29590 238867 29876 240625
rect 25347 234188 25481 237330
rect 32789 237766 34043 240890
rect 34931 237766 36169 240890
rect 32789 236455 33518 237766
rect 32789 234583 33147 236455
rect 22452 226484 22668 226499
rect 22344 225995 22668 226484
rect 21636 225706 22668 225995
rect 21636 225359 22884 225706
rect 21520 224776 22884 225359
rect 23753 224943 24039 229763
rect 27796 226892 27846 227507
rect 27796 225562 27964 226892
rect 27532 224943 27964 225562
rect 28396 224943 28682 229503
rect 35384 225716 36169 237766
rect 681431 238434 682216 250484
rect 688918 246697 689204 251257
rect 689636 250638 690068 251257
rect 689636 249308 689804 250638
rect 689754 248693 689804 249308
rect 693561 246437 693847 251257
rect 694716 250841 696080 251424
rect 694716 250494 695964 250841
rect 694932 250205 695964 250494
rect 694932 249716 695256 250205
rect 694932 249701 695148 249716
rect 684453 239745 684811 241617
rect 684082 238434 684811 239745
rect 681431 235310 682669 238434
rect 683557 235310 684811 238434
rect 692119 238870 692253 242012
rect 687724 235575 688010 237333
rect 690639 235575 690809 237333
rect 692119 235575 692355 238870
rect 687724 235552 692355 235575
rect 694233 235552 694469 242012
rect 696449 238870 696633 242012
rect 696347 235552 696633 238870
rect 687724 235266 696633 235552
rect 703733 242192 705676 251483
rect 703733 235312 705677 242192
rect 706576 250123 713395 251483
rect 706576 235674 706938 250123
rect 711303 249897 713395 250123
rect 711303 238006 711695 249897
rect 712309 238006 713395 249897
rect 711303 235674 713395 238006
rect 706576 235313 713395 235674
rect 706576 235312 711646 235313
rect 21520 224717 22303 224776
rect 23753 224657 28682 224943
rect 38135 224717 38867 225422
rect 678733 205578 679465 206283
rect 688918 206057 693847 206343
rect 695297 206224 696080 206283
rect 5954 197687 11024 197688
rect 4205 197326 11024 197687
rect 4205 194994 6297 197326
rect 4205 183103 5291 194994
rect 5905 183103 6297 194994
rect 4205 182877 6297 183103
rect 10662 182877 11024 197326
rect 4205 181517 11024 182877
rect 11923 190808 13867 197688
rect 11924 181517 13867 190808
rect 20967 197448 29876 197734
rect 20967 194130 21253 197448
rect 20967 190988 21151 194130
rect 23131 190988 23367 197448
rect 25245 197425 29876 197448
rect 25245 194130 25481 197425
rect 26791 195667 26961 197425
rect 29590 195667 29876 197425
rect 25347 190988 25481 194130
rect 32789 194566 34043 197690
rect 34931 194566 36169 197690
rect 32789 193255 33518 194566
rect 32789 191383 33147 193255
rect 22452 183284 22668 183299
rect 22344 182795 22668 183284
rect 21636 182506 22668 182795
rect 21636 182159 22884 182506
rect 21520 181576 22884 182159
rect 23753 181743 24039 186563
rect 27796 183692 27846 184307
rect 27796 182362 27964 183692
rect 27532 181743 27964 182362
rect 28396 181743 28682 186303
rect 35384 182516 36169 194566
rect 681431 193234 682216 205284
rect 688918 201497 689204 206057
rect 689636 205438 690068 206057
rect 689636 204108 689804 205438
rect 689754 203493 689804 204108
rect 693561 201237 693847 206057
rect 694716 205641 696080 206224
rect 694716 205294 695964 205641
rect 694932 205005 695964 205294
rect 694932 204516 695256 205005
rect 694932 204501 695148 204516
rect 684453 194545 684811 196417
rect 684082 193234 684811 194545
rect 681431 190110 682669 193234
rect 683557 190110 684811 193234
rect 692119 193670 692253 196812
rect 687724 190375 688010 192133
rect 690639 190375 690809 192133
rect 692119 190375 692355 193670
rect 687724 190352 692355 190375
rect 694233 190352 694469 196812
rect 696449 193670 696633 196812
rect 696347 190352 696633 193670
rect 687724 190066 696633 190352
rect 703733 196992 705676 206283
rect 703733 190112 705677 196992
rect 706576 204923 713395 206283
rect 706576 190474 706938 204923
rect 711303 204697 713395 204923
rect 711303 192806 711695 204697
rect 712309 192806 713395 204697
rect 711303 190474 713395 192806
rect 706576 190113 713395 190474
rect 706576 190112 711646 190113
rect 21520 181517 22303 181576
rect 23753 181457 28682 181743
rect 38135 181517 38867 182222
rect 678733 160578 679465 161283
rect 688918 161057 693847 161343
rect 695297 161224 696080 161283
rect 681431 148234 682216 160284
rect 688918 156497 689204 161057
rect 689636 160438 690068 161057
rect 689636 159108 689804 160438
rect 689754 158493 689804 159108
rect 693561 156237 693847 161057
rect 694716 160641 696080 161224
rect 694716 160294 695964 160641
rect 694932 160005 695964 160294
rect 694932 159516 695256 160005
rect 694932 159501 695148 159516
rect 684453 149545 684811 151417
rect 684082 148234 684811 149545
rect 681431 145110 682669 148234
rect 683557 145110 684811 148234
rect 692119 148670 692253 151812
rect 687724 145375 688010 147133
rect 690639 145375 690809 147133
rect 692119 145375 692355 148670
rect 687724 145352 692355 145375
rect 694233 145352 694469 151812
rect 696449 148670 696633 151812
rect 696347 145352 696633 148670
rect 687724 145066 696633 145352
rect 703733 151992 705676 161283
rect 703733 145112 705677 151992
rect 706576 159923 713395 161283
rect 706576 145474 706938 159923
rect 711303 159697 713395 159923
rect 711303 147806 711695 159697
rect 712309 147806 713395 159697
rect 711303 145474 713395 147806
rect 706576 145113 713395 145474
rect 706576 145112 711646 145113
rect 39559 112572 39863 124393
rect 678733 115378 679465 116083
rect 688918 115857 693847 116143
rect 695297 116024 696080 116083
rect 681431 103034 682216 115084
rect 688918 111297 689204 115857
rect 689636 115238 690068 115857
rect 689636 113908 689804 115238
rect 689754 113293 689804 113908
rect 693561 111037 693847 115857
rect 694716 115441 696080 116024
rect 694716 115094 695964 115441
rect 694932 114805 695964 115094
rect 694932 114316 695256 114805
rect 694932 114301 695148 114316
rect 684453 104345 684811 106217
rect 684082 103034 684811 104345
rect 681431 99910 682669 103034
rect 683557 99910 684811 103034
rect 692119 103470 692253 106612
rect 687724 100175 688010 101933
rect 690639 100175 690809 101933
rect 692119 100175 692355 103470
rect 687724 100152 692355 100175
rect 694233 100152 694469 106612
rect 696449 103470 696633 106612
rect 696347 100152 696633 103470
rect 687724 99866 696633 100152
rect 703733 106792 705676 116083
rect 703733 99912 705677 106792
rect 706576 114723 713395 116083
rect 706576 100274 706938 114723
rect 711303 114497 713395 114723
rect 711303 102606 711695 114497
rect 712309 102606 713395 114497
rect 711303 100274 713395 102606
rect 706576 99913 713395 100274
rect 706576 99912 711646 99913
rect 79607 39559 91428 39863
rect 569807 39559 581628 39863
rect 623607 39559 635428 39863
rect 201778 38135 202483 38867
rect 310378 38135 311083 38867
rect 365178 38135 365883 38867
rect 419978 38135 420683 38867
rect 474778 38135 475483 38867
rect 529578 38135 530283 38867
rect 186310 35384 201484 36169
rect 294910 35384 310084 36169
rect 349710 35384 364884 36169
rect 404510 35384 419684 36169
rect 459310 35384 474484 36169
rect 514110 35384 529284 36169
rect 186310 34931 189434 35384
rect 294910 34931 298034 35384
rect 349710 34931 352834 35384
rect 404510 34931 407634 35384
rect 459310 34931 462434 35384
rect 514110 34931 517234 35384
rect 186310 33518 189434 34043
rect 294910 33518 298034 34043
rect 349710 33518 352834 34043
rect 404510 33518 407634 34043
rect 459310 33518 462434 34043
rect 514110 33518 517234 34043
rect 186310 33147 190745 33518
rect 294910 33147 299345 33518
rect 349710 33147 354145 33518
rect 404510 33147 408945 33518
rect 459310 33147 463745 33518
rect 514110 33147 518545 33518
rect 186310 32789 192617 33147
rect 294910 32789 301217 33147
rect 349710 32789 356017 33147
rect 404510 32789 410817 33147
rect 459310 32789 465617 33147
rect 514110 32789 520417 33147
rect 186266 29590 188333 29876
rect 294866 29590 296933 29876
rect 349666 29590 351733 29876
rect 404466 29590 406533 29876
rect 459266 29590 461333 29876
rect 514066 29590 516133 29876
rect 186266 26961 186575 29590
rect 197697 28396 202543 28682
rect 202257 27964 202543 28396
rect 200308 27846 202543 27964
rect 199693 27796 202543 27846
rect 201638 27532 202543 27796
rect 186266 26791 188333 26961
rect 186266 25481 186575 26791
rect 186266 25347 193012 25481
rect 186266 25245 189870 25347
rect 186266 23367 186552 25245
rect 202257 24039 202543 27532
rect 197437 23753 202543 24039
rect 294866 26961 295175 29590
rect 306297 28396 311143 28682
rect 310857 27964 311143 28396
rect 308908 27846 311143 27964
rect 308293 27796 311143 27846
rect 310238 27532 311143 27796
rect 294866 26791 296933 26961
rect 294866 25481 295175 26791
rect 294866 25347 301612 25481
rect 294866 25245 298470 25347
rect 294866 23367 295152 25245
rect 310857 24039 311143 27532
rect 306037 23753 311143 24039
rect 349666 26961 349975 29590
rect 361097 28396 365943 28682
rect 365657 27964 365943 28396
rect 363708 27846 365943 27964
rect 363093 27796 365943 27846
rect 365038 27532 365943 27796
rect 349666 26791 351733 26961
rect 349666 25481 349975 26791
rect 349666 25347 356412 25481
rect 349666 25245 353270 25347
rect 349666 23367 349952 25245
rect 365657 24039 365943 27532
rect 360837 23753 365943 24039
rect 404466 26961 404775 29590
rect 415897 28396 420743 28682
rect 420457 27964 420743 28396
rect 418508 27846 420743 27964
rect 417893 27796 420743 27846
rect 419838 27532 420743 27796
rect 404466 26791 406533 26961
rect 404466 25481 404775 26791
rect 404466 25347 411212 25481
rect 404466 25245 408070 25347
rect 404466 23367 404752 25245
rect 420457 24039 420743 27532
rect 415637 23753 420743 24039
rect 459266 26961 459575 29590
rect 470697 28396 475543 28682
rect 475257 27964 475543 28396
rect 473308 27846 475543 27964
rect 472693 27796 475543 27846
rect 474638 27532 475543 27796
rect 459266 26791 461333 26961
rect 459266 25481 459575 26791
rect 459266 25347 466012 25481
rect 459266 25245 462870 25347
rect 459266 23367 459552 25245
rect 475257 24039 475543 27532
rect 470437 23753 475543 24039
rect 514066 26961 514375 29590
rect 525497 28396 530343 28682
rect 530057 27964 530343 28396
rect 528108 27846 530343 27964
rect 527493 27796 530343 27846
rect 529438 27532 530343 27796
rect 514066 26791 516133 26961
rect 514066 25481 514375 26791
rect 514066 25347 520812 25481
rect 514066 25245 517670 25347
rect 514066 23367 514352 25245
rect 530057 24039 530343 27532
rect 525237 23753 530343 24039
rect 186266 23131 193012 23367
rect 294866 23131 301612 23367
rect 349666 23131 356412 23367
rect 404466 23131 411212 23367
rect 459266 23131 466012 23367
rect 514066 23131 520812 23367
rect 186266 21253 186552 23131
rect 201494 22668 202424 22884
rect 200701 22452 202424 22668
rect 200716 22344 202424 22452
rect 201205 22303 202424 22344
rect 201205 21636 202483 22303
rect 201841 21520 202483 21636
rect 186266 21151 189870 21253
rect 186266 20967 193012 21151
rect 294866 21253 295152 23131
rect 310094 22668 311024 22884
rect 309301 22452 311024 22668
rect 309316 22344 311024 22452
rect 309805 22303 311024 22344
rect 309805 21636 311083 22303
rect 310441 21520 311083 21636
rect 294866 21151 298470 21253
rect 294866 20967 301612 21151
rect 349666 21253 349952 23131
rect 364894 22668 365824 22884
rect 364101 22452 365824 22668
rect 364116 22344 365824 22452
rect 364605 22303 365824 22344
rect 364605 21636 365883 22303
rect 365241 21520 365883 21636
rect 349666 21151 353270 21253
rect 349666 20967 356412 21151
rect 404466 21253 404752 23131
rect 419694 22668 420624 22884
rect 418901 22452 420624 22668
rect 418916 22344 420624 22452
rect 419405 22303 420624 22344
rect 419405 21636 420683 22303
rect 420041 21520 420683 21636
rect 404466 21151 408070 21253
rect 404466 20967 411212 21151
rect 459266 21253 459552 23131
rect 474494 22668 475424 22884
rect 473701 22452 475424 22668
rect 473716 22344 475424 22452
rect 474205 22303 475424 22344
rect 474205 21636 475483 22303
rect 474841 21520 475483 21636
rect 459266 21151 462870 21253
rect 459266 20967 466012 21151
rect 514066 21253 514352 23131
rect 529294 22668 530224 22884
rect 528501 22452 530224 22668
rect 528516 22344 530224 22452
rect 529005 22303 530224 22344
rect 529005 21636 530283 22303
rect 529641 21520 530283 21636
rect 514066 21151 517670 21253
rect 514066 20967 520812 21151
rect 132534 11924 147666 13867
rect 186312 11924 202483 13867
rect 294912 11924 311083 13867
rect 349712 11924 365883 13867
rect 404512 11924 420683 13867
rect 459312 11924 475483 13867
rect 514112 11924 530283 13867
rect 186312 11923 193192 11924
rect 294912 11923 301792 11924
rect 349712 11923 356592 11924
rect 404512 11923 411392 11924
rect 459312 11923 466192 11924
rect 514112 11923 520992 11924
rect 132476 10662 147703 11024
rect 132476 6297 132981 10662
rect 147265 6297 147703 10662
rect 132476 5958 147703 6297
rect 186312 10662 202483 11024
rect 186312 6297 186674 10662
rect 201123 6297 202483 10662
rect 186312 5954 202483 6297
rect 294912 10662 311083 11024
rect 294912 6297 295274 10662
rect 309723 6297 311083 10662
rect 294912 5954 311083 6297
rect 349712 10662 365883 11024
rect 349712 6297 350074 10662
rect 364523 6297 365883 10662
rect 349712 5954 365883 6297
rect 404512 10662 420683 11024
rect 404512 6297 404874 10662
rect 419323 6297 420683 10662
rect 404512 5954 420683 6297
rect 459312 10662 475483 11024
rect 459312 6297 459674 10662
rect 474123 6297 475483 10662
rect 459312 5954 475483 6297
rect 514112 10662 530283 11024
rect 514112 6297 514474 10662
rect 528923 6297 530283 10662
rect 514112 5954 530283 6297
rect 186313 5905 202483 5954
rect 186313 5291 189006 5905
rect 200897 5291 202483 5905
rect 186313 4205 202483 5291
rect 294913 5905 311083 5954
rect 294913 5291 297606 5905
rect 309497 5291 311083 5905
rect 294913 4205 311083 5291
rect 349713 5905 365883 5954
rect 349713 5291 352406 5905
rect 364297 5291 365883 5905
rect 349713 4205 365883 5291
rect 404513 5905 420683 5954
rect 404513 5291 407206 5905
rect 419097 5291 420683 5905
rect 404513 4205 420683 5291
rect 459313 5905 475483 5954
rect 459313 5291 462006 5905
rect 473897 5291 475483 5905
rect 459313 4205 475483 5291
rect 514113 5905 530283 5954
rect 514113 5291 516806 5905
rect 528697 5291 530283 5905
rect 514113 4205 530283 5291
<< pwell >>
rect 231099 997787 232657 1002358
rect 282699 997787 284257 1002358
rect 677787 965343 682358 966901
rect 35242 870499 39813 872057
rect 696187 877357 703671 878443
rect 696187 876540 696851 877357
rect 696591 870523 696851 876540
rect 697993 877253 703671 877357
rect 697993 870523 698310 877253
rect 696591 869232 697197 870523
rect 696591 869082 696652 869232
rect 696795 863046 697197 869232
rect 697764 867824 698310 870523
rect 697504 863046 698310 867824
rect 696795 862827 698310 863046
rect 702627 870351 703671 877253
rect 702627 865018 703463 870351
rect 702627 862827 703671 865018
rect 696795 862342 703671 862827
rect 705737 862342 706513 878458
rect 677787 831143 682358 832701
rect 11087 784342 11863 800458
rect 13929 799973 20805 800458
rect 13929 797782 14973 799973
rect 14137 792449 14973 797782
rect 13929 785547 14973 792449
rect 19290 799754 20805 799973
rect 19290 794976 20096 799754
rect 19290 792277 19836 794976
rect 20403 793568 20805 799754
rect 20948 793568 21009 793718
rect 20403 792277 21009 793568
rect 19290 785547 19607 792277
rect 13929 785443 19607 785547
rect 20749 786260 21009 792277
rect 20749 785443 21413 786260
rect 13929 784357 21413 785443
rect 696187 788157 703671 789243
rect 696187 787340 696851 788157
rect 696591 781323 696851 787340
rect 697993 788053 703671 788157
rect 697993 781323 698310 788053
rect 696591 780032 697197 781323
rect 696591 779882 696652 780032
rect 696795 773846 697197 780032
rect 697764 778624 698310 781323
rect 697504 773846 698310 778624
rect 696795 773627 698310 773846
rect 702627 781151 703671 788053
rect 702627 775818 703463 781151
rect 702627 773627 703671 775818
rect 696795 773142 703671 773627
rect 705737 773142 706513 789258
rect 11087 741142 11863 757258
rect 13929 756773 20805 757258
rect 13929 754582 14973 756773
rect 14137 749249 14973 754582
rect 13929 742347 14973 749249
rect 19290 756554 20805 756773
rect 19290 751776 20096 756554
rect 19290 749077 19836 751776
rect 20403 750368 20805 756554
rect 20948 750368 21009 750518
rect 20403 749077 21009 750368
rect 19290 742347 19607 749077
rect 13929 742243 19607 742347
rect 20749 743060 21009 749077
rect 20749 742243 21413 743060
rect 13929 741157 21413 742243
rect 696187 743157 703671 744243
rect 696187 742340 696851 743157
rect 696591 736323 696851 742340
rect 697993 743053 703671 743157
rect 697993 736323 698310 743053
rect 696591 735032 697197 736323
rect 696591 734882 696652 735032
rect 696795 728846 697197 735032
rect 697764 733624 698310 736323
rect 697504 728846 698310 733624
rect 696795 728627 698310 728846
rect 702627 736151 703671 743053
rect 702627 730818 703463 736151
rect 702627 728627 703671 730818
rect 696795 728142 703671 728627
rect 705737 728142 706513 744258
rect 11087 697942 11863 714058
rect 13929 713573 20805 714058
rect 13929 711382 14973 713573
rect 14137 706049 14973 711382
rect 13929 699147 14973 706049
rect 19290 713354 20805 713573
rect 19290 708576 20096 713354
rect 19290 705877 19836 708576
rect 20403 707168 20805 713354
rect 20948 707168 21009 707318
rect 20403 705877 21009 707168
rect 19290 699147 19607 705877
rect 13929 699043 19607 699147
rect 20749 699860 21009 705877
rect 20749 699043 21413 699860
rect 13929 697957 21413 699043
rect 696187 698157 703671 699243
rect 696187 697340 696851 698157
rect 696591 691323 696851 697340
rect 697993 698053 703671 698157
rect 697993 691323 698310 698053
rect 696591 690032 697197 691323
rect 696591 689882 696652 690032
rect 696795 683846 697197 690032
rect 697764 688624 698310 691323
rect 697504 683846 698310 688624
rect 696795 683627 698310 683846
rect 702627 691151 703671 698053
rect 702627 685818 703463 691151
rect 702627 683627 703671 685818
rect 696795 683142 703671 683627
rect 705737 683142 706513 699258
rect 11087 654742 11863 670858
rect 13929 670373 20805 670858
rect 13929 668182 14973 670373
rect 14137 662849 14973 668182
rect 13929 655947 14973 662849
rect 19290 670154 20805 670373
rect 19290 665376 20096 670154
rect 19290 662677 19836 665376
rect 20403 663968 20805 670154
rect 20948 663968 21009 664118
rect 20403 662677 21009 663968
rect 19290 655947 19607 662677
rect 13929 655843 19607 655947
rect 20749 656660 21009 662677
rect 20749 655843 21413 656660
rect 13929 654757 21413 655843
rect 696187 652957 703671 654043
rect 696187 652140 696851 652957
rect 696591 646123 696851 652140
rect 697993 652853 703671 652957
rect 697993 646123 698310 652853
rect 696591 644832 697197 646123
rect 696591 644682 696652 644832
rect 696795 638646 697197 644832
rect 697764 643424 698310 646123
rect 697504 638646 698310 643424
rect 696795 638427 698310 638646
rect 702627 645951 703671 652853
rect 702627 640618 703463 645951
rect 702627 638427 703671 640618
rect 696795 637942 703671 638427
rect 705737 637942 706513 654058
rect 11087 611542 11863 627658
rect 13929 627173 20805 627658
rect 13929 624982 14973 627173
rect 14137 619649 14973 624982
rect 13929 612747 14973 619649
rect 19290 626954 20805 627173
rect 19290 622176 20096 626954
rect 19290 619477 19836 622176
rect 20403 620768 20805 626954
rect 20948 620768 21009 620918
rect 20403 619477 21009 620768
rect 19290 612747 19607 619477
rect 13929 612643 19607 612747
rect 20749 613460 21009 619477
rect 20749 612643 21413 613460
rect 13929 611557 21413 612643
rect 696187 607957 703671 609043
rect 696187 607140 696851 607957
rect 696591 601123 696851 607140
rect 697993 607853 703671 607957
rect 697993 601123 698310 607853
rect 696591 599832 697197 601123
rect 696591 599682 696652 599832
rect 696795 593646 697197 599832
rect 697764 598424 698310 601123
rect 697504 593646 698310 598424
rect 696795 593427 698310 593646
rect 702627 600951 703671 607853
rect 702627 595618 703463 600951
rect 702627 593427 703671 595618
rect 696795 592942 703671 593427
rect 705737 592942 706513 609058
rect 11087 568342 11863 584458
rect 13929 583973 20805 584458
rect 13929 581782 14973 583973
rect 14137 576449 14973 581782
rect 13929 569547 14973 576449
rect 19290 583754 20805 583973
rect 19290 578976 20096 583754
rect 19290 576277 19836 578976
rect 20403 577568 20805 583754
rect 20948 577568 21009 577718
rect 20403 576277 21009 577568
rect 19290 569547 19607 576277
rect 13929 569443 19607 569547
rect 20749 570260 21009 576277
rect 20749 569443 21413 570260
rect 13929 568357 21413 569443
rect 696187 562757 703671 563843
rect 696187 561940 696851 562757
rect 696591 555923 696851 561940
rect 697993 562653 703671 562757
rect 697993 555923 698310 562653
rect 696591 554632 697197 555923
rect 696591 554482 696652 554632
rect 696795 548446 697197 554632
rect 697764 553224 698310 555923
rect 697504 548446 698310 553224
rect 696795 548227 698310 548446
rect 702627 555751 703671 562653
rect 702627 550418 703463 555751
rect 702627 548227 703671 550418
rect 696795 547742 703671 548227
rect 705737 547742 706513 563858
rect 11087 525142 11863 541258
rect 13929 540773 20805 541258
rect 13929 538582 14973 540773
rect 14137 533249 14973 538582
rect 13929 526347 14973 533249
rect 19290 540554 20805 540773
rect 19290 535776 20096 540554
rect 19290 533077 19836 535776
rect 20403 534368 20805 540554
rect 20948 534368 21009 534518
rect 20403 533077 21009 534368
rect 19290 526347 19607 533077
rect 13929 526243 19607 526347
rect 20749 527060 21009 533077
rect 20749 526243 21413 527060
rect 13929 525157 21413 526243
rect 677787 516543 682358 518101
rect 35242 483699 39813 485257
rect 11087 397542 11863 413658
rect 13929 413173 20805 413658
rect 13929 410982 14973 413173
rect 14137 405649 14973 410982
rect 13929 398747 14973 405649
rect 19290 412954 20805 413173
rect 19290 408176 20096 412954
rect 19290 405477 19836 408176
rect 20403 406768 20805 412954
rect 20948 406768 21009 406918
rect 20403 405477 21009 406768
rect 19290 398747 19607 405477
rect 13929 398643 19607 398747
rect 20749 399460 21009 405477
rect 20749 398643 21413 399460
rect 13929 397557 21413 398643
rect 696187 385557 703671 386643
rect 696187 384740 696851 385557
rect 696591 378723 696851 384740
rect 697993 385453 703671 385557
rect 697993 378723 698310 385453
rect 696591 377432 697197 378723
rect 696591 377282 696652 377432
rect 11087 354342 11863 370458
rect 13929 369973 20805 370458
rect 13929 367782 14973 369973
rect 14137 362449 14973 367782
rect 13929 355547 14973 362449
rect 19290 369754 20805 369973
rect 19290 364976 20096 369754
rect 19290 362277 19836 364976
rect 20403 363568 20805 369754
rect 696795 371246 697197 377432
rect 697764 376024 698310 378723
rect 697504 371246 698310 376024
rect 696795 371027 698310 371246
rect 702627 378551 703671 385453
rect 702627 373218 703463 378551
rect 702627 371027 703671 373218
rect 696795 370542 703671 371027
rect 705737 370542 706513 386658
rect 20948 363568 21009 363718
rect 20403 362277 21009 363568
rect 19290 355547 19607 362277
rect 13929 355443 19607 355547
rect 20749 356260 21009 362277
rect 20749 355443 21413 356260
rect 13929 354357 21413 355443
rect 696187 340357 703671 341443
rect 696187 339540 696851 340357
rect 696591 333523 696851 339540
rect 697993 340253 703671 340357
rect 697993 333523 698310 340253
rect 696591 332232 697197 333523
rect 696591 332082 696652 332232
rect 11087 311142 11863 327258
rect 13929 326773 20805 327258
rect 13929 324582 14973 326773
rect 14137 319249 14973 324582
rect 13929 312347 14973 319249
rect 19290 326554 20805 326773
rect 19290 321776 20096 326554
rect 19290 319077 19836 321776
rect 20403 320368 20805 326554
rect 696795 326046 697197 332232
rect 697764 330824 698310 333523
rect 697504 326046 698310 330824
rect 696795 325827 698310 326046
rect 702627 333351 703671 340253
rect 702627 328018 703463 333351
rect 702627 325827 703671 328018
rect 696795 325342 703671 325827
rect 705737 325342 706513 341458
rect 20948 320368 21009 320518
rect 20403 319077 21009 320368
rect 19290 312347 19607 319077
rect 13929 312243 19607 312347
rect 20749 313060 21009 319077
rect 20749 312243 21413 313060
rect 13929 311157 21413 312243
rect 11087 267942 11863 284058
rect 13929 283573 20805 284058
rect 13929 281382 14973 283573
rect 14137 276049 14973 281382
rect 13929 269147 14973 276049
rect 19290 283354 20805 283573
rect 19290 278576 20096 283354
rect 19290 275877 19836 278576
rect 20403 277168 20805 283354
rect 20948 277168 21009 277318
rect 20403 275877 21009 277168
rect 19290 269147 19607 275877
rect 13929 269043 19607 269147
rect 20749 269860 21009 275877
rect 20749 269043 21413 269860
rect 13929 267957 21413 269043
rect 696187 295357 703671 296443
rect 696187 294540 696851 295357
rect 696591 288523 696851 294540
rect 697993 295253 703671 295357
rect 697993 288523 698310 295253
rect 696591 287232 697197 288523
rect 696591 287082 696652 287232
rect 696795 281046 697197 287232
rect 697764 285824 698310 288523
rect 697504 281046 698310 285824
rect 696795 280827 698310 281046
rect 702627 288351 703671 295253
rect 702627 283018 703463 288351
rect 702627 280827 703671 283018
rect 696795 280342 703671 280827
rect 705737 280342 706513 296458
rect 11087 224742 11863 240858
rect 13929 240373 20805 240858
rect 13929 238182 14973 240373
rect 14137 232849 14973 238182
rect 13929 225947 14973 232849
rect 19290 240154 20805 240373
rect 19290 235376 20096 240154
rect 19290 232677 19836 235376
rect 20403 233968 20805 240154
rect 20948 233968 21009 234118
rect 20403 232677 21009 233968
rect 19290 225947 19607 232677
rect 13929 225843 19607 225947
rect 20749 226660 21009 232677
rect 20749 225843 21413 226660
rect 13929 224757 21413 225843
rect 696187 250357 703671 251443
rect 696187 249540 696851 250357
rect 696591 243523 696851 249540
rect 697993 250253 703671 250357
rect 697993 243523 698310 250253
rect 696591 242232 697197 243523
rect 696591 242082 696652 242232
rect 696795 236046 697197 242232
rect 697764 240824 698310 243523
rect 697504 236046 698310 240824
rect 696795 235827 698310 236046
rect 702627 243351 703671 250253
rect 702627 238018 703463 243351
rect 702627 235827 703671 238018
rect 696795 235342 703671 235827
rect 705737 235342 706513 251458
rect 11087 181542 11863 197658
rect 13929 197173 20805 197658
rect 13929 194982 14973 197173
rect 14137 189649 14973 194982
rect 13929 182747 14973 189649
rect 19290 196954 20805 197173
rect 19290 192176 20096 196954
rect 19290 189477 19836 192176
rect 20403 190768 20805 196954
rect 20948 190768 21009 190918
rect 20403 189477 21009 190768
rect 19290 182747 19607 189477
rect 13929 182643 19607 182747
rect 20749 183460 21009 189477
rect 20749 182643 21413 183460
rect 13929 181557 21413 182643
rect 696187 205157 703671 206243
rect 696187 204340 696851 205157
rect 696591 198323 696851 204340
rect 697993 205053 703671 205157
rect 697993 198323 698310 205053
rect 696591 197032 697197 198323
rect 696591 196882 696652 197032
rect 696795 190846 697197 197032
rect 697764 195624 698310 198323
rect 697504 190846 698310 195624
rect 696795 190627 698310 190846
rect 702627 198151 703671 205053
rect 702627 192818 703463 198151
rect 702627 190627 703671 192818
rect 696795 190142 703671 190627
rect 705737 190142 706513 206258
rect 696187 160157 703671 161243
rect 696187 159340 696851 160157
rect 696591 153323 696851 159340
rect 697993 160053 703671 160157
rect 697993 153323 698310 160053
rect 696591 152032 697197 153323
rect 696591 151882 696652 152032
rect 696795 145846 697197 152032
rect 697764 150624 698310 153323
rect 697504 145846 698310 150624
rect 696795 145627 698310 145846
rect 702627 153151 703671 160053
rect 702627 147818 703463 153151
rect 702627 145627 703671 147818
rect 696795 145142 703671 145627
rect 705737 145142 706513 161258
rect 35242 110899 39813 112457
rect 696187 114957 703671 116043
rect 696187 114140 696851 114957
rect 696591 108123 696851 114140
rect 697993 114853 703671 114957
rect 697993 108123 698310 114853
rect 696591 106832 697197 108123
rect 696591 106682 696652 106832
rect 696795 100646 697197 106832
rect 697764 105424 698310 108123
rect 697504 100646 698310 105424
rect 696795 100427 698310 100646
rect 702627 107951 703671 114853
rect 702627 102618 703463 107951
rect 702627 100427 703671 102618
rect 696795 99942 703671 100427
rect 705737 99942 706513 116058
rect 635543 35242 637101 39813
rect 200540 21009 202443 21413
rect 193082 20948 202443 21009
rect 309140 21009 311043 21413
rect 301682 20948 311043 21009
rect 363940 21009 365843 21413
rect 356482 20948 365843 21009
rect 418740 21009 420643 21413
rect 411282 20948 420643 21009
rect 473540 21009 475443 21413
rect 466082 20948 475443 21009
rect 528340 21009 530243 21413
rect 520882 20948 530243 21009
rect 193232 20805 202443 20948
rect 301832 20805 311043 20948
rect 356632 20805 365843 20948
rect 411432 20805 420643 20948
rect 466232 20805 475443 20948
rect 521032 20805 530243 20948
rect 186342 20749 202443 20805
rect 135906 20653 147626 20654
rect 132574 20401 147626 20653
rect 132574 20154 133214 20401
rect 135906 20154 147626 20401
rect 132574 19495 147626 20154
rect 132574 15173 132888 19495
rect 147313 15173 147626 19495
rect 132574 14137 147626 15173
rect 132574 13929 135218 14137
rect 139250 13929 147626 14137
rect 186342 20403 194523 20749
rect 186342 20096 187046 20403
rect 186342 19836 191824 20096
rect 186342 19607 194523 19836
rect 201357 19607 202443 20749
rect 186342 19290 202443 19607
rect 186342 14973 186827 19290
rect 201253 14973 202443 19290
rect 186342 14137 202443 14973
rect 186342 13929 189018 14137
rect 194351 13929 202443 14137
rect 294942 20749 311043 20805
rect 294942 20403 303123 20749
rect 294942 20096 295646 20403
rect 294942 19836 300424 20096
rect 294942 19607 303123 19836
rect 309957 19607 311043 20749
rect 294942 19290 311043 19607
rect 294942 14973 295427 19290
rect 309853 14973 311043 19290
rect 294942 14137 311043 14973
rect 294942 13929 297618 14137
rect 302951 13929 311043 14137
rect 349742 20749 365843 20805
rect 349742 20403 357923 20749
rect 349742 20096 350446 20403
rect 349742 19836 355224 20096
rect 349742 19607 357923 19836
rect 364757 19607 365843 20749
rect 349742 19290 365843 19607
rect 349742 14973 350227 19290
rect 364653 14973 365843 19290
rect 349742 14137 365843 14973
rect 349742 13929 352418 14137
rect 357751 13929 365843 14137
rect 404542 20749 420643 20805
rect 404542 20403 412723 20749
rect 404542 20096 405246 20403
rect 404542 19836 410024 20096
rect 404542 19607 412723 19836
rect 419557 19607 420643 20749
rect 404542 19290 420643 19607
rect 404542 14973 405027 19290
rect 419453 14973 420643 19290
rect 404542 14137 420643 14973
rect 404542 13929 407218 14137
rect 412551 13929 420643 14137
rect 459342 20749 475443 20805
rect 459342 20403 467523 20749
rect 459342 20096 460046 20403
rect 459342 19836 464824 20096
rect 459342 19607 467523 19836
rect 474357 19607 475443 20749
rect 459342 19290 475443 19607
rect 459342 14973 459827 19290
rect 474253 14973 475443 19290
rect 459342 14137 475443 14973
rect 459342 13929 462018 14137
rect 467351 13929 475443 14137
rect 514142 20749 530243 20805
rect 514142 20403 522323 20749
rect 514142 20096 514846 20403
rect 514142 19836 519624 20096
rect 514142 19607 522323 19836
rect 529157 19607 530243 20749
rect 514142 19290 530243 19607
rect 514142 14973 514627 19290
rect 529053 14973 530243 19290
rect 514142 14137 530243 14973
rect 514142 13929 516818 14137
rect 522151 13929 530243 14137
rect 132542 11087 147658 11863
rect 186342 11087 202458 11863
rect 294942 11087 311058 11863
rect 349742 11087 365858 11863
rect 404542 11087 420658 11863
rect 459342 11087 475458 11863
rect 514142 11087 530258 11863
<< obsli1 >>
rect 76781 1007253 90609 1033820
rect 128181 1007253 142009 1033820
rect 179581 1007253 193409 1033820
rect 230522 998007 244971 1037539
rect 282122 998007 296571 1037539
rect 333614 998007 347955 1037539
rect 384381 1007253 398209 1033820
rect 473381 1007253 487209 1033820
rect 524781 1007253 538609 1033820
rect 575814 998007 590155 1037539
rect 626581 1007253 640409 1033820
rect 230522 997813 232631 998007
rect 232807 997984 233009 998007
rect 244346 997984 244536 998007
rect 232807 997794 244536 997984
rect 282122 997813 284231 998007
rect 284407 997984 284609 998007
rect 295946 997984 296136 998007
rect 284407 997794 296136 997984
rect 335813 997978 336009 998007
rect 347352 997978 347530 998007
rect 335813 997800 347530 997978
rect 578013 997978 578209 998007
rect 589552 997978 589730 998007
rect 578013 997800 589730 997978
rect 3780 954781 30347 968609
rect 677813 965369 717539 967478
rect 678007 965193 717539 965369
rect 677794 964991 717539 965193
rect 677794 953654 677984 964991
rect 678007 953654 717539 964991
rect 677794 953464 717539 953654
rect 678007 953029 717539 953464
rect 44 912048 39396 926951
rect 678204 907649 717556 922552
rect 61 883936 39593 884371
rect 61 883746 39806 883936
rect 61 872409 39593 883746
rect 39616 872409 39806 883746
rect 696779 878417 703644 878423
rect 703855 878417 705630 878423
rect 678799 878400 679399 878417
rect 689044 878400 693721 878417
rect 695363 878400 696014 878417
rect 696213 878400 703645 878417
rect 703799 878400 705630 878417
rect 705763 878400 706487 878432
rect 706631 878417 711618 878423
rect 706631 878400 713329 878417
rect 61 872207 39806 872409
rect 61 872031 39593 872207
rect 61 869922 39787 872031
rect 677646 862400 717541 878400
rect 681497 862376 682603 862400
rect 683623 862376 684745 862400
rect 687850 862383 696516 862400
rect 696821 862368 703645 862400
rect 703799 862383 705611 862400
rect 705763 862368 706487 862400
rect 706643 862379 713329 862400
rect 61 841730 39593 842155
rect 61 841552 39800 841730
rect 61 830209 39593 841552
rect 39622 830209 39800 841552
rect 677813 831169 717539 833278
rect 678007 830993 717539 831169
rect 61 830013 39800 830209
rect 677794 830791 717539 830993
rect 61 827814 39593 830013
rect 677794 819454 677984 830791
rect 678007 819454 717539 830791
rect 677794 819264 717539 819454
rect 678007 818829 717539 819264
rect 4271 800400 10957 800421
rect 11113 800400 11837 800432
rect 11989 800400 13801 800417
rect 13955 800400 20779 800432
rect 21084 800400 29750 800417
rect 32855 800400 33977 800424
rect 34997 800400 36103 800424
rect 59 784400 39954 800400
rect 696779 789217 703644 789223
rect 703855 789217 705630 789223
rect 678799 789200 679399 789217
rect 689044 789200 693721 789217
rect 695363 789200 696014 789217
rect 696213 789200 703645 789217
rect 703799 789200 705630 789217
rect 705763 789200 706487 789232
rect 706631 789217 711618 789223
rect 706631 789200 713329 789217
rect 4271 784383 10969 784400
rect 5982 784377 10969 784383
rect 11113 784368 11837 784400
rect 11970 784383 13801 784400
rect 13955 784383 21387 784400
rect 21586 784383 22237 784400
rect 23879 784383 28556 784400
rect 38201 784383 38801 784400
rect 11970 784377 13745 784383
rect 13956 784377 20821 784383
rect 677646 773200 717541 789200
rect 681497 773176 682603 773200
rect 683623 773176 684745 773200
rect 687850 773183 696516 773200
rect 696821 773168 703645 773200
rect 703799 773183 705611 773200
rect 705763 773168 706487 773200
rect 706643 773179 713329 773200
rect 4271 757200 10957 757221
rect 11113 757200 11837 757232
rect 11989 757200 13801 757217
rect 13955 757200 20779 757232
rect 21084 757200 29750 757217
rect 32855 757200 33977 757224
rect 34997 757200 36103 757224
rect 59 741200 39954 757200
rect 696779 744217 703644 744223
rect 703855 744217 705630 744223
rect 678799 744200 679399 744217
rect 689044 744200 693721 744217
rect 695363 744200 696014 744217
rect 696213 744200 703645 744217
rect 703799 744200 705630 744217
rect 705763 744200 706487 744232
rect 706631 744217 711618 744223
rect 706631 744200 713329 744217
rect 4271 741183 10969 741200
rect 5982 741177 10969 741183
rect 11113 741168 11837 741200
rect 11970 741183 13801 741200
rect 13955 741183 21387 741200
rect 21586 741183 22237 741200
rect 23879 741183 28556 741200
rect 38201 741183 38801 741200
rect 11970 741177 13745 741183
rect 13956 741177 20821 741183
rect 677646 728200 717541 744200
rect 681497 728176 682603 728200
rect 683623 728176 684745 728200
rect 687850 728183 696516 728200
rect 696821 728168 703645 728200
rect 703799 728183 705611 728200
rect 705763 728168 706487 728200
rect 706643 728179 713329 728200
rect 4271 714000 10957 714021
rect 11113 714000 11837 714032
rect 11989 714000 13801 714017
rect 13955 714000 20779 714032
rect 21084 714000 29750 714017
rect 32855 714000 33977 714024
rect 34997 714000 36103 714024
rect 59 698000 39954 714000
rect 696779 699217 703644 699223
rect 703855 699217 705630 699223
rect 678799 699200 679399 699217
rect 689044 699200 693721 699217
rect 695363 699200 696014 699217
rect 696213 699200 703645 699217
rect 703799 699200 705630 699217
rect 705763 699200 706487 699232
rect 706631 699217 711618 699223
rect 706631 699200 713329 699217
rect 4271 697983 10969 698000
rect 5982 697977 10969 697983
rect 11113 697968 11837 698000
rect 11970 697983 13801 698000
rect 13955 697983 21387 698000
rect 21586 697983 22237 698000
rect 23879 697983 28556 698000
rect 38201 697983 38801 698000
rect 11970 697977 13745 697983
rect 13956 697977 20821 697983
rect 677646 683200 717541 699200
rect 681497 683176 682603 683200
rect 683623 683176 684745 683200
rect 687850 683183 696516 683200
rect 696821 683168 703645 683200
rect 703799 683183 705611 683200
rect 705763 683168 706487 683200
rect 706643 683179 713329 683200
rect 4271 670800 10957 670821
rect 11113 670800 11837 670832
rect 11989 670800 13801 670817
rect 13955 670800 20779 670832
rect 21084 670800 29750 670817
rect 32855 670800 33977 670824
rect 34997 670800 36103 670824
rect 59 654800 39954 670800
rect 4271 654783 10969 654800
rect 5982 654777 10969 654783
rect 11113 654768 11837 654800
rect 11970 654783 13801 654800
rect 13955 654783 21387 654800
rect 21586 654783 22237 654800
rect 23879 654783 28556 654800
rect 38201 654783 38801 654800
rect 11970 654777 13745 654783
rect 13956 654777 20821 654783
rect 696779 654017 703644 654023
rect 703855 654017 705630 654023
rect 678799 654000 679399 654017
rect 689044 654000 693721 654017
rect 695363 654000 696014 654017
rect 696213 654000 703645 654017
rect 703799 654000 705630 654017
rect 705763 654000 706487 654032
rect 706631 654017 711618 654023
rect 706631 654000 713329 654017
rect 677646 638000 717541 654000
rect 681497 637976 682603 638000
rect 683623 637976 684745 638000
rect 687850 637983 696516 638000
rect 696821 637968 703645 638000
rect 703799 637983 705611 638000
rect 705763 637968 706487 638000
rect 706643 637979 713329 638000
rect 4271 627600 10957 627621
rect 11113 627600 11837 627632
rect 11989 627600 13801 627617
rect 13955 627600 20779 627632
rect 21084 627600 29750 627617
rect 32855 627600 33977 627624
rect 34997 627600 36103 627624
rect 59 611600 39954 627600
rect 4271 611583 10969 611600
rect 5982 611577 10969 611583
rect 11113 611568 11837 611600
rect 11970 611583 13801 611600
rect 13955 611583 21387 611600
rect 21586 611583 22237 611600
rect 23879 611583 28556 611600
rect 38201 611583 38801 611600
rect 11970 611577 13745 611583
rect 13956 611577 20821 611583
rect 696779 609017 703644 609023
rect 703855 609017 705630 609023
rect 678799 609000 679399 609017
rect 689044 609000 693721 609017
rect 695363 609000 696014 609017
rect 696213 609000 703645 609017
rect 703799 609000 705630 609017
rect 705763 609000 706487 609032
rect 706631 609017 711618 609023
rect 706631 609000 713329 609017
rect 677646 593000 717541 609000
rect 681497 592976 682603 593000
rect 683623 592976 684745 593000
rect 687850 592983 696516 593000
rect 696821 592968 703645 593000
rect 703799 592983 705611 593000
rect 705763 592968 706487 593000
rect 706643 592979 713329 593000
rect 4271 584400 10957 584421
rect 11113 584400 11837 584432
rect 11989 584400 13801 584417
rect 13955 584400 20779 584432
rect 21084 584400 29750 584417
rect 32855 584400 33977 584424
rect 34997 584400 36103 584424
rect 59 568400 39954 584400
rect 4271 568383 10969 568400
rect 5982 568377 10969 568383
rect 11113 568368 11837 568400
rect 11970 568383 13801 568400
rect 13955 568383 21387 568400
rect 21586 568383 22237 568400
rect 23879 568383 28556 568400
rect 38201 568383 38801 568400
rect 11970 568377 13745 568383
rect 13956 568377 20821 568383
rect 696779 563817 703644 563823
rect 703855 563817 705630 563823
rect 678799 563800 679399 563817
rect 689044 563800 693721 563817
rect 695363 563800 696014 563817
rect 696213 563800 703645 563817
rect 703799 563800 705630 563817
rect 705763 563800 706487 563832
rect 706631 563817 711618 563823
rect 706631 563800 713329 563817
rect 677646 547800 717541 563800
rect 681497 547776 682603 547800
rect 683623 547776 684745 547800
rect 687850 547783 696516 547800
rect 696821 547768 703645 547800
rect 703799 547783 705611 547800
rect 705763 547768 706487 547800
rect 706643 547779 713329 547800
rect 4271 541200 10957 541221
rect 11113 541200 11837 541232
rect 11989 541200 13801 541217
rect 13955 541200 20779 541232
rect 21084 541200 29750 541217
rect 32855 541200 33977 541224
rect 34997 541200 36103 541224
rect 59 525200 39954 541200
rect 4271 525183 10969 525200
rect 5982 525177 10969 525183
rect 11113 525168 11837 525200
rect 11970 525183 13801 525200
rect 13955 525183 21387 525200
rect 21586 525183 22237 525200
rect 23879 525183 28556 525200
rect 38201 525183 38801 525200
rect 11970 525177 13745 525183
rect 13956 525177 20821 525183
rect 677813 516569 717539 518678
rect 678007 516393 717539 516569
rect 677794 516191 717539 516393
rect 677794 504854 677984 516191
rect 678007 504854 717539 516191
rect 677794 504664 717539 504854
rect 678007 504229 717539 504664
rect 61 497136 39593 497571
rect 61 496946 39806 497136
rect 61 485609 39593 496946
rect 39616 485609 39806 496946
rect 61 485407 39806 485609
rect 61 485231 39593 485407
rect 61 483122 39787 485231
rect 678204 459849 717556 474752
rect 44 440848 39396 455751
rect 678007 428187 717539 430386
rect 677800 427991 717539 428187
rect 677800 416648 677978 427991
rect 678007 416648 717539 427991
rect 677800 416470 717539 416648
rect 678007 416045 717539 416470
rect 4271 413600 10957 413621
rect 11113 413600 11837 413632
rect 11989 413600 13801 413617
rect 13955 413600 20779 413632
rect 21084 413600 29750 413617
rect 32855 413600 33977 413624
rect 34997 413600 36103 413624
rect 59 397600 39954 413600
rect 4271 397583 10969 397600
rect 5982 397577 10969 397583
rect 11113 397568 11837 397600
rect 11970 397583 13801 397600
rect 13955 397583 21387 397600
rect 21586 397583 22237 397600
rect 23879 397583 28556 397600
rect 38201 397583 38801 397600
rect 11970 397577 13745 397583
rect 13956 397577 20821 397583
rect 696779 386617 703644 386623
rect 703855 386617 705630 386623
rect 678799 386600 679399 386617
rect 689044 386600 693721 386617
rect 695363 386600 696014 386617
rect 696213 386600 703645 386617
rect 703799 386600 705630 386617
rect 705763 386600 706487 386632
rect 706631 386617 711618 386623
rect 706631 386600 713329 386617
rect 677646 370600 717541 386600
rect 681497 370576 682603 370600
rect 683623 370576 684745 370600
rect 687850 370583 696516 370600
rect 696821 370568 703645 370600
rect 703799 370583 705611 370600
rect 705763 370568 706487 370600
rect 706643 370579 713329 370600
rect 4271 370400 10957 370421
rect 11113 370400 11837 370432
rect 11989 370400 13801 370417
rect 13955 370400 20779 370432
rect 21084 370400 29750 370417
rect 32855 370400 33977 370424
rect 34997 370400 36103 370424
rect 59 354400 39954 370400
rect 4271 354383 10969 354400
rect 5982 354377 10969 354383
rect 11113 354368 11837 354400
rect 11970 354383 13801 354400
rect 13955 354383 21387 354400
rect 21586 354383 22237 354400
rect 23879 354383 28556 354400
rect 38201 354383 38801 354400
rect 11970 354377 13745 354383
rect 13956 354377 20821 354383
rect 696779 341417 703644 341423
rect 703855 341417 705630 341423
rect 678799 341400 679399 341417
rect 689044 341400 693721 341417
rect 695363 341400 696014 341417
rect 696213 341400 703645 341417
rect 703799 341400 705630 341417
rect 705763 341400 706487 341432
rect 706631 341417 711618 341423
rect 706631 341400 713329 341417
rect 4271 327200 10957 327221
rect 11113 327200 11837 327232
rect 11989 327200 13801 327217
rect 13955 327200 20779 327232
rect 21084 327200 29750 327217
rect 32855 327200 33977 327224
rect 34997 327200 36103 327224
rect 59 311200 39954 327200
rect 677646 325400 717541 341400
rect 681497 325376 682603 325400
rect 683623 325376 684745 325400
rect 687850 325383 696516 325400
rect 696821 325368 703645 325400
rect 703799 325383 705611 325400
rect 705763 325368 706487 325400
rect 706643 325379 713329 325400
rect 4271 311183 10969 311200
rect 5982 311177 10969 311183
rect 11113 311168 11837 311200
rect 11970 311183 13801 311200
rect 13955 311183 21387 311200
rect 21586 311183 22237 311200
rect 23879 311183 28556 311200
rect 38201 311183 38801 311200
rect 11970 311177 13745 311183
rect 13956 311177 20821 311183
rect 696779 296417 703644 296423
rect 703855 296417 705630 296423
rect 678799 296400 679399 296417
rect 689044 296400 693721 296417
rect 695363 296400 696014 296417
rect 696213 296400 703645 296417
rect 703799 296400 705630 296417
rect 705763 296400 706487 296432
rect 706631 296417 711618 296423
rect 706631 296400 713329 296417
rect 4271 284000 10957 284021
rect 11113 284000 11837 284032
rect 11989 284000 13801 284017
rect 13955 284000 20779 284032
rect 21084 284000 29750 284017
rect 32855 284000 33977 284024
rect 34997 284000 36103 284024
rect 59 268000 39954 284000
rect 677646 280400 717541 296400
rect 681497 280376 682603 280400
rect 683623 280376 684745 280400
rect 687850 280383 696516 280400
rect 696821 280368 703645 280400
rect 703799 280383 705611 280400
rect 705763 280368 706487 280400
rect 706643 280379 713329 280400
rect 4271 267983 10969 268000
rect 5982 267977 10969 267983
rect 11113 267968 11837 268000
rect 11970 267983 13801 268000
rect 13955 267983 21387 268000
rect 21586 267983 22237 268000
rect 23879 267983 28556 268000
rect 38201 267983 38801 268000
rect 11970 267977 13745 267983
rect 13956 267977 20821 267983
rect 696779 251417 703644 251423
rect 703855 251417 705630 251423
rect 678799 251400 679399 251417
rect 689044 251400 693721 251417
rect 695363 251400 696014 251417
rect 696213 251400 703645 251417
rect 703799 251400 705630 251417
rect 705763 251400 706487 251432
rect 706631 251417 711618 251423
rect 706631 251400 713329 251417
rect 4271 240800 10957 240821
rect 11113 240800 11837 240832
rect 11989 240800 13801 240817
rect 13955 240800 20779 240832
rect 21084 240800 29750 240817
rect 32855 240800 33977 240824
rect 34997 240800 36103 240824
rect 59 224800 39954 240800
rect 677646 235400 717541 251400
rect 681497 235376 682603 235400
rect 683623 235376 684745 235400
rect 687850 235383 696516 235400
rect 696821 235368 703645 235400
rect 703799 235383 705611 235400
rect 705763 235368 706487 235400
rect 706643 235379 713329 235400
rect 4271 224783 10969 224800
rect 5982 224777 10969 224783
rect 11113 224768 11837 224800
rect 11970 224783 13801 224800
rect 13955 224783 21387 224800
rect 21586 224783 22237 224800
rect 23879 224783 28556 224800
rect 38201 224783 38801 224800
rect 11970 224777 13745 224783
rect 13956 224777 20821 224783
rect 696779 206217 703644 206223
rect 703855 206217 705630 206223
rect 678799 206200 679399 206217
rect 689044 206200 693721 206217
rect 695363 206200 696014 206217
rect 696213 206200 703645 206217
rect 703799 206200 705630 206217
rect 705763 206200 706487 206232
rect 706631 206217 711618 206223
rect 706631 206200 713329 206217
rect 4271 197600 10957 197621
rect 11113 197600 11837 197632
rect 11989 197600 13801 197617
rect 13955 197600 20779 197632
rect 21084 197600 29750 197617
rect 32855 197600 33977 197624
rect 34997 197600 36103 197624
rect 59 181600 39954 197600
rect 677646 190200 717541 206200
rect 681497 190176 682603 190200
rect 683623 190176 684745 190200
rect 687850 190183 696516 190200
rect 696821 190168 703645 190200
rect 703799 190183 705611 190200
rect 705763 190168 706487 190200
rect 706643 190179 713329 190200
rect 4271 181583 10969 181600
rect 5982 181577 10969 181583
rect 11113 181568 11837 181600
rect 11970 181583 13801 181600
rect 13955 181583 21387 181600
rect 21586 181583 22237 181600
rect 23879 181583 28556 181600
rect 38201 181583 38801 181600
rect 11970 181577 13745 181583
rect 13956 181577 20821 181583
rect 696779 161217 703644 161223
rect 703855 161217 705630 161223
rect 678799 161200 679399 161217
rect 689044 161200 693721 161217
rect 695363 161200 696014 161217
rect 696213 161200 703645 161217
rect 703799 161200 705630 161217
rect 705763 161200 706487 161232
rect 706631 161217 711618 161223
rect 706631 161200 713329 161217
rect 677646 145200 717541 161200
rect 681497 145176 682603 145200
rect 683623 145176 684745 145200
rect 687850 145183 696516 145200
rect 696821 145168 703645 145200
rect 703799 145183 705611 145200
rect 705763 145168 706487 145200
rect 706643 145179 713329 145200
rect 61 124336 39593 124771
rect 61 124146 39806 124336
rect 61 112809 39593 124146
rect 39616 112809 39806 124146
rect 696779 116017 703644 116023
rect 703855 116017 705630 116023
rect 678799 116000 679399 116017
rect 689044 116000 693721 116017
rect 695363 116000 696014 116017
rect 696213 116000 703645 116017
rect 703799 116000 705630 116017
rect 705763 116000 706487 116032
rect 706631 116017 711618 116023
rect 706631 116000 713329 116017
rect 61 112607 39806 112809
rect 61 112431 39593 112607
rect 61 110322 39787 112431
rect 677646 100000 717541 116000
rect 681497 99976 682603 100000
rect 683623 99976 684745 100000
rect 687850 99983 696516 100000
rect 696821 99968 703645 100000
rect 703799 99983 705611 100000
rect 705763 99968 706487 100000
rect 706643 99979 713329 100000
rect 44 68048 39396 82951
rect 79670 39622 91387 39800
rect 79670 39593 79848 39622
rect 91191 39593 91387 39622
rect 79245 61 93586 39593
rect 132600 19721 147600 39963
rect 186400 38801 202400 39954
rect 186400 38201 202417 38801
rect 186400 36103 202400 38201
rect 186376 34997 202400 36103
rect 186400 33977 202400 34997
rect 186376 32855 202400 33977
rect 186400 29750 202400 32855
rect 186383 28556 202400 29750
rect 186383 23879 202417 28556
rect 186383 22237 202400 23879
rect 186383 21586 202417 22237
rect 186383 21387 202400 21586
rect 186383 21084 202417 21387
rect 186400 20821 202417 21084
rect 186400 20779 202423 20821
rect 132600 13955 147653 19721
rect 186368 13956 202423 20779
rect 186368 13955 202417 13956
rect 132600 11837 147600 13955
rect 186400 13801 202400 13955
rect 186383 13745 202417 13801
rect 186383 11989 202423 13745
rect 186400 11970 202423 11989
rect 186400 11837 202400 11970
rect 132568 11113 147632 11837
rect 186368 11113 202432 11837
rect 132600 156 147600 11113
rect 186400 10969 202400 11113
rect 186400 10957 202423 10969
rect 186379 5982 202423 10957
rect 186379 4271 202417 5982
rect 186400 59 202400 4271
rect 241249 44 256152 39396
rect 295000 38801 311000 39954
rect 349800 38801 365800 39954
rect 404600 38801 420600 39954
rect 459400 38801 475400 39954
rect 514200 38801 530200 39954
rect 569870 39622 581587 39800
rect 569870 39593 570048 39622
rect 581391 39593 581587 39622
rect 623664 39616 635393 39806
rect 623664 39593 623854 39616
rect 635191 39593 635393 39616
rect 635569 39593 637678 39787
rect 295000 38201 311017 38801
rect 349800 38201 365817 38801
rect 404600 38201 420617 38801
rect 459400 38201 475417 38801
rect 514200 38201 530217 38801
rect 295000 36103 311000 38201
rect 349800 36103 365800 38201
rect 404600 36103 420600 38201
rect 459400 36103 475400 38201
rect 514200 36103 530200 38201
rect 294976 34997 311000 36103
rect 349776 34997 365800 36103
rect 404576 34997 420600 36103
rect 459376 34997 475400 36103
rect 514176 34997 530200 36103
rect 295000 33977 311000 34997
rect 349800 33977 365800 34997
rect 404600 33977 420600 34997
rect 459400 33977 475400 34997
rect 514200 33977 530200 34997
rect 294976 32855 311000 33977
rect 349776 32855 365800 33977
rect 404576 32855 420600 33977
rect 459376 32855 475400 33977
rect 514176 32855 530200 33977
rect 295000 29750 311000 32855
rect 349800 29750 365800 32855
rect 404600 29750 420600 32855
rect 459400 29750 475400 32855
rect 514200 29750 530200 32855
rect 294983 28556 311000 29750
rect 349783 28556 365800 29750
rect 404583 28556 420600 29750
rect 459383 28556 475400 29750
rect 514183 28556 530200 29750
rect 294983 23879 311017 28556
rect 349783 23879 365817 28556
rect 404583 23879 420617 28556
rect 459383 23879 475417 28556
rect 514183 23879 530217 28556
rect 294983 22237 311000 23879
rect 349783 22237 365800 23879
rect 404583 22237 420600 23879
rect 459383 22237 475400 23879
rect 514183 22237 530200 23879
rect 294983 21586 311017 22237
rect 349783 21586 365817 22237
rect 404583 21586 420617 22237
rect 459383 21586 475417 22237
rect 514183 21586 530217 22237
rect 294983 21387 311000 21586
rect 349783 21387 365800 21586
rect 404583 21387 420600 21586
rect 459383 21387 475400 21586
rect 514183 21387 530200 21586
rect 294983 21084 311017 21387
rect 349783 21084 365817 21387
rect 404583 21084 420617 21387
rect 459383 21084 475417 21387
rect 514183 21084 530217 21387
rect 295000 20821 311017 21084
rect 349800 20821 365817 21084
rect 404600 20821 420617 21084
rect 459400 20821 475417 21084
rect 514200 20821 530217 21084
rect 295000 20779 311023 20821
rect 349800 20779 365823 20821
rect 404600 20779 420623 20821
rect 459400 20779 475423 20821
rect 514200 20779 530223 20821
rect 294968 13956 311023 20779
rect 349768 13956 365823 20779
rect 404568 13956 420623 20779
rect 459368 13956 475423 20779
rect 514168 13956 530223 20779
rect 294968 13955 311017 13956
rect 349768 13955 365817 13956
rect 404568 13955 420617 13956
rect 459368 13955 475417 13956
rect 514168 13955 530217 13956
rect 295000 13801 311000 13955
rect 349800 13801 365800 13955
rect 404600 13801 420600 13955
rect 459400 13801 475400 13955
rect 514200 13801 530200 13955
rect 294983 13745 311017 13801
rect 349783 13745 365817 13801
rect 404583 13745 420617 13801
rect 459383 13745 475417 13801
rect 514183 13745 530217 13801
rect 294983 11989 311023 13745
rect 349783 11989 365823 13745
rect 404583 11989 420623 13745
rect 459383 11989 475423 13745
rect 514183 11989 530223 13745
rect 295000 11970 311023 11989
rect 349800 11970 365823 11989
rect 404600 11970 420623 11989
rect 459400 11970 475423 11989
rect 514200 11970 530223 11989
rect 295000 11837 311000 11970
rect 349800 11837 365800 11970
rect 404600 11837 420600 11970
rect 459400 11837 475400 11970
rect 514200 11837 530200 11970
rect 294968 11113 311032 11837
rect 349768 11113 365832 11837
rect 404568 11113 420632 11837
rect 459368 11113 475432 11837
rect 514168 11113 530232 11837
rect 295000 10969 311000 11113
rect 349800 10969 365800 11113
rect 404600 10969 420600 11113
rect 459400 10969 475400 11113
rect 514200 10969 530200 11113
rect 295000 10957 311023 10969
rect 349800 10957 365823 10969
rect 404600 10957 420623 10969
rect 459400 10957 475423 10969
rect 514200 10957 530223 10969
rect 294979 5982 311023 10957
rect 349779 5982 365823 10957
rect 404579 5982 420623 10957
rect 459379 5982 475423 10957
rect 514179 5982 530223 10957
rect 294979 4271 311017 5982
rect 349779 4271 365817 5982
rect 404579 4271 420617 5982
rect 459379 4271 475417 5982
rect 514179 4271 530217 5982
rect 295000 59 311000 4271
rect 349800 59 365800 4271
rect 404600 59 420600 4271
rect 459400 59 475400 4271
rect 514200 59 530200 4271
rect 569445 61 583786 39593
rect 623229 61 637678 39593
<< metal1 >>
rect 673730 870816 673736 870868
rect 673788 870856 673794 870868
rect 675386 870856 675392 870868
rect 673788 870828 675392 870856
rect 673788 870816 673794 870828
rect 675386 870816 675392 870828
rect 675444 870816 675450 870868
rect 42242 787244 42248 787296
rect 42300 787284 42306 787296
rect 42426 787284 42432 787296
rect 42300 787256 42432 787284
rect 42300 787244 42306 787256
rect 42426 787244 42432 787256
rect 42484 787244 42490 787296
rect 673730 785952 673736 786004
rect 673788 785992 673794 786004
rect 675202 785992 675208 786004
rect 673788 785964 675208 785992
rect 673788 785952 673794 785964
rect 675202 785952 675208 785964
rect 675260 785992 675266 786004
rect 675386 785992 675392 786004
rect 675260 785964 675392 785992
rect 675260 785952 675266 785964
rect 675386 785952 675392 785964
rect 675444 785952 675450 786004
rect 673730 781600 673736 781652
rect 673788 781640 673794 781652
rect 675202 781640 675208 781652
rect 673788 781612 675208 781640
rect 673788 781600 673794 781612
rect 675202 781600 675208 781612
rect 675260 781640 675266 781652
rect 675386 781640 675392 781652
rect 675260 781612 675392 781640
rect 675260 781600 675266 781612
rect 675386 781600 675392 781612
rect 675444 781600 675450 781652
rect 673730 740936 673736 740988
rect 673788 740976 673794 740988
rect 675202 740976 675208 740988
rect 673788 740948 675208 740976
rect 673788 740936 673794 740948
rect 675202 740936 675208 740948
rect 675260 740976 675266 740988
rect 675386 740976 675392 740988
rect 675260 740948 675392 740976
rect 675260 740936 675266 740948
rect 675386 740936 675392 740948
rect 675444 740936 675450 740988
rect 673730 736992 673736 737044
rect 673788 737032 673794 737044
rect 675202 737032 675208 737044
rect 673788 737004 675208 737032
rect 673788 736992 673794 737004
rect 675202 736992 675208 737004
rect 675260 737032 675266 737044
rect 675386 737032 675392 737044
rect 675260 737004 675392 737032
rect 675260 736992 675266 737004
rect 675386 736992 675392 737004
rect 675444 736992 675450 737044
rect 673730 695920 673736 695972
rect 673788 695960 673794 695972
rect 675202 695960 675208 695972
rect 673788 695932 675208 695960
rect 673788 695920 673794 695932
rect 675202 695920 675208 695932
rect 675260 695960 675266 695972
rect 675386 695960 675392 695972
rect 675260 695932 675392 695960
rect 675260 695920 675266 695932
rect 675386 695920 675392 695932
rect 675444 695920 675450 695972
rect 673730 692044 673736 692096
rect 673788 692084 673794 692096
rect 675202 692084 675208 692096
rect 673788 692056 675208 692084
rect 673788 692044 673794 692056
rect 675202 692044 675208 692056
rect 675260 692084 675266 692096
rect 675386 692084 675392 692096
rect 675260 692056 675392 692084
rect 675260 692044 675266 692056
rect 675386 692044 675392 692056
rect 675444 692044 675450 692096
rect 673730 651108 673736 651160
rect 673788 651148 673794 651160
rect 675386 651148 675392 651160
rect 673788 651120 675392 651148
rect 673788 651108 673794 651120
rect 675386 651108 675392 651120
rect 675444 651108 675450 651160
rect 673730 646416 673736 646468
rect 673788 646456 673794 646468
rect 675386 646456 675392 646468
rect 673788 646428 675392 646456
rect 673788 646416 673794 646428
rect 675386 646416 675392 646428
rect 675444 646416 675450 646468
rect 673730 605752 673736 605804
rect 673788 605792 673794 605804
rect 675202 605792 675208 605804
rect 673788 605764 675208 605792
rect 673788 605752 673794 605764
rect 675202 605752 675208 605764
rect 675260 605792 675266 605804
rect 675386 605792 675392 605804
rect 675260 605764 675392 605792
rect 675260 605752 675266 605764
rect 675386 605752 675392 605764
rect 675444 605752 675450 605804
rect 673730 601808 673736 601860
rect 673788 601848 673794 601860
rect 675202 601848 675208 601860
rect 673788 601820 675208 601848
rect 673788 601808 673794 601820
rect 675202 601808 675208 601820
rect 675260 601848 675266 601860
rect 675386 601848 675392 601860
rect 675260 601820 675392 601848
rect 675260 601808 675266 601820
rect 675386 601808 675392 601820
rect 675444 601808 675450 601860
rect 673730 561076 673736 561128
rect 673788 561116 673794 561128
rect 675202 561116 675208 561128
rect 673788 561088 675208 561116
rect 673788 561076 673794 561088
rect 675202 561076 675208 561088
rect 675260 561076 675266 561128
rect 673638 556588 673644 556640
rect 673696 556628 673702 556640
rect 675202 556628 675208 556640
rect 673696 556600 675208 556628
rect 673696 556588 673702 556600
rect 675202 556588 675208 556600
rect 675260 556628 675266 556640
rect 675386 556628 675392 556640
rect 675260 556600 675392 556628
rect 675260 556588 675266 556600
rect 675386 556588 675392 556600
rect 675444 556588 675450 556640
rect 673638 384276 673644 384328
rect 673696 384316 673702 384328
rect 675386 384316 675392 384328
rect 673696 384288 675392 384316
rect 673696 384276 673702 384288
rect 675386 384276 675392 384288
rect 675444 384276 675450 384328
rect 673638 379040 673644 379092
rect 673696 379080 673702 379092
rect 675386 379080 675392 379092
rect 673696 379052 675392 379080
rect 673696 379040 673702 379052
rect 675386 379040 675392 379052
rect 675444 379040 675450 379092
rect 673638 338784 673644 338836
rect 673696 338824 673702 338836
rect 675386 338824 675392 338836
rect 673696 338796 675392 338824
rect 673696 338784 673702 338796
rect 675386 338784 675392 338796
rect 675444 338784 675450 338836
rect 673822 334228 673828 334280
rect 673880 334268 673886 334280
rect 675386 334268 675392 334280
rect 673880 334240 675392 334268
rect 673880 334228 673886 334240
rect 675386 334228 675392 334240
rect 675444 334228 675450 334280
rect 673822 294652 673828 294704
rect 673880 294692 673886 294704
rect 675294 294692 675300 294704
rect 673880 294664 675300 294692
rect 673880 294652 673886 294664
rect 675294 294652 675300 294664
rect 675352 294652 675358 294704
rect 673638 288804 673644 288856
rect 673696 288844 673702 288856
rect 675386 288844 675392 288856
rect 673696 288816 675392 288844
rect 673696 288804 673702 288816
rect 675386 288804 675392 288816
rect 675444 288804 675450 288856
rect 673638 249092 673644 249144
rect 673696 249132 673702 249144
rect 675386 249132 675392 249144
rect 673696 249104 675392 249132
rect 673696 249092 673702 249104
rect 675386 249092 675392 249104
rect 675444 249092 675450 249144
rect 673822 243788 673828 243840
rect 673880 243828 673886 243840
rect 675386 243828 675392 243840
rect 673880 243800 675392 243828
rect 673880 243788 673886 243800
rect 675386 243788 675392 243800
rect 675444 243788 675450 243840
rect 673822 203464 673828 203516
rect 673880 203504 673886 203516
rect 675294 203504 675300 203516
rect 673880 203476 675300 203504
rect 673880 203464 673886 203476
rect 675294 203464 675300 203476
rect 675352 203464 675358 203516
rect 673730 199044 673736 199096
rect 673788 199084 673794 199096
rect 675386 199084 675392 199096
rect 673788 199056 675392 199084
rect 673788 199044 673794 199056
rect 675386 199044 675392 199056
rect 675444 199044 675450 199096
rect 41782 189116 41788 189168
rect 41840 189156 41846 189168
rect 42426 189156 42432 189168
rect 41840 189128 42432 189156
rect 41840 189116 41846 189128
rect 42426 189116 42432 189128
rect 42484 189116 42490 189168
rect 673730 158584 673736 158636
rect 673788 158624 673794 158636
rect 675386 158624 675392 158636
rect 673788 158596 675392 158624
rect 673788 158584 673794 158596
rect 675386 158584 675392 158596
rect 675444 158584 675450 158636
rect 673638 154096 673644 154148
rect 673696 154136 673702 154148
rect 675294 154136 675300 154148
rect 673696 154108 675300 154136
rect 673696 154096 673702 154108
rect 675294 154096 675300 154108
rect 675352 154096 675358 154148
rect 673638 113704 673644 113756
rect 673696 113744 673702 113756
rect 675386 113744 675392 113756
rect 673696 113716 675392 113744
rect 673696 113704 673702 113716
rect 675386 113704 675392 113716
rect 675444 113704 675450 113756
rect 673638 108400 673644 108452
rect 673696 108440 673702 108452
rect 675386 108440 675392 108452
rect 673696 108412 675392 108440
rect 673696 108400 673702 108412
rect 675386 108400 675392 108412
rect 675444 108400 675450 108452
rect 673638 46968 673644 46980
rect 52454 46860 52460 46912
rect 52512 46900 52518 46912
rect 143534 46900 143540 46912
rect 52512 46872 143540 46900
rect 52512 46860 52518 46872
rect 143534 46860 143540 46872
rect 143592 46860 143598 46912
rect 527468 46940 673644 46968
rect 527468 46912 527496 46940
rect 673638 46928 673644 46940
rect 673696 46928 673702 46980
rect 527450 46860 527456 46912
rect 527508 46860 527514 46912
rect 468294 44384 468300 44396
rect 358722 44316 358728 44328
rect 349908 44288 358728 44316
rect 303890 44248 303896 44260
rect 206986 44220 303896 44248
rect 143534 44140 143540 44192
rect 143592 44180 143598 44192
rect 145098 44180 145104 44192
rect 143592 44152 145104 44180
rect 143592 44140 143598 44152
rect 145098 44140 145104 44152
rect 145156 44180 145162 44192
rect 195330 44180 195336 44192
rect 145156 44152 195336 44180
rect 145156 44140 145162 44152
rect 195330 44140 195336 44152
rect 195388 44180 195394 44192
rect 199654 44180 199660 44192
rect 195388 44152 199660 44180
rect 195388 44140 195394 44152
rect 199654 44140 199660 44152
rect 199712 44180 199718 44192
rect 206986 44180 207014 44220
rect 303890 44208 303896 44220
rect 303948 44248 303954 44260
rect 308214 44248 308220 44260
rect 303948 44220 308220 44248
rect 303948 44208 303954 44220
rect 308214 44208 308220 44220
rect 308272 44248 308278 44260
rect 349908 44248 349936 44288
rect 358722 44276 358728 44288
rect 358780 44316 358786 44328
rect 363046 44316 363052 44328
rect 358780 44288 363052 44316
rect 358780 44276 358786 44288
rect 363046 44276 363052 44288
rect 363104 44316 363110 44328
rect 417896 44356 468300 44384
rect 363104 44288 363368 44316
rect 363104 44276 363110 44288
rect 363340 44248 363368 44288
rect 417896 44260 417924 44356
rect 468294 44344 468300 44356
rect 468352 44384 468358 44396
rect 472618 44384 472624 44396
rect 468352 44356 472624 44384
rect 468352 44344 468358 44356
rect 472618 44344 472624 44356
rect 472676 44384 472682 44396
rect 472676 44356 477494 44384
rect 472676 44344 472682 44356
rect 477466 44316 477494 44356
rect 477466 44288 523172 44316
rect 413554 44248 413560 44260
rect 308272 44220 349936 44248
rect 363340 44220 413560 44248
rect 308272 44208 308278 44220
rect 199712 44152 207014 44180
rect 199712 44140 199718 44152
rect 413554 44208 413560 44220
rect 413612 44248 413618 44260
rect 417878 44248 417884 44260
rect 413612 44220 417884 44248
rect 413612 44208 413618 44220
rect 417878 44208 417884 44220
rect 417936 44208 417942 44260
rect 523144 44192 523172 44288
rect 523126 44140 523132 44192
rect 523184 44180 523190 44192
rect 527450 44180 527456 44192
rect 523184 44152 527456 44180
rect 523184 44140 523190 44152
rect 527450 44140 527456 44152
rect 527508 44140 527514 44192
rect 409322 41760 409328 41812
rect 409380 41800 409386 41812
rect 412358 41800 412364 41812
rect 409380 41772 412364 41800
rect 409380 41760 409386 41772
rect 412358 41760 412364 41772
rect 412416 41800 412422 41812
rect 415210 41800 415216 41812
rect 412416 41772 415216 41800
rect 412416 41760 412422 41772
rect 415210 41760 415216 41772
rect 415268 41760 415274 41812
rect 464154 41760 464160 41812
rect 464212 41800 464218 41812
rect 467190 41800 467196 41812
rect 464212 41772 467196 41800
rect 464212 41760 464218 41772
rect 467190 41760 467196 41772
rect 467248 41800 467254 41812
rect 470042 41800 470048 41812
rect 467248 41772 470048 41800
rect 467248 41760 467254 41772
rect 470042 41760 470048 41772
rect 470100 41760 470106 41812
<< via1 >>
rect 673736 870816 673788 870868
rect 675392 870816 675444 870868
rect 42248 787244 42300 787296
rect 42432 787244 42484 787296
rect 673736 785952 673788 786004
rect 675208 785952 675260 786004
rect 675392 785952 675444 786004
rect 673736 781600 673788 781652
rect 675208 781600 675260 781652
rect 675392 781600 675444 781652
rect 673736 740936 673788 740988
rect 675208 740936 675260 740988
rect 675392 740936 675444 740988
rect 673736 736992 673788 737044
rect 675208 736992 675260 737044
rect 675392 736992 675444 737044
rect 673736 695920 673788 695972
rect 675208 695920 675260 695972
rect 675392 695920 675444 695972
rect 673736 692044 673788 692096
rect 675208 692044 675260 692096
rect 675392 692044 675444 692096
rect 673736 651108 673788 651160
rect 675392 651108 675444 651160
rect 673736 646416 673788 646468
rect 675392 646416 675444 646468
rect 673736 605752 673788 605804
rect 675208 605752 675260 605804
rect 675392 605752 675444 605804
rect 673736 601808 673788 601860
rect 675208 601808 675260 601860
rect 675392 601808 675444 601860
rect 673736 561076 673788 561128
rect 675208 561076 675260 561128
rect 673644 556588 673696 556640
rect 675208 556588 675260 556640
rect 675392 556588 675444 556640
rect 673644 384276 673696 384328
rect 675392 384276 675444 384328
rect 673644 379040 673696 379092
rect 675392 379040 675444 379092
rect 673644 338784 673696 338836
rect 675392 338784 675444 338836
rect 673828 334228 673880 334280
rect 675392 334228 675444 334280
rect 673828 294652 673880 294704
rect 675300 294652 675352 294704
rect 673644 288804 673696 288856
rect 675392 288804 675444 288856
rect 673644 249092 673696 249144
rect 675392 249092 675444 249144
rect 673828 243788 673880 243840
rect 675392 243788 675444 243840
rect 673828 203464 673880 203516
rect 675300 203464 675352 203516
rect 673736 199044 673788 199096
rect 675392 199044 675444 199096
rect 41788 189116 41840 189168
rect 42432 189116 42484 189168
rect 673736 158584 673788 158636
rect 675392 158584 675444 158636
rect 673644 154096 673696 154148
rect 675300 154096 675352 154148
rect 673644 113704 673696 113756
rect 675392 113704 675444 113756
rect 673644 108400 673696 108452
rect 675392 108400 675444 108452
rect 52460 46860 52512 46912
rect 143540 46860 143592 46912
rect 673644 46928 673696 46980
rect 527456 46860 527508 46912
rect 143540 44140 143592 44192
rect 145104 44140 145156 44192
rect 195336 44140 195388 44192
rect 199660 44140 199712 44192
rect 303896 44208 303948 44260
rect 308220 44208 308272 44260
rect 358728 44276 358780 44328
rect 363052 44276 363104 44328
rect 468300 44344 468352 44396
rect 472624 44344 472676 44396
rect 413560 44208 413612 44260
rect 417884 44208 417936 44260
rect 523132 44140 523184 44192
rect 527456 44140 527508 44192
rect 409328 41760 409380 41812
rect 412364 41760 412416 41812
rect 415216 41760 415268 41812
rect 464160 41760 464212 41812
rect 467196 41760 467248 41812
rect 470048 41760 470100 41812
<< obsm1 >>
rect 77050 1006851 90288 1007371
rect 128450 1006851 141688 1007371
rect 179850 1006851 193088 1007371
rect 230437 998007 244983 1037545
rect 282037 998007 296583 1037545
rect 333437 998007 348124 1037545
rect 384650 1006851 397888 1007371
rect 473650 1006851 486888 1007371
rect 525050 1006851 538288 1007371
rect 575637 998007 590324 1037545
rect 626850 1006851 640088 1007371
rect 231125 997826 232171 998007
rect 232807 997984 233070 998007
tri 233070 997984 233093 998007 sw
tri 244285 997984 244308 998007 se
rect 244308 997984 244536 998007
rect 232807 997794 244536 997984
rect 282725 997826 283771 998007
rect 284407 997984 284670 998007
tri 284670 997984 284693 998007 sw
tri 295885 997984 295908 998007 se
rect 295908 997984 296136 998007
rect 284407 997794 296136 997984
rect 335807 997984 336070 998007
tri 336070 997984 336093 998007 sw
tri 347285 997984 347308 998007 se
rect 347308 997984 347536 998007
rect 335807 997794 347536 997984
rect 578007 997984 578270 998007
tri 578270 997984 578293 998007 sw
tri 589485 997984 589508 998007 se
rect 589508 997984 589736 998007
rect 578007 997794 589736 997984
rect 585042 996384 585106 996396
rect 674742 996384 674806 996396
rect 585042 996356 674806 996384
rect 585042 996344 585106 996356
rect 674742 996344 674806 996356
rect 356054 990876 356118 990888
rect 673546 990876 673610 990888
rect 356054 990848 673610 990876
rect 356054 990836 356118 990848
rect 673546 990836 673610 990848
rect 42242 990196 42306 990208
rect 42242 990168 52454 990196
rect 42242 990156 42306 990168
rect 44910 990088 44974 990140
rect 52426 990128 52454 990168
rect 343634 990128 343698 990140
rect 356054 990128 356118 990140
rect 52426 990100 356118 990128
rect 343634 990088 343698 990100
rect 356054 990088 356118 990100
rect 44928 990060 44956 990088
rect 673454 990060 673518 990072
rect 44928 990032 673518 990060
rect 673454 990020 673518 990032
rect 30229 955050 30749 968288
rect 678007 966875 717545 967563
rect 677826 965829 717545 966875
rect 678007 965193 717545 965829
rect 677794 964930 717545 965193
rect 677794 953692 677984 964930
tri 677984 964907 678007 964930 nw
tri 677984 953692 678007 953715 sw
rect 678007 953692 717545 964930
rect 677794 953464 717545 953692
rect 678007 953017 717545 953464
rect 24523 928387 40977 929187
tri 40977 928387 41777 929187 sw
rect 24523 927240 41777 928387
rect 32 923313 39593 927000
rect 39756 923313 41777 927240
rect 32 916185 41777 923313
rect 678007 919269 717568 922576
rect 678000 918415 717568 919269
rect 32 915331 39600 916185
rect 32 912024 39593 915331
rect 675823 911287 717568 918415
rect 675823 907360 677844 911287
rect 678007 907600 717568 911287
rect 675823 906213 693077 907360
tri 675823 905413 676623 906213 ne
rect 676623 905413 693077 906213
rect 55 883936 39593 884383
rect 55 883708 39806 883936
rect 55 872470 39593 883708
tri 39593 883685 39616 883708 ne
tri 39593 872470 39616 872493 se
rect 39616 872470 39806 883708
rect 689038 878400 693727 878423
rect 695550 878400 695896 878429
rect 696779 878400 703644 878423
rect 703855 878400 711618 878423
rect 673546 874528 673610 874540
rect 675386 874528 675450 874540
rect 673546 874500 675450 874528
rect 673546 874488 673610 874500
rect 675386 874488 675450 874500
rect 55 872207 39806 872470
rect 673454 872420 673518 872432
rect 673638 872420 673702 872432
rect 675386 872420 675450 872432
rect 673454 872392 675450 872420
rect 673454 872380 673518 872392
rect 673638 872380 673702 872392
rect 675386 872380 675450 872392
rect 55 871571 39593 872207
rect 55 870525 39774 871571
rect 55 869837 39593 870525
rect 673822 870176 673886 870188
rect 675386 870176 675450 870188
rect 673822 870148 675450 870176
rect 673822 870136 673886 870148
rect 675386 870136 675450 870148
rect 673454 864260 673518 864272
rect 675386 864260 675450 864272
rect 673454 864232 675450 864260
rect 673454 864220 673518 864232
rect 675386 864220 675450 864232
rect 673822 863240 673886 863252
rect 675386 863240 675450 863252
rect 673822 863212 675450 863240
rect 673822 863200 673886 863212
rect 675386 863200 675450 863212
rect 676231 862400 717600 878400
rect 681497 862377 682603 862400
rect 683624 862377 684745 862400
rect 687844 862388 696516 862400
rect 687844 862377 692186 862388
tri 692186 862377 692197 862388 nw
rect 696779 862371 703644 862400
rect 703855 862371 711618 862400
rect 713380 862396 713795 862400
rect 55 841736 39593 842324
rect 55 841508 39806 841736
rect 55 830270 39593 841508
tri 39593 841485 39616 841508 ne
tri 39593 830270 39616 830293 se
rect 39616 830270 39806 841508
rect 678007 832675 717545 833363
rect 677826 831629 717545 832675
rect 678007 830993 717545 831629
rect 55 830007 39806 830270
rect 677794 830730 717545 830993
rect 55 827637 39593 830007
rect 677794 819492 677984 830730
tri 677984 830707 678007 830730 nw
tri 677984 819492 678007 819515 sw
rect 678007 819492 717545 830730
rect 677794 819264 717545 819492
rect 678007 818817 717545 819264
rect 675294 818360 675358 818372
rect 677594 818360 677658 818372
rect 675294 818332 677658 818360
rect 675294 818320 675358 818332
rect 677594 818320 677658 818332
rect 3805 800400 4220 800404
rect 5982 800400 13745 800429
rect 13956 800400 20821 800429
tri 25403 800412 25414 800423 se
rect 25414 800412 29756 800423
rect 21084 800400 29756 800412
rect 32855 800400 33976 800423
rect 34997 800400 36103 800423
rect 0 784400 41369 800400
rect 41782 797756 41846 797768
rect 42610 797756 42674 797768
rect 41782 797728 42674 797756
rect 41782 797716 41846 797728
rect 42610 797716 42674 797728
rect 41782 791364 41846 791376
rect 42426 791364 42490 791376
rect 41782 791336 42490 791364
rect 41782 791324 41846 791336
rect 42426 791324 42490 791336
rect 689038 789200 693727 789223
rect 695550 789200 695896 789229
rect 696779 789200 703644 789223
rect 703855 789200 711618 789223
rect 41782 788304 41846 788316
rect 42334 788304 42398 788316
rect 41782 788276 42398 788304
rect 41782 788264 41846 788276
rect 42334 788264 42398 788276
rect 41782 787244 41846 787296
rect 41800 787080 41828 787244
rect 42242 787080 42306 787092
rect 41800 787052 42306 787080
rect 42242 787040 42306 787052
rect 42334 787012 42398 787024
rect 42518 787012 42582 787024
rect 42334 786984 42582 787012
rect 42334 786972 42398 786984
rect 42518 786972 42582 786984
rect 673546 785720 673610 785732
rect 675386 785720 675450 785732
rect 673546 785692 675450 785720
rect 673546 785680 673610 785692
rect 675386 785680 675450 785692
rect 5982 784377 13745 784400
rect 13956 784377 20821 784400
rect 21704 784371 22050 784400
rect 23873 784377 28562 784400
rect 673638 782320 673702 782332
rect 675386 782320 675450 782332
rect 673638 782292 675450 782320
rect 673638 782280 673702 782292
rect 675386 782280 675450 782292
rect 675202 781028 675266 781040
rect 675386 781028 675450 781040
rect 675202 781000 675450 781028
rect 675202 780988 675266 781000
rect 675386 780988 675450 781000
rect 673454 775860 673518 775872
rect 675386 775860 675450 775872
rect 673454 775832 675450 775860
rect 673454 775820 673518 775832
rect 675386 775820 675450 775832
rect 676231 773200 717600 789200
rect 681497 773177 682603 773200
rect 683624 773177 684745 773200
rect 687844 773188 696516 773200
rect 687844 773177 692186 773188
tri 692186 773177 692197 773188 nw
rect 696779 773171 703644 773200
rect 703855 773171 711618 773200
rect 713380 773196 713795 773200
rect 42242 757636 42306 757648
rect 42794 757636 42858 757648
rect 42242 757608 42858 757636
rect 42242 757596 42306 757608
rect 42794 757596 42858 757608
rect 42334 757568 42398 757580
rect 42702 757568 42766 757580
rect 42334 757540 42766 757568
rect 42334 757528 42398 757540
rect 42702 757528 42766 757540
rect 3805 757200 4220 757204
rect 5982 757200 13745 757229
rect 13956 757200 20821 757229
tri 25403 757212 25414 757223 se
rect 25414 757212 29756 757223
rect 21084 757200 29756 757212
rect 32855 757200 33976 757223
rect 34997 757200 36103 757223
rect 0 741200 41369 757200
rect 41782 755460 41846 755472
rect 42610 755460 42674 755472
rect 41782 755432 42674 755460
rect 41782 755420 41846 755432
rect 42610 755420 42674 755432
rect 41782 747708 41846 747720
rect 42702 747708 42766 747720
rect 41782 747680 42766 747708
rect 41782 747668 41846 747680
rect 42702 747668 42766 747680
rect 689038 744200 693727 744223
rect 695550 744200 695896 744229
rect 696779 744200 703644 744223
rect 703855 744200 711618 744223
rect 41782 744036 41846 744048
rect 42794 744036 42858 744048
rect 41782 744008 42858 744036
rect 41782 743996 41846 744008
rect 42794 743996 42858 744008
rect 5982 741177 13745 741200
rect 13956 741177 20821 741200
rect 21704 741171 22050 741200
rect 23873 741177 28562 741200
rect 673546 740364 673610 740376
rect 673822 740364 673886 740376
rect 675386 740364 675450 740376
rect 673546 740336 675450 740364
rect 673546 740324 673610 740336
rect 673822 740324 673886 740336
rect 675386 740324 675450 740336
rect 673638 738120 673702 738132
rect 675386 738120 675450 738132
rect 673638 738092 675450 738120
rect 673638 738080 673702 738092
rect 675386 738080 675450 738092
rect 673454 730912 673518 730924
rect 674006 730912 674070 730924
rect 675386 730912 675450 730924
rect 673454 730884 675450 730912
rect 673454 730872 673518 730884
rect 674006 730872 674070 730884
rect 675386 730872 675450 730884
rect 676231 728200 717600 744200
rect 681497 728177 682603 728200
rect 683624 728177 684745 728200
rect 687844 728188 696516 728200
rect 687844 728177 692186 728188
tri 692186 728177 692197 728188 nw
rect 696779 728171 703644 728200
rect 703855 728171 711618 728200
rect 713380 728196 713795 728200
rect 3805 714000 4220 714004
rect 5982 714000 13745 714029
rect 13956 714000 20821 714029
tri 25403 714012 25414 714023 se
rect 25414 714012 29756 714023
rect 21084 714000 29756 714012
rect 32855 714000 33976 714023
rect 34997 714000 36103 714023
rect 0 698000 41369 714000
rect 41782 712280 41846 712292
rect 42610 712280 42674 712292
rect 41782 712252 42674 712280
rect 41782 712240 41846 712252
rect 42610 712240 42674 712252
rect 41782 703984 41846 703996
rect 42426 703984 42490 703996
rect 42702 703984 42766 703996
rect 41782 703956 42766 703984
rect 41782 703944 41846 703956
rect 42426 703944 42490 703956
rect 42702 703944 42766 703956
rect 41782 700856 41846 700868
rect 42610 700856 42674 700868
rect 41782 700828 42674 700856
rect 41782 700816 41846 700828
rect 42610 700816 42674 700828
rect 689038 699200 693727 699223
rect 695550 699200 695896 699229
rect 696779 699200 703644 699223
rect 703855 699200 711618 699223
rect 5982 697977 13745 698000
rect 13956 697977 20821 698000
rect 21704 697971 22050 698000
rect 23873 697977 28562 698000
rect 673454 695348 673518 695360
rect 673822 695348 673886 695360
rect 675386 695348 675450 695360
rect 673454 695320 675450 695348
rect 673454 695308 673518 695320
rect 673822 695308 673886 695320
rect 675386 695308 675450 695320
rect 673914 692288 673978 692300
rect 675386 692288 675450 692300
rect 673914 692260 675450 692288
rect 673914 692248 673978 692260
rect 675386 692248 675450 692260
rect 673546 685216 673610 685228
rect 674006 685216 674070 685228
rect 675386 685216 675450 685228
rect 673546 685188 675450 685216
rect 673546 685176 673610 685188
rect 674006 685176 674070 685188
rect 675386 685176 675450 685188
rect 676231 683200 717600 699200
rect 681497 683177 682603 683200
rect 683624 683177 684745 683200
rect 687844 683188 696516 683200
rect 687844 683177 692186 683188
tri 692186 683177 692197 683188 nw
rect 696779 683171 703644 683200
rect 703855 683171 711618 683200
rect 713380 683196 713795 683200
rect 3805 670800 4220 670804
rect 5982 670800 13745 670829
rect 13956 670800 20821 670829
tri 25403 670812 25414 670823 se
rect 25414 670812 29756 670823
rect 21084 670800 29756 670812
rect 32855 670800 33976 670823
rect 34997 670800 36103 670823
rect 0 654800 41369 670800
rect 41782 668148 41846 668160
rect 42518 668148 42582 668160
rect 41782 668120 42582 668148
rect 41782 668108 41846 668120
rect 42518 668108 42582 668120
rect 41782 661076 41846 661088
rect 42426 661076 42490 661088
rect 41782 661048 42490 661076
rect 41782 661036 41846 661048
rect 42426 661036 42490 661048
rect 41782 658696 41846 658708
rect 42610 658696 42674 658708
rect 41782 658668 42674 658696
rect 41782 658656 41846 658668
rect 42610 658656 42674 658668
rect 5982 654777 13745 654800
rect 13956 654777 20821 654800
rect 21704 654771 22050 654800
rect 23873 654777 28562 654800
rect 689038 654000 693727 654023
rect 695550 654000 695896 654029
rect 696779 654000 703644 654023
rect 703855 654000 711618 654023
rect 673454 650536 673518 650548
rect 675386 650536 675450 650548
rect 673454 650508 675450 650536
rect 673454 650496 673518 650508
rect 675386 650496 675450 650508
rect 673454 647204 673518 647216
rect 673638 647204 673702 647216
rect 673454 647176 673702 647204
rect 673454 647164 673518 647176
rect 673638 647164 673702 647176
rect 673454 647068 673518 647080
rect 673914 647068 673978 647080
rect 675386 647068 675450 647080
rect 673454 647040 675450 647068
rect 673454 647028 673518 647040
rect 673914 647028 673978 647040
rect 675386 647028 675450 647040
rect 675202 645776 675266 645788
rect 675386 645776 675450 645788
rect 675202 645748 675450 645776
rect 675202 645736 675266 645748
rect 675386 645736 675450 645748
rect 673546 640676 673610 640688
rect 675386 640676 675450 640688
rect 673546 640648 675450 640676
rect 673546 640636 673610 640648
rect 675386 640636 675450 640648
rect 676231 638000 717600 654000
rect 681497 637977 682603 638000
rect 683624 637977 684745 638000
rect 687844 637988 696516 638000
rect 687844 637977 692186 637988
tri 692186 637977 692197 637988 nw
rect 696779 637971 703644 638000
rect 703855 637971 711618 638000
rect 713380 637996 713795 638000
rect 3805 627600 4220 627604
rect 5982 627600 13745 627629
rect 13956 627600 20821 627629
tri 25403 627612 25414 627623 se
rect 25414 627612 29756 627623
rect 21084 627600 29756 627612
rect 32855 627600 33976 627623
rect 34997 627600 36103 627623
rect 0 611600 41369 627600
rect 41782 624968 41846 624980
rect 42518 624968 42582 624980
rect 41782 624940 42582 624968
rect 41782 624928 41846 624940
rect 42518 624928 42582 624940
rect 41782 618508 41846 618520
rect 42426 618508 42490 618520
rect 41782 618480 42490 618508
rect 41782 618468 41846 618480
rect 42426 618468 42490 618480
rect 41782 615516 41846 615528
rect 42610 615516 42674 615528
rect 41782 615488 42674 615516
rect 41782 615476 41846 615488
rect 42610 615476 42674 615488
rect 5982 611577 13745 611600
rect 13956 611577 20821 611600
rect 21704 611571 22050 611600
rect 23873 611577 28562 611600
rect 689038 609000 693727 609023
rect 695550 609000 695896 609029
rect 696779 609000 703644 609023
rect 703855 609000 711618 609023
rect 673638 605112 673702 605124
rect 675386 605112 675450 605124
rect 673638 605084 675450 605112
rect 673638 605072 673702 605084
rect 675386 605072 675450 605084
rect 42518 603168 42582 603220
rect 42536 603016 42564 603168
rect 42518 602964 42582 603016
rect 673454 602936 673518 602948
rect 675386 602936 675450 602948
rect 673454 602908 675450 602936
rect 673454 602896 673518 602908
rect 675386 602896 675450 602908
rect 673546 595048 673610 595060
rect 675386 595048 675450 595060
rect 673546 595020 675450 595048
rect 673546 595008 673610 595020
rect 675386 595008 675450 595020
rect 676231 593000 717600 609000
rect 681497 592977 682603 593000
rect 683624 592977 684745 593000
rect 687844 592988 696516 593000
rect 687844 592977 692186 592988
tri 692186 592977 692197 592988 nw
rect 696779 592971 703644 593000
rect 703855 592971 711618 593000
rect 713380 592996 713795 593000
rect 3805 584400 4220 584404
rect 5982 584400 13745 584429
rect 13956 584400 20821 584429
tri 25403 584412 25414 584423 se
rect 25414 584412 29756 584423
rect 21084 584400 29756 584412
rect 32855 584400 33976 584423
rect 34997 584400 36103 584423
rect 0 568400 41369 584400
rect 41782 581720 41846 581732
rect 42426 581720 42490 581732
rect 41782 581692 42490 581720
rect 41782 581680 41846 581692
rect 42426 581680 42490 581692
rect 41782 575260 41846 575272
rect 42702 575260 42766 575272
rect 41782 575232 42766 575260
rect 41782 575220 41846 575232
rect 42702 575220 42766 575232
rect 41782 572268 41846 572280
rect 42518 572268 42582 572280
rect 42794 572268 42858 572280
rect 41782 572240 42858 572268
rect 41782 572228 41846 572240
rect 42518 572228 42582 572240
rect 42794 572228 42858 572240
rect 42242 571180 42306 571192
rect 42426 571180 42490 571192
rect 42242 571152 42490 571180
rect 42242 571140 42306 571152
rect 42426 571140 42490 571152
rect 5982 568377 13745 568400
rect 13956 568377 20821 568400
rect 21704 568371 22050 568400
rect 23873 568377 28562 568400
rect 689038 563800 693727 563823
rect 695550 563800 695896 563829
rect 696779 563800 703644 563823
rect 703855 563800 711618 563823
rect 673638 560980 673702 560992
rect 675386 560980 675450 560992
rect 673638 560952 675450 560980
rect 673638 560940 673702 560952
rect 675386 560940 675450 560952
rect 673454 557852 673518 557864
rect 675386 557852 675450 557864
rect 673454 557824 675450 557852
rect 673454 557812 673518 557824
rect 675386 557812 675450 557824
rect 675202 555608 675266 555620
rect 675386 555608 675450 555620
rect 675202 555580 675450 555608
rect 675202 555568 675266 555580
rect 675386 555568 675450 555580
rect 673546 550508 673610 550520
rect 675386 550508 675450 550520
rect 673546 550480 675450 550508
rect 673546 550468 673610 550480
rect 675386 550468 675450 550480
rect 676231 547800 717600 563800
rect 681497 547777 682603 547800
rect 683624 547777 684745 547800
rect 687844 547788 696516 547800
rect 687844 547777 692186 547788
tri 692186 547777 692197 547788 nw
rect 696779 547771 703644 547800
rect 703855 547771 711618 547800
rect 713380 547796 713795 547800
rect 42242 543096 42306 543108
rect 42426 543096 42490 543108
rect 42242 543068 42490 543096
rect 42242 543056 42306 543068
rect 42426 543056 42490 543068
rect 3805 541200 4220 541204
rect 5982 541200 13745 541229
rect 13956 541200 20821 541229
tri 25403 541212 25414 541223 se
rect 25414 541212 29756 541223
rect 21084 541200 29756 541212
rect 32855 541200 33976 541223
rect 34997 541200 36103 541223
rect 0 525200 41369 541200
rect 41782 539492 41846 539504
rect 42426 539492 42490 539504
rect 42794 539492 42858 539504
rect 41782 539464 42858 539492
rect 41782 539452 41846 539464
rect 42426 539452 42490 539464
rect 42794 539452 42858 539464
rect 41782 531196 41846 531208
rect 42426 531196 42490 531208
rect 41782 531168 42490 531196
rect 41782 531156 41846 531168
rect 42426 531156 42490 531168
rect 41782 528068 41846 528080
rect 42334 528068 42398 528080
rect 42702 528068 42766 528080
rect 41782 528040 42766 528068
rect 41782 528028 41846 528040
rect 42334 528028 42398 528040
rect 42702 528028 42766 528040
rect 5982 525177 13745 525200
rect 13956 525177 20821 525200
rect 21704 525171 22050 525200
rect 23873 525177 28562 525200
rect 678007 518075 717545 518763
rect 677826 517029 717545 518075
rect 678007 516393 717545 517029
rect 677794 516130 717545 516393
rect 675294 513788 675358 513800
rect 677686 513788 677750 513800
rect 675294 513760 677750 513788
rect 675294 513748 675358 513760
rect 677686 513748 677750 513760
rect 677794 504892 677984 516130
tri 677984 516107 678007 516130 nw
tri 677984 504892 678007 504915 sw
rect 678007 504892 717545 516130
rect 677794 504664 717545 504892
rect 678007 504217 717545 504664
rect 55 497136 39593 497583
rect 55 496908 39806 497136
rect 55 485670 39593 496908
tri 39593 496885 39616 496908 ne
tri 39593 485670 39616 485693 se
rect 39616 485670 39806 496908
rect 55 485407 39806 485670
rect 55 484771 39593 485407
rect 55 483725 39774 484771
rect 55 483037 39593 483725
rect 678007 471469 717568 474776
rect 678000 470615 717568 471469
rect 675823 463487 717568 470615
rect 675823 459560 677844 463487
rect 678007 459800 717568 463487
rect 675823 458413 693077 459560
tri 675823 457987 676249 458413 ne
rect 676249 457987 693077 458413
rect 24523 457187 40977 457987
tri 40977 457187 41777 457987 sw
tri 676249 457613 676623 457987 ne
rect 676623 457613 693077 457987
rect 24523 456040 41777 457187
rect 32 452113 39593 455800
rect 39756 452113 41777 456040
rect 32 444985 41777 452113
rect 32 444131 39600 444985
rect 32 440824 39593 444131
rect 678007 428193 717545 430563
rect 677794 427930 717545 428193
rect 674742 427836 674806 427848
rect 677502 427836 677566 427848
rect 674742 427808 677566 427836
rect 674742 427796 674806 427808
rect 677502 427796 677566 427808
rect 677794 416692 677984 427930
tri 677984 427907 678007 427930 nw
tri 677984 416692 678007 416715 sw
rect 678007 416692 717545 427930
rect 677794 416464 717545 416692
rect 678007 415876 717545 416464
rect 3805 413600 4220 413604
rect 5982 413600 13745 413629
rect 13956 413600 20821 413629
tri 25403 413612 25414 413623 se
rect 25414 413612 29756 413623
rect 21084 413600 29756 413612
rect 32855 413600 33976 413623
rect 34997 413600 36103 413623
rect 0 397600 41369 413600
rect 41782 410972 41846 410984
rect 42518 410972 42582 410984
rect 42794 410972 42858 410984
rect 41782 410944 42858 410972
rect 41782 410932 41846 410944
rect 42518 410932 42582 410944
rect 42794 410932 42858 410944
rect 41782 404512 41846 404524
rect 42426 404512 42490 404524
rect 42610 404512 42674 404524
rect 41782 404484 42674 404512
rect 41782 404472 41846 404484
rect 42426 404472 42490 404484
rect 42610 404472 42674 404484
rect 41782 400840 41846 400852
rect 42702 400840 42766 400852
rect 41782 400812 42766 400840
rect 41782 400800 41846 400812
rect 42702 400800 42766 400812
rect 5982 397577 13745 397600
rect 13956 397577 20821 397600
rect 21704 397571 22050 397600
rect 23873 397577 28562 397600
rect 689038 386600 693727 386623
rect 695550 386600 695896 386629
rect 696779 386600 703644 386623
rect 703855 386600 711618 386623
rect 673546 382752 673610 382764
rect 675386 382752 675450 382764
rect 673546 382724 675450 382752
rect 673546 382712 673610 382724
rect 675386 382712 675450 382724
rect 673730 379692 673794 379704
rect 675386 379692 675450 379704
rect 673730 379664 675450 379692
rect 673730 379652 673794 379664
rect 675386 379652 675450 379664
rect 673454 372348 673518 372360
rect 673914 372348 673978 372360
rect 675386 372348 675450 372360
rect 673454 372320 675450 372348
rect 673454 372308 673518 372320
rect 673914 372308 673978 372320
rect 675386 372308 675450 372320
rect 676231 370600 717600 386600
rect 681497 370577 682603 370600
rect 683624 370577 684745 370600
rect 687844 370588 696516 370600
rect 687844 370577 692186 370588
tri 692186 370577 692197 370588 nw
rect 696779 370571 703644 370600
rect 703855 370571 711618 370600
rect 713380 370596 713795 370600
rect 3805 370400 4220 370404
rect 5982 370400 13745 370429
rect 13956 370400 20821 370429
tri 25403 370412 25414 370423 se
rect 25414 370412 29756 370423
rect 21084 370400 29756 370412
rect 32855 370400 33976 370423
rect 34997 370400 36103 370423
rect 0 354400 41369 370400
rect 41782 369560 41846 369572
rect 42334 369560 42398 369572
rect 41782 369532 42398 369560
rect 41782 369520 41846 369532
rect 42334 369520 42398 369532
rect 41782 368676 41846 368688
rect 42518 368676 42582 368688
rect 41782 368648 42582 368676
rect 41782 368636 41846 368648
rect 42518 368636 42582 368648
rect 41782 362624 41846 362636
rect 42334 362624 42398 362636
rect 41782 362596 42398 362624
rect 41782 362584 41846 362596
rect 42334 362584 42398 362596
rect 41782 360720 41846 360732
rect 42610 360720 42674 360732
rect 41782 360692 42674 360720
rect 41782 360680 41846 360692
rect 42610 360680 42674 360692
rect 41782 357252 41846 357264
rect 42518 357252 42582 357264
rect 42702 357252 42766 357264
rect 41782 357224 42766 357252
rect 41782 357212 41846 357224
rect 42518 357212 42582 357224
rect 42702 357212 42766 357224
rect 5982 354377 13745 354400
rect 13956 354377 20821 354400
rect 21704 354371 22050 354400
rect 23873 354377 28562 354400
rect 689038 341400 693727 341423
rect 695550 341400 695896 341429
rect 696779 341400 703644 341423
rect 703855 341400 711618 341423
rect 673546 337532 673610 337544
rect 675386 337532 675450 337544
rect 673546 337504 675450 337532
rect 673546 337492 673610 337504
rect 675386 337492 675450 337504
rect 673730 334472 673794 334484
rect 674006 334472 674070 334484
rect 675386 334472 675450 334484
rect 673730 334444 675450 334472
rect 673730 334432 673794 334444
rect 674006 334432 674070 334444
rect 675386 334432 675450 334444
rect 673914 328080 673978 328092
rect 675386 328080 675450 328092
rect 673914 328052 675450 328080
rect 673914 328040 673978 328052
rect 675386 328040 675450 328052
rect 3805 327200 4220 327204
rect 5982 327200 13745 327229
rect 13956 327200 20821 327229
tri 25403 327212 25414 327223 se
rect 25414 327212 29756 327223
rect 21084 327200 29756 327212
rect 32855 327200 33976 327223
rect 34997 327200 36103 327223
rect 0 311200 41369 327200
rect 41782 325496 41846 325508
rect 42426 325496 42490 325508
rect 42794 325496 42858 325508
rect 41782 325468 42858 325496
rect 41782 325456 41846 325468
rect 42426 325456 42490 325468
rect 42794 325456 42858 325468
rect 676231 325400 717600 341400
rect 681497 325377 682603 325400
rect 683624 325377 684745 325400
rect 687844 325388 696516 325400
rect 687844 325377 692186 325388
tri 692186 325377 692197 325388 nw
rect 696779 325371 703644 325400
rect 703855 325371 711618 325400
rect 713380 325396 713795 325400
rect 41782 317200 41846 317212
rect 42610 317200 42674 317212
rect 41782 317172 42674 317200
rect 41782 317160 41846 317172
rect 42610 317160 42674 317172
rect 41782 314072 41846 314084
rect 42518 314072 42582 314084
rect 42702 314072 42766 314084
rect 41782 314044 42766 314072
rect 41782 314032 41846 314044
rect 42518 314032 42582 314044
rect 42702 314032 42766 314044
rect 5982 311177 13745 311200
rect 13956 311177 20821 311200
rect 21704 311171 22050 311200
rect 23873 311177 28562 311200
rect 689038 296400 693727 296423
rect 695550 296400 695896 296429
rect 696779 296400 703644 296423
rect 703855 296400 711618 296423
rect 673454 293196 673518 293208
rect 675386 293196 675450 293208
rect 673454 293168 675450 293196
rect 673454 293156 673518 293168
rect 675386 293156 675450 293168
rect 673546 289524 673610 289536
rect 674006 289524 674070 289536
rect 675386 289524 675450 289536
rect 673546 289496 675450 289524
rect 673546 289484 673610 289496
rect 674006 289484 674070 289496
rect 675386 289484 675450 289496
rect 3805 284000 4220 284004
rect 5982 284000 13745 284029
rect 13956 284000 20821 284029
tri 25403 284012 25414 284023 se
rect 25414 284012 29756 284023
rect 21084 284000 29756 284012
rect 32855 284000 33976 284023
rect 34997 284000 36103 284023
rect 0 268000 41369 284000
rect 673914 283064 673978 283076
rect 675386 283064 675450 283076
rect 673914 283036 675450 283064
rect 673914 283024 673978 283036
rect 675386 283024 675450 283036
rect 41782 281364 41846 281376
rect 42426 281364 42490 281376
rect 42794 281364 42858 281376
rect 41782 281336 42858 281364
rect 41782 281324 41846 281336
rect 42426 281324 42490 281336
rect 42794 281324 42858 281336
rect 676231 280400 717600 296400
rect 681497 280377 682603 280400
rect 683624 280377 684745 280400
rect 687844 280388 696516 280400
rect 687844 280377 692186 280388
tri 692186 280377 692197 280388 nw
rect 696779 280371 703644 280400
rect 703855 280371 711618 280400
rect 713380 280396 713795 280400
rect 41782 274564 41846 274576
rect 42610 274564 42674 274576
rect 41782 274536 42674 274564
rect 41782 274524 41846 274536
rect 42610 274524 42674 274536
rect 41782 271912 41846 271924
rect 42702 271912 42766 271924
rect 41782 271884 42766 271912
rect 41782 271872 41846 271884
rect 42702 271872 42766 271884
rect 5982 267977 13745 268000
rect 13956 267977 20821 268000
rect 21704 267971 22050 268000
rect 23873 267977 28562 268000
rect 689038 251400 693727 251423
rect 695550 251400 695896 251429
rect 696779 251400 703644 251423
rect 703855 251400 711618 251423
rect 673454 248588 673518 248600
rect 674006 248588 674070 248600
rect 675386 248588 675450 248600
rect 673454 248560 675450 248588
rect 673454 248548 673518 248560
rect 674006 248548 674070 248560
rect 675386 248548 675450 248560
rect 673546 244916 673610 244928
rect 675386 244916 675450 244928
rect 673546 244888 675450 244916
rect 673546 244876 673610 244888
rect 675386 244876 675450 244888
rect 3805 240800 4220 240804
rect 5982 240800 13745 240829
rect 13956 240800 20821 240829
tri 25403 240812 25414 240823 se
rect 25414 240812 29756 240823
rect 21084 240800 29756 240812
rect 32855 240800 33976 240823
rect 34997 240800 36103 240823
rect 0 224800 41369 240800
rect 41782 238116 41846 238128
rect 42426 238116 42490 238128
rect 41782 238088 42490 238116
rect 41782 238076 41846 238088
rect 42426 238076 42490 238088
rect 673914 237708 673978 237720
rect 675386 237708 675450 237720
rect 673914 237680 675450 237708
rect 673914 237668 673978 237680
rect 675386 237668 675450 237680
rect 676231 235400 717600 251400
rect 681497 235377 682603 235400
rect 683624 235377 684745 235400
rect 687844 235388 696516 235400
rect 687844 235377 692186 235388
tri 692186 235377 692197 235388 nw
rect 696779 235371 703644 235400
rect 703855 235371 711618 235400
rect 713380 235396 713795 235400
rect 41782 231724 41846 231736
rect 42518 231724 42582 231736
rect 41782 231696 42582 231724
rect 41782 231684 41846 231696
rect 42518 231684 42582 231696
rect 41782 228664 41846 228676
rect 42610 228664 42674 228676
rect 41782 228636 42674 228664
rect 41782 228624 41846 228636
rect 42610 228624 42674 228636
rect 42242 227508 42306 227520
rect 42518 227508 42582 227520
rect 42242 227480 42582 227508
rect 42242 227468 42306 227480
rect 42518 227468 42582 227480
rect 5982 224777 13745 224800
rect 13956 224777 20821 224800
rect 21704 224771 22050 224800
rect 23873 224777 28562 224800
rect 689038 206200 693727 206223
rect 695550 206200 695896 206229
rect 696779 206200 703644 206223
rect 703855 206200 711618 206223
rect 674006 202348 674070 202360
rect 675386 202348 675450 202360
rect 674006 202320 675450 202348
rect 674006 202308 674070 202320
rect 675386 202308 675450 202320
rect 673546 199288 673610 199300
rect 675386 199288 675450 199300
rect 673546 199260 675450 199288
rect 673546 199248 673610 199260
rect 675386 199248 675450 199260
rect 3805 197600 4220 197604
rect 5982 197600 13745 197629
rect 13956 197600 20821 197629
tri 25403 197612 25414 197623 se
rect 25414 197612 29756 197623
rect 21084 197600 29756 197612
rect 32855 197600 33976 197623
rect 34997 197600 36103 197623
rect 0 181600 41369 197600
rect 41782 195888 41846 195900
rect 42518 195888 42582 195900
rect 41782 195860 42582 195888
rect 41782 195848 41846 195860
rect 42518 195848 42582 195860
rect 673914 191944 673978 191956
rect 675386 191944 675450 191956
rect 673914 191916 675450 191944
rect 673914 191904 673978 191916
rect 675386 191904 675450 191916
rect 676231 190200 717600 206200
rect 681497 190177 682603 190200
rect 683624 190177 684745 190200
rect 687844 190188 696516 190200
rect 687844 190177 692186 190188
tri 692186 190177 692197 190188 nw
rect 696779 190171 703644 190200
rect 703855 190171 711618 190200
rect 713380 190196 713795 190200
rect 41966 187592 42030 187604
rect 42518 187592 42582 187604
rect 41966 187564 42582 187592
rect 41966 187552 42030 187564
rect 42518 187552 42582 187564
rect 41782 184464 41846 184476
rect 42610 184464 42674 184476
rect 41782 184436 42674 184464
rect 41782 184424 41846 184436
rect 42260 184204 42288 184436
rect 42610 184424 42674 184436
rect 42242 184152 42306 184204
rect 5982 181577 13745 181600
rect 13956 181577 20821 181600
rect 21704 181571 22050 181600
rect 23873 181577 28562 181600
rect 689038 161200 693727 161223
rect 695550 161200 695896 161229
rect 696779 161200 703644 161223
rect 703855 161200 711618 161223
rect 673454 158352 673518 158364
rect 674006 158352 674070 158364
rect 675386 158352 675450 158364
rect 673454 158324 675450 158352
rect 673454 158312 673518 158324
rect 674006 158312 674070 158324
rect 675386 158312 675450 158324
rect 673546 155224 673610 155236
rect 675386 155224 675450 155236
rect 673546 155196 675450 155224
rect 673546 155184 673610 155196
rect 675386 155184 675450 155196
rect 673730 146928 673794 146940
rect 673914 146928 673978 146940
rect 675386 146928 675450 146940
rect 673730 146900 675450 146928
rect 673730 146888 673794 146900
rect 673914 146888 673978 146900
rect 675386 146888 675450 146900
rect 676231 145200 717600 161200
rect 681497 145177 682603 145200
rect 683624 145177 684745 145200
rect 687844 145188 696516 145200
rect 687844 145177 692186 145188
tri 692186 145177 692197 145188 nw
rect 696779 145171 703644 145200
rect 703855 145171 711618 145200
rect 713380 145196 713795 145200
rect 55 124336 39593 124783
rect 55 124108 39806 124336
rect 55 112870 39593 124108
tri 39593 124085 39616 124108 ne
tri 39593 112870 39616 112893 se
rect 39616 112870 39806 124108
rect 42518 121496 42582 121508
rect 44174 121496 44238 121508
rect 42518 121468 44238 121496
rect 42518 121456 42582 121468
rect 44174 121456 44238 121468
rect 689038 116000 693727 116023
rect 695550 116000 695896 116029
rect 696779 116000 703644 116023
rect 703855 116000 711618 116023
rect 673454 113200 673518 113212
rect 675386 113200 675450 113212
rect 673454 113172 675450 113200
rect 673454 113160 673518 113172
rect 675386 113160 675450 113172
rect 55 112607 39806 112870
rect 55 111971 39593 112607
rect 55 110925 39774 111971
rect 55 110237 39593 110925
rect 673546 109528 673610 109540
rect 675386 109528 675450 109540
rect 673546 109500 675450 109528
rect 673546 109488 673610 109500
rect 675386 109488 675450 109500
rect 673730 101708 673794 101720
rect 675386 101708 675450 101720
rect 673730 101680 675450 101708
rect 673730 101668 673794 101680
rect 675386 101668 675450 101680
rect 676231 100000 717600 116000
rect 681497 99977 682603 100000
rect 683624 99977 684745 100000
rect 687844 99988 696516 100000
rect 687844 99977 692186 99988
tri 692186 99977 692197 99988 nw
rect 696779 99971 703644 100000
rect 703855 99971 711618 100000
rect 713380 99996 713795 100000
rect 31928 85187 32702 85239
rect 31928 84387 40900 85187
tri 40900 84387 41700 85187 sw
rect 31928 83240 41700 84387
rect 31928 83049 32702 83240
rect 32 79313 39593 83000
rect 39756 79313 41700 83240
rect 42426 82872 42490 82884
rect 44174 82872 44238 82884
rect 42426 82844 44238 82872
rect 42426 82832 42490 82844
rect 44174 82832 44238 82844
rect 32 72099 41700 79313
rect 32 71331 39600 72099
rect 39796 71731 41700 72099
tri 39796 71331 40196 71731 ne
rect 40196 71331 41300 71731
tri 41300 71331 41700 71731 nw
rect 32 68024 39593 71331
rect 44818 46968 44882 46980
rect 44818 46940 187694 46968
rect 44818 46928 44882 46940
rect 149072 46912 149100 46940
rect 149054 46860 149118 46912
rect 187666 46900 187694 46940
rect 200868 46940 297772 46968
rect 200868 46912 200896 46940
rect 188522 46900 188586 46912
rect 187666 46872 188586 46900
rect 188522 46860 188586 46872
rect 200850 46860 200914 46912
rect 240888 46900 240916 46940
rect 297744 46912 297772 46940
rect 309428 46940 352604 46968
rect 309428 46912 309456 46940
rect 352576 46912 352604 46940
rect 364260 46940 407436 46968
rect 364260 46912 364288 46940
rect 407408 46912 407436 46940
rect 419092 46940 462176 46968
rect 419092 46912 419120 46940
rect 462148 46912 462176 46940
rect 473832 46940 517008 46968
rect 473832 46912 473860 46940
rect 516980 46912 517008 46940
rect 256234 46900 256298 46912
rect 240888 46872 256298 46900
rect 256234 46860 256298 46872
rect 297726 46860 297790 46912
rect 309410 46860 309474 46912
rect 352558 46860 352622 46912
rect 364242 46860 364306 46912
rect 407390 46860 407454 46912
rect 419074 46860 419138 46912
rect 462130 46860 462194 46912
rect 473814 46860 473878 46912
rect 516962 46860 517026 46912
rect 42242 45608 42306 45620
rect 140958 45608 141022 45620
rect 42242 45580 141022 45608
rect 42242 45568 42306 45580
rect 140958 45568 141022 45580
rect 523770 45608 523834 45620
rect 673546 45608 673610 45620
rect 523770 45580 673610 45608
rect 523770 45568 523834 45580
rect 673546 45568 673610 45580
rect 44910 45540 44974 45552
rect 195974 45540 196038 45552
rect 44910 45512 196038 45540
rect 44910 45500 44974 45512
rect 195974 45500 196038 45512
rect 518710 45540 518774 45552
rect 673730 45540 673794 45552
rect 518710 45512 673794 45540
rect 518710 45500 518774 45512
rect 673730 45500 673794 45512
rect 195974 44452 196038 44464
rect 304534 44452 304598 44464
rect 306282 44452 306346 44464
rect 195974 44424 306346 44452
rect 195974 44412 196038 44424
rect 304534 44412 304598 44424
rect 306282 44412 306346 44424
rect 406746 44452 406810 44464
rect 461486 44452 461550 44464
rect 406746 44424 461550 44452
rect 406746 44412 406810 44424
rect 461486 44412 461550 44424
rect 468938 44452 469002 44464
rect 523770 44452 523834 44464
rect 468938 44424 523834 44452
rect 468938 44412 469002 44424
rect 523770 44412 523834 44424
rect 351914 44384 351978 44396
rect 354398 44384 354462 44396
rect 360562 44384 360626 44396
rect 322906 44356 380894 44384
rect 188522 44316 188586 44328
rect 192846 44316 192910 44328
rect 201494 44316 201558 44328
rect 297082 44316 297146 44328
rect 299566 44316 299630 44328
rect 305730 44316 305794 44328
rect 322906 44316 322934 44356
rect 351914 44344 351978 44356
rect 354398 44344 354462 44356
rect 360562 44344 360626 44356
rect 188522 44288 322934 44316
rect 188522 44276 188586 44288
rect 192846 44276 192910 44288
rect 201494 44276 201558 44288
rect 297082 44276 297146 44288
rect 299566 44276 299630 44288
rect 305730 44276 305794 44288
rect 186682 44248 186746 44260
rect 194686 44248 194750 44260
rect 186682 44220 194750 44248
rect 186682 44208 186746 44220
rect 194686 44208 194750 44220
rect 380866 44316 380894 44356
rect 406746 44316 406810 44328
rect 380866 44288 406810 44316
rect 359366 44248 359430 44260
rect 406746 44276 406810 44288
rect 468938 44316 469002 44328
rect 419506 44288 469002 44316
rect 350000 44220 361574 44248
rect 295242 44180 295306 44192
rect 303246 44180 303310 44192
rect 295242 44152 303310 44180
rect 295242 44140 295306 44152
rect 303246 44140 303310 44152
rect 306282 44180 306346 44192
rect 350000 44180 350028 44220
rect 359366 44208 359430 44220
rect 306282 44152 350028 44180
rect 350074 44180 350138 44192
rect 358078 44180 358142 44192
rect 350074 44152 358142 44180
rect 361546 44180 361574 44220
rect 414198 44180 414262 44192
rect 419506 44180 419534 44288
rect 468938 44276 469002 44288
rect 461486 44248 461550 44260
rect 516318 44248 516382 44260
rect 518710 44248 518774 44260
rect 461486 44220 518774 44248
rect 461486 44208 461550 44220
rect 516318 44208 516382 44220
rect 518710 44208 518774 44220
rect 361546 44152 419534 44180
rect 306282 44140 306346 44152
rect 350074 44140 350138 44152
rect 358078 44140 358142 44152
rect 414198 44140 414262 44152
rect 579890 42752 579954 42764
rect 673454 42752 673518 42764
rect 579890 42724 673518 42752
rect 579890 42712 579954 42724
rect 673454 42712 673518 42724
rect 189258 41936 189322 41948
rect 191098 41936 191162 41948
rect 192294 41936 192358 41948
rect 193582 41936 193646 41948
rect 196434 41936 196498 41948
rect 189258 41908 196498 41936
rect 189258 41896 189322 41908
rect 191098 41896 191162 41908
rect 192294 41896 192358 41908
rect 193582 41896 193646 41908
rect 196434 41896 196498 41908
rect 198458 41936 198522 41948
rect 200114 41936 200178 41948
rect 198458 41908 200178 41936
rect 198458 41896 198522 41908
rect 200114 41896 200178 41908
rect 297910 41936 297974 41948
rect 300670 41936 300734 41948
rect 297910 41908 300734 41936
rect 297910 41896 297974 41908
rect 300670 41896 300734 41908
rect 302234 41936 302298 41948
rect 305270 41936 305334 41948
rect 306558 41936 306622 41948
rect 308674 41936 308738 41948
rect 302234 41908 308738 41936
rect 302234 41896 302298 41908
rect 305270 41896 305334 41908
rect 306558 41896 306622 41908
rect 308674 41896 308738 41908
rect 352650 41936 352714 41948
rect 355502 41936 355566 41948
rect 352650 41908 355566 41936
rect 352650 41896 352714 41908
rect 355502 41896 355566 41908
rect 356974 41936 357038 41948
rect 359826 41936 359890 41948
rect 361114 41936 361178 41948
rect 363506 41936 363570 41948
rect 356974 41908 363570 41936
rect 356974 41896 357038 41908
rect 359826 41896 359890 41908
rect 361114 41896 361178 41908
rect 363506 41896 363570 41908
rect 407482 41936 407546 41948
rect 410242 41936 410306 41948
rect 411530 41936 411594 41948
rect 414566 41936 414630 41948
rect 415854 41936 415918 41948
rect 418246 41936 418310 41948
rect 407482 41908 418310 41936
rect 407482 41896 407546 41908
rect 410242 41896 410306 41908
rect 411530 41896 411594 41908
rect 414566 41896 414630 41908
rect 415854 41896 415918 41908
rect 418246 41896 418310 41908
rect 462314 41936 462378 41948
rect 465074 41936 465138 41948
rect 466362 41936 466426 41948
rect 469398 41936 469462 41948
rect 470686 41936 470750 41948
rect 473078 41936 473142 41948
rect 462314 41908 473142 41936
rect 462314 41896 462378 41908
rect 465074 41896 465138 41908
rect 466362 41896 466426 41908
rect 469398 41896 469462 41908
rect 470686 41896 470750 41908
rect 473078 41896 473142 41908
rect 517054 41936 517118 41948
rect 519906 41936 519970 41948
rect 521194 41936 521258 41948
rect 524230 41936 524294 41948
rect 525518 41936 525582 41948
rect 527910 41936 527974 41948
rect 517054 41908 527974 41936
rect 517054 41896 517118 41908
rect 519906 41896 519970 41908
rect 521194 41896 521258 41908
rect 524230 41896 524294 41908
rect 525518 41896 525582 41908
rect 527910 41896 527974 41908
rect 147122 41868 147186 41880
rect 568850 41868 568914 41880
rect 579890 41868 579954 41880
rect 147122 41840 579954 41868
rect 147122 41828 147186 41840
rect 568850 41828 568914 41840
rect 579890 41828 579954 41840
rect 198918 41800 198982 41812
rect 307754 41800 307818 41812
rect 362494 41800 362558 41812
rect 168346 41772 380894 41800
rect 93762 41528 93826 41540
rect 168346 41528 168374 41772
rect 198918 41760 198982 41772
rect 307754 41760 307818 41772
rect 362494 41760 362558 41772
rect 93762 41500 168374 41528
rect 93762 41488 93826 41500
tri 239482 41369 239813 41700 se
rect 239813 41369 252469 41700
rect 135162 40236 135226 40248
rect 143534 40236 143598 40248
rect 135162 40208 143598 40236
rect 135162 40196 135226 40208
rect 143534 40196 143598 40208
rect 140990 40100 141054 40112
rect 143066 40100 143130 40112
rect 144546 40100 144610 40112
rect 147122 40100 147186 40112
rect 140990 40072 147186 40100
rect 140990 40060 141054 40072
rect 142586 40000 142614 40072
rect 143066 40060 143130 40072
rect 144546 40060 144610 40072
rect 147122 40060 147186 40072
rect 132600 39878 140940 39963
rect 140996 39934 141048 40000
rect 141104 39878 141313 39963
rect 141369 39934 141499 40000
rect 141555 39878 141898 39963
rect 141954 39934 142084 40000
rect 142140 39878 142517 39963
rect 79664 39616 91393 39806
rect 79664 39593 79892 39616
tri 79892 39593 79915 39616 nw
tri 91107 39593 91130 39616 ne
rect 91130 39593 91393 39616
rect 79076 55 93763 39593
rect 132600 37949 142517 39878
rect 142573 38005 142619 40000
rect 142675 39878 143012 39963
rect 143068 39934 143128 40000
rect 143184 39878 144517 39963
rect 144573 39934 144689 40000
rect 144745 39878 145035 39963
rect 145091 39934 145143 40000
rect 145199 39878 147600 39963
rect 142675 37949 147600 39878
rect 132600 20821 147600 37949
rect 186400 36103 202400 41369
rect 186377 34997 202400 36103
rect 186400 33976 202400 34997
rect 186377 32855 202400 33976
rect 186400 29756 202400 32855
tri 239013 40900 239482 41369 se
rect 239482 41300 252469 41369
tri 252469 41300 252869 41700 sw
rect 380866 41528 380894 41772
rect 417326 41800 417390 41812
rect 417252 41772 417390 41800
rect 417252 41528 417280 41772
rect 417326 41760 417390 41772
rect 472158 41800 472222 41812
rect 526714 41800 526778 41812
rect 472084 41772 472222 41800
rect 472084 41528 472112 41772
rect 472158 41760 472222 41772
rect 516106 41772 526778 41800
rect 516106 41528 516134 41772
rect 526714 41760 526778 41772
rect 380866 41500 516134 41528
rect 239482 40900 252869 41300
rect 239013 40196 252869 40900
rect 239013 39796 252469 40196
tri 252469 39796 252869 40196 nw
rect 239013 39756 252101 39796
rect 239013 32702 240960 39756
rect 244887 39600 252101 39756
rect 244887 39593 252869 39600
rect 238961 31928 241151 32702
rect 186377 28562 202400 29756
rect 186377 25414 202423 28562
tri 186377 25403 186388 25414 ne
rect 186388 23873 202423 25414
rect 186388 22050 202400 23873
rect 186388 21704 202429 22050
rect 186388 21084 202400 21704
rect 186400 20821 202400 21084
rect 132571 13956 147629 20821
rect 186371 13956 202423 20821
rect 132600 13745 147600 13956
rect 186400 13745 202400 13956
rect 132571 5982 147629 13745
rect 186371 5982 202423 13745
rect 132600 158 147600 5982
rect 186400 4220 202400 5982
rect 186396 3805 202400 4220
rect 186400 0 202400 3805
rect 241200 32 256176 39593
rect 295000 36103 311000 41369
rect 349800 36103 365800 41369
rect 404600 36103 420600 41369
rect 459400 36103 475400 41369
rect 514200 36103 530200 41369
rect 569864 39616 581593 39806
rect 569864 39593 570092 39616
tri 570092 39593 570115 39616 nw
tri 581307 39593 581330 39616 ne
rect 581330 39593 581593 39616
rect 623664 39616 635393 39806
rect 623664 39593 623892 39616
tri 623892 39593 623915 39616 nw
tri 635107 39593 635130 39616 ne
rect 635130 39593 635393 39616
rect 636029 39593 637075 39774
rect 294977 34997 311000 36103
rect 349777 34997 365800 36103
rect 404577 34997 420600 36103
rect 459377 34997 475400 36103
rect 514177 34997 530200 36103
rect 295000 33976 311000 34997
rect 349800 33976 365800 34997
rect 404600 33976 420600 34997
rect 459400 33976 475400 34997
rect 514200 33976 530200 34997
rect 294977 32855 311000 33976
rect 349777 32855 365800 33976
rect 404577 32855 420600 33976
rect 459377 32855 475400 33976
rect 514177 32855 530200 33976
rect 295000 29756 311000 32855
rect 349800 29756 365800 32855
rect 404600 29756 420600 32855
rect 459400 29756 475400 32855
rect 514200 29756 530200 32855
rect 294977 28562 311000 29756
rect 349777 28562 365800 29756
rect 404577 28562 420600 29756
rect 459377 28562 475400 29756
rect 514177 28562 530200 29756
rect 294977 25414 311023 28562
tri 294977 25403 294988 25414 ne
rect 294988 23873 311023 25414
rect 349777 25414 365823 28562
tri 349777 25403 349788 25414 ne
rect 349788 23873 365823 25414
rect 404577 25414 420623 28562
tri 404577 25403 404588 25414 ne
rect 404588 23873 420623 25414
rect 459377 25414 475423 28562
tri 459377 25403 459388 25414 ne
rect 459388 23873 475423 25414
rect 514177 25414 530223 28562
tri 514177 25403 514188 25414 ne
rect 514188 23873 530223 25414
rect 294988 22050 311000 23873
rect 349788 22050 365800 23873
rect 404588 22050 420600 23873
rect 459388 22050 475400 23873
rect 514188 22050 530200 23873
rect 294988 21704 311029 22050
rect 349788 21704 365829 22050
rect 404588 21704 420629 22050
rect 459388 21704 475429 22050
rect 514188 21704 530229 22050
rect 294988 21084 311000 21704
rect 349788 21084 365800 21704
rect 404588 21084 420600 21704
rect 459388 21084 475400 21704
rect 514188 21084 530200 21704
rect 295000 20821 311000 21084
rect 349800 20821 365800 21084
rect 404600 20821 420600 21084
rect 459400 20821 475400 21084
rect 514200 20821 530200 21084
rect 294971 13956 311023 20821
rect 349771 13956 365823 20821
rect 404571 13956 420623 20821
rect 459371 13956 475423 20821
rect 514171 13956 530223 20821
rect 295000 13745 311000 13956
rect 349800 13745 365800 13956
rect 404600 13745 420600 13956
rect 459400 13745 475400 13956
rect 514200 13745 530200 13956
rect 294971 5982 311023 13745
rect 349771 5982 365823 13745
rect 404571 5982 420623 13745
rect 459371 5982 475423 13745
rect 514171 5982 530223 13745
rect 295000 4220 311000 5982
rect 349800 4220 365800 5982
rect 404600 4220 420600 5982
rect 459400 4220 475400 5982
rect 514200 4220 530200 5982
rect 294996 3805 311000 4220
rect 349796 3805 365800 4220
rect 404596 3805 420600 4220
rect 459396 3805 475400 4220
rect 514196 3805 530200 4220
rect 295000 0 311000 3805
rect 349800 0 365800 3805
rect 404600 0 420600 3805
rect 459400 0 475400 3805
rect 514200 0 530200 3805
rect 569276 55 583963 39593
rect 623217 55 637763 39593
<< metal2 >>
rect 230499 997600 235279 998011
rect 240478 997600 245258 1002732
rect 282099 997600 286879 998011
rect 292078 997600 296858 1002732
rect 41713 799417 42193 799473
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 795093 42193 795149
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 41713 791466 42193 791469
rect 41713 791438 42288 791466
rect 41713 791413 42193 791438
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 42260 787302 42288 791438
rect 42248 787296 42300 787302
rect 41892 787244 42248 787250
rect 41892 787238 42300 787244
rect 42432 787296 42484 787302
rect 42432 787238 42484 787244
rect 41892 787222 42288 787238
rect 41892 787145 41920 787222
rect 41713 787089 42193 787145
rect 41722 787086 41920 787089
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 41713 784697 42193 784753
rect 41713 756217 42193 756273
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751893 42193 751949
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 41713 748213 42193 748269
rect 41892 747974 41920 748213
rect 42444 747974 42472 787238
rect 41892 747946 42472 747974
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 41713 743889 42193 743945
rect 41800 743730 41828 743889
rect 42260 743730 42288 747946
rect 41800 743702 42288 743730
rect 41713 743337 42193 743393
rect 41713 742693 42193 742749
rect 41713 742049 42193 742105
rect 41713 741497 42193 741553
rect 42260 728654 42288 743702
rect 42260 728626 42380 728654
rect 41713 713017 42193 713073
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708693 42193 708749
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 41713 705013 42193 705069
rect 41892 704970 41920 705013
rect 42352 704970 42380 728626
rect 41892 704942 42380 704970
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 41722 700745 41920 700754
rect 41713 700689 42193 700745
rect 41892 700618 41920 700689
rect 42260 700618 42288 704942
rect 41892 700590 42288 700618
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 41713 698297 42193 698353
rect 42260 690014 42288 700590
rect 42260 689986 42380 690014
rect 41713 669817 42193 669873
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 665493 42193 665549
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 42352 661994 42380 689986
rect 41800 661966 42380 661994
rect 41800 661869 41828 661966
rect 41713 661813 42193 661869
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 42260 657642 42288 661966
rect 673736 870868 673788 870874
rect 673736 870810 673788 870816
rect 673748 786010 673776 870810
rect 673736 786004 673788 786010
rect 673736 785946 673788 785952
rect 673736 781652 673788 781658
rect 673736 781594 673788 781600
rect 673748 740994 673776 781594
rect 673736 740988 673788 740994
rect 673736 740930 673788 740936
rect 41892 657614 42288 657642
rect 41892 657545 41920 657614
rect 41713 657489 42193 657545
rect 41722 657478 41920 657489
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 41713 655097 42193 655153
rect 42260 651374 42288 657614
rect 42260 651346 42380 651374
rect 41713 626617 42193 626673
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 622293 42193 622349
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 42352 618746 42380 651346
rect 41800 618718 42380 618746
rect 41800 618669 41828 618718
rect 41713 618613 42193 618669
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41713 614331 42193 614345
rect 42260 614331 42288 618718
rect 41713 614303 42288 614331
rect 41713 614289 42193 614303
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 42260 612734 42288 614303
rect 42260 612706 42380 612734
rect 41713 612449 42193 612505
rect 41713 611897 42193 611953
rect 41713 583417 42193 583473
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 579093 42193 579149
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 41713 575455 42193 575469
rect 42352 575455 42380 612706
rect 673736 737044 673788 737050
rect 673736 736986 673788 736992
rect 673748 695978 673776 736986
rect 673736 695972 673788 695978
rect 673736 695914 673788 695920
rect 673736 692096 673788 692102
rect 673736 692038 673788 692044
rect 41713 575427 42380 575455
rect 41713 575413 42193 575427
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 42260 571282 42288 575427
rect 41800 571254 42380 571282
rect 41800 571146 41828 571254
rect 41722 571145 41828 571146
rect 41713 571089 42193 571145
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 41713 568697 42193 568753
rect 41713 540217 42193 540273
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535893 42193 535949
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 41713 532213 42193 532269
rect 41892 532114 41920 532213
rect 42352 532114 42380 571254
rect 41892 532086 42380 532114
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 41713 527917 42193 527945
rect 41708 527898 42193 527917
rect 42260 527898 42288 532086
rect 673748 651166 673776 692038
rect 673736 651160 673788 651166
rect 673736 651102 673788 651108
rect 673748 646474 673776 651102
rect 673736 646468 673788 646474
rect 673736 646410 673788 646416
rect 673748 605810 673776 646410
rect 673736 605804 673788 605810
rect 673736 605746 673788 605752
rect 673736 601860 673788 601866
rect 673736 601802 673788 601808
rect 673748 561134 673776 601802
rect 673736 561128 673788 561134
rect 673736 561070 673788 561076
rect 673644 556640 673696 556646
rect 673644 556582 673696 556588
rect 41708 527870 42288 527898
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 41713 525497 42193 525553
rect 42260 419534 42288 527870
rect 42260 419506 42380 419534
rect 41713 412617 42193 412673
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 408293 42193 408349
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 42352 405226 42380 419506
rect 41800 405198 42380 405226
rect 41800 404682 41828 405198
rect 41722 404669 41828 404682
rect 41713 404613 42193 404669
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41713 400330 42193 400345
rect 42260 400330 42288 405198
rect 41713 400302 42288 400330
rect 41713 400289 42193 400302
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 41713 397897 42193 397953
rect 41713 369417 42193 369473
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 365093 42193 365149
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 41713 361434 42193 361469
rect 42260 361434 42288 400302
rect 41713 361413 42288 361434
rect 41722 361406 42288 361413
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41713 357089 42193 357145
rect 41984 356674 42012 357089
rect 42260 356674 42288 361406
rect 41984 356646 42288 356674
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 41713 354697 42193 354753
rect 42260 332602 42288 356646
rect 42260 332574 42380 332602
rect 41713 326217 42193 326273
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321893 42193 321949
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 41713 318255 42193 318269
rect 42352 318255 42380 332574
rect 41713 318227 42380 318255
rect 41713 318213 42193 318227
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 41713 313889 42193 313945
rect 41800 313834 41828 313889
rect 42260 313834 42288 318227
rect 673656 384334 673684 556582
rect 677600 962721 678011 967501
rect 677600 952742 682732 957522
rect 675407 878047 675887 878103
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675407 875697 675887 875711
rect 675312 875669 675887 875697
rect 675312 871373 675340 875669
rect 675407 875655 675887 875669
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 871373 675887 871387
rect 675312 871345 675887 871373
rect 675404 871331 675887 871345
rect 675404 870874 675432 871331
rect 675392 870868 675444 870874
rect 675392 870810 675444 870816
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867651 675887 867707
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675407 863327 675887 863383
rect 675407 788847 675887 788903
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 675407 786483 675887 786511
rect 675404 786455 675887 786483
rect 675404 786010 675432 786455
rect 675208 786004 675260 786010
rect 675208 785946 675260 785952
rect 675392 786004 675444 786010
rect 675392 785946 675444 785952
rect 675220 781658 675248 785946
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 782159 675887 782187
rect 675404 782131 675887 782159
rect 675404 781658 675432 782131
rect 675208 781652 675260 781658
rect 675208 781594 675260 781600
rect 675392 781652 675444 781658
rect 675392 781594 675444 781600
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 778451 675887 778507
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675407 774127 675887 774183
rect 675407 743847 675887 743903
rect 675407 743295 675887 743351
rect 675407 742651 675887 742707
rect 675407 742007 675887 742063
rect 675407 741483 675887 741511
rect 675404 741455 675887 741483
rect 675404 740994 675432 741455
rect 675208 740988 675260 740994
rect 675208 740930 675260 740936
rect 675392 740988 675444 740994
rect 675392 740930 675444 740936
rect 675220 737050 675248 740930
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 737159 675887 737187
rect 675404 737131 675887 737159
rect 675404 737050 675432 737131
rect 675208 737044 675260 737050
rect 675208 736986 675260 736992
rect 675392 737044 675444 737050
rect 675392 736986 675444 736992
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 733451 675887 733507
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675407 729127 675887 729183
rect 675407 698847 675887 698903
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675407 696483 675887 696511
rect 675404 696455 675887 696483
rect 675404 695978 675432 696455
rect 675208 695972 675260 695978
rect 675208 695914 675260 695920
rect 675392 695972 675444 695978
rect 675392 695914 675444 695920
rect 675220 692102 675248 695914
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 692172 675887 692187
rect 675404 692131 675887 692172
rect 675404 692102 675432 692131
rect 675208 692096 675260 692102
rect 675208 692038 675260 692044
rect 675392 692096 675444 692102
rect 675392 692038 675444 692044
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 688451 675887 688507
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675407 684127 675887 684183
rect 675407 653647 675887 653703
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 675407 651283 675887 651311
rect 675404 651255 675887 651283
rect 675404 651166 675432 651255
rect 675392 651160 675444 651166
rect 675392 651102 675444 651108
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 646959 675887 646987
rect 675404 646931 675887 646959
rect 675404 646474 675432 646931
rect 675392 646468 675444 646474
rect 675392 646410 675444 646416
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 643251 675887 643307
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675407 638927 675887 638983
rect 675407 608647 675887 608703
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 675407 606283 675887 606311
rect 675404 606255 675887 606283
rect 675404 605810 675432 606255
rect 675208 605804 675260 605810
rect 675208 605746 675260 605752
rect 675392 605804 675444 605810
rect 675392 605746 675444 605752
rect 675220 601866 675248 605746
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 601959 675887 601987
rect 675404 601931 675887 601959
rect 675404 601866 675432 601931
rect 675208 601860 675260 601866
rect 675208 601802 675260 601808
rect 675392 601860 675444 601866
rect 675392 601802 675444 601808
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 598251 675887 598307
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675407 593927 675887 593983
rect 675407 563447 675887 563503
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 675220 561134 675248 561165
rect 675208 561128 675260 561134
rect 675407 561082 675887 561111
rect 675260 561076 675887 561082
rect 675208 561070 675887 561076
rect 675220 561055 675887 561070
rect 675220 561054 675418 561055
rect 675220 556646 675248 561054
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675407 556759 675887 556787
rect 675404 556731 675887 556759
rect 675404 556646 675432 556731
rect 675208 556640 675260 556646
rect 675208 556582 675260 556588
rect 675392 556640 675444 556646
rect 675392 556582 675444 556588
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 553051 675887 553107
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675407 548727 675887 548783
rect 675407 386247 675887 386303
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 673644 384328 673696 384334
rect 673644 384270 673696 384276
rect 675392 384328 675444 384334
rect 675392 384270 675444 384276
rect 675404 384010 675432 384270
rect 675312 383982 675432 384010
rect 673644 379092 673696 379098
rect 673644 379034 673696 379040
rect 673656 338842 673684 379034
rect 673644 338836 673696 338842
rect 673644 338778 673696 338784
rect 41800 313806 42288 313834
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 41713 311497 42193 311553
rect 42260 303614 42288 313806
rect 42260 303586 42380 303614
rect 41713 283017 42193 283073
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278693 42193 278749
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 42352 275210 42380 303586
rect 41800 275182 42380 275210
rect 41800 275074 41828 275182
rect 41722 275069 41828 275074
rect 41713 275013 42193 275069
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 42260 270858 42288 275182
rect 41892 270830 42288 270858
rect 41892 270745 41920 270830
rect 41713 270689 42193 270745
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 41713 268297 42193 268353
rect 42260 264974 42288 270830
rect 42260 264946 42380 264974
rect 41713 239817 42193 239873
rect 41713 237977 42193 238033
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 41713 231855 42193 231869
rect 42352 231855 42380 264946
rect 41713 231827 42380 231855
rect 41713 231813 42193 231827
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 42260 227610 42288 231827
rect 41800 227582 42380 227610
rect 41800 227545 41828 227582
rect 41713 227489 42193 227545
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 41713 225097 42193 225153
rect 42352 197554 42380 227582
rect 675312 379573 675340 383982
rect 675404 383911 675432 383982
rect 675404 383860 675887 383911
rect 675407 383855 675887 383860
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675407 379573 675887 379587
rect 675312 379545 675887 379573
rect 675404 379531 675887 379545
rect 675404 379098 675432 379531
rect 675392 379092 675444 379098
rect 675392 379034 675444 379040
rect 673828 334280 673880 334286
rect 673828 334222 673880 334228
rect 673840 294710 673868 334222
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675407 371527 675887 371583
rect 675407 341047 675887 341103
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675392 338836 675444 338842
rect 675392 338778 675444 338784
rect 675404 338711 675432 338778
rect 675404 338655 675887 338711
rect 675404 338178 675432 338655
rect 675312 338150 675432 338178
rect 673828 294704 673880 294710
rect 673828 294646 673880 294652
rect 673644 288856 673696 288862
rect 673644 288798 673696 288804
rect 673656 249150 673684 288798
rect 675312 334370 675340 338150
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 334370 675887 334387
rect 675312 334342 675887 334370
rect 675404 334331 675887 334342
rect 675404 334286 675432 334331
rect 675392 334280 675444 334286
rect 675392 334222 675444 334228
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675407 326327 675887 326383
rect 675407 296047 675887 296103
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675300 294704 675352 294710
rect 675300 294646 675352 294652
rect 675312 293706 675340 294646
rect 675407 294207 675887 294263
rect 675407 293706 675887 293711
rect 675312 293678 675887 293706
rect 675312 289354 675340 293678
rect 675407 293655 675887 293678
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 289354 675887 289387
rect 675312 289331 675887 289354
rect 675312 289326 675432 289331
rect 675404 288862 675432 289326
rect 675392 288856 675444 288862
rect 675392 288798 675444 288804
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 675407 281327 675887 281383
rect 673644 249144 673696 249150
rect 673644 249086 673696 249092
rect 42352 197526 42472 197554
rect 41713 196617 42193 196673
rect 41713 194777 42193 194833
rect 41713 192937 42193 192993
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 41788 189168 41840 189174
rect 41788 189110 41840 189116
rect 41800 188669 41828 189110
rect 41713 188613 42193 188669
rect 42444 189174 42472 197526
rect 42432 189168 42484 189174
rect 42432 189110 42484 189116
rect 42444 188034 42472 189110
rect 42260 188006 42472 188034
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 41713 184331 42193 184345
rect 42260 184331 42288 188006
rect 41713 184303 42380 184331
rect 41713 184289 42193 184303
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 41713 181897 42193 181953
rect 42352 47025 42380 184303
rect 673828 243840 673880 243846
rect 673828 243782 673880 243788
rect 673840 203522 673868 243782
rect 675407 251047 675887 251103
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675392 249144 675444 249150
rect 675392 249086 675444 249092
rect 675404 248711 675432 249086
rect 675404 248690 675887 248711
rect 675312 248662 675887 248690
rect 673828 203516 673880 203522
rect 673828 203458 673880 203464
rect 673736 199096 673788 199102
rect 673736 199038 673788 199044
rect 673748 158642 673776 199038
rect 675312 244373 675340 248662
rect 675407 248655 675887 248662
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 244373 675887 244387
rect 675312 244345 675887 244373
rect 675404 244331 675887 244345
rect 675404 243846 675432 244331
rect 675392 243840 675444 243846
rect 675392 243782 675444 243788
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 675407 238167 675887 238223
rect 675407 236327 675887 236383
rect 675407 205847 675887 205903
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 675312 203522 675340 203580
rect 675300 203516 675352 203522
rect 675407 203497 675887 203511
rect 675352 203469 675887 203497
rect 675300 203458 675352 203464
rect 673736 158636 673788 158642
rect 673736 158578 673788 158584
rect 42338 47016 42394 47025
rect 42338 46951 42394 46960
rect 52460 46912 52512 46918
rect 52458 46880 52460 46889
rect 143540 46912 143592 46918
rect 52512 46880 52514 46889
rect 143540 46854 143592 46860
rect 527456 46912 527508 46918
rect 527456 46854 527508 46860
rect 52458 46815 52514 46824
rect 143552 44198 143580 46854
rect 143540 44192 143592 44198
rect 143540 44134 143592 44140
rect 145104 44192 145156 44198
rect 145104 44134 145156 44140
rect 145116 40202 145144 44134
rect 145103 40174 145144 40202
rect 145103 40000 145131 40174
rect 195336 44192 195388 44198
rect 195336 44134 195388 44140
rect 195348 42193 195376 44134
rect 199660 44192 199712 44198
rect 199660 44134 199712 44140
rect 199672 42193 199700 44134
rect 187327 41713 187383 42193
rect 194043 41713 194099 42193
rect 195331 41713 195387 42193
rect 199655 41713 199711 42193
rect 145091 39706 145143 40000
rect 303896 44260 303948 44266
rect 303896 44202 303948 44208
rect 303908 42193 303936 44202
rect 308220 44260 308272 44266
rect 308220 44202 308272 44208
rect 308232 42193 308260 44202
rect 358728 44328 358780 44334
rect 358728 44270 358780 44276
rect 358740 42193 358768 44270
rect 363052 44328 363104 44334
rect 363052 44270 363104 44276
rect 363064 42193 363092 44270
rect 411074 44432 411130 44441
rect 411074 44367 411130 44376
rect 411088 42193 411116 44367
rect 413560 44260 413612 44266
rect 413560 44202 413612 44208
rect 417884 44260 417936 44266
rect 417884 44202 417936 44208
rect 413572 42193 413600 44202
rect 417896 42193 417924 44202
rect 419722 44432 419778 44441
rect 419722 44367 419778 44376
rect 419736 42193 419764 44367
rect 465814 44432 465870 44441
rect 465814 44367 465870 44376
rect 468300 44396 468352 44402
rect 465828 42193 465856 44367
rect 468300 44338 468352 44344
rect 468312 42193 468340 44338
rect 472624 44396 472676 44402
rect 472624 44338 472676 44344
rect 472636 42193 472664 44338
rect 474462 44432 474518 44441
rect 474462 44367 474518 44376
rect 474476 42193 474504 44367
rect 518806 44296 518862 44305
rect 518806 44231 518862 44240
rect 518820 42193 518848 44231
rect 523132 44192 523184 44198
rect 523132 44134 523184 44140
rect 523144 42193 523172 44134
rect 524970 44296 525026 44305
rect 524970 44231 525026 44240
rect 524984 42193 525012 44231
rect 527468 44198 527496 46854
rect 527456 44192 527508 44198
rect 527456 44134 527508 44140
rect 527468 42193 527496 44134
rect 673644 154148 673696 154154
rect 673644 154090 673696 154096
rect 673656 113762 673684 154090
rect 675312 199186 675340 203458
rect 675407 203455 675887 203469
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 199186 675887 199187
rect 675312 199158 675887 199186
rect 675404 199131 675887 199158
rect 675404 199102 675432 199131
rect 675392 199096 675444 199102
rect 675392 199038 675444 199044
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 675407 194807 675887 194863
rect 675407 192967 675887 193023
rect 675407 191127 675887 191183
rect 675407 160847 675887 160903
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675392 158636 675444 158642
rect 675392 158578 675444 158584
rect 675404 158522 675432 158578
rect 675312 158511 675432 158522
rect 675312 158494 675887 158511
rect 675312 154170 675340 158494
rect 675407 158455 675887 158494
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 154170 675887 154187
rect 675312 154154 675887 154170
rect 675300 154148 675887 154154
rect 675352 154142 675887 154148
rect 675407 154131 675887 154142
rect 675300 154090 675352 154096
rect 675312 154059 675340 154090
rect 673644 113756 673696 113762
rect 673644 113698 673696 113704
rect 673644 108452 673696 108458
rect 673644 108394 673696 108400
rect 673656 46986 673684 108394
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675407 146127 675887 146183
rect 675407 115647 675887 115703
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675392 113756 675444 113762
rect 675392 113698 675444 113704
rect 675404 113311 675432 113698
rect 675404 113297 675887 113311
rect 675312 113269 675887 113297
rect 675312 108973 675340 113269
rect 675407 113255 675887 113269
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675407 108973 675887 108987
rect 675312 108945 675887 108973
rect 675404 108931 675887 108945
rect 675404 108458 675432 108931
rect 675392 108452 675444 108458
rect 675392 108394 675444 108400
rect 673644 46980 673696 46986
rect 673644 46922 673696 46928
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675407 100927 675887 100983
rect 302643 41713 302699 42193
rect 303908 41806 303987 42193
rect 303931 41713 303987 41806
rect 306967 41713 307023 42193
rect 308232 41806 308311 42193
rect 308255 41713 308311 41806
rect 310095 41713 310151 42193
rect 357443 41713 357499 42193
rect 358731 41713 358787 42193
rect 361767 41713 361823 42193
rect 363055 41713 363111 42193
rect 364895 41713 364951 42193
rect 405527 41713 405583 42193
rect 409207 41834 409263 42193
rect 409207 41818 409368 41834
rect 409207 41812 409380 41818
rect 409207 41806 409328 41812
rect 409207 41713 409263 41806
rect 409328 41754 409380 41760
rect 411047 41820 411116 42193
rect 411047 41713 411103 41820
rect 412243 41834 412299 42193
rect 412243 41818 412404 41834
rect 413531 41820 413600 42193
rect 415371 41834 415427 42193
rect 412243 41812 412416 41818
rect 412243 41806 412364 41812
rect 412243 41713 412299 41806
rect 412364 41754 412416 41760
rect 413531 41713 413587 41820
rect 415228 41818 415427 41834
rect 415216 41812 415427 41818
rect 415268 41806 415427 41812
rect 415216 41754 415268 41760
rect 415371 41713 415427 41806
rect 416567 41713 416623 42193
rect 417855 41820 417924 42193
rect 419695 41820 419764 42193
rect 417855 41713 417911 41820
rect 419695 41713 419751 41820
rect 460327 41713 460383 42193
rect 464007 41834 464063 42193
rect 464007 41818 464200 41834
rect 464007 41812 464212 41818
rect 464007 41806 464160 41812
rect 464007 41713 464063 41806
rect 464160 41754 464212 41760
rect 465828 41806 465903 42193
rect 465847 41713 465903 41806
rect 467043 41834 467099 42193
rect 467043 41818 467236 41834
rect 467043 41812 467248 41818
rect 467043 41806 467196 41812
rect 467043 41713 467099 41806
rect 468312 41806 468387 42193
rect 470171 41834 470227 42193
rect 470060 41818 470227 41834
rect 467196 41754 467248 41760
rect 468331 41713 468387 41806
rect 470048 41812 470227 41818
rect 470100 41806 470227 41812
rect 470048 41754 470100 41760
rect 470171 41713 470227 41806
rect 471367 41713 471423 42193
rect 472636 41806 472711 42193
rect 474476 41806 474551 42193
rect 472655 41713 472711 41806
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 518807 41713 518863 42193
rect 520647 41713 520703 42193
rect 521843 41713 521899 42193
rect 523131 41713 523187 42193
rect 524971 41713 525027 42193
rect 526167 41713 526223 42193
rect 527455 41713 527511 42193
rect 529295 41713 529351 42193
<< via2 >>
rect 42338 46960 42394 47016
rect 52458 46860 52460 46880
rect 52460 46860 52512 46880
rect 52512 46860 52514 46880
rect 52458 46824 52514 46860
rect 411074 44376 411130 44432
rect 419722 44376 419778 44432
rect 465814 44376 465870 44432
rect 474462 44376 474518 44432
rect 518806 44240 518862 44296
rect 524970 44240 525026 44296
<< obsm2 >>
rect 77050 1006851 90288 1007371
rect 128450 1006851 141688 1007371
rect 179850 1006851 193088 1007371
rect 230453 1002788 245258 1036615
rect 282053 1002788 296858 1036615
rect 230453 998067 240422 1002788
rect 235335 998007 240422 998067
rect 235579 997600 235979 997984
rect 282053 998067 292022 1002788
rect 286935 998007 292022 998067
rect 287179 997600 287579 997984
rect 333453 998007 348258 1036615
rect 384650 1006851 397888 1007371
rect 473650 1006851 486888 1007371
rect 525050 1006851 538288 1007371
rect 575653 998007 590458 1036615
rect 626850 1006851 640088 1007371
rect 333499 997600 338279 998007
rect 338579 997600 338979 997984
rect 343478 997600 348258 998007
rect 575699 997600 580479 998007
rect 580779 997600 581179 997984
rect 585678 997600 590458 998007
rect 585046 997455 585102 997529
rect 343638 997047 343694 997121
rect 42248 990150 42300 990214
rect 30229 955050 30749 968288
rect 7 927240 30281 929187
rect 30753 927000 31683 929228
rect 32033 927240 34915 929187
rect 7 926940 39593 927000
rect 7 922819 39600 926940
rect 7 922707 39593 922819
rect 7 916185 39600 922707
rect 7 916099 39593 916185
rect 7 912100 39600 916099
rect 7 912000 39593 912100
rect 30760 909805 31690 912000
rect 985 879878 40000 884658
rect 985 874679 39593 879878
rect 39616 874979 40000 875379
rect 985 869899 40000 874679
rect 985 869853 39593 869899
rect 985 837678 40000 842458
rect 985 832479 39593 837678
rect 39616 832779 40000 833179
rect 985 827699 40000 832479
rect 985 827653 39593 827699
rect 0 800173 41713 800383
rect 0 800005 41657 800173
rect 42260 800170 42288 990150
rect 343652 990146 343680 997047
rect 585060 996402 585088 997455
rect 585048 996338 585100 996402
rect 674748 996338 674800 996402
rect 356060 990830 356112 990894
rect 673552 990830 673604 990894
rect 356072 990146 356100 990830
rect 44916 990082 44968 990146
rect 343640 990082 343692 990146
rect 356060 990082 356112 990146
rect 44928 888734 44956 990082
rect 673460 990014 673512 990078
rect 44836 888706 44956 888734
rect 44836 870097 44864 888706
rect 673472 872438 673500 990014
rect 673564 874546 673592 990830
rect 673552 874482 673604 874546
rect 673460 872374 673512 872438
rect 42338 870023 42394 870097
rect 44822 870023 44878 870097
rect 42352 805934 42380 870023
rect 673460 864214 673512 864278
rect 42352 805906 42472 805934
rect 42260 800142 42380 800170
rect 41713 800103 42193 800117
rect 41713 800075 42288 800103
rect 41713 800061 42193 800075
rect 0 799529 41713 800005
rect 0 799361 41657 799529
rect 0 798885 41713 799361
rect 0 798717 41657 798885
rect 41713 798773 42193 798829
rect 0 798333 41713 798717
rect 0 798165 41657 798333
rect 41713 798221 42193 798277
rect 0 797689 41713 798165
rect 41800 797774 41828 798221
rect 41788 797710 41840 797774
rect 0 797521 41657 797689
rect 0 797045 41713 797521
rect 0 796877 41657 797045
rect 0 796493 41713 796877
rect 0 796325 41657 796493
rect 41713 796381 42193 796437
rect 0 795849 41713 796325
rect 0 795681 41657 795849
rect 0 795205 41713 795681
rect 0 795037 41657 795205
rect 0 794653 41713 795037
rect 0 794485 41657 794653
rect 0 794009 41713 794485
rect 0 793841 41657 794009
rect 0 793365 41713 793841
rect 0 793197 41657 793365
rect 0 792813 41713 793197
rect 0 792645 41657 792813
rect 0 792169 41713 792645
rect 42260 792282 42288 800075
rect 41892 792254 42288 792282
rect 0 792001 41657 792169
rect 41892 792113 41920 792254
rect 41713 792057 42193 792113
rect 0 791525 41713 792001
rect 0 791357 41657 791525
rect 0 790881 41713 791357
rect 41788 791318 41840 791382
rect 0 790713 41657 790881
rect 41800 790825 41828 791318
rect 41713 790769 42193 790825
rect 41722 790758 41828 790769
rect 0 790329 41713 790713
rect 0 790161 41657 790329
rect 0 789685 41713 790161
rect 0 789517 41657 789685
rect 0 789041 41713 789517
rect 0 788873 41657 789041
rect 0 788489 41713 788873
rect 0 788321 41657 788489
rect 0 787845 41713 788321
rect 41788 788258 41840 788322
rect 0 787677 41657 787845
rect 41800 787794 41828 788258
rect 41722 787789 41828 787794
rect 41713 787733 42193 787789
rect 0 787201 41713 787677
rect 41800 787302 41828 787733
rect 42352 788322 42380 800142
rect 42444 791382 42472 805906
rect 42616 797710 42668 797774
rect 42432 791318 42484 791382
rect 42340 788258 42392 788322
rect 42444 787386 42472 791318
rect 42444 787358 42564 787386
rect 41788 787238 41840 787302
rect 0 787033 41657 787201
rect 42248 787034 42300 787098
rect 0 786649 41713 787033
rect 0 786481 41657 786649
rect 0 786005 41713 786481
rect 0 785837 41657 786005
rect 0 785361 41713 785837
rect 0 785193 41657 785361
rect 0 784809 41713 785193
rect 0 784641 41657 784809
rect 0 784442 41713 784641
rect 42260 757654 42288 787034
rect 42340 786966 42392 787030
rect 42248 757590 42300 757654
rect 42352 757586 42380 786966
rect 42340 757522 42392 757586
rect 0 756973 41713 757183
rect 0 756805 41657 756973
rect 41722 756917 42288 756922
rect 41713 756894 42288 756917
rect 41713 756861 42193 756894
rect 0 756329 41713 756805
rect 0 756161 41657 756329
rect 0 755685 41713 756161
rect 0 755517 41657 755685
rect 41713 755573 42193 755629
rect 0 755133 41713 755517
rect 41788 755414 41840 755478
rect 0 754965 41657 755133
rect 41800 755077 41828 755414
rect 41713 755021 42193 755077
rect 0 754489 41713 754965
rect 0 754321 41657 754489
rect 0 753845 41713 754321
rect 0 753677 41657 753845
rect 0 753293 41713 753677
rect 0 753125 41657 753293
rect 41713 753181 42193 753237
rect 0 752649 41713 753125
rect 0 752481 41657 752649
rect 0 752005 41713 752481
rect 0 751837 41657 752005
rect 0 751453 41713 751837
rect 0 751285 41657 751453
rect 0 750809 41713 751285
rect 0 750641 41657 750809
rect 0 750165 41713 750641
rect 0 749997 41657 750165
rect 0 749613 41713 749997
rect 0 749445 41657 749613
rect 0 748969 41713 749445
rect 42260 749034 42288 756894
rect 41800 749006 42288 749034
rect 0 748801 41657 748969
rect 41800 748913 41828 749006
rect 41713 748857 42193 748913
rect 0 748325 41713 748801
rect 0 748157 41657 748325
rect 0 747681 41713 748157
rect 42536 787030 42564 787358
rect 42524 786966 42576 787030
rect 42628 755478 42656 797710
rect 673472 775878 673500 864214
rect 673564 785738 673592 874482
rect 673644 872374 673696 872438
rect 673552 785674 673604 785738
rect 673460 775814 673512 775878
rect 42800 757590 42852 757654
rect 42708 757522 42760 757586
rect 42616 755414 42668 755478
rect 0 747513 41657 747681
rect 41788 747662 41840 747726
rect 41800 747625 41828 747662
rect 41713 747569 42193 747625
rect 0 747129 41713 747513
rect 0 746961 41657 747129
rect 0 746485 41713 746961
rect 0 746317 41657 746485
rect 0 745841 41713 746317
rect 0 745673 41657 745841
rect 0 745289 41713 745673
rect 0 745121 41657 745289
rect 0 744645 41713 745121
rect 0 744477 41657 744645
rect 41713 744533 42193 744589
rect 0 744001 41713 744477
rect 41800 744054 41828 744533
rect 0 743833 41657 744001
rect 41788 743990 41840 744054
rect 0 743449 41713 743833
rect 0 743281 41657 743449
rect 0 742805 41713 743281
rect 0 742637 41657 742805
rect 0 742161 41713 742637
rect 0 741993 41657 742161
rect 0 741609 41713 741993
rect 0 741441 41657 741609
rect 0 741242 41713 741441
rect 0 713773 41713 713983
rect 0 713605 41657 713773
rect 41713 713703 42193 713717
rect 41713 713675 42288 713703
rect 41713 713661 42193 713675
rect 0 713129 41713 713605
rect 0 712961 41657 713129
rect 0 712485 41713 712961
rect 0 712317 41657 712485
rect 41713 712373 42193 712429
rect 0 711933 41713 712317
rect 41788 712234 41840 712298
rect 0 711765 41657 711933
rect 41800 711877 41828 712234
rect 41713 711821 42193 711877
rect 0 711289 41713 711765
rect 0 711121 41657 711289
rect 0 710645 41713 711121
rect 0 710477 41657 710645
rect 0 710093 41713 710477
rect 0 709925 41657 710093
rect 41713 709981 42193 710037
rect 0 709449 41713 709925
rect 0 709281 41657 709449
rect 0 708805 41713 709281
rect 0 708637 41657 708805
rect 0 708253 41713 708637
rect 0 708085 41657 708253
rect 0 707609 41713 708085
rect 0 707441 41657 707609
rect 0 706965 41713 707441
rect 0 706797 41657 706965
rect 0 706413 41713 706797
rect 0 706245 41657 706413
rect 0 705769 41713 706245
rect 42260 706194 42288 713675
rect 41892 706166 42288 706194
rect 0 705601 41657 705769
rect 41892 705713 41920 706166
rect 41713 705657 42193 705713
rect 0 705125 41713 705601
rect 0 704957 41657 705125
rect 42628 712298 42656 755414
rect 42720 747726 42748 757522
rect 42708 747662 42760 747726
rect 42616 712234 42668 712298
rect 42628 709334 42656 712234
rect 0 704481 41713 704957
rect 42536 709306 42656 709334
rect 0 704313 41657 704481
rect 41722 704425 41828 704426
rect 41713 704369 42193 704425
rect 0 703929 41713 704313
rect 41800 704002 41828 704369
rect 41788 703938 41840 704002
rect 0 703761 41657 703929
rect 0 703285 41713 703761
rect 0 703117 41657 703285
rect 0 702641 41713 703117
rect 0 702473 41657 702641
rect 0 702089 41713 702473
rect 0 701921 41657 702089
rect 0 701445 41713 701921
rect 0 701277 41657 701445
rect 41713 701333 42193 701389
rect 0 700801 41713 701277
rect 41800 700874 41828 701333
rect 41788 700810 41840 700874
rect 0 700633 41657 700801
rect 0 700249 41713 700633
rect 42432 703938 42484 704002
rect 0 700081 41657 700249
rect 0 699605 41713 700081
rect 0 699437 41657 699605
rect 0 698961 41713 699437
rect 0 698793 41657 698961
rect 0 698409 41713 698793
rect 0 698241 41657 698409
rect 0 698042 41713 698241
rect 0 670573 41713 670783
rect 0 670405 41657 670573
rect 41713 670503 42193 670517
rect 41713 670475 42288 670503
rect 41713 670461 42193 670475
rect 0 669929 41713 670405
rect 0 669761 41657 669929
rect 0 669285 41713 669761
rect 0 669117 41657 669285
rect 41713 669173 42193 669229
rect 0 668733 41713 669117
rect 0 668565 41657 668733
rect 41713 668621 42193 668677
rect 0 668089 41713 668565
rect 41800 668166 41828 668621
rect 41788 668102 41840 668166
rect 0 667921 41657 668089
rect 0 667445 41713 667921
rect 0 667277 41657 667445
rect 0 666893 41713 667277
rect 0 666725 41657 666893
rect 41713 666781 42193 666837
rect 0 666249 41713 666725
rect 0 666081 41657 666249
rect 0 665605 41713 666081
rect 0 665437 41657 665605
rect 0 665053 41713 665437
rect 0 664885 41657 665053
rect 0 664409 41713 664885
rect 0 664241 41657 664409
rect 0 663765 41713 664241
rect 0 663597 41657 663765
rect 0 663213 41713 663597
rect 0 663045 41657 663213
rect 0 662569 41713 663045
rect 0 662401 41657 662569
rect 42260 662538 42288 670475
rect 41708 662510 42288 662538
rect 41708 662485 42193 662510
rect 41713 662457 42193 662485
rect 0 661925 41713 662401
rect 0 661757 41657 661925
rect 0 661281 41713 661757
rect 0 661113 41657 661281
rect 41713 661169 42193 661225
rect 0 660729 41713 661113
rect 41800 661094 41828 661169
rect 41788 661030 41840 661094
rect 0 660561 41657 660729
rect 0 660085 41713 660561
rect 0 659917 41657 660085
rect 0 659441 41713 659917
rect 0 659273 41657 659441
rect 0 658889 41713 659273
rect 0 658721 41657 658889
rect 0 658245 41713 658721
rect 41788 658650 41840 658714
rect 0 658077 41657 658245
rect 41800 658189 41828 658650
rect 41713 658133 42193 658189
rect 0 657601 41713 658077
rect 42444 661094 42472 703938
rect 42536 668166 42564 709306
rect 42720 704002 42748 747662
rect 42812 744054 42840 757590
rect 42800 743990 42852 744054
rect 42708 703938 42760 704002
rect 42812 700890 42840 743990
rect 673472 730930 673500 775814
rect 673564 740382 673592 785674
rect 673656 782338 673684 872374
rect 673828 870130 673880 870194
rect 673840 863258 673868 870130
rect 673828 863194 673880 863258
rect 673644 782274 673696 782338
rect 673552 740318 673604 740382
rect 673656 738138 673684 782274
rect 673828 740318 673880 740382
rect 673644 738074 673696 738138
rect 673460 730866 673512 730930
rect 42628 700874 42840 700890
rect 42616 700862 42840 700874
rect 42616 700810 42668 700862
rect 42524 668102 42576 668166
rect 42432 661030 42484 661094
rect 0 657433 41657 657601
rect 0 657049 41713 657433
rect 0 656881 41657 657049
rect 0 656405 41713 656881
rect 0 656237 41657 656405
rect 0 655761 41713 656237
rect 0 655593 41657 655761
rect 0 655209 41713 655593
rect 0 655041 41657 655209
rect 0 654842 41713 655041
rect 0 627373 41713 627583
rect 0 627205 41657 627373
rect 41713 627314 42193 627317
rect 41713 627286 42288 627314
rect 41713 627261 42193 627286
rect 0 626729 41713 627205
rect 0 626561 41657 626729
rect 0 626085 41713 626561
rect 0 625917 41657 626085
rect 41713 625973 42193 626029
rect 0 625533 41713 625917
rect 0 625365 41657 625533
rect 41713 625421 42193 625477
rect 0 624889 41713 625365
rect 41800 624986 41828 625421
rect 41788 624922 41840 624986
rect 0 624721 41657 624889
rect 0 624245 41713 624721
rect 0 624077 41657 624245
rect 0 623693 41713 624077
rect 0 623525 41657 623693
rect 41713 623581 42193 623637
rect 0 623049 41713 623525
rect 0 622881 41657 623049
rect 0 622405 41713 622881
rect 0 622237 41657 622405
rect 0 621853 41713 622237
rect 0 621685 41657 621853
rect 0 621209 41713 621685
rect 0 621041 41657 621209
rect 0 620565 41713 621041
rect 0 620397 41657 620565
rect 0 620013 41713 620397
rect 0 619845 41657 620013
rect 0 619369 41713 619845
rect 42260 619426 42288 627286
rect 41800 619398 42288 619426
rect 0 619201 41657 619369
rect 41800 619313 41828 619398
rect 41713 619257 42193 619313
rect 0 618725 41713 619201
rect 0 618557 41657 618725
rect 0 618081 41713 618557
rect 41788 618462 41840 618526
rect 0 617913 41657 618081
rect 41800 618025 41828 618462
rect 41713 617969 42193 618025
rect 0 617529 41713 617913
rect 0 617361 41657 617529
rect 0 616885 41713 617361
rect 0 616717 41657 616885
rect 0 616241 41713 616717
rect 0 616073 41657 616241
rect 0 615689 41713 616073
rect 0 615521 41657 615689
rect 0 615045 41713 615521
rect 41788 615470 41840 615534
rect 0 614877 41657 615045
rect 41800 614989 41828 615470
rect 41713 614933 42193 614989
rect 0 614401 41713 614877
rect 0 614233 41657 614401
rect 42444 618526 42472 661030
rect 42536 624986 42564 668102
rect 42628 658714 42656 700810
rect 673460 695302 673512 695366
rect 42616 658650 42668 658714
rect 42524 624922 42576 624986
rect 42432 618462 42484 618526
rect 0 613849 41713 614233
rect 0 613681 41657 613849
rect 0 613205 41713 613681
rect 0 613037 41657 613205
rect 0 612561 41713 613037
rect 0 612393 41657 612561
rect 0 612009 41713 612393
rect 0 611841 41657 612009
rect 0 611642 41713 611841
rect 0 584173 41713 584383
rect 0 584005 41657 584173
rect 41713 584103 42193 584117
rect 41713 584075 42288 584103
rect 41713 584061 42193 584075
rect 0 583529 41713 584005
rect 0 583361 41657 583529
rect 0 582885 41713 583361
rect 0 582717 41657 582885
rect 41713 582773 42193 582829
rect 0 582333 41713 582717
rect 0 582165 41657 582333
rect 41713 582221 42193 582277
rect 0 581689 41713 582165
rect 41800 581738 41828 582221
rect 0 581521 41657 581689
rect 41788 581674 41840 581738
rect 0 581045 41713 581521
rect 0 580877 41657 581045
rect 0 580493 41713 580877
rect 0 580325 41657 580493
rect 41713 580381 42193 580437
rect 0 579849 41713 580325
rect 0 579681 41657 579849
rect 0 579205 41713 579681
rect 0 579037 41657 579205
rect 0 578653 41713 579037
rect 0 578485 41657 578653
rect 0 578009 41713 578485
rect 0 577841 41657 578009
rect 0 577365 41713 577841
rect 0 577197 41657 577365
rect 0 576813 41713 577197
rect 0 576645 41657 576813
rect 0 576169 41713 576645
rect 42260 576178 42288 584075
rect 0 576001 41657 576169
rect 41800 576150 42288 576178
rect 41800 576113 41828 576150
rect 41713 576057 42193 576113
rect 0 575525 41713 576001
rect 0 575357 41657 575525
rect 42444 603106 42472 618462
rect 42536 603226 42564 624922
rect 42628 615534 42656 658650
rect 673472 650554 673500 695302
rect 673656 692322 673684 738074
rect 673840 695366 673868 740318
rect 674012 730866 674064 730930
rect 673828 695302 673880 695366
rect 673656 692306 673960 692322
rect 673656 692294 673972 692306
rect 673920 692242 673972 692294
rect 673552 685170 673604 685234
rect 673460 650490 673512 650554
rect 673472 647222 673500 650490
rect 673460 647158 673512 647222
rect 673460 647022 673512 647086
rect 42616 615470 42668 615534
rect 42628 612734 42656 615470
rect 42628 612706 42840 612734
rect 42524 603162 42576 603226
rect 42444 603078 42656 603106
rect 42524 602958 42576 603022
rect 42536 585134 42564 602958
rect 42628 593414 42656 603078
rect 42628 593386 42748 593414
rect 42444 585106 42564 585134
rect 42444 581738 42472 585106
rect 42432 581674 42484 581738
rect 0 574881 41713 575357
rect 41788 575214 41840 575278
rect 0 574713 41657 574881
rect 41800 574825 41828 575214
rect 41713 574769 42193 574825
rect 0 574329 41713 574713
rect 0 574161 41657 574329
rect 0 573685 41713 574161
rect 0 573517 41657 573685
rect 0 573041 41713 573517
rect 0 572873 41657 573041
rect 0 572489 41713 572873
rect 0 572321 41657 572489
rect 0 571845 41713 572321
rect 41788 572222 41840 572286
rect 0 571677 41657 571845
rect 41800 571789 41828 572222
rect 41713 571733 42193 571789
rect 0 571201 41713 571677
rect 0 571033 41657 571201
rect 42248 571134 42300 571198
rect 0 570649 41713 571033
rect 0 570481 41657 570649
rect 0 570005 41713 570481
rect 0 569837 41657 570005
rect 0 569361 41713 569837
rect 0 569193 41657 569361
rect 0 568809 41713 569193
rect 0 568641 41657 568809
rect 0 568442 41713 568641
rect 42260 543114 42288 571134
rect 42248 543050 42300 543114
rect 0 540973 41713 541183
rect 0 540805 41657 540973
rect 41713 540903 42193 540917
rect 41713 540875 42288 540903
rect 41713 540861 42193 540875
rect 0 540329 41713 540805
rect 0 540161 41657 540329
rect 0 539685 41713 540161
rect 0 539517 41657 539685
rect 41713 539573 42193 539629
rect 0 539133 41713 539517
rect 41788 539446 41840 539510
rect 0 538965 41657 539133
rect 41800 539077 41828 539446
rect 41713 539021 42193 539077
rect 0 538489 41713 538965
rect 0 538321 41657 538489
rect 0 537845 41713 538321
rect 0 537677 41657 537845
rect 0 537293 41713 537677
rect 0 537125 41657 537293
rect 41713 537181 42193 537237
rect 0 536649 41713 537125
rect 0 536481 41657 536649
rect 0 536005 41713 536481
rect 0 535837 41657 536005
rect 0 535453 41713 535837
rect 0 535285 41657 535453
rect 0 534809 41713 535285
rect 0 534641 41657 534809
rect 0 534165 41713 534641
rect 0 533997 41657 534165
rect 0 533613 41713 533997
rect 0 533445 41657 533613
rect 0 532969 41713 533445
rect 42260 533066 42288 540875
rect 41800 533038 42288 533066
rect 0 532801 41657 532969
rect 41800 532913 41828 533038
rect 41713 532857 42193 532913
rect 0 532325 41713 532801
rect 0 532157 41657 532325
rect 0 531681 41713 532157
rect 42444 571198 42472 581674
rect 42720 575278 42748 593386
rect 42708 575214 42760 575278
rect 42524 572222 42576 572286
rect 42432 571134 42484 571198
rect 42432 543050 42484 543114
rect 42444 539510 42472 543050
rect 42432 539446 42484 539510
rect 0 531513 41657 531681
rect 41713 531569 42193 531625
rect 0 531129 41713 531513
rect 41800 531214 41828 531569
rect 41788 531150 41840 531214
rect 0 530961 41657 531129
rect 0 530485 41713 530961
rect 0 530317 41657 530485
rect 0 529841 41713 530317
rect 0 529673 41657 529841
rect 0 529289 41713 529673
rect 0 529121 41657 529289
rect 0 528645 41713 529121
rect 0 528477 41657 528645
rect 41713 528533 42193 528589
rect 0 528001 41713 528477
rect 41800 528086 41828 528533
rect 41788 528022 41840 528086
rect 0 527833 41657 528001
rect 42536 531434 42564 572222
rect 42720 554774 42748 575214
rect 42812 572286 42840 612706
rect 673472 602954 673500 647022
rect 673564 640694 673592 685170
rect 673644 647158 673696 647222
rect 673552 640630 673604 640694
rect 673460 602890 673512 602954
rect 42800 572222 42852 572286
rect 673472 557870 673500 602890
rect 673564 595066 673592 640630
rect 673656 605130 673684 647158
rect 673932 647086 673960 692242
rect 674024 685234 674052 730866
rect 674012 685170 674064 685234
rect 673920 647022 673972 647086
rect 673644 605066 673696 605130
rect 673552 595002 673604 595066
rect 673460 557806 673512 557870
rect 42352 531406 42564 531434
rect 42628 554746 42748 554774
rect 42352 528086 42380 531406
rect 42628 531298 42656 554746
rect 673564 550526 673592 595002
rect 673656 560998 673684 605066
rect 673644 560934 673696 560998
rect 673552 550462 673604 550526
rect 673564 546494 673592 550462
rect 673472 546466 673592 546494
rect 42800 539446 42852 539510
rect 42444 531270 42656 531298
rect 42444 531214 42472 531270
rect 42432 531150 42484 531214
rect 42340 528022 42392 528086
rect 0 527449 41713 527833
rect 0 527281 41657 527449
rect 0 526805 41713 527281
rect 0 526637 41657 526805
rect 0 526161 41713 526637
rect 0 525993 41657 526161
rect 0 525609 41713 525993
rect 0 525441 41657 525609
rect 0 525242 41713 525441
rect 985 493078 40000 497858
rect 985 487879 39593 493078
rect 39616 488179 40000 488579
rect 985 483099 40000 487879
rect 985 483053 39593 483099
rect 7 456040 30281 457987
rect 30753 455800 31683 458028
rect 32033 456040 34915 457987
rect 7 455740 39593 455800
rect 7 451619 39600 455740
rect 7 451507 39593 451619
rect 7 444985 39600 451507
rect 7 444899 39593 444985
rect 7 440900 39600 444899
rect 7 440800 39593 440900
rect 30760 438605 31690 440800
rect 0 413373 41713 413583
rect 0 413205 41657 413373
rect 41713 413303 42193 413317
rect 41713 413275 42288 413303
rect 41713 413261 42193 413275
rect 0 412729 41713 413205
rect 0 412561 41657 412729
rect 0 412085 41713 412561
rect 0 411917 41657 412085
rect 41713 411973 42193 412029
rect 0 411533 41713 411917
rect 0 411365 41657 411533
rect 41722 411477 41828 411482
rect 41713 411421 42193 411477
rect 0 410889 41713 411365
rect 41800 410990 41828 411421
rect 41788 410926 41840 410990
rect 0 410721 41657 410889
rect 0 410245 41713 410721
rect 0 410077 41657 410245
rect 0 409693 41713 410077
rect 0 409525 41657 409693
rect 41713 409581 42193 409637
rect 0 409049 41713 409525
rect 0 408881 41657 409049
rect 0 408405 41713 408881
rect 0 408237 41657 408405
rect 0 407853 41713 408237
rect 0 407685 41657 407853
rect 0 407209 41713 407685
rect 0 407041 41657 407209
rect 0 406565 41713 407041
rect 0 406397 41657 406565
rect 0 406013 41713 406397
rect 0 405845 41657 406013
rect 0 405369 41713 405845
rect 42260 405498 42288 413275
rect 41800 405470 42288 405498
rect 0 405201 41657 405369
rect 41800 405313 41828 405470
rect 41713 405257 42193 405313
rect 0 404725 41713 405201
rect 0 404557 41657 404725
rect 0 404081 41713 404557
rect 41788 404466 41840 404530
rect 0 403913 41657 404081
rect 41800 404025 41828 404466
rect 41713 403969 42193 404025
rect 0 403529 41713 403913
rect 0 403361 41657 403529
rect 0 402885 41713 403361
rect 0 402717 41657 402885
rect 0 402241 41713 402717
rect 0 402073 41657 402241
rect 0 401689 41713 402073
rect 0 401521 41657 401689
rect 0 401045 41713 401521
rect 0 400877 41657 401045
rect 41713 400933 42193 400989
rect 0 400401 41713 400877
rect 41800 400858 41828 400933
rect 41788 400794 41840 400858
rect 0 400233 41657 400401
rect 42444 404530 42472 531150
rect 42708 528022 42760 528086
rect 42524 410926 42576 410990
rect 42432 404466 42484 404530
rect 0 399849 41713 400233
rect 0 399681 41657 399849
rect 0 399205 41713 399681
rect 0 399037 41657 399205
rect 0 398561 41713 399037
rect 0 398393 41657 398561
rect 0 398009 41713 398393
rect 0 397841 41657 398009
rect 0 397642 41713 397841
rect 0 370173 41713 370383
rect 0 370005 41657 370173
rect 41713 370061 42193 370117
rect 0 369529 41713 370005
rect 41800 369578 41828 370061
rect 0 369361 41657 369529
rect 41788 369514 41840 369578
rect 0 368885 41713 369361
rect 0 368717 41657 368885
rect 41713 368773 42193 368829
rect 0 368333 41713 368717
rect 41788 368630 41840 368694
rect 0 368165 41657 368333
rect 41800 368277 41828 368630
rect 41713 368221 42193 368277
rect 0 367689 41713 368165
rect 0 367521 41657 367689
rect 0 367045 41713 367521
rect 0 366877 41657 367045
rect 0 366493 41713 366877
rect 0 366325 41657 366493
rect 41713 366381 42193 366437
rect 0 365849 41713 366325
rect 0 365681 41657 365849
rect 0 365205 41713 365681
rect 0 365037 41657 365205
rect 0 364653 41713 365037
rect 0 364485 41657 364653
rect 0 364009 41713 364485
rect 0 363841 41657 364009
rect 0 363365 41713 363841
rect 0 363197 41657 363365
rect 0 362813 41713 363197
rect 0 362645 41657 362813
rect 0 362169 41713 362645
rect 41788 362578 41840 362642
rect 0 362001 41657 362169
rect 41800 362114 41828 362578
rect 41722 362113 41828 362114
rect 41713 362057 42193 362113
rect 0 361525 41713 362001
rect 0 361357 41657 361525
rect 42340 369514 42392 369578
rect 42352 362642 42380 369514
rect 42536 368694 42564 410926
rect 42616 404466 42668 404530
rect 42524 368630 42576 368694
rect 42340 362578 42392 362642
rect 42536 361574 42564 368630
rect 0 360881 41713 361357
rect 0 360713 41657 360881
rect 41713 360769 42193 360825
rect 41800 360738 41828 360769
rect 0 360329 41713 360713
rect 41788 360674 41840 360738
rect 0 360161 41657 360329
rect 0 359685 41713 360161
rect 0 359517 41657 359685
rect 0 359041 41713 359517
rect 0 358873 41657 359041
rect 0 358489 41713 358873
rect 0 358321 41657 358489
rect 0 357845 41713 358321
rect 0 357677 41657 357845
rect 41713 357733 42193 357789
rect 0 357201 41713 357677
rect 41800 357270 41828 357733
rect 41788 357206 41840 357270
rect 0 357033 41657 357201
rect 0 356649 41713 357033
rect 0 356481 41657 356649
rect 0 356005 41713 356481
rect 0 355837 41657 356005
rect 0 355361 41713 355837
rect 0 355193 41657 355361
rect 0 354809 41713 355193
rect 0 354641 41657 354809
rect 0 354442 41713 354641
rect 42352 361546 42564 361574
rect 42352 342254 42380 361546
rect 42628 360738 42656 404466
rect 42720 400858 42748 528022
rect 42812 410990 42840 539446
rect 42800 410926 42852 410990
rect 42708 400794 42760 400858
rect 42616 360674 42668 360738
rect 42524 357206 42576 357270
rect 42352 342226 42472 342254
rect 0 326973 41713 327183
rect 0 326805 41657 326973
rect 41713 326861 42193 326917
rect 0 326329 41713 326805
rect 41892 326754 41920 326861
rect 41892 326726 42288 326754
rect 0 326161 41657 326329
rect 0 325685 41713 326161
rect 0 325517 41657 325685
rect 41713 325573 42193 325629
rect 0 325133 41713 325517
rect 41788 325450 41840 325514
rect 0 324965 41657 325133
rect 41800 325077 41828 325450
rect 41713 325021 42193 325077
rect 0 324489 41713 324965
rect 0 324321 41657 324489
rect 0 323845 41713 324321
rect 0 323677 41657 323845
rect 0 323293 41713 323677
rect 0 323125 41657 323293
rect 41713 323181 42193 323237
rect 0 322649 41713 323125
rect 0 322481 41657 322649
rect 0 322005 41713 322481
rect 0 321837 41657 322005
rect 0 321453 41713 321837
rect 0 321285 41657 321453
rect 0 320809 41713 321285
rect 0 320641 41657 320809
rect 0 320165 41713 320641
rect 0 319997 41657 320165
rect 0 319613 41713 319997
rect 0 319445 41657 319613
rect 0 318969 41713 319445
rect 0 318801 41657 318969
rect 41713 318899 42193 318913
rect 42260 318899 42288 326726
rect 41713 318871 42288 318899
rect 41713 318857 42193 318871
rect 0 318325 41713 318801
rect 0 318157 41657 318325
rect 42444 325514 42472 342226
rect 42432 325450 42484 325514
rect 0 317681 41713 318157
rect 0 317513 41657 317681
rect 41713 317569 42193 317625
rect 0 317129 41713 317513
rect 41800 317218 41828 317569
rect 41788 317154 41840 317218
rect 0 316961 41657 317129
rect 0 316485 41713 316961
rect 0 316317 41657 316485
rect 0 315841 41713 316317
rect 0 315673 41657 315841
rect 0 315289 41713 315673
rect 0 315121 41657 315289
rect 0 314645 41713 315121
rect 0 314477 41657 314645
rect 41713 314533 42193 314589
rect 0 314001 41713 314477
rect 41800 314090 41828 314533
rect 41788 314026 41840 314090
rect 0 313833 41657 314001
rect 42536 314090 42564 357206
rect 42628 317218 42656 360674
rect 42720 357270 42748 400794
rect 673472 372366 673500 546466
rect 674760 427854 674788 996338
rect 678067 962665 716615 967547
rect 677600 962021 677984 962421
rect 678007 957578 716615 962665
rect 682788 952742 716615 957578
rect 685910 922600 686840 924795
rect 678007 922500 717593 922600
rect 678000 918501 717593 922500
rect 678007 918415 717593 918501
rect 678000 911893 717593 918415
rect 678007 911781 717593 911893
rect 678000 907660 717593 911781
rect 678007 907600 717593 907660
rect 682685 905413 685567 907360
rect 685917 905372 686847 907600
rect 687319 905413 717593 907360
rect 675887 878159 717600 878358
rect 675943 877991 717600 878159
rect 675887 877607 717600 877991
rect 675943 877439 717600 877607
rect 675887 876963 717600 877439
rect 675943 876795 717600 876963
rect 675887 876319 717600 876795
rect 675943 876151 717600 876319
rect 675887 875767 717600 876151
rect 675943 875599 717600 875767
rect 675887 875123 717600 875599
rect 675407 875039 675887 875067
rect 675404 875011 675887 875039
rect 675404 874546 675432 875011
rect 675943 874955 717600 875123
rect 675392 874482 675444 874546
rect 675887 874479 717600 874955
rect 675943 874311 717600 874479
rect 675887 873927 717600 874311
rect 675943 873759 717600 873927
rect 675887 873283 717600 873759
rect 675943 873115 717600 873283
rect 675887 872639 717600 873115
rect 675943 872471 717600 872639
rect 675392 872374 675444 872438
rect 675404 872031 675432 872374
rect 675887 872087 717600 872471
rect 675404 872003 675887 872031
rect 675407 871975 675887 872003
rect 675943 871919 717600 872087
rect 675887 871443 717600 871919
rect 675943 871275 717600 871443
rect 675887 870799 717600 871275
rect 675407 870740 675887 870743
rect 675404 870687 675887 870740
rect 675404 870194 675432 870687
rect 675943 870631 717600 870799
rect 675392 870130 675444 870194
rect 675887 870155 717600 870631
rect 675943 869987 717600 870155
rect 675887 869603 717600 869987
rect 675943 869435 717600 869603
rect 675887 868959 717600 869435
rect 675943 868791 717600 868959
rect 675887 868315 717600 868791
rect 675943 868147 717600 868315
rect 675887 867763 717600 868147
rect 675943 867595 717600 867763
rect 675887 867119 717600 867595
rect 675943 866951 717600 867119
rect 675887 866475 717600 866951
rect 675407 866363 675887 866419
rect 675943 866307 717600 866475
rect 675887 865923 717600 866307
rect 675943 865755 717600 865923
rect 675887 865279 717600 865755
rect 675943 865111 717600 865279
rect 675887 864635 717600 865111
rect 675407 864551 675887 864579
rect 675404 864523 675887 864551
rect 675404 864278 675432 864523
rect 675943 864467 717600 864635
rect 675392 864214 675444 864278
rect 675887 864083 717600 864467
rect 675407 863971 675887 864027
rect 675943 863915 717600 864083
rect 675887 863439 717600 863915
rect 675943 863271 717600 863439
rect 675392 863194 675444 863258
rect 675404 862739 675432 863194
rect 675887 862795 717600 863271
rect 675404 862716 675887 862739
rect 675407 862683 675887 862716
rect 675943 862627 717600 862795
rect 675887 862417 717600 862627
rect 678007 833301 716615 833347
rect 677600 828521 716615 833301
rect 677600 827821 677984 828221
rect 678007 823322 716615 828521
rect 677600 818542 716615 823322
rect 675300 818314 675352 818378
rect 677598 818343 677654 818417
rect 677600 818314 677652 818343
rect 675312 786614 675340 818314
rect 675887 788959 717600 789158
rect 675943 788791 717600 788959
rect 675887 788407 717600 788791
rect 675943 788239 717600 788407
rect 675887 787763 717600 788239
rect 675943 787595 717600 787763
rect 675887 787119 717600 787595
rect 675943 786951 717600 787119
rect 675128 786586 675340 786614
rect 675128 728906 675156 786586
rect 675887 786567 717600 786951
rect 675943 786399 717600 786567
rect 675887 785923 717600 786399
rect 675407 785839 675887 785867
rect 675404 785811 675887 785839
rect 675404 785738 675432 785811
rect 675943 785755 717600 785923
rect 675392 785674 675444 785738
rect 675887 785279 717600 785755
rect 675943 785111 717600 785279
rect 675887 784727 717600 785111
rect 675943 784559 717600 784727
rect 675887 784083 717600 784559
rect 675943 783915 717600 784083
rect 675887 783439 717600 783915
rect 675943 783271 717600 783439
rect 675887 782887 717600 783271
rect 675407 782803 675887 782831
rect 675404 782775 675887 782803
rect 675404 782338 675432 782775
rect 675943 782719 717600 782887
rect 675392 782274 675444 782338
rect 675887 782243 717600 782719
rect 675943 782075 717600 782243
rect 675887 781599 717600 782075
rect 675407 781524 675887 781543
rect 675404 781487 675887 781524
rect 675404 781046 675432 781487
rect 675943 781431 717600 781599
rect 675208 780982 675260 781046
rect 675392 780982 675444 781046
rect 675220 773514 675248 780982
rect 675887 780955 717600 781431
rect 675943 780787 717600 780955
rect 675887 780403 717600 780787
rect 675943 780235 717600 780403
rect 675887 779759 717600 780235
rect 675943 779591 717600 779759
rect 675887 779115 717600 779591
rect 675943 778947 717600 779115
rect 675887 778563 717600 778947
rect 675943 778395 717600 778563
rect 675887 777919 717600 778395
rect 675943 777751 717600 777919
rect 675887 777275 717600 777751
rect 675407 777163 675887 777219
rect 675943 777107 717600 777275
rect 675887 776723 717600 777107
rect 675943 776555 717600 776723
rect 675887 776079 717600 776555
rect 675943 775911 717600 776079
rect 675392 775814 675444 775878
rect 675404 775379 675432 775814
rect 675887 775435 717600 775911
rect 675404 775351 675887 775379
rect 675407 775323 675887 775351
rect 675943 775267 717600 775435
rect 675887 774883 717600 775267
rect 675407 774771 675887 774827
rect 675943 774715 717600 774883
rect 675887 774239 717600 774715
rect 675943 774071 717600 774239
rect 675887 773595 717600 774071
rect 675407 773514 675887 773539
rect 675220 773486 675887 773514
rect 675407 773483 675887 773486
rect 675943 773427 717600 773595
rect 675887 773217 717600 773427
rect 675887 743959 717600 744158
rect 675943 743791 717600 743959
rect 675887 743407 717600 743791
rect 675943 743239 717600 743407
rect 675887 742763 717600 743239
rect 675943 742595 717600 742763
rect 675887 742119 717600 742595
rect 675943 741951 717600 742119
rect 675887 741567 717600 741951
rect 675943 741399 717600 741567
rect 675887 740923 717600 741399
rect 675407 740860 675887 740867
rect 675404 740811 675887 740860
rect 675404 740382 675432 740811
rect 675943 740755 717600 740923
rect 675392 740318 675444 740382
rect 675887 740279 717600 740755
rect 675943 740111 717600 740279
rect 675887 739727 717600 740111
rect 675943 739559 717600 739727
rect 675887 739083 717600 739559
rect 675943 738915 717600 739083
rect 675887 738439 717600 738915
rect 675943 738271 717600 738439
rect 675392 738074 675444 738138
rect 675404 737831 675432 738074
rect 675887 737887 717600 738271
rect 675404 737803 675887 737831
rect 675407 737775 675887 737803
rect 675943 737719 717600 737887
rect 675887 737243 717600 737719
rect 675943 737075 717600 737243
rect 675887 736599 717600 737075
rect 675407 736522 675887 736543
rect 675312 736494 675887 736522
rect 675312 729042 675340 736494
rect 675407 736487 675887 736494
rect 675943 736431 717600 736599
rect 675887 735955 717600 736431
rect 675943 735787 717600 735955
rect 675887 735403 717600 735787
rect 675943 735235 717600 735403
rect 675887 734759 717600 735235
rect 675943 734591 717600 734759
rect 675887 734115 717600 734591
rect 675943 733947 717600 734115
rect 675887 733563 717600 733947
rect 675943 733395 717600 733563
rect 675887 732919 717600 733395
rect 675943 732751 717600 732919
rect 675887 732275 717600 732751
rect 675407 732163 675887 732219
rect 675943 732107 717600 732275
rect 675887 731723 717600 732107
rect 675943 731555 717600 731723
rect 675887 731079 717600 731555
rect 675392 730866 675444 730930
rect 675943 730911 717600 731079
rect 675404 730379 675432 730866
rect 675887 730435 717600 730911
rect 675404 730351 675887 730379
rect 675407 730323 675887 730351
rect 675943 730267 717600 730435
rect 675887 729883 717600 730267
rect 675407 729771 675887 729827
rect 675943 729715 717600 729883
rect 675887 729239 717600 729715
rect 675943 729071 717600 729239
rect 675312 729014 675432 729042
rect 675128 728878 675340 728906
rect 675312 701054 675340 728878
rect 675404 728539 675432 729014
rect 675887 728595 717600 729071
rect 675404 728484 675887 728539
rect 675407 728483 675887 728484
rect 675943 728427 717600 728595
rect 675887 728217 717600 728427
rect 675128 701026 675340 701054
rect 675128 681734 675156 701026
rect 675887 698959 717600 699158
rect 675943 698791 717600 698959
rect 675887 698407 717600 698791
rect 675943 698239 717600 698407
rect 675887 697763 717600 698239
rect 675943 697595 717600 697763
rect 675887 697119 717600 697595
rect 675943 696951 717600 697119
rect 675887 696567 717600 696951
rect 675943 696399 717600 696567
rect 675887 695923 717600 696399
rect 675407 695844 675887 695867
rect 675404 695811 675887 695844
rect 675404 695366 675432 695811
rect 675943 695755 717600 695923
rect 675392 695302 675444 695366
rect 675887 695279 717600 695755
rect 675943 695111 717600 695279
rect 675887 694727 717600 695111
rect 675943 694559 717600 694727
rect 675887 694083 717600 694559
rect 675943 693915 717600 694083
rect 675887 693439 717600 693915
rect 675943 693271 717600 693439
rect 675887 692887 717600 693271
rect 675407 692803 675887 692831
rect 675404 692775 675887 692803
rect 675404 692306 675432 692775
rect 675943 692719 717600 692887
rect 675392 692242 675444 692306
rect 675887 692243 717600 692719
rect 675943 692075 717600 692243
rect 675312 691614 675432 691642
rect 675312 683525 675340 691614
rect 675404 691543 675432 691614
rect 675887 691599 717600 692075
rect 675404 691492 675887 691543
rect 675407 691487 675887 691492
rect 675943 691431 717600 691599
rect 675887 690955 717600 691431
rect 675943 690787 717600 690955
rect 675887 690403 717600 690787
rect 675943 690235 717600 690403
rect 675887 689759 717600 690235
rect 675943 689591 717600 689759
rect 675887 689115 717600 689591
rect 675943 688947 717600 689115
rect 675887 688563 717600 688947
rect 675943 688395 717600 688563
rect 675887 687919 717600 688395
rect 675943 687751 717600 687919
rect 675887 687275 717600 687751
rect 675407 687163 675887 687219
rect 675943 687107 717600 687275
rect 675887 686723 717600 687107
rect 675943 686555 717600 686723
rect 675887 686079 717600 686555
rect 675943 685911 717600 686079
rect 675887 685435 717600 685911
rect 675407 685372 675887 685379
rect 675404 685323 675887 685372
rect 675404 685234 675432 685323
rect 675943 685267 717600 685435
rect 675392 685170 675444 685234
rect 675887 684883 717600 685267
rect 675407 684771 675887 684827
rect 675943 684715 717600 684883
rect 675887 684239 717600 684715
rect 675943 684071 717600 684239
rect 675887 683595 717600 684071
rect 675407 683525 675887 683539
rect 675312 683497 675887 683525
rect 675407 683483 675887 683497
rect 675943 683427 717600 683595
rect 675887 683217 717600 683427
rect 675128 681706 675340 681734
rect 675312 651374 675340 681706
rect 675887 653759 717600 653958
rect 675943 653591 717600 653759
rect 675887 653207 717600 653591
rect 675943 653039 717600 653207
rect 675887 652563 717600 653039
rect 675943 652395 717600 652563
rect 675887 651919 717600 652395
rect 675943 651751 717600 651919
rect 675128 651346 675340 651374
rect 675887 651367 717600 651751
rect 675128 632054 675156 651346
rect 675943 651199 717600 651367
rect 675887 650723 717600 651199
rect 675407 650639 675887 650667
rect 675404 650611 675887 650639
rect 675404 650554 675432 650611
rect 675943 650555 717600 650723
rect 675392 650490 675444 650554
rect 675887 650079 717600 650555
rect 675943 649911 717600 650079
rect 675887 649527 717600 649911
rect 675943 649359 717600 649527
rect 675887 648883 717600 649359
rect 675943 648715 717600 648883
rect 675887 648239 717600 648715
rect 675943 648071 717600 648239
rect 675887 647687 717600 648071
rect 675407 647603 675887 647631
rect 675404 647575 675887 647603
rect 675404 647086 675432 647575
rect 675943 647519 717600 647687
rect 675392 647022 675444 647086
rect 675887 647043 717600 647519
rect 675943 646875 717600 647043
rect 675887 646399 717600 646875
rect 675407 646340 675887 646343
rect 675404 646287 675887 646340
rect 675404 645794 675432 646287
rect 675943 646231 717600 646399
rect 675208 645730 675260 645794
rect 675392 645730 675444 645794
rect 675887 645755 717600 646231
rect 675220 638330 675248 645730
rect 675943 645587 717600 645755
rect 675887 645203 717600 645587
rect 675943 645035 717600 645203
rect 675887 644559 717600 645035
rect 675943 644391 717600 644559
rect 675887 643915 717600 644391
rect 675943 643747 717600 643915
rect 675887 643363 717600 643747
rect 675943 643195 717600 643363
rect 675887 642719 717600 643195
rect 675943 642551 717600 642719
rect 675887 642075 717600 642551
rect 675407 641963 675887 642019
rect 675943 641907 717600 642075
rect 675887 641523 717600 641907
rect 675943 641355 717600 641523
rect 675887 640879 717600 641355
rect 675943 640711 717600 640879
rect 675392 640630 675444 640694
rect 675404 640179 675432 640630
rect 675887 640235 717600 640711
rect 675404 640151 675887 640179
rect 675407 640123 675887 640151
rect 675943 640067 717600 640235
rect 675887 639683 717600 640067
rect 675407 639571 675887 639627
rect 675943 639515 717600 639683
rect 675887 639039 717600 639515
rect 675943 638871 717600 639039
rect 675887 638395 717600 638871
rect 675407 638330 675887 638339
rect 675220 638302 675887 638330
rect 675407 638283 675887 638302
rect 675943 638227 717600 638395
rect 675887 638017 717600 638227
rect 675128 632026 675340 632054
rect 675312 612734 675340 632026
rect 675128 612706 675340 612734
rect 675128 593722 675156 612706
rect 675887 608759 717600 608958
rect 675943 608591 717600 608759
rect 675887 608207 717600 608591
rect 675943 608039 717600 608207
rect 675887 607563 717600 608039
rect 675943 607395 717600 607563
rect 675887 606919 717600 607395
rect 675943 606751 717600 606919
rect 675887 606367 717600 606751
rect 675943 606199 717600 606367
rect 675887 605723 717600 606199
rect 675407 605639 675887 605667
rect 675404 605611 675887 605639
rect 675404 605130 675432 605611
rect 675943 605555 717600 605723
rect 675392 605066 675444 605130
rect 675887 605079 717600 605555
rect 675943 604911 717600 605079
rect 675887 604527 717600 604911
rect 675943 604359 717600 604527
rect 675887 603883 717600 604359
rect 675943 603715 717600 603883
rect 675887 603239 717600 603715
rect 675943 603071 717600 603239
rect 675392 602890 675444 602954
rect 675404 602631 675432 602890
rect 675887 602687 717600 603071
rect 675404 602603 675887 602631
rect 675407 602575 675887 602603
rect 675943 602519 717600 602687
rect 675887 602043 717600 602519
rect 675943 601875 717600 602043
rect 675887 601399 717600 601875
rect 675407 601338 675887 601343
rect 675312 601310 675887 601338
rect 675312 593858 675340 601310
rect 675407 601287 675887 601310
rect 675943 601231 717600 601399
rect 675887 600755 717600 601231
rect 675943 600587 717600 600755
rect 675887 600203 717600 600587
rect 675943 600035 717600 600203
rect 675887 599559 717600 600035
rect 675943 599391 717600 599559
rect 675887 598915 717600 599391
rect 675943 598747 717600 598915
rect 675887 598363 717600 598747
rect 675943 598195 717600 598363
rect 675887 597719 717600 598195
rect 675943 597551 717600 597719
rect 675887 597075 717600 597551
rect 675407 596963 675887 597019
rect 675943 596907 717600 597075
rect 675887 596523 717600 596907
rect 675943 596355 717600 596523
rect 675887 595879 717600 596355
rect 675943 595711 717600 595879
rect 675887 595235 717600 595711
rect 675407 595151 675887 595179
rect 675404 595123 675887 595151
rect 675404 595066 675432 595123
rect 675943 595067 717600 595235
rect 675392 595002 675444 595066
rect 675887 594683 717600 595067
rect 675407 594571 675887 594627
rect 675943 594515 717600 594683
rect 675887 594039 717600 594515
rect 675943 593871 717600 594039
rect 675312 593830 675432 593858
rect 675128 593694 675340 593722
rect 675312 574094 675340 593694
rect 675404 593339 675432 593830
rect 675887 593395 717600 593871
rect 675404 593300 675887 593339
rect 675407 593283 675887 593300
rect 675943 593227 717600 593395
rect 675887 593017 717600 593227
rect 675128 574066 675340 574094
rect 675128 546494 675156 574066
rect 675887 563559 717600 563758
rect 675943 563391 717600 563559
rect 675887 563007 717600 563391
rect 675943 562839 717600 563007
rect 675887 562363 717600 562839
rect 675943 562195 717600 562363
rect 675887 561719 717600 562195
rect 675943 561551 717600 561719
rect 675887 561167 717600 561551
rect 675943 560999 717600 561167
rect 675392 560934 675444 560998
rect 675404 560467 675432 560934
rect 675887 560523 717600 560999
rect 675404 560439 675887 560467
rect 675407 560411 675887 560439
rect 675943 560355 717600 560523
rect 675887 559879 717600 560355
rect 675943 559711 717600 559879
rect 675887 559327 717600 559711
rect 675943 559159 717600 559327
rect 675887 558683 717600 559159
rect 675943 558515 717600 558683
rect 675887 558039 717600 558515
rect 675943 557871 717600 558039
rect 675392 557806 675444 557870
rect 675404 557431 675432 557806
rect 675887 557487 717600 557871
rect 675404 557396 675887 557431
rect 675407 557375 675887 557396
rect 675943 557319 717600 557487
rect 675887 556843 717600 557319
rect 675943 556675 717600 556843
rect 675887 556199 717600 556675
rect 675407 556115 675887 556143
rect 675404 556087 675887 556115
rect 675404 555626 675432 556087
rect 675943 556031 717600 556199
rect 675208 555562 675260 555626
rect 675392 555562 675444 555626
rect 675220 548125 675248 555562
rect 675887 555555 717600 556031
rect 675943 555387 717600 555555
rect 675887 555003 717600 555387
rect 675943 554835 717600 555003
rect 675887 554359 717600 554835
rect 675943 554191 717600 554359
rect 675887 553715 717600 554191
rect 675943 553547 717600 553715
rect 675887 553163 717600 553547
rect 675943 552995 717600 553163
rect 675887 552519 717600 552995
rect 675943 552351 717600 552519
rect 675887 551875 717600 552351
rect 675407 551763 675887 551819
rect 675943 551707 717600 551875
rect 675887 551323 717600 551707
rect 675943 551155 717600 551323
rect 675887 550679 717600 551155
rect 675392 550462 675444 550526
rect 675943 550511 717600 550679
rect 675404 549979 675432 550462
rect 675887 550035 717600 550511
rect 675404 549951 675887 549979
rect 675407 549923 675887 549951
rect 675943 549867 717600 550035
rect 675887 549483 717600 549867
rect 675407 549371 675887 549427
rect 675943 549315 717600 549483
rect 675887 548839 717600 549315
rect 675943 548671 717600 548839
rect 675887 548195 717600 548671
rect 675407 548125 675887 548139
rect 675220 548097 675887 548125
rect 675407 548083 675887 548097
rect 675943 548027 717600 548195
rect 675887 547817 717600 548027
rect 675128 546466 675340 546494
rect 675312 513806 675340 546466
rect 678007 518701 716615 518747
rect 677600 513921 716615 518701
rect 675300 513742 675352 513806
rect 677692 513777 677744 513806
rect 677690 513703 677746 513777
rect 677600 513221 677984 513621
rect 678007 508722 716615 513921
rect 677600 503942 716615 508722
rect 685910 474800 686840 476995
rect 678007 474700 717593 474800
rect 678000 470701 717593 474700
rect 678007 470615 717593 470701
rect 678000 464093 717593 470615
rect 678007 463981 717593 464093
rect 678000 459860 717593 463981
rect 678007 459800 717593 459860
rect 682685 457613 685567 459560
rect 685917 457572 686847 459800
rect 687319 457613 717593 459560
rect 678007 430501 716615 430547
rect 674748 427790 674800 427854
rect 677508 427790 677560 427854
rect 677520 425649 677548 427790
rect 677600 425721 716615 430501
rect 677506 425575 677562 425649
rect 677600 425021 677984 425421
rect 678007 420522 716615 425721
rect 677600 415742 716615 420522
rect 675887 386359 717600 386558
rect 675943 386191 717600 386359
rect 675887 385807 717600 386191
rect 675943 385639 717600 385807
rect 675887 385163 717600 385639
rect 675943 384995 717600 385163
rect 675887 384519 717600 384995
rect 675943 384351 717600 384519
rect 673552 382706 673604 382770
rect 673460 372302 673512 372366
rect 42708 357206 42760 357270
rect 673564 337550 673592 382706
rect 673736 379646 673788 379710
rect 673552 337486 673604 337550
rect 42800 325450 42852 325514
rect 42616 317154 42668 317218
rect 42524 314026 42576 314090
rect 0 313449 41713 313833
rect 0 313281 41657 313449
rect 0 312805 41713 313281
rect 0 312637 41657 312805
rect 0 312161 41713 312637
rect 0 311993 41657 312161
rect 0 311609 41713 311993
rect 0 311441 41657 311609
rect 0 311242 41713 311441
rect 0 283773 41713 283983
rect 0 283605 41657 283773
rect 41713 283703 42193 283717
rect 41713 283675 42288 283703
rect 41713 283661 42193 283675
rect 0 283129 41713 283605
rect 0 282961 41657 283129
rect 0 282485 41713 282961
rect 0 282317 41657 282485
rect 41713 282373 42193 282429
rect 0 281933 41713 282317
rect 0 281765 41657 281933
rect 41713 281821 42193 281877
rect 0 281289 41713 281765
rect 41800 281382 41828 281821
rect 41788 281318 41840 281382
rect 0 281121 41657 281289
rect 0 280645 41713 281121
rect 0 280477 41657 280645
rect 0 280093 41713 280477
rect 0 279925 41657 280093
rect 41713 279981 42193 280037
rect 0 279449 41713 279925
rect 0 279281 41657 279449
rect 0 278805 41713 279281
rect 0 278637 41657 278805
rect 0 278253 41713 278637
rect 0 278085 41657 278253
rect 0 277609 41713 278085
rect 0 277441 41657 277609
rect 0 276965 41713 277441
rect 0 276797 41657 276965
rect 0 276413 41713 276797
rect 0 276245 41657 276413
rect 0 275769 41713 276245
rect 0 275601 41657 275769
rect 41713 275699 42193 275713
rect 42260 275699 42288 283675
rect 41713 275671 42288 275699
rect 41713 275657 42193 275671
rect 0 275125 41713 275601
rect 42432 281318 42484 281382
rect 0 274957 41657 275125
rect 0 274481 41713 274957
rect 41788 274518 41840 274582
rect 0 274313 41657 274481
rect 41800 274425 41828 274518
rect 41713 274369 42193 274425
rect 41722 274366 41828 274369
rect 0 273929 41713 274313
rect 0 273761 41657 273929
rect 0 273285 41713 273761
rect 0 273117 41657 273285
rect 0 272641 41713 273117
rect 0 272473 41657 272641
rect 0 272089 41713 272473
rect 0 271921 41657 272089
rect 0 271445 41713 271921
rect 41788 271866 41840 271930
rect 0 271277 41657 271445
rect 41800 271402 41828 271866
rect 41722 271389 41828 271402
rect 41713 271333 42193 271389
rect 0 270801 41713 271277
rect 0 270633 41657 270801
rect 0 270249 41713 270633
rect 0 270081 41657 270249
rect 0 269605 41713 270081
rect 0 269437 41657 269605
rect 0 268961 41713 269437
rect 0 268793 41657 268961
rect 0 268409 41713 268793
rect 0 268241 41657 268409
rect 0 268042 41713 268241
rect 0 240573 41713 240783
rect 0 240405 41657 240573
rect 41722 240517 42288 240530
rect 41713 240502 42288 240517
rect 41713 240461 42193 240502
rect 0 239929 41713 240405
rect 0 239761 41657 239929
rect 0 239285 41713 239761
rect 0 239117 41657 239285
rect 41713 239173 42193 239229
rect 0 238733 41713 239117
rect 0 238565 41657 238733
rect 41713 238621 42193 238677
rect 0 238089 41713 238565
rect 41800 238134 41828 238621
rect 0 237921 41657 238089
rect 41788 238070 41840 238134
rect 0 237445 41713 237921
rect 0 237277 41657 237445
rect 41713 237333 42193 237389
rect 0 236893 41713 237277
rect 0 236725 41657 236893
rect 41713 236781 42193 236837
rect 0 236249 41713 236725
rect 0 236081 41657 236249
rect 0 235605 41713 236081
rect 0 235437 41657 235605
rect 41713 235493 42193 235549
rect 0 235053 41713 235437
rect 0 234885 41657 235053
rect 0 234409 41713 234885
rect 0 234241 41657 234409
rect 0 233765 41713 234241
rect 0 233597 41657 233765
rect 0 233213 41713 233597
rect 0 233045 41657 233213
rect 0 232569 41713 233045
rect 42260 232642 42288 240502
rect 41800 232614 42288 232642
rect 0 232401 41657 232569
rect 41800 232513 41828 232614
rect 41713 232457 42193 232513
rect 0 231925 41713 232401
rect 0 231757 41657 231925
rect 42444 238134 42472 281318
rect 42628 274582 42656 317154
rect 42708 314026 42760 314090
rect 42616 274530 42668 274582
rect 42536 274518 42668 274530
rect 42536 274502 42656 274518
rect 42432 238070 42484 238134
rect 0 231281 41713 231757
rect 41788 231678 41840 231742
rect 0 231113 41657 231281
rect 41800 231225 41828 231678
rect 41713 231169 42193 231225
rect 0 230729 41713 231113
rect 0 230561 41657 230729
rect 0 230085 41713 230561
rect 0 229917 41657 230085
rect 0 229441 41713 229917
rect 0 229273 41657 229441
rect 0 228889 41713 229273
rect 0 228721 41657 228889
rect 0 228245 41713 228721
rect 41788 228618 41840 228682
rect 0 228077 41657 228245
rect 41800 228189 41828 228618
rect 41713 228133 42193 228189
rect 41722 228126 41828 228133
rect 0 227601 41713 228077
rect 0 227433 41657 227601
rect 42248 227462 42300 227526
rect 0 227049 41713 227433
rect 0 226881 41657 227049
rect 0 226405 41713 226881
rect 0 226237 41657 226405
rect 0 225761 41713 226237
rect 0 225593 41657 225761
rect 0 225209 41713 225593
rect 0 225041 41657 225209
rect 0 224842 41713 225041
rect 0 197373 41713 197583
rect 42260 197418 42288 227462
rect 42444 226334 42472 238070
rect 42536 231742 42564 274502
rect 42720 271930 42748 314026
rect 42812 281382 42840 325450
rect 673564 295334 673592 337486
rect 673748 334490 673776 379646
rect 675887 383967 717600 384351
rect 675943 383799 717600 383967
rect 675887 383323 717600 383799
rect 675407 383239 675887 383267
rect 675404 383211 675887 383239
rect 675404 382770 675432 383211
rect 675943 383155 717600 383323
rect 675392 382706 675444 382770
rect 675887 382679 717600 383155
rect 675943 382511 717600 382679
rect 675887 382127 717600 382511
rect 675943 381959 717600 382127
rect 675887 381483 717600 381959
rect 675943 381315 717600 381483
rect 675887 380839 717600 381315
rect 675943 380671 717600 380839
rect 675887 380287 717600 380671
rect 675407 380188 675887 380231
rect 675404 380175 675887 380188
rect 675404 379710 675432 380175
rect 675943 380119 717600 380287
rect 675392 379646 675444 379710
rect 675887 379643 717600 380119
rect 675943 379475 717600 379643
rect 675887 378999 717600 379475
rect 675407 378929 675887 378943
rect 675312 378901 675887 378929
rect 673920 372302 673972 372366
rect 673736 334426 673788 334490
rect 673472 295306 673592 295334
rect 673472 293214 673500 295306
rect 673932 328098 673960 372302
rect 675312 370925 675340 378901
rect 675407 378887 675887 378901
rect 675943 378831 717600 378999
rect 675887 378355 717600 378831
rect 675943 378187 717600 378355
rect 675887 377803 717600 378187
rect 675943 377635 717600 377803
rect 675887 377159 717600 377635
rect 675943 376991 717600 377159
rect 675887 376515 717600 376991
rect 675943 376347 717600 376515
rect 675887 375963 717600 376347
rect 675407 375851 675887 375907
rect 675943 375795 717600 375963
rect 675887 375319 717600 375795
rect 675943 375151 717600 375319
rect 675887 374675 717600 375151
rect 675407 374563 675887 374619
rect 675943 374507 717600 374675
rect 675887 374123 717600 374507
rect 675407 374011 675887 374067
rect 675943 373955 717600 374123
rect 675887 373479 717600 373955
rect 675943 373311 717600 373479
rect 675887 372835 717600 373311
rect 675407 372751 675887 372779
rect 675404 372723 675887 372751
rect 675404 372366 675432 372723
rect 675943 372667 717600 372835
rect 675392 372302 675444 372366
rect 675887 372283 717600 372667
rect 675407 372171 675887 372227
rect 675943 372115 717600 372283
rect 675887 371639 717600 372115
rect 675943 371471 717600 371639
rect 675887 370995 717600 371471
rect 675407 370925 675887 370939
rect 675312 370897 675887 370925
rect 675407 370883 675887 370897
rect 675943 370827 717600 370995
rect 675887 370617 717600 370827
rect 675887 341159 717600 341358
rect 675943 340991 717600 341159
rect 675887 340607 717600 340991
rect 675943 340439 717600 340607
rect 675887 339963 717600 340439
rect 675943 339795 717600 339963
rect 675887 339319 717600 339795
rect 675943 339151 717600 339319
rect 675887 338767 717600 339151
rect 675943 338599 717600 338767
rect 674012 334426 674064 334490
rect 673920 328034 673972 328098
rect 673460 293150 673512 293214
rect 42800 281318 42852 281382
rect 42708 271866 42760 271930
rect 42720 245654 42748 271866
rect 673472 248606 673500 293150
rect 673552 289478 673604 289542
rect 673460 248542 673512 248606
rect 42628 245626 42748 245654
rect 42524 231678 42576 231742
rect 42536 227526 42564 231678
rect 42628 228682 42656 245626
rect 673564 244934 673592 289478
rect 673932 283082 673960 328034
rect 674024 289542 674052 334426
rect 675887 338123 717600 338599
rect 675407 338028 675887 338067
rect 675404 338011 675887 338028
rect 675404 337550 675432 338011
rect 675943 337955 717600 338123
rect 675392 337486 675444 337550
rect 675887 337479 717600 337955
rect 675943 337311 717600 337479
rect 675887 336927 717600 337311
rect 675943 336759 717600 336927
rect 675887 336283 717600 336759
rect 675943 336115 717600 336283
rect 675887 335639 717600 336115
rect 675943 335471 717600 335639
rect 675887 335087 717600 335471
rect 675407 335003 675887 335031
rect 675404 334975 675887 335003
rect 675404 334490 675432 334975
rect 675943 334919 717600 335087
rect 675392 334426 675444 334490
rect 675887 334443 717600 334919
rect 675943 334275 717600 334443
rect 675887 333799 717600 334275
rect 675407 333729 675887 333743
rect 675312 333701 675887 333729
rect 675312 325725 675340 333701
rect 675407 333687 675887 333701
rect 675943 333631 717600 333799
rect 675887 333155 717600 333631
rect 675943 332987 717600 333155
rect 675887 332603 717600 332987
rect 675943 332435 717600 332603
rect 675887 331959 717600 332435
rect 675943 331791 717600 331959
rect 675887 331315 717600 331791
rect 675943 331147 717600 331315
rect 675887 330763 717600 331147
rect 675407 330651 675887 330707
rect 675943 330595 717600 330763
rect 675887 330119 717600 330595
rect 675943 329951 717600 330119
rect 675887 329475 717600 329951
rect 675407 329363 675887 329419
rect 675943 329307 717600 329475
rect 675887 328923 717600 329307
rect 675407 328811 675887 328867
rect 675943 328755 717600 328923
rect 675887 328279 717600 328755
rect 675943 328111 717600 328279
rect 675392 328034 675444 328098
rect 675404 327579 675432 328034
rect 675887 327635 717600 328111
rect 675404 327556 675887 327579
rect 675407 327523 675887 327556
rect 675943 327467 717600 327635
rect 675887 327083 717600 327467
rect 675407 326971 675887 327027
rect 675943 326915 717600 327083
rect 675887 326439 717600 326915
rect 675943 326271 717600 326439
rect 675887 325795 717600 326271
rect 675407 325725 675887 325739
rect 675312 325697 675887 325725
rect 675407 325683 675887 325697
rect 675943 325627 717600 325795
rect 675887 325417 717600 325627
rect 675887 296159 717600 296358
rect 675943 295991 717600 296159
rect 675887 295607 717600 295991
rect 675943 295439 717600 295607
rect 675887 294963 717600 295439
rect 675943 294795 717600 294963
rect 675887 294319 717600 294795
rect 675943 294151 717600 294319
rect 675887 293767 717600 294151
rect 674012 289478 674064 289542
rect 675943 293599 717600 293767
rect 675392 293150 675444 293214
rect 675404 293067 675432 293150
rect 675887 293123 717600 293599
rect 675404 293012 675887 293067
rect 675407 293011 675887 293012
rect 675943 292955 717600 293123
rect 675887 292479 717600 292955
rect 675943 292311 717600 292479
rect 675887 291927 717600 292311
rect 675943 291759 717600 291927
rect 675887 291283 717600 291759
rect 675943 291115 717600 291283
rect 675887 290639 717600 291115
rect 675943 290471 717600 290639
rect 675887 290087 717600 290471
rect 675407 290020 675887 290031
rect 675404 289975 675887 290020
rect 675404 289542 675432 289975
rect 675943 289919 717600 290087
rect 675392 289478 675444 289542
rect 675887 289443 717600 289919
rect 675943 289275 717600 289443
rect 675887 288799 717600 289275
rect 675407 288729 675887 288743
rect 675312 288701 675887 288729
rect 673920 283018 673972 283082
rect 673932 276014 673960 283018
rect 675312 280725 675340 288701
rect 675407 288687 675887 288701
rect 675943 288631 717600 288799
rect 675887 288155 717600 288631
rect 675943 287987 717600 288155
rect 675887 287603 717600 287987
rect 675943 287435 717600 287603
rect 675887 286959 717600 287435
rect 675943 286791 717600 286959
rect 675887 286315 717600 286791
rect 675943 286147 717600 286315
rect 675887 285763 717600 286147
rect 675407 285651 675887 285707
rect 675943 285595 717600 285763
rect 675887 285119 717600 285595
rect 675943 284951 717600 285119
rect 675887 284475 717600 284951
rect 675407 284363 675887 284419
rect 675943 284307 717600 284475
rect 675887 283923 717600 284307
rect 675407 283811 675887 283867
rect 675943 283755 717600 283923
rect 675887 283279 717600 283755
rect 675943 283111 717600 283279
rect 675392 283018 675444 283082
rect 675404 282579 675432 283018
rect 675887 282635 717600 283111
rect 675404 282540 675887 282579
rect 675407 282523 675887 282540
rect 675943 282467 717600 282635
rect 675887 282083 717600 282467
rect 675407 281971 675887 282027
rect 675943 281915 717600 282083
rect 675887 281439 717600 281915
rect 675943 281271 717600 281439
rect 675887 280795 717600 281271
rect 675407 280725 675887 280739
rect 675312 280697 675887 280725
rect 675407 280683 675887 280697
rect 675943 280627 717600 280795
rect 675887 280417 717600 280627
rect 673748 275986 673960 276014
rect 673748 264974 673776 275986
rect 673748 264946 673960 264974
rect 673552 244870 673604 244934
rect 42616 228618 42668 228682
rect 42524 227462 42576 227526
rect 42444 226306 42564 226334
rect 42260 197390 42380 197418
rect 0 197205 41657 197373
rect 41713 197282 42193 197317
rect 41713 197261 42288 197282
rect 41722 197254 42288 197261
rect 0 196729 41713 197205
rect 0 196561 41657 196729
rect 0 196085 41713 196561
rect 0 195917 41657 196085
rect 41713 195973 42193 196029
rect 0 195533 41713 195917
rect 41788 195842 41840 195906
rect 0 195365 41657 195533
rect 41800 195477 41828 195842
rect 41713 195421 42193 195477
rect 0 194889 41713 195365
rect 0 194721 41657 194889
rect 0 194245 41713 194721
rect 0 194077 41657 194245
rect 41713 194133 42193 194189
rect 0 193693 41713 194077
rect 0 193525 41657 193693
rect 41713 193581 42193 193637
rect 0 193049 41713 193525
rect 0 192881 41657 193049
rect 0 192405 41713 192881
rect 0 192237 41657 192405
rect 41713 192293 42193 192349
rect 0 191853 41713 192237
rect 0 191685 41657 191853
rect 0 191209 41713 191685
rect 0 191041 41657 191209
rect 0 190565 41713 191041
rect 0 190397 41657 190565
rect 0 190013 41713 190397
rect 0 189845 41657 190013
rect 0 189369 41713 189845
rect 42260 189394 42288 197254
rect 0 189201 41657 189369
rect 41892 189366 42288 189394
rect 41892 189313 41920 189366
rect 41713 189257 42193 189313
rect 0 188725 41713 189201
rect 0 188557 41657 188725
rect 0 188081 41713 188557
rect 42352 188170 42380 197390
rect 42536 195906 42564 226306
rect 42524 195842 42576 195906
rect 41892 188142 42380 188170
rect 0 187913 41657 188081
rect 41892 188034 41920 188142
rect 41722 188025 41920 188034
rect 41984 188025 42012 188142
rect 41713 187969 42193 188025
rect 0 187529 41713 187913
rect 41984 187610 42012 187969
rect 41972 187546 42024 187610
rect 0 187361 41657 187529
rect 0 186885 41713 187361
rect 0 186717 41657 186885
rect 0 186241 41713 186717
rect 0 186073 41657 186241
rect 0 185689 41713 186073
rect 0 185521 41657 185689
rect 0 185045 41713 185521
rect 0 184877 41657 185045
rect 41713 184933 42193 184989
rect 0 184401 41713 184877
rect 41800 184482 41828 184933
rect 41788 184418 41840 184482
rect 0 184233 41657 184401
rect 42536 187694 42564 195842
rect 42444 187666 42564 187694
rect 0 183849 41713 184233
rect 42248 184146 42300 184210
rect 0 183681 41657 183849
rect 0 183205 41713 183681
rect 0 183037 41657 183205
rect 0 182561 41713 183037
rect 0 182393 41657 182561
rect 0 182009 41713 182393
rect 0 181841 41657 182009
rect 0 181642 41713 181841
rect 985 120278 40000 125058
rect 985 115079 39593 120278
rect 39616 115379 40000 115779
rect 985 110299 40000 115079
rect 985 110253 39593 110299
rect 30753 83000 31683 85228
rect 31928 83049 32702 85239
rect 714 82940 39593 83000
rect 714 78819 39600 82940
rect 714 78707 39593 78819
rect 714 72185 39600 78707
rect 714 72099 39593 72185
rect 714 68100 39600 72099
rect 714 68098 39593 68100
rect 42260 45626 42288 184146
rect 42444 82890 42472 187666
rect 42524 187546 42576 187610
rect 42536 121514 42564 187546
rect 42628 184482 42656 228618
rect 673564 199306 673592 244870
rect 673932 237726 673960 264946
rect 675887 251159 717600 251358
rect 675943 250991 717600 251159
rect 675887 250607 717600 250991
rect 675943 250439 717600 250607
rect 675887 249963 717600 250439
rect 675943 249795 717600 249963
rect 675887 249319 717600 249795
rect 675943 249151 717600 249319
rect 675887 248767 717600 249151
rect 674012 248542 674064 248606
rect 673920 237662 673972 237726
rect 673552 199242 673604 199306
rect 42616 184418 42668 184482
rect 673460 158306 673512 158370
rect 42524 121450 42576 121514
rect 44180 121450 44232 121514
rect 44192 110537 44220 121450
rect 673472 113218 673500 158306
rect 673564 155242 673592 199242
rect 673932 191962 673960 237662
rect 674024 202366 674052 248542
rect 675392 248542 675444 248606
rect 675943 248599 717600 248767
rect 675404 248067 675432 248542
rect 675887 248123 717600 248599
rect 675404 248039 675887 248067
rect 675407 248011 675887 248039
rect 675943 247955 717600 248123
rect 675887 247479 717600 247955
rect 675943 247311 717600 247479
rect 675887 246927 717600 247311
rect 675943 246759 717600 246927
rect 675887 246283 717600 246759
rect 675943 246115 717600 246283
rect 675887 245639 717600 246115
rect 675943 245471 717600 245639
rect 675887 245087 717600 245471
rect 675407 245004 675887 245031
rect 675404 244975 675887 245004
rect 675404 244934 675432 244975
rect 675392 244870 675444 244934
rect 675943 244919 717600 245087
rect 675887 244443 717600 244919
rect 675943 244275 717600 244443
rect 675887 243799 717600 244275
rect 675407 243729 675887 243743
rect 675312 243701 675887 243729
rect 675312 235725 675340 243701
rect 675407 243687 675887 243701
rect 675943 243631 717600 243799
rect 675887 243155 717600 243631
rect 675943 242987 717600 243155
rect 675887 242603 717600 242987
rect 675943 242435 717600 242603
rect 675887 241959 717600 242435
rect 675943 241791 717600 241959
rect 675887 241315 717600 241791
rect 675943 241147 717600 241315
rect 675887 240763 717600 241147
rect 675407 240651 675887 240707
rect 675943 240595 717600 240763
rect 675887 240119 717600 240595
rect 675943 239951 717600 240119
rect 675887 239475 717600 239951
rect 675407 239363 675887 239419
rect 675943 239307 717600 239475
rect 675887 238923 717600 239307
rect 675407 238811 675887 238867
rect 675943 238755 717600 238923
rect 675887 238279 717600 238755
rect 675943 238111 717600 238279
rect 675392 237662 675444 237726
rect 675404 237579 675432 237662
rect 675887 237635 717600 238111
rect 675404 237524 675887 237579
rect 675407 237523 675887 237524
rect 675943 237467 717600 237635
rect 675887 237083 717600 237467
rect 675407 236971 675887 237027
rect 675943 236915 717600 237083
rect 675887 236439 717600 236915
rect 675943 236271 717600 236439
rect 675887 235795 717600 236271
rect 675407 235725 675887 235739
rect 675312 235697 675887 235725
rect 675407 235683 675887 235697
rect 675943 235627 717600 235795
rect 675887 235417 717600 235627
rect 675887 205959 717600 206158
rect 675943 205791 717600 205959
rect 675887 205407 717600 205791
rect 675943 205239 717600 205407
rect 675887 204763 717600 205239
rect 675943 204595 717600 204763
rect 675887 204119 717600 204595
rect 675943 203951 717600 204119
rect 675887 203567 717600 203951
rect 674012 202302 674064 202366
rect 673920 191898 673972 191962
rect 673552 155178 673604 155242
rect 673460 113154 673512 113218
rect 44178 110463 44234 110537
rect 44822 110463 44878 110537
rect 44836 110414 44864 110463
rect 44836 110386 44956 110414
rect 42432 82826 42484 82890
rect 44180 82826 44232 82890
rect 44192 71913 44220 82826
rect 44178 71839 44234 71913
rect 44822 71839 44878 71913
rect 44836 46986 44864 71839
rect 44824 46922 44876 46986
rect 42248 45562 42300 45626
rect 44928 45558 44956 110386
rect 149060 46854 149112 46918
rect 188528 46854 188580 46918
rect 200856 46854 200908 46918
rect 256240 46854 256292 46918
rect 297732 46854 297784 46918
rect 309416 46854 309468 46918
rect 352564 46854 352616 46918
rect 364248 46854 364300 46918
rect 407396 46854 407448 46918
rect 419080 46854 419132 46918
rect 462136 46854 462188 46918
rect 473820 46854 473872 46918
rect 516968 46854 517020 46918
rect 140964 45562 141016 45626
rect 44916 45494 44968 45558
rect 93768 41482 93820 41546
rect 93780 40225 93808 41482
rect 135168 40225 135220 40254
rect 93766 40151 93822 40225
rect 135166 40151 135222 40225
rect 140976 40202 141004 45562
rect 143540 40225 143592 40254
rect 140976 40174 141036 40202
rect 141008 40118 141036 40174
rect 143078 40151 143134 40225
rect 143538 40151 143594 40225
rect 147128 41822 147180 41886
rect 143084 40118 143112 40151
rect 140996 40054 141048 40118
rect 143072 40054 143124 40118
rect 144552 40054 144604 40118
rect 141008 40000 141036 40054
rect 143084 40000 143112 40054
rect 144564 40000 144592 40054
rect 147140 40118 147168 41822
rect 149072 40361 149100 46854
rect 188540 44334 188568 46854
rect 195980 45494 196032 45558
rect 195992 44470 196020 45494
rect 195980 44406 196032 44470
rect 188528 44270 188580 44334
rect 192852 44270 192904 44334
rect 186688 44202 186740 44266
rect 186700 42193 186728 44202
rect 188540 42193 188568 44270
rect 192864 42193 192892 44270
rect 194692 44202 194744 44266
rect 194704 42193 194732 44202
rect 195992 42193 196020 44406
rect 200868 42193 200896 46854
rect 201500 44270 201552 44334
rect 201512 42193 201540 44270
rect 186683 41713 186739 42193
rect 187971 41713 188027 42193
rect 188523 41713 188579 42193
rect 189167 41834 189223 42193
rect 189264 41890 189316 41954
rect 189276 41834 189304 41890
rect 189167 41806 189304 41834
rect 189167 41713 189223 41806
rect 189811 41713 189867 42193
rect 190363 41713 190419 42193
rect 191007 41834 191063 42193
rect 191104 41890 191156 41954
rect 191116 41834 191144 41890
rect 191007 41806 191144 41834
rect 191007 41713 191063 41806
rect 191651 41713 191707 42193
rect 192203 41834 192259 42193
rect 192300 41890 192352 41954
rect 192312 41834 192340 41890
rect 192203 41806 192340 41834
rect 192203 41713 192259 41806
rect 192847 41713 192903 42193
rect 193491 41834 193547 42193
rect 193588 41890 193640 41954
rect 193600 41834 193628 41890
rect 193491 41806 193628 41834
rect 193491 41713 193547 41806
rect 194687 41713 194743 42193
rect 195975 41713 196031 42193
rect 196440 41890 196492 41954
rect 196452 41834 196480 41890
rect 196527 41834 196583 42193
rect 197171 41834 197227 42193
rect 197815 41834 197871 42193
rect 198367 41834 198423 42193
rect 198464 41890 198516 41954
rect 198476 41834 198504 41890
rect 199011 41834 199067 42193
rect 196452 41806 198504 41834
rect 198936 41818 199067 41834
rect 198924 41806 199067 41818
rect 196527 41713 196583 41806
rect 197171 41713 197227 41806
rect 197815 41713 197871 41806
rect 198367 41713 198423 41806
rect 198924 41754 198976 41806
rect 199011 41713 199067 41806
rect 200120 41890 200172 41954
rect 200132 41834 200160 41890
rect 200207 41834 200263 42193
rect 200851 41834 200907 42193
rect 200132 41806 200907 41834
rect 200207 41713 200263 41806
rect 200851 41713 200907 41806
rect 201495 41713 201551 42193
rect 202047 41713 202103 42193
rect 186417 41657 186627 41713
rect 186795 41657 187271 41713
rect 187439 41657 187915 41713
rect 188083 41657 188467 41713
rect 188635 41657 189111 41713
rect 189279 41657 189755 41713
rect 189923 41657 190307 41713
rect 190475 41657 190951 41713
rect 191119 41657 191595 41713
rect 191763 41657 192147 41713
rect 192315 41657 192791 41713
rect 192959 41657 193435 41713
rect 193603 41657 193987 41713
rect 194155 41657 194631 41713
rect 194799 41657 195275 41713
rect 195443 41657 195919 41713
rect 196087 41657 196471 41713
rect 196639 41657 197115 41713
rect 197283 41657 197759 41713
rect 197927 41657 198311 41713
rect 198479 41657 198955 41713
rect 199123 41657 199599 41713
rect 199767 41657 200151 41713
rect 200319 41657 200795 41713
rect 200963 41657 201439 41713
rect 201607 41657 201991 41713
rect 202159 41657 202358 41713
rect 149058 40287 149114 40361
rect 147128 40054 147180 40118
rect 78942 39593 83722 40000
rect 88221 39616 88621 40000
rect 88921 39593 93701 40000
rect 132617 39878 132897 40000
rect 132953 39934 133157 40000
rect 133213 39878 140940 40000
rect 132617 39816 140940 39878
rect 140996 39872 141048 40000
rect 141104 39878 141313 40000
rect 141369 39934 141499 40000
rect 141555 39878 141611 40000
rect 141667 39934 141813 40000
rect 141869 39878 141898 40000
rect 141954 39934 142084 40000
rect 142140 39878 143012 40000
rect 141104 39816 143012 39878
rect 78942 985 93747 39593
rect 132617 39204 143012 39816
rect 132617 39147 142955 39204
rect 143068 39151 143128 40000
rect 143184 39662 143299 40000
rect 143355 39718 143585 40000
rect 143641 39831 143762 40000
rect 143818 39887 144151 40000
rect 144207 39831 144517 40000
rect 144564 39916 144689 40000
rect 143641 39747 144517 39831
rect 144573 39803 144689 39916
rect 144745 39747 145035 40000
rect 143641 39662 145035 39747
rect 145199 39878 145765 40000
rect 145821 39934 145915 40000
rect 145971 39878 147532 40000
rect 143184 39650 145035 39662
rect 145199 39650 147532 39878
rect 143184 39369 147532 39650
rect 143184 39297 144495 39369
rect 145520 39341 147532 39369
rect 143184 39243 144441 39297
rect 144551 39285 145464 39313
rect 144551 39271 145530 39285
rect 145586 39275 147532 39341
rect 144551 39261 145436 39271
rect 143184 39207 144367 39243
rect 144551 39241 144623 39261
rect 144625 39241 144645 39261
rect 145414 39247 145461 39261
rect 145464 39247 145530 39271
rect 143244 39169 144367 39207
rect 144497 39233 144551 39241
rect 144571 39233 144625 39241
rect 144497 39205 144625 39233
rect 145414 39219 145530 39247
rect 145414 39214 145461 39219
rect 144497 39187 144551 39205
rect 144571 39187 144625 39205
rect 143068 39148 143188 39151
rect 132617 39076 141720 39147
rect 143011 39091 143188 39148
rect 143244 39147 144345 39169
rect 144423 39113 144571 39187
rect 144701 39185 145358 39205
rect 144681 39158 145358 39185
rect 145461 39191 145525 39214
rect 145530 39191 145599 39219
rect 145655 39206 147532 39275
rect 145461 39163 145599 39191
rect 144681 39131 145405 39158
rect 145461 39150 145525 39163
rect 145530 39150 145599 39163
rect 144401 39091 144497 39113
rect 132617 39010 141654 39076
rect 141776 39063 144497 39091
rect 141776 39049 141847 39063
rect 143068 39049 143128 39063
rect 144423 39049 144497 39063
rect 144627 39094 145405 39131
rect 145525 39135 145591 39150
rect 145599 39135 145653 39150
rect 144627 39057 145469 39094
rect 145525 39085 145653 39135
rect 145525 39084 145591 39085
rect 141776 39039 144497 39049
rect 141776 39020 141847 39039
rect 141850 39020 141869 39039
rect 144553 39028 145469 39057
rect 141710 39011 141776 39020
rect 141784 39011 141850 39020
rect 132617 37861 141628 39010
rect 141710 38969 141850 39011
rect 144553 38983 145545 39028
rect 141710 38954 141776 38969
rect 141784 38954 141850 38969
rect 141925 38964 145545 38983
rect 141684 38928 141710 38954
rect 141736 38928 141784 38954
rect 141684 38906 141784 38928
rect 132617 37823 141590 37861
rect 132617 36927 141538 37823
rect 141684 37805 141736 38906
rect 141906 38898 145545 38964
rect 141840 38850 145545 38898
rect 141646 37783 141736 37805
rect 141646 37767 141684 37783
rect 141720 37767 141736 37783
rect 141792 38284 145545 38850
rect 141792 38216 145477 38284
rect 145601 38228 145653 39085
rect 141792 38176 145437 38216
rect 145533 38178 145653 38228
rect 141792 38110 145371 38176
rect 145533 38160 145601 38178
rect 145607 38160 145653 38178
rect 145493 38150 145533 38160
rect 145567 38150 145607 38160
rect 145493 38136 145607 38150
rect 145493 38120 145533 38136
rect 145567 38120 145607 38136
rect 141594 37693 141720 37767
rect 141792 37711 145319 38110
rect 145427 38108 145493 38120
rect 145501 38108 145567 38120
rect 145427 38080 145567 38108
rect 145709 38104 147532 39206
rect 145427 38054 145493 38080
rect 145501 38054 145567 38080
rect 145663 38064 147532 38104
rect 132617 36860 141471 36927
rect 141594 36871 141646 37693
rect 141776 37637 145319 37711
rect 132617 35845 141419 36860
rect 141527 36821 141646 36871
rect 141527 36804 141594 36821
rect 141601 36804 141646 36821
rect 141475 36730 141601 36804
rect 141702 36748 145319 37637
rect 141475 35901 141527 36730
rect 141657 36674 145319 36748
rect 141583 35845 145319 36674
rect 132617 34484 145319 35845
rect 145375 37980 145501 38054
rect 145623 37998 147532 38064
rect 145375 34678 145427 37980
rect 145557 37924 147532 37998
rect 145483 34734 147532 37924
rect 145375 34540 145470 34678
rect 132617 34469 145362 34484
rect 132617 33839 145319 34469
rect 145418 34413 145470 34540
rect 145375 34371 145470 34413
rect 145375 34370 145418 34371
rect 145375 34275 145470 34370
rect 132617 33810 145290 33839
rect 132617 33765 145245 33810
rect 145375 33783 145427 34275
rect 145526 34219 147532 34734
rect 132617 32852 145240 33765
rect 145346 33754 145427 33783
rect 145301 33747 145346 33754
rect 145375 33747 145427 33754
rect 145301 33733 145427 33747
rect 145301 33709 145346 33733
rect 145375 33709 145427 33733
rect 145296 33704 145301 33709
rect 145348 33704 145375 33709
rect 145296 33682 145375 33704
rect 132617 32688 145114 32852
rect 145296 32796 145348 33682
rect 145483 33653 147532 34219
rect 145431 33626 147532 33653
rect 145170 32744 145348 32796
rect 145404 32688 147532 33626
rect 132617 158 147532 32688
rect 186417 0 202358 41657
rect 241260 39593 245381 39600
rect 245493 39593 252015 39600
rect 252101 39593 256100 39600
rect 238961 31928 241151 32702
rect 241200 31683 256100 39593
rect 256252 39545 256280 46854
rect 297088 44270 297140 44334
rect 295248 44134 295300 44198
rect 295260 42193 295288 44134
rect 297100 42193 297128 44270
rect 297744 42193 297772 46854
rect 304540 44406 304592 44470
rect 306288 44406 306340 44470
rect 299572 44270 299624 44334
rect 299584 42193 299612 44270
rect 303252 44134 303304 44198
rect 303264 42193 303292 44134
rect 304552 42193 304580 44406
rect 305736 44270 305788 44334
rect 305748 42193 305776 44270
rect 306300 44198 306328 44406
rect 306288 44134 306340 44198
rect 309428 42193 309456 46854
rect 351920 44338 351972 44402
rect 350080 44134 350132 44198
rect 350092 42193 350120 44134
rect 351932 42193 351960 44338
rect 352576 42193 352604 46854
rect 354404 44338 354456 44402
rect 360568 44338 360620 44402
rect 354416 42193 354444 44338
rect 358084 44134 358136 44198
rect 358096 42193 358124 44134
rect 359372 44202 359424 44266
rect 359384 42193 359412 44202
rect 360580 42193 360608 44338
rect 364260 42193 364288 46854
rect 406752 44406 406804 44470
rect 406764 44334 406792 44406
rect 404910 44231 404966 44305
rect 406752 44270 406804 44334
rect 404924 42193 404952 44231
rect 406764 42193 406792 44270
rect 407408 42193 407436 46854
rect 412914 44231 412970 44305
rect 412928 42193 412956 44231
rect 414204 44134 414256 44198
rect 414216 42193 414244 44134
rect 419092 42193 419120 46854
rect 461492 44406 461544 44470
rect 459650 44231 459706 44305
rect 461504 44266 461532 44406
rect 459664 42193 459692 44231
rect 461492 44202 461544 44266
rect 461504 42193 461532 44202
rect 462148 42193 462176 46854
rect 468944 44406 468996 44470
rect 467654 44231 467710 44305
rect 467668 42193 467696 44231
rect 468956 44334 468984 44406
rect 468944 44270 468996 44334
rect 468956 42193 468984 44270
rect 473832 42193 473860 46854
rect 514482 44231 514538 44305
rect 514496 42193 514524 44231
rect 516324 44202 516376 44266
rect 516336 42193 516364 44202
rect 516980 42193 517008 46854
rect 523776 45562 523828 45626
rect 518716 45494 518768 45558
rect 518728 44266 518756 45494
rect 523788 44470 523816 45562
rect 522486 44367 522542 44441
rect 523776 44406 523828 44470
rect 518716 44202 518768 44266
rect 522500 42193 522528 44367
rect 523788 42193 523816 44406
rect 673472 42770 673500 113154
rect 673564 109546 673592 155178
rect 673932 146946 673960 191898
rect 674024 158370 674052 202302
rect 675943 203399 717600 203567
rect 675887 202923 717600 203399
rect 675407 202844 675887 202867
rect 675404 202811 675887 202844
rect 675404 202366 675432 202811
rect 675943 202755 717600 202923
rect 675392 202302 675444 202366
rect 675887 202279 717600 202755
rect 675943 202111 717600 202279
rect 675887 201727 717600 202111
rect 675943 201559 717600 201727
rect 675887 201083 717600 201559
rect 675943 200915 717600 201083
rect 675887 200439 717600 200915
rect 675943 200271 717600 200439
rect 675887 199887 717600 200271
rect 675407 199803 675887 199831
rect 675404 199775 675887 199803
rect 675404 199306 675432 199775
rect 675943 199719 717600 199887
rect 675392 199242 675444 199306
rect 675887 199243 717600 199719
rect 675943 199075 717600 199243
rect 675312 198614 675432 198642
rect 675312 190525 675340 198614
rect 675404 198543 675432 198614
rect 675887 198599 717600 199075
rect 675404 198492 675887 198543
rect 675407 198487 675887 198492
rect 675943 198431 717600 198599
rect 675887 197955 717600 198431
rect 675943 197787 717600 197955
rect 675887 197403 717600 197787
rect 675943 197235 717600 197403
rect 675887 196759 717600 197235
rect 675943 196591 717600 196759
rect 675887 196115 717600 196591
rect 675943 195947 717600 196115
rect 675887 195563 717600 195947
rect 675407 195451 675887 195507
rect 675943 195395 717600 195563
rect 675887 194919 717600 195395
rect 675943 194751 717600 194919
rect 675887 194275 717600 194751
rect 675407 194163 675887 194219
rect 675943 194107 717600 194275
rect 675887 193723 717600 194107
rect 675407 193611 675887 193667
rect 675943 193555 717600 193723
rect 675887 193079 717600 193555
rect 675943 192911 717600 193079
rect 675887 192435 717600 192911
rect 675407 192372 675887 192379
rect 675404 192323 675887 192372
rect 675404 191962 675432 192323
rect 675943 192267 717600 192435
rect 675392 191898 675444 191962
rect 675887 191883 717600 192267
rect 675407 191771 675887 191827
rect 675943 191715 717600 191883
rect 675887 191239 717600 191715
rect 675943 191071 717600 191239
rect 675887 190595 717600 191071
rect 675407 190525 675887 190539
rect 675312 190497 675887 190525
rect 675407 190483 675887 190497
rect 675943 190427 717600 190595
rect 675887 190217 717600 190427
rect 675887 160959 717600 161158
rect 675943 160791 717600 160959
rect 675887 160407 717600 160791
rect 675943 160239 717600 160407
rect 675887 159763 717600 160239
rect 675943 159595 717600 159763
rect 675887 159119 717600 159595
rect 675943 158951 717600 159119
rect 675887 158567 717600 158951
rect 674012 158306 674064 158370
rect 675943 158399 717600 158567
rect 675392 158306 675444 158370
rect 675404 157867 675432 158306
rect 675887 157923 717600 158399
rect 675404 157828 675887 157867
rect 675407 157811 675887 157828
rect 675943 157755 717600 157923
rect 675887 157279 717600 157755
rect 675943 157111 717600 157279
rect 675887 156727 717600 157111
rect 675943 156559 717600 156727
rect 675887 156083 717600 156559
rect 675943 155915 717600 156083
rect 675887 155439 717600 155915
rect 675943 155271 717600 155439
rect 675392 155178 675444 155242
rect 675404 154831 675432 155178
rect 675887 154887 717600 155271
rect 675404 154803 675887 154831
rect 675407 154775 675887 154803
rect 675943 154719 717600 154887
rect 675887 154243 717600 154719
rect 675943 154075 717600 154243
rect 675887 153599 717600 154075
rect 675407 153529 675887 153543
rect 675312 153501 675887 153529
rect 673736 146882 673788 146946
rect 673920 146882 673972 146946
rect 673552 109482 673604 109546
rect 673564 45626 673592 109482
rect 673748 101726 673776 146882
rect 675312 145525 675340 153501
rect 675407 153487 675887 153501
rect 675943 153431 717600 153599
rect 675887 152955 717600 153431
rect 675943 152787 717600 152955
rect 675887 152403 717600 152787
rect 675943 152235 717600 152403
rect 675887 151759 717600 152235
rect 675943 151591 717600 151759
rect 675887 151115 717600 151591
rect 675943 150947 717600 151115
rect 675887 150563 717600 150947
rect 675407 150451 675887 150507
rect 675943 150395 717600 150563
rect 675887 149919 717600 150395
rect 675943 149751 717600 149919
rect 675887 149275 717600 149751
rect 675407 149163 675887 149219
rect 675943 149107 717600 149275
rect 675887 148723 717600 149107
rect 675407 148611 675887 148667
rect 675943 148555 717600 148723
rect 675887 148079 717600 148555
rect 675943 147911 717600 148079
rect 675887 147435 717600 147911
rect 675407 147356 675887 147379
rect 675404 147323 675887 147356
rect 675404 146946 675432 147323
rect 675943 147267 717600 147435
rect 675392 146882 675444 146946
rect 675887 146883 717600 147267
rect 675407 146771 675887 146827
rect 675943 146715 717600 146883
rect 675887 146239 717600 146715
rect 675943 146071 717600 146239
rect 675887 145595 717600 146071
rect 675407 145525 675887 145539
rect 675312 145497 675887 145525
rect 675407 145483 675887 145497
rect 675943 145427 717600 145595
rect 675887 145217 717600 145427
rect 675887 115759 717600 115958
rect 675943 115591 717600 115759
rect 675887 115207 717600 115591
rect 675943 115039 717600 115207
rect 675887 114563 717600 115039
rect 675943 114395 717600 114563
rect 675887 113919 717600 114395
rect 675943 113751 717600 113919
rect 675887 113367 717600 113751
rect 675392 113154 675444 113218
rect 675943 113199 717600 113367
rect 675404 112667 675432 113154
rect 675887 112723 717600 113199
rect 675404 112639 675887 112667
rect 675407 112611 675887 112639
rect 675943 112555 717600 112723
rect 675887 112079 717600 112555
rect 675943 111911 717600 112079
rect 675887 111527 717600 111911
rect 675943 111359 717600 111527
rect 675887 110883 717600 111359
rect 675943 110715 717600 110883
rect 675887 110239 717600 110715
rect 675943 110071 717600 110239
rect 675887 109687 717600 110071
rect 675407 109603 675887 109631
rect 675404 109575 675887 109603
rect 675404 109546 675432 109575
rect 675392 109482 675444 109546
rect 675943 109519 717600 109687
rect 675887 109043 717600 109519
rect 675943 108875 717600 109043
rect 675887 108399 717600 108875
rect 675407 108338 675887 108343
rect 675312 108310 675887 108338
rect 673736 101662 673788 101726
rect 673552 45562 673604 45626
rect 673748 45558 673776 101662
rect 675312 100314 675340 108310
rect 675407 108287 675887 108310
rect 675943 108231 717600 108399
rect 675887 107755 717600 108231
rect 675943 107587 717600 107755
rect 675887 107203 717600 107587
rect 675943 107035 717600 107203
rect 675887 106559 717600 107035
rect 675943 106391 717600 106559
rect 675887 105915 717600 106391
rect 675943 105747 717600 105915
rect 675887 105363 717600 105747
rect 675407 105251 675887 105307
rect 675943 105195 717600 105363
rect 675887 104719 717600 105195
rect 675943 104551 717600 104719
rect 675887 104075 717600 104551
rect 675407 103963 675887 104019
rect 675943 103907 717600 104075
rect 675887 103523 717600 103907
rect 675407 103411 675887 103467
rect 675943 103355 717600 103523
rect 675887 102879 717600 103355
rect 675943 102711 717600 102879
rect 675887 102235 717600 102711
rect 675407 102151 675887 102179
rect 675404 102123 675887 102151
rect 675404 101726 675432 102123
rect 675943 102067 717600 102235
rect 675392 101662 675444 101726
rect 675887 101683 717600 102067
rect 675407 101571 675887 101627
rect 675943 101515 717600 101683
rect 675887 101039 717600 101515
rect 675943 100871 717600 101039
rect 675887 100395 717600 100871
rect 675407 100314 675887 100339
rect 675312 100286 675887 100314
rect 675407 100283 675887 100286
rect 675943 100227 717600 100395
rect 675887 100017 717600 100227
rect 673736 45494 673788 45558
rect 579896 42706 579948 42770
rect 673460 42706 673512 42770
rect 295260 41806 295339 42193
rect 295283 41713 295339 41806
rect 295927 41713 295983 42193
rect 296571 41713 296627 42193
rect 297100 41806 297179 42193
rect 297744 41834 297823 42193
rect 297916 41890 297968 41954
rect 297928 41834 297956 41890
rect 297744 41806 297956 41834
rect 297123 41713 297179 41806
rect 297767 41713 297823 41806
rect 298411 41713 298467 42193
rect 298963 41713 299019 42193
rect 299584 41806 299663 42193
rect 299607 41713 299663 41806
rect 300251 41713 300307 42193
rect 300676 41890 300728 41954
rect 300688 41834 300716 41890
rect 300803 41834 300859 42193
rect 301447 41834 301503 42193
rect 302091 41834 302147 42193
rect 302240 41890 302292 41954
rect 302252 41834 302280 41890
rect 300688 41806 302280 41834
rect 300803 41713 300859 41806
rect 301447 41713 301503 41806
rect 302091 41713 302147 41806
rect 303264 41806 303343 42193
rect 304552 41806 304631 42193
rect 303287 41713 303343 41806
rect 304575 41713 304631 41806
rect 305127 41834 305183 42193
rect 305276 41890 305328 41954
rect 305288 41834 305316 41890
rect 305127 41806 305316 41834
rect 305748 41806 305827 42193
rect 305127 41713 305183 41806
rect 305771 41713 305827 41806
rect 306415 41834 306471 42193
rect 306564 41890 306616 41954
rect 306576 41834 306604 41890
rect 306415 41806 306604 41834
rect 306415 41713 306471 41806
rect 307611 41834 307667 42193
rect 307611 41818 307800 41834
rect 307611 41806 307812 41818
rect 308680 41890 308732 41954
rect 308692 41834 308720 41890
rect 308807 41834 308863 42193
rect 309428 41834 309507 42193
rect 308692 41806 309507 41834
rect 307611 41713 307667 41806
rect 307760 41754 307812 41806
rect 308807 41713 308863 41806
rect 309451 41713 309507 41806
rect 310647 41713 310703 42193
rect 350083 41713 350139 42193
rect 350727 41713 350783 42193
rect 351371 41713 351427 42193
rect 351923 41713 351979 42193
rect 352567 41970 352623 42193
rect 352567 41954 352696 41970
rect 352567 41942 352708 41954
rect 352567 41713 352623 41942
rect 352656 41890 352708 41942
rect 353211 41713 353267 42193
rect 353763 41713 353819 42193
rect 354407 41713 354463 42193
rect 355051 41713 355107 42193
rect 355508 41890 355560 41954
rect 355520 41834 355548 41890
rect 355603 41834 355659 42193
rect 356247 41834 356303 42193
rect 356891 41834 356947 42193
rect 356980 41890 357032 41954
rect 356992 41834 357020 41890
rect 355520 41806 357020 41834
rect 355603 41713 355659 41806
rect 356247 41713 356303 41806
rect 356891 41713 356947 41806
rect 358087 41713 358143 42193
rect 359375 41713 359431 42193
rect 359832 41890 359884 41954
rect 359844 41834 359872 41890
rect 359927 41834 359983 42193
rect 359844 41806 359983 41834
rect 359927 41713 359983 41806
rect 360571 41713 360627 42193
rect 361120 41890 361172 41954
rect 361132 41834 361160 41890
rect 361215 41834 361271 42193
rect 361132 41806 361271 41834
rect 361215 41713 361271 41806
rect 362411 41834 362467 42193
rect 362411 41818 362540 41834
rect 362411 41806 362552 41818
rect 362411 41713 362467 41806
rect 362500 41754 362552 41806
rect 363512 41890 363564 41954
rect 363524 41834 363552 41890
rect 363607 41834 363663 42193
rect 364251 41834 364307 42193
rect 363524 41806 364307 41834
rect 363607 41713 363663 41806
rect 364251 41713 364307 41806
rect 365447 41713 365503 42193
rect 404883 41820 404952 42193
rect 404883 41713 404939 41820
rect 406171 41713 406227 42193
rect 406723 41820 406792 42193
rect 407367 41970 407436 42193
rect 407367 41954 407528 41970
rect 407367 41942 407540 41954
rect 407367 41820 407436 41942
rect 407488 41890 407540 41942
rect 406723 41713 406779 41820
rect 407367 41713 407423 41820
rect 408011 41713 408067 42193
rect 408563 41713 408619 42193
rect 409851 41713 409907 42193
rect 410248 41890 410300 41954
rect 410260 41834 410288 41890
rect 410403 41834 410459 42193
rect 410260 41806 410459 41834
rect 410403 41713 410459 41806
rect 411536 41890 411588 41954
rect 411548 41834 411576 41890
rect 411691 41834 411747 42193
rect 411548 41806 411747 41834
rect 411691 41713 411747 41806
rect 412887 41820 412956 42193
rect 414175 41820 414244 42193
rect 414572 41890 414624 41954
rect 414584 41834 414612 41890
rect 414727 41834 414783 42193
rect 415860 41890 415912 41954
rect 412887 41713 412943 41820
rect 414175 41713 414231 41820
rect 414584 41806 414783 41834
rect 414727 41713 414783 41806
rect 415872 41834 415900 41890
rect 416015 41834 416071 42193
rect 415872 41806 416071 41834
rect 416015 41713 416071 41806
rect 417211 41834 417267 42193
rect 417211 41818 417372 41834
rect 418252 41890 418304 41954
rect 418264 41834 418292 41890
rect 418407 41834 418463 42193
rect 419051 41834 419120 42193
rect 418264 41820 419120 41834
rect 417211 41806 417384 41818
rect 417211 41713 417267 41806
rect 417332 41754 417384 41806
rect 418264 41806 419107 41820
rect 418407 41713 418463 41806
rect 419051 41713 419107 41806
rect 420247 41713 420303 42193
rect 459664 41806 459739 42193
rect 459683 41713 459739 41806
rect 460971 41713 461027 42193
rect 461504 41806 461579 42193
rect 462148 41834 462223 42193
rect 462320 41890 462372 41954
rect 462332 41834 462360 41890
rect 462148 41806 462360 41834
rect 461523 41713 461579 41806
rect 462167 41713 462223 41806
rect 462811 41713 462867 42193
rect 463363 41713 463419 42193
rect 464651 41713 464707 42193
rect 465080 41890 465132 41954
rect 465092 41834 465120 41890
rect 465203 41834 465259 42193
rect 465092 41806 465259 41834
rect 466368 41890 466420 41954
rect 466380 41834 466408 41890
rect 466491 41834 466547 42193
rect 466380 41806 466547 41834
rect 465203 41713 465259 41806
rect 466491 41713 466547 41806
rect 467668 41806 467743 42193
rect 468956 41806 469031 42193
rect 469404 41890 469456 41954
rect 469416 41834 469444 41890
rect 469527 41834 469583 42193
rect 470692 41890 470744 41954
rect 469416 41806 469583 41834
rect 467687 41713 467743 41806
rect 468975 41713 469031 41806
rect 469527 41713 469583 41806
rect 470704 41834 470732 41890
rect 470815 41834 470871 42193
rect 470704 41806 470871 41834
rect 470815 41713 470871 41806
rect 472011 41834 472067 42193
rect 472011 41818 472204 41834
rect 472011 41806 472216 41818
rect 473084 41890 473136 41954
rect 473096 41834 473124 41890
rect 473207 41834 473263 42193
rect 473832 41834 473907 42193
rect 473096 41806 473907 41834
rect 472011 41713 472067 41806
rect 472164 41754 472216 41806
rect 473207 41713 473263 41806
rect 473851 41713 473907 41806
rect 475047 41713 475103 42193
rect 514483 41713 514539 42193
rect 515771 41713 515827 42193
rect 516323 41713 516379 42193
rect 516967 41970 517023 42193
rect 516967 41954 517100 41970
rect 516967 41942 517112 41954
rect 516967 41713 517023 41942
rect 517060 41890 517112 41942
rect 517611 41713 517667 42193
rect 518163 41713 518219 42193
rect 519451 41713 519507 42193
rect 519912 41890 519964 41954
rect 519924 41834 519952 41890
rect 520003 41834 520059 42193
rect 519924 41806 520059 41834
rect 520003 41713 520059 41806
rect 521200 41890 521252 41954
rect 521212 41834 521240 41890
rect 521291 41834 521347 42193
rect 521212 41806 521347 41834
rect 521291 41713 521347 41806
rect 522487 41713 522543 42193
rect 523775 41713 523831 42193
rect 524236 41890 524288 41954
rect 524248 41834 524276 41890
rect 524327 41834 524383 42193
rect 524248 41806 524383 41834
rect 524327 41713 524383 41806
rect 525524 41890 525576 41954
rect 525536 41834 525564 41890
rect 525615 41834 525671 42193
rect 525536 41806 525671 41834
rect 525615 41713 525671 41806
rect 526811 41834 526867 42193
rect 526732 41818 526867 41834
rect 526720 41806 526867 41818
rect 526720 41754 526772 41806
rect 526811 41713 526867 41806
rect 527916 41890 527968 41954
rect 527928 41834 527956 41890
rect 528007 41834 528063 42193
rect 528651 41834 528707 42193
rect 527928 41806 528707 41834
rect 528007 41713 528063 41806
rect 528651 41713 528707 41806
rect 529847 41713 529903 42193
rect 579908 41886 579936 42706
rect 568856 41822 568908 41886
rect 579896 41822 579948 41886
rect 295017 41657 295227 41713
rect 295395 41657 295871 41713
rect 296039 41657 296515 41713
rect 296683 41657 297067 41713
rect 297235 41657 297711 41713
rect 297879 41657 298355 41713
rect 298523 41657 298907 41713
rect 299075 41657 299551 41713
rect 299719 41657 300195 41713
rect 300363 41657 300747 41713
rect 300915 41657 301391 41713
rect 301559 41657 302035 41713
rect 302203 41657 302587 41713
rect 302755 41657 303231 41713
rect 303399 41657 303875 41713
rect 304043 41657 304519 41713
rect 304687 41657 305071 41713
rect 305239 41657 305715 41713
rect 305883 41657 306359 41713
rect 306527 41657 306911 41713
rect 307079 41657 307555 41713
rect 307723 41657 308199 41713
rect 308367 41657 308751 41713
rect 308919 41657 309395 41713
rect 309563 41657 310039 41713
rect 310207 41657 310591 41713
rect 310759 41657 310958 41713
rect 256238 39471 256294 39545
rect 238972 30753 256100 31683
rect 241200 714 256100 30753
rect 295017 0 310958 41657
rect 349817 41657 350027 41713
rect 350195 41657 350671 41713
rect 350839 41657 351315 41713
rect 351483 41657 351867 41713
rect 352035 41657 352511 41713
rect 352679 41657 353155 41713
rect 353323 41657 353707 41713
rect 353875 41657 354351 41713
rect 354519 41657 354995 41713
rect 355163 41657 355547 41713
rect 355715 41657 356191 41713
rect 356359 41657 356835 41713
rect 357003 41657 357387 41713
rect 357555 41657 358031 41713
rect 358199 41657 358675 41713
rect 358843 41657 359319 41713
rect 359487 41657 359871 41713
rect 360039 41657 360515 41713
rect 360683 41657 361159 41713
rect 361327 41657 361711 41713
rect 361879 41657 362355 41713
rect 362523 41657 362999 41713
rect 363167 41657 363551 41713
rect 363719 41657 364195 41713
rect 364363 41657 364839 41713
rect 365007 41657 365391 41713
rect 365559 41657 365758 41713
rect 349817 0 365758 41657
rect 404617 41657 404827 41713
rect 404995 41657 405471 41713
rect 405639 41657 406115 41713
rect 406283 41657 406667 41713
rect 406835 41657 407311 41713
rect 407479 41657 407955 41713
rect 408123 41657 408507 41713
rect 408675 41657 409151 41713
rect 409319 41657 409795 41713
rect 409963 41657 410347 41713
rect 410515 41657 410991 41713
rect 411159 41657 411635 41713
rect 411803 41657 412187 41713
rect 412355 41657 412831 41713
rect 412999 41657 413475 41713
rect 413643 41657 414119 41713
rect 414287 41657 414671 41713
rect 414839 41657 415315 41713
rect 415483 41657 415959 41713
rect 416127 41657 416511 41713
rect 416679 41657 417155 41713
rect 417323 41657 417799 41713
rect 417967 41657 418351 41713
rect 418519 41657 418995 41713
rect 419163 41657 419639 41713
rect 419807 41657 420191 41713
rect 420359 41657 420558 41713
rect 404617 0 420558 41657
rect 459417 41657 459627 41713
rect 459795 41657 460271 41713
rect 460439 41657 460915 41713
rect 461083 41657 461467 41713
rect 461635 41657 462111 41713
rect 462279 41657 462755 41713
rect 462923 41657 463307 41713
rect 463475 41657 463951 41713
rect 464119 41657 464595 41713
rect 464763 41657 465147 41713
rect 465315 41657 465791 41713
rect 465959 41657 466435 41713
rect 466603 41657 466987 41713
rect 467155 41657 467631 41713
rect 467799 41657 468275 41713
rect 468443 41657 468919 41713
rect 469087 41657 469471 41713
rect 469639 41657 470115 41713
rect 470283 41657 470759 41713
rect 470927 41657 471311 41713
rect 471479 41657 471955 41713
rect 472123 41657 472599 41713
rect 472767 41657 473151 41713
rect 473319 41657 473795 41713
rect 473963 41657 474439 41713
rect 474607 41657 474991 41713
rect 475159 41657 475358 41713
rect 459417 0 475358 41657
rect 514217 41657 514427 41713
rect 514595 41657 515071 41713
rect 515239 41657 515715 41713
rect 515883 41657 516267 41713
rect 516435 41657 516911 41713
rect 517079 41657 517555 41713
rect 517723 41657 518107 41713
rect 518275 41657 518751 41713
rect 518919 41657 519395 41713
rect 519563 41657 519947 41713
rect 520115 41657 520591 41713
rect 520759 41657 521235 41713
rect 521403 41657 521787 41713
rect 521955 41657 522431 41713
rect 522599 41657 523075 41713
rect 523243 41657 523719 41713
rect 523887 41657 524271 41713
rect 524439 41657 524915 41713
rect 525083 41657 525559 41713
rect 525727 41657 526111 41713
rect 526279 41657 526755 41713
rect 526923 41657 527399 41713
rect 527567 41657 527951 41713
rect 528119 41657 528595 41713
rect 528763 41657 529239 41713
rect 529407 41657 529791 41713
rect 529959 41657 530158 41713
rect 514217 0 530158 41657
rect 568868 39681 568896 41822
rect 568854 39607 568910 39681
rect 569142 39593 573922 40000
rect 578421 39616 578821 40000
rect 579121 39593 583901 40000
rect 622942 39593 627722 40000
rect 632221 39616 632621 40000
rect 632921 39593 637701 40000
rect 569142 985 583947 39593
rect 622942 985 637747 39593
<< metal3 >>
rect 81144 997600 86144 1014070
rect 132544 997600 137544 1014070
rect 183944 997600 188944 1014070
rect 240478 997600 254800 1000737
rect 292078 997600 306400 1000737
rect 388744 997600 393744 1014070
rect 477744 997600 482744 1014070
rect 529144 997600 534144 1014070
rect 630944 997600 635944 1014070
rect 23530 959144 40000 964144
rect 677600 943200 680737 957522
rect 678000 469900 685920 474700
rect 31680 440900 39600 445700
rect 42333 47018 42399 47021
rect 42333 47016 44834 47018
rect 42333 46960 42338 47016
rect 42394 46960 44834 47016
rect 42333 46958 44834 46960
rect 42333 46955 42399 46958
rect 44774 46882 44834 46958
rect 52453 46882 52519 46885
rect 44774 46880 52519 46882
rect 44774 46824 52458 46880
rect 52514 46824 52519 46880
rect 44774 46822 52519 46824
rect 52453 46819 52519 46822
rect 411069 44434 411135 44437
rect 419717 44434 419783 44437
rect 411069 44432 419783 44434
rect 411069 44376 411074 44432
rect 411130 44376 419722 44432
rect 419778 44376 419783 44432
rect 411069 44374 419783 44376
rect 411069 44371 411135 44374
rect 419717 44371 419783 44374
rect 465809 44434 465875 44437
rect 474457 44434 474523 44437
rect 465809 44432 474523 44434
rect 465809 44376 465814 44432
rect 465870 44376 474462 44432
rect 474518 44376 474523 44432
rect 465809 44374 474523 44376
rect 465809 44371 465875 44374
rect 474457 44371 474523 44374
rect 518801 44298 518867 44301
rect 524965 44298 525031 44301
rect 518801 44296 525031 44298
rect 518801 44240 518806 44296
rect 518862 44240 524970 44296
rect 525026 44240 525031 44296
rect 518801 44238 525031 44240
rect 518801 44235 518867 44238
rect 524965 44235 525031 44238
rect 141667 38031 141813 40000
rect 141667 37971 141873 38031
rect 141667 37911 141820 37971
rect 141873 37911 141966 37971
rect 141667 37818 141966 37911
rect 141820 37046 141966 37818
<< obsm3 >>
rect 76291 1014150 91050 1032263
rect 76291 1000581 81064 1014150
rect 86224 1000581 91050 1014150
rect 127691 1014150 142450 1032263
rect 127691 1000581 132464 1014150
rect 137624 1000581 142450 1014150
rect 179091 1014150 193850 1032263
rect 179091 1000581 183864 1014150
rect 189024 1000581 193850 1014150
rect 221000 1000817 254800 1037600
rect 272600 1000817 306400 1037600
rect 333448 1002850 348258 1037600
rect 383891 1014150 398650 1032263
rect 221000 997600 235279 1000737
rect 235359 999946 240398 1000817
rect 235359 998225 237898 999946
rect 235359 998145 235499 998225
rect 237859 998145 237898 998225
rect 235579 997600 237779 998145
rect 237978 997600 240178 999866
rect 240258 998145 240398 999946
rect 272600 997600 286879 1000737
rect 286959 999946 291998 1000817
rect 286959 998225 289498 999946
rect 286959 998145 287099 998225
rect 289459 998145 289498 998225
rect 287179 997600 289379 998145
rect 289578 997600 291778 999866
rect 291858 998145 291998 999946
rect 333499 997600 338279 1002770
rect 338359 998007 343398 1002850
rect 338579 997600 340779 998007
rect 340978 997600 343178 998007
rect 343478 997600 348258 1002770
rect 383891 1000581 388664 1014150
rect 393824 1000581 398650 1014150
rect 472891 1014150 487650 1032263
rect 472891 1000581 477664 1014150
rect 482824 1000581 487650 1014150
rect 524291 1014150 539050 1032263
rect 524291 1000581 529064 1014150
rect 534224 1000581 539050 1014150
rect 575648 1005032 590458 1036620
rect 626091 1014150 640850 1032263
rect 575648 1004183 585598 1005032
rect 575699 997600 580479 1004103
rect 580559 998007 585598 1004183
rect 580779 997600 582979 998007
rect 583178 997600 585378 998007
rect 585678 997600 590458 1004952
rect 626091 1000581 630864 1014150
rect 636024 1000581 640850 1014150
rect 343590 997117 343650 997600
rect 585041 997522 585107 997525
rect 585734 997522 585794 997600
rect 585041 997462 585794 997522
rect 585041 997459 585107 997462
rect 343590 997054 343699 997117
rect 343633 997051 343699 997054
rect 5337 964224 37019 969050
rect 5337 959064 23450 964224
rect 677600 962721 680737 977000
rect 680817 962641 717600 977000
rect 678145 962501 717600 962641
rect 677600 960221 678145 962421
rect 678225 960141 717600 962501
rect 678145 960102 717600 960141
rect 5337 954291 37019 959064
rect 677600 957822 679866 960022
rect 679946 957742 717600 960102
rect 678145 957602 717600 957742
rect 680817 943200 717600 957602
rect 7 927240 4850 929187
rect 30753 927121 31683 929228
rect 33910 927240 34840 929187
rect 7 922071 38140 927000
rect 38220 922151 39600 926940
rect 685910 922779 686840 924795
rect 678007 922580 717593 922600
rect 7 921851 39593 922071
rect 7 919676 39600 921851
rect 7 919376 39593 919676
rect 7 917200 39600 919376
rect 678000 917700 679380 922500
rect 679460 917620 717593 922580
rect 678007 917400 717593 917620
rect 7 916980 39593 917200
rect 7 912020 38140 916980
rect 38220 912100 39600 916900
rect 678000 915224 717593 917400
rect 678007 914924 717593 915224
rect 678000 912749 717593 914924
rect 678007 912529 717593 912749
rect 7 912000 39593 912020
rect 30760 909805 31690 911821
rect 678000 907660 679380 912449
rect 679460 907600 717593 912529
rect 682760 905413 683690 907360
rect 685917 905372 686847 907479
rect 712750 905413 717593 907360
rect 0 879798 35960 884658
rect 36040 879878 40000 884658
rect 0 879578 39593 879798
rect 0 877378 40000 879578
rect 0 877179 39593 877378
rect 0 874979 40000 877179
rect 0 874759 39593 874979
rect 0 869848 35960 874759
rect 36040 870090 40000 874679
rect 42333 870090 42399 870093
rect 44817 870090 44883 870093
rect 36040 870030 44883 870090
rect 36040 869899 40000 870030
rect 42333 870027 42399 870030
rect 44817 870027 44883 870030
rect 677338 862486 717600 878338
rect 980 837598 32568 842458
rect 32648 837678 40000 842458
rect 980 837378 39593 837598
rect 980 835178 40000 837378
rect 980 834979 39593 835178
rect 980 832779 40000 834979
rect 980 832559 39593 832779
rect 980 827648 33417 832559
rect 33497 827699 40000 832479
rect 677600 828521 680592 833301
rect 680672 828441 717600 833352
rect 678007 828221 717600 828441
rect 677600 826021 717600 828221
rect 678007 825822 717600 826021
rect 677600 823622 717600 825822
rect 678007 823402 717600 823622
rect 677600 818542 680592 823322
rect 680672 818542 717600 823402
rect 677593 818410 677659 818413
rect 677734 818410 677794 818542
rect 677593 818350 677794 818410
rect 677593 818347 677659 818350
rect 0 784462 40262 800314
rect 677338 773286 717600 789138
rect 0 741262 40262 757114
rect 677338 728286 717600 744138
rect 0 698062 40262 713914
rect 677338 683286 717600 699138
rect 0 654862 40262 670714
rect 677338 638086 717600 653938
rect 0 611662 40262 627514
rect 677338 593086 717600 608938
rect 0 568462 40262 584314
rect 677338 547886 717600 563738
rect 0 525262 40262 541114
rect 677600 513921 680592 518701
rect 677734 513773 677794 513921
rect 680672 513841 717600 518752
rect 677685 513710 677794 513773
rect 677685 513707 677751 513710
rect 678007 513621 717600 513841
rect 677600 511421 717600 513621
rect 678007 511222 717600 511421
rect 677600 509022 717600 511222
rect 678007 508802 717600 509022
rect 677600 503942 680592 508722
rect 680672 503942 717600 508802
rect 0 492998 36928 497858
rect 37008 493078 40000 497858
rect 0 492778 39593 492998
rect 0 490578 40000 492778
rect 0 490379 39593 490578
rect 0 488179 40000 490379
rect 0 487959 39593 488179
rect 0 483048 36928 487959
rect 37008 483099 40000 487879
rect 685910 474979 686840 476995
rect 678007 474780 717593 474800
rect 686000 469820 717593 474780
rect 678007 469600 717593 469820
rect 678000 467424 717593 469600
rect 678007 467124 717593 467424
rect 678000 464949 717593 467124
rect 678007 464729 717593 464949
rect 678000 459860 685920 464649
rect 686000 459800 717593 464729
rect 7 456040 4850 457987
rect 30753 455921 31683 458028
rect 33910 456040 34840 457987
rect 682760 457613 683690 459560
rect 685917 457572 686847 459679
rect 712750 457613 717593 459560
rect 7 450871 31600 455800
rect 31680 450951 39600 455740
rect 7 450651 39593 450871
rect 7 448476 39600 450651
rect 7 448176 39593 448476
rect 7 446000 39600 448176
rect 7 445780 39593 446000
rect 7 440820 31600 445780
rect 7 440800 39593 440820
rect 30760 438605 31690 440621
rect 677600 425721 684103 430501
rect 677501 425642 677567 425645
rect 677734 425642 677794 425721
rect 677501 425582 677794 425642
rect 684183 425641 716620 430552
rect 677501 425579 677567 425582
rect 678007 425421 716620 425641
rect 677600 423221 716620 425421
rect 678007 423022 716620 423221
rect 677600 420822 716620 423022
rect 678007 420602 716620 420822
rect 677600 415742 684952 420522
rect 685032 415742 716620 420602
rect 0 397662 40262 413514
rect 677338 370686 717600 386538
rect 0 354462 40262 370314
rect 0 311262 40262 327114
rect 677338 325486 717600 341338
rect 0 268062 40262 283914
rect 677338 280486 717600 296338
rect 0 224862 40262 240714
rect 677338 235486 717600 251338
rect 0 181662 40262 197514
rect 677338 190286 717600 206138
rect 677338 145286 717600 161138
rect 0 120198 35960 125058
rect 36040 120278 40000 125058
rect 0 119978 39593 120198
rect 0 117778 40000 119978
rect 0 117579 39593 117778
rect 0 115379 40000 117579
rect 0 115159 39593 115379
rect 0 110248 35960 115159
rect 36040 110530 40000 115079
rect 44173 110530 44239 110533
rect 44817 110530 44883 110533
rect 36040 110470 44883 110530
rect 36040 110299 40000 110470
rect 44173 110467 44239 110470
rect 44817 110467 44883 110470
rect 677338 100086 717600 115938
rect 30753 83121 31683 85228
rect 31961 83088 32654 85228
rect 879 78071 38140 83000
rect 38220 78151 39600 82940
rect 879 77851 39593 78071
rect 879 75676 39600 77851
rect 879 75376 39593 75676
rect 879 73200 39600 75376
rect 879 72980 39593 73200
rect 879 68098 38140 72980
rect 38220 71906 39600 72900
rect 44173 71906 44239 71909
rect 44817 71906 44883 71909
rect 38220 71846 44883 71906
rect 38220 68100 39600 71846
rect 44173 71843 44239 71846
rect 44817 71843 44883 71846
rect 522481 44434 522547 44437
rect 516090 44374 522547 44434
rect 404905 44298 404971 44301
rect 412909 44298 412975 44301
rect 404905 44238 412975 44298
rect 404905 44235 404971 44238
rect 412909 44235 412975 44238
rect 459645 44298 459711 44301
rect 467649 44298 467715 44301
rect 459645 44238 467715 44298
rect 459645 44235 459711 44238
rect 467649 44235 467715 44238
rect 514477 44298 514543 44301
rect 516090 44298 516150 44374
rect 522481 44371 522547 44374
rect 514477 44238 516150 44298
rect 514477 44235 514543 44238
rect 149053 40354 149119 40357
rect 145838 40294 149119 40354
rect 93761 40218 93827 40221
rect 135161 40218 135227 40221
rect 91142 40158 93827 40218
rect 91142 40000 91202 40158
rect 93761 40155 93827 40158
rect 133094 40158 135227 40218
rect 133094 40000 133154 40158
rect 135161 40155 135227 40158
rect 143073 40218 143139 40221
rect 143533 40218 143599 40221
rect 143073 40158 143458 40218
rect 143073 40155 143139 40158
rect 143398 40000 143458 40158
rect 143533 40158 144010 40218
rect 143533 40155 143599 40158
rect 143950 40000 144010 40158
rect 145838 40014 145898 40294
rect 149053 40291 149119 40294
rect 145820 40000 145898 40014
rect 47600 32953 51202 36017
rect 51600 32953 55202 36017
rect 55600 32953 59202 36017
rect 59600 32953 63202 36017
rect 63600 32953 67202 36017
rect 67600 32953 71202 36017
rect 78942 32648 83722 40000
rect 84022 39593 86222 40000
rect 86421 39593 88621 40000
rect 83802 33417 88841 39593
rect 88921 33497 93701 40000
rect 83802 32568 93752 33417
rect 101400 32953 105002 36017
rect 105400 32953 109002 36017
rect 109400 32953 113002 36017
rect 113400 32953 117002 36017
rect 117400 32953 121002 36017
rect 121400 32953 125002 36017
rect 78942 980 93752 32568
rect 132660 30216 132868 39875
rect 132660 26680 132735 30216
rect 132948 30136 133162 40000
rect 132815 27080 133162 30136
rect 133242 37738 141587 39875
rect 141893 38746 143275 39875
rect 141893 38453 142982 38746
rect 143355 38666 143585 40000
rect 141893 38397 142926 38453
rect 141893 38111 142710 38397
rect 143062 38390 143585 38666
rect 143062 38373 143375 38390
rect 143388 38373 143585 38390
rect 143665 39293 143738 39875
rect 143818 39373 144151 40000
rect 144231 39293 145736 39875
rect 143006 38360 143062 38373
rect 143079 38360 143388 38373
rect 143006 38330 143388 38360
rect 143006 38317 143315 38330
rect 143332 38317 143388 38330
rect 141953 38051 142710 38111
rect 133242 36966 141740 37738
rect 142046 37467 142710 38051
rect 142790 38300 143006 38317
rect 143019 38300 143332 38317
rect 142790 38004 143332 38300
rect 143665 38293 145736 39293
rect 143468 38237 145736 38293
rect 142790 37547 143019 38004
rect 143412 37924 145736 38237
rect 143099 37467 145736 37924
rect 142046 36966 145736 37467
rect 133242 36603 145736 36966
rect 145816 36843 145920 40000
rect 146000 36923 147407 39875
rect 146042 36881 147407 36923
rect 145816 36801 145962 36843
rect 145816 36711 146052 36801
rect 146132 36791 147407 36881
rect 145816 36683 145934 36711
rect 145936 36683 146142 36711
rect 146222 36701 147407 36791
rect 145934 36621 146142 36683
rect 133242 36511 145854 36603
rect 145934 36591 146245 36621
rect 133242 36396 145946 36511
rect 146026 36476 146245 36591
rect 133242 33821 146061 36396
rect 133242 33704 145944 33821
rect 146141 33741 146245 36476
rect 133242 33561 145801 33704
rect 146024 33639 146245 33741
rect 146024 33624 146155 33639
rect 146170 33624 146245 33639
rect 145881 33609 146024 33624
rect 146027 33609 146170 33624
rect 133242 33444 145684 33561
rect 145881 33489 146170 33609
rect 146325 33544 147407 36701
rect 145881 33481 146024 33489
rect 146027 33481 146170 33489
rect 145764 33459 145881 33481
rect 145889 33459 146027 33481
rect 133242 33401 145641 33444
rect 133242 33095 143065 33401
rect 145764 33369 146027 33459
rect 146250 33401 147407 33544
rect 145764 33364 145885 33369
rect 145910 33364 146027 33369
rect 145721 33339 145764 33364
rect 145769 33339 145910 33364
rect 145721 33321 145910 33339
rect 143145 33261 145910 33321
rect 146107 33284 147407 33401
rect 143145 33260 145777 33261
rect 145806 33260 145910 33261
rect 143145 33175 145806 33260
rect 145990 33180 147407 33284
rect 145886 33095 147407 33180
rect 133242 27160 147407 33095
rect 155200 32953 158802 36017
rect 159200 32953 162802 36017
rect 163200 32953 166802 36017
rect 167200 32953 170802 36017
rect 171200 32953 174802 36017
rect 175200 32953 178802 36017
rect 132815 26760 133482 27080
rect 133562 26840 147407 27160
rect 132660 26360 133082 26680
rect 133162 26480 133762 26760
rect 133842 26560 147407 26840
rect 133162 26450 133949 26480
rect 133162 26440 133482 26450
rect 133502 26440 133949 26450
rect 132660 26103 133402 26360
rect 133482 26293 133949 26440
rect 134029 26373 147407 26560
rect 133482 26270 133942 26293
rect 133949 26270 134122 26293
rect 133482 26210 134122 26270
rect 133482 26183 133739 26210
rect 133742 26183 134122 26210
rect 134202 26200 147407 26373
rect 133739 26120 134122 26183
rect 132660 25913 133659 26103
rect 133739 26000 134392 26120
rect 133739 25993 133929 26000
rect 133952 25993 134392 26000
rect 132660 25720 133849 25913
rect 133929 25850 134392 25993
rect 134472 25930 147407 26200
rect 133929 25820 134628 25850
rect 133929 25800 134122 25820
rect 134132 25800 134628 25820
rect 132660 25478 134042 25720
rect 134122 25584 134628 25800
rect 134122 25558 134364 25584
rect 134368 25558 134628 25584
rect 134364 25520 134628 25558
rect 132660 25440 134284 25478
rect 132660 20991 134322 25440
rect 134402 21071 134628 25520
rect 134708 20991 147407 25930
rect 132660 0 147407 20991
rect 186486 0 202338 40262
rect 210000 32953 213602 36017
rect 214000 32953 217602 36017
rect 218000 32953 221602 36017
rect 222000 32953 225602 36017
rect 226000 32953 229602 36017
rect 230000 32953 233602 36017
rect 238972 31961 241112 32654
rect 238972 30753 241079 31683
rect 241260 31680 246049 39600
rect 246349 39593 248524 39600
rect 248824 39593 251000 39600
rect 246129 31600 251220 39593
rect 251300 39538 256100 39600
rect 256233 39538 256299 39541
rect 251300 39478 256299 39538
rect 251300 31680 256100 39478
rect 256233 39475 256299 39478
rect 263800 32953 267402 36017
rect 267800 32953 271402 36017
rect 271800 32953 275402 36017
rect 275800 32953 279402 36017
rect 279800 32953 283402 36017
rect 283800 32953 287402 36017
rect 241200 879 256100 31600
rect 295086 0 310938 40262
rect 318600 32953 322202 36017
rect 322600 32953 326202 36017
rect 326600 32953 330202 36017
rect 330600 32953 334202 36017
rect 334600 32953 338202 36017
rect 338600 32953 342202 36017
rect 349886 0 365738 40262
rect 373400 32953 377002 36017
rect 377400 32953 381002 36017
rect 381400 32953 385002 36017
rect 385400 32953 389002 36017
rect 389400 32953 393002 36017
rect 393400 32953 397002 36017
rect 404686 0 420538 40262
rect 428200 32953 431802 36017
rect 432200 32953 435802 36017
rect 436200 32953 439802 36017
rect 440200 32953 443802 36017
rect 444200 32953 447802 36017
rect 448200 32953 451802 36017
rect 459486 0 475338 40262
rect 483000 32953 486602 36017
rect 487000 32953 490602 36017
rect 491000 32953 494602 36017
rect 495000 32953 498602 36017
rect 499000 32953 502602 36017
rect 503000 32953 506602 36017
rect 514286 0 530138 40262
rect 568849 39674 568915 39677
rect 569142 39674 573922 40000
rect 568849 39614 573922 39674
rect 568849 39611 568915 39614
rect 537800 32953 541402 36017
rect 541800 32953 545402 36017
rect 545800 32953 549402 36017
rect 549800 32953 553402 36017
rect 553800 32953 557402 36017
rect 557800 32953 561402 36017
rect 569142 34830 573922 39614
rect 574222 39593 576422 40000
rect 576621 39593 578821 40000
rect 574002 34750 579041 39593
rect 579121 34830 583901 40000
rect 622942 37008 627722 40000
rect 628022 39593 630222 40000
rect 630421 39593 632621 40000
rect 627802 36928 632841 39593
rect 632921 37008 637701 40000
rect 569142 0 583952 34750
rect 591600 32953 595202 36017
rect 595600 32953 599202 36017
rect 599600 32953 603202 36017
rect 603600 32953 607202 36017
rect 607600 32953 611202 36017
rect 611600 32953 615202 36017
rect 622942 0 637752 36928
rect 645400 32953 649002 36017
rect 649400 32953 653002 36017
rect 653400 32953 657002 36017
rect 657400 32953 661002 36017
rect 661400 32953 665002 36017
rect 665400 32953 669002 36017
<< metal4 >>
rect 7 455800 4843 456093
rect 0 455546 4843 455800
rect 28653 407018 28719 525722
rect 32933 455546 33623 483254
rect 36323 455607 37013 483193
rect 37293 455546 38223 483254
rect 38503 455546 39593 483254
rect 679377 430346 680307 460054
rect 680587 430407 681277 459993
rect 688881 430346 688947 554382
rect 93607 36323 132793 37013
rect 93546 31674 132854 31683
rect 93546 30762 132869 31674
rect 93546 30753 132854 30762
rect 93546 28653 192982 28719
<< obsm4 >>
rect 0 1032677 40466 1037600
rect 40546 1032757 76454 1037600
rect 0 1016680 40549 1032677
rect 40800 1016680 76200 1032757
rect 76534 1032677 90866 1037600
rect 90946 1032757 127854 1037600
rect 76393 1016680 91007 1032677
rect 91200 1016680 127600 1032757
rect 127934 1032677 142266 1037600
rect 142346 1032757 179254 1037600
rect 127793 1016680 142407 1032677
rect 142600 1016680 179000 1032757
rect 179334 1032677 193666 1037600
rect 193746 1032757 230641 1037600
rect 179193 1016680 193807 1032677
rect 194000 1016680 221000 1032757
rect 230721 1032677 246097 1037600
rect 246177 1032757 282241 1037600
rect 230448 1016680 246177 1032677
rect 254800 1016680 272600 1032757
rect 282321 1032677 297697 1037600
rect 297777 1032757 333654 1037600
rect 282048 1016680 297777 1032677
rect 306400 1016680 333400 1032757
rect 333734 1032677 348066 1037600
rect 348146 1032757 384054 1037600
rect 333593 1016680 348207 1032677
rect 348400 1016680 381800 1032757
rect 382800 1016680 383800 1032757
rect 384134 1032677 398466 1037600
rect 398546 1032757 473054 1037600
rect 383993 1016680 398607 1032677
rect 398800 1016680 472800 1032757
rect 473134 1032677 487466 1037600
rect 487546 1032757 524454 1037600
rect 472993 1016680 487607 1032677
rect 487800 1016680 524200 1032757
rect 524534 1032677 538866 1037600
rect 538946 1032757 575854 1037600
rect 524393 1016680 539007 1032677
rect 539200 1016680 575600 1032757
rect 575934 1032677 590266 1037600
rect 590346 1032757 626254 1037600
rect 575793 1016680 590407 1032677
rect 590600 1016680 626000 1032757
rect 626334 1032677 640666 1037600
rect 640746 1032757 677887 1037600
rect 641000 1032677 677600 1032757
rect 677967 1032677 717600 1037600
rect 626193 1016680 640807 1032677
rect 641000 1016680 717600 1032677
rect 0 1011527 40349 1016680
rect 40429 1011607 76454 1016600
rect 76534 1011527 90866 1016680
rect 90946 1011607 127854 1016600
rect 127934 1011527 142266 1016680
rect 142346 1011607 179254 1016600
rect 179334 1011527 193666 1016680
rect 193746 1011607 230543 1016600
rect 230623 1011527 246097 1016680
rect 246177 1011607 282143 1016600
rect 282223 1011527 297697 1016680
rect 297777 1011607 333654 1016600
rect 333734 1011527 348066 1016680
rect 348146 1011607 384054 1016600
rect 384134 1011527 398466 1016680
rect 398546 1011607 473054 1016600
rect 473134 1011527 487466 1016680
rect 487546 1011607 524454 1016600
rect 524534 1011527 538866 1016680
rect 538946 1011607 575854 1016600
rect 575934 1011527 590266 1016680
rect 590346 1011607 626254 1016600
rect 626334 1011527 640666 1016680
rect 640746 1011607 678129 1016600
rect 678209 1011527 717600 1016680
rect 0 1011387 40549 1011527
rect 40800 1011387 76200 1011527
rect 76393 1011387 91007 1011527
rect 91200 1011387 127600 1011527
rect 127793 1011387 142407 1011527
rect 142600 1011387 179000 1011527
rect 179193 1011387 193807 1011527
rect 194000 1011387 221000 1011527
rect 230448 1011387 246177 1011527
rect 254800 1011387 272600 1011527
rect 282048 1011387 297777 1011527
rect 306400 1011387 333400 1011527
rect 333593 1011387 348207 1011527
rect 348400 1011387 381800 1011527
rect 382800 1011387 383800 1011527
rect 383993 1011387 398607 1011527
rect 398800 1011387 472800 1011527
rect 472993 1011387 487607 1011527
rect 487800 1011387 524200 1011527
rect 524393 1011387 539007 1011527
rect 539200 1011387 575600 1011527
rect 575793 1011387 590407 1011527
rect 590600 1011387 626000 1011527
rect 626193 1011387 640807 1011527
rect 641000 1011387 717600 1011527
rect 0 1010337 40466 1011387
rect 40546 1010417 76454 1011307
rect 76534 1010337 90866 1011387
rect 90946 1010417 127854 1011307
rect 127934 1010337 142266 1011387
rect 142346 1010417 179254 1011307
rect 179334 1010337 193666 1011387
rect 193746 1010417 230543 1011307
rect 230623 1010337 246097 1011387
rect 246177 1010417 282143 1011307
rect 282223 1010337 297697 1011387
rect 297777 1010417 333654 1011307
rect 333734 1010337 348066 1011387
rect 348146 1010417 384054 1011307
rect 384134 1010337 398466 1011387
rect 398546 1010417 473054 1011307
rect 473134 1010337 487466 1011387
rect 487546 1010417 524454 1011307
rect 524534 1010337 538866 1011387
rect 538946 1010417 575854 1011307
rect 575934 1010337 590266 1011387
rect 590346 1010417 626254 1011307
rect 626334 1010337 640666 1011387
rect 640746 1010417 677896 1011307
rect 677976 1010337 717600 1011387
rect 0 1010217 40549 1010337
rect 40800 1010217 76200 1010337
rect 76393 1010217 91007 1010337
rect 91200 1010217 127600 1010337
rect 127793 1010217 142407 1010337
rect 142600 1010217 179000 1010337
rect 179193 1010217 193807 1010337
rect 194000 1010217 221000 1010337
rect 230448 1010217 246177 1010337
rect 254800 1010217 272600 1010337
rect 282048 1010217 297777 1010337
rect 306400 1010217 333400 1010337
rect 333593 1010217 348207 1010337
rect 348400 1010217 381800 1010337
rect 382800 1010217 383800 1010337
rect 383993 1010217 398607 1010337
rect 398800 1010217 472800 1010337
rect 472993 1010217 487607 1010337
rect 487800 1010217 524200 1010337
rect 524393 1010217 539007 1010337
rect 539200 1010217 575600 1010337
rect 575793 1010217 590407 1010337
rect 590600 1010217 626000 1010337
rect 626193 1010217 640807 1010337
rect 641000 1010217 717600 1010337
rect 0 1009167 40466 1010217
rect 40546 1009247 76454 1010137
rect 76534 1009167 90866 1010217
rect 90946 1009247 127854 1010137
rect 127934 1009167 142266 1010217
rect 142346 1009247 179254 1010137
rect 179334 1009167 193666 1010217
rect 193746 1009247 230543 1010137
rect 230623 1009167 246097 1010217
rect 246177 1009247 282143 1010137
rect 282223 1009167 297697 1010217
rect 297777 1009247 333654 1010137
rect 333734 1009167 348066 1010217
rect 348146 1009247 384054 1010137
rect 384134 1009167 398466 1010217
rect 398546 1009247 473054 1010137
rect 473134 1009167 487466 1010217
rect 487546 1009247 524454 1010137
rect 524534 1009167 538866 1010217
rect 538946 1009247 575854 1010137
rect 575934 1009167 590266 1010217
rect 590346 1009247 626254 1010137
rect 626334 1009167 640666 1010217
rect 640746 1009247 677925 1010137
rect 678005 1009167 717600 1010217
rect 0 1009027 40549 1009167
rect 40800 1009027 76200 1009167
rect 76393 1009027 91007 1009167
rect 91200 1009027 127600 1009167
rect 127793 1009027 142407 1009167
rect 142600 1009027 179000 1009167
rect 179193 1009027 193807 1009167
rect 194000 1009027 221000 1009167
rect 230448 1009027 246177 1009167
rect 254800 1009027 272600 1009167
rect 282048 1009027 297777 1009167
rect 306400 1009027 333400 1009167
rect 333593 1009027 348207 1009167
rect 348400 1009027 381800 1009167
rect 382800 1009027 383800 1009167
rect 383993 1009027 398607 1009167
rect 398800 1009027 472800 1009167
rect 472993 1009027 487607 1009167
rect 487800 1009027 524200 1009167
rect 524393 1009027 539007 1009167
rect 539200 1009027 575600 1009167
rect 575793 1009027 590407 1009167
rect 590600 1009027 626000 1009167
rect 626193 1009027 640807 1009167
rect 641000 1009027 717600 1009167
rect 0 1008801 35285 1009027
rect 35365 1008881 381800 1008947
rect 382800 1008881 575854 1008947
rect 575934 1008901 590266 1009027
rect 590346 1008881 682235 1008947
rect 0 1008145 35338 1008801
rect 35418 1008225 682182 1008821
rect 682315 1008801 717600 1009027
rect 0 1007849 36409 1008145
rect 36489 1007929 76454 1008165
rect 76534 1007949 90866 1008145
rect 90946 1007929 127854 1008165
rect 127934 1007949 142266 1008145
rect 142346 1007929 179254 1008165
rect 179334 1007949 193666 1008145
rect 193746 1007929 230448 1008165
rect 230528 1007949 246097 1008145
rect 246177 1007929 282048 1008165
rect 282128 1007949 297697 1008145
rect 297777 1007929 333654 1008165
rect 333734 1007949 348066 1008145
rect 348146 1007929 381800 1008165
rect 382800 1007929 384054 1008165
rect 384134 1007949 398466 1008145
rect 398546 1007929 473054 1008165
rect 473134 1007949 487466 1008145
rect 487546 1007929 524454 1008165
rect 524534 1007949 538866 1008145
rect 538946 1007929 575854 1008165
rect 575934 1007949 590266 1008145
rect 590346 1007929 626254 1008165
rect 626334 1007949 640666 1008145
rect 640746 1007929 681910 1008165
rect 682262 1008145 717600 1008801
rect 0 1007293 36545 1007849
rect 0 1007067 36005 1007293
rect 36625 1007273 681787 1007869
rect 681990 1007849 717600 1008145
rect 36085 1007147 381800 1007213
rect 382800 1007147 575854 1007213
rect 575934 1007067 590266 1007193
rect 590346 1007147 681515 1007213
rect 681867 1007193 717600 1007849
rect 681595 1007067 717600 1007193
rect 0 1006927 40549 1007067
rect 76393 1006927 91007 1007067
rect 127793 1006927 142407 1007067
rect 179193 1006927 193807 1007067
rect 230448 1006927 246177 1007067
rect 282048 1006927 297777 1007067
rect 333593 1006927 348207 1007067
rect 383993 1006927 398607 1007067
rect 472993 1006927 487607 1007067
rect 524393 1006927 539007 1007067
rect 575793 1006927 590407 1007067
rect 626193 1006927 640807 1007067
rect 677600 1006927 717600 1007067
rect 0 1005837 40466 1006927
rect 40546 1005917 76454 1006847
rect 76534 1005837 90866 1006927
rect 90946 1005917 127854 1006847
rect 127934 1005837 142266 1006927
rect 142346 1005917 179254 1006847
rect 179334 1005837 193666 1006927
rect 193746 1005917 230450 1006847
rect 230530 1005837 246097 1006927
rect 246177 1005917 282050 1006847
rect 282130 1005837 297697 1006927
rect 297777 1005917 333654 1006847
rect 333734 1005837 348066 1006927
rect 348146 1005917 382800 1006847
rect 383800 1005917 384054 1006847
rect 384134 1005837 398466 1006927
rect 398546 1005917 473054 1006847
rect 473134 1005837 487466 1006927
rect 487546 1005917 524454 1006847
rect 524534 1005837 538866 1006927
rect 538946 1005917 575854 1006847
rect 575934 1005837 590266 1006927
rect 590346 1005917 626254 1006847
rect 626334 1005837 640666 1006927
rect 640746 1005917 677895 1006847
rect 677975 1005837 717600 1006927
rect 0 1005717 40549 1005837
rect 76393 1005717 91007 1005837
rect 127793 1005717 142407 1005837
rect 179193 1005717 193807 1005837
rect 230448 1005717 246177 1005837
rect 282048 1005717 297777 1005837
rect 333593 1005717 348207 1005837
rect 383993 1005717 398607 1005837
rect 472993 1005717 487607 1005837
rect 524393 1005717 539007 1005837
rect 575793 1005717 590407 1005837
rect 626193 1005717 640807 1005837
rect 677600 1005717 717600 1005837
rect 0 1004867 40466 1005717
rect 40546 1004947 76454 1005637
rect 76534 1004867 90866 1005717
rect 90946 1004947 127854 1005637
rect 127934 1004867 142266 1005717
rect 142346 1004947 179254 1005637
rect 179334 1004867 193666 1005717
rect 193746 1004947 230543 1005637
rect 230623 1004867 246097 1005717
rect 246177 1004947 282143 1005637
rect 282223 1004867 297697 1005717
rect 297777 1004947 333654 1005637
rect 333734 1004867 348066 1005717
rect 348146 1004947 381800 1005637
rect 382800 1004947 384054 1005637
rect 384134 1004867 398466 1005717
rect 398546 1004947 473054 1005637
rect 473134 1004867 487466 1005717
rect 487546 1004947 524454 1005637
rect 524534 1004867 538866 1005717
rect 538946 1004947 575854 1005637
rect 575934 1004867 590266 1005717
rect 590346 1004947 626254 1005637
rect 626334 1004867 640666 1005717
rect 640746 1004947 677867 1005637
rect 677947 1004867 717600 1005717
rect 0 1004747 40549 1004867
rect 76393 1004747 91007 1004867
rect 127793 1004747 142407 1004867
rect 179193 1004747 193807 1004867
rect 230448 1004747 246177 1004867
rect 282048 1004747 297777 1004867
rect 333593 1004747 348207 1004867
rect 383993 1004747 398607 1004867
rect 472993 1004747 487607 1004867
rect 524393 1004747 539007 1004867
rect 575793 1004747 590407 1004867
rect 626193 1004747 640807 1004867
rect 677600 1004747 717600 1004867
rect 0 1003897 40466 1004747
rect 40546 1003977 76454 1004667
rect 76534 1003897 90866 1004747
rect 90946 1003977 127854 1004667
rect 127934 1003897 142266 1004747
rect 142346 1003977 179254 1004667
rect 179334 1003897 193666 1004747
rect 193746 1003977 230543 1004667
rect 230623 1003897 246097 1004747
rect 246177 1003977 282143 1004667
rect 282223 1003897 297697 1004747
rect 297777 1003977 333654 1004667
rect 333734 1003897 348066 1004747
rect 348146 1003977 384054 1004667
rect 384134 1003897 398466 1004747
rect 398546 1003977 473054 1004667
rect 473134 1003897 487466 1004747
rect 487546 1003977 524454 1004667
rect 524534 1003897 538866 1004747
rect 538946 1003977 575854 1004667
rect 575934 1003897 590266 1004747
rect 590346 1003977 626254 1004667
rect 626334 1003897 640666 1004747
rect 640746 1003977 677877 1004667
rect 677957 1003897 717600 1004747
rect 0 1003777 40549 1003897
rect 76393 1003777 91007 1003897
rect 127793 1003777 142407 1003897
rect 179193 1003777 193807 1003897
rect 230448 1003777 246177 1003897
rect 282048 1003777 297777 1003897
rect 333593 1003777 348207 1003897
rect 383993 1003777 398607 1003897
rect 472993 1003777 487607 1003897
rect 524393 1003777 539007 1003897
rect 575793 1003777 590407 1003897
rect 626193 1003777 640807 1003897
rect 677600 1003777 717600 1003897
rect 0 1002687 40466 1003777
rect 40546 1002767 76454 1003697
rect 76534 1002687 90866 1003777
rect 90946 1002767 127854 1003697
rect 127934 1002687 142266 1003777
rect 142346 1002767 179254 1003697
rect 179334 1002687 193666 1003777
rect 193746 1002767 230543 1003697
rect 230623 1002687 246097 1003777
rect 246177 1002767 282143 1003697
rect 282223 1002687 297697 1003777
rect 297777 1002767 333654 1003697
rect 333734 1002687 348066 1003777
rect 348146 1002767 384054 1003697
rect 384134 1002687 398466 1003777
rect 398546 1002767 473054 1003697
rect 473134 1002687 487466 1003777
rect 487546 1002767 524454 1003697
rect 524534 1002687 538866 1003777
rect 538946 1002767 575854 1003697
rect 575934 1002687 590266 1003777
rect 590346 1002767 626254 1003697
rect 626334 1002687 640666 1003777
rect 640746 1002767 677920 1003697
rect 678000 1002687 717600 1003777
rect 0 1002567 40549 1002687
rect 76393 1002567 91007 1002687
rect 127793 1002567 142407 1002687
rect 179193 1002567 193807 1002687
rect 230448 1002567 246177 1002687
rect 282048 1002567 297777 1002687
rect 333593 1002567 348207 1002687
rect 383993 1002567 398607 1002687
rect 472993 1002567 487607 1002687
rect 524393 1002567 539007 1002687
rect 575793 1002567 590407 1002687
rect 626193 1002567 640807 1002687
rect 677600 1002567 717600 1002687
rect 0 1002315 40466 1002567
rect 0 998209 28573 1002315
rect 28799 1002262 40466 1002315
rect 0 997967 20920 998209
rect 0 997600 4843 997887
rect 4923 997600 20920 997967
rect 0 969200 20920 997600
rect 0 968946 4843 969200
rect 4923 968866 20920 969007
rect 21000 968946 25993 998129
rect 26073 998005 28573 998209
rect 26073 997976 27383 998005
rect 26073 969200 26213 997976
rect 26073 968866 26213 969007
rect 26293 968946 27183 997896
rect 27263 969200 27383 997976
rect 27263 968866 27383 969007
rect 27463 968946 28353 997925
rect 28433 969200 28573 998005
rect 28433 968866 28573 969007
rect 0 954534 28573 968866
rect 0 954200 4843 954454
rect 4923 954393 20920 954534
rect 0 927000 20920 954200
rect 0 926957 4850 927000
rect 0 926746 4843 926957
rect 4923 926666 20920 927000
rect 21000 926746 25993 954454
rect 26073 954393 26213 954534
rect 26073 926666 26213 954200
rect 26293 926746 27183 954454
rect 27263 954393 27383 954534
rect 27263 926666 27383 954200
rect 27463 926746 28353 954454
rect 28433 954393 28573 954534
rect 28433 926666 28573 954200
rect 0 912334 28573 926666
rect 0 912000 4843 912254
rect 4923 912000 20920 912334
rect 0 884800 20920 912000
rect 0 884546 4843 884800
rect 4923 884466 20920 884607
rect 21000 884546 25993 912254
rect 26073 884800 26213 912334
rect 26073 884466 26213 884607
rect 26293 884546 27183 912254
rect 27263 884800 27383 912334
rect 27263 884466 27383 884607
rect 27463 884546 28353 912254
rect 28433 884800 28573 912334
rect 28433 884466 28573 884607
rect 0 870134 28573 884466
rect 0 869800 4843 870054
rect 4923 869993 20920 870134
rect 0 842600 20920 869800
rect 0 842346 4843 842600
rect 4923 842266 20920 842407
rect 21000 842346 25993 870054
rect 26073 869993 26213 870134
rect 26073 842600 26213 869800
rect 26073 842266 26213 842407
rect 26293 842346 27183 870054
rect 27263 869993 27383 870134
rect 27263 842600 27383 869800
rect 27263 842266 27383 842407
rect 27463 842346 28353 870054
rect 28433 869993 28573 870134
rect 28433 842600 28573 869800
rect 28433 842266 28573 842407
rect 28653 842346 28719 1002235
rect 0 827934 28699 842266
rect 0 827600 4843 827854
rect 4923 827793 20920 827934
rect 0 800400 20920 827600
rect 0 800146 4843 800400
rect 4923 800066 20920 800194
rect 21000 800146 25993 827854
rect 26073 827793 26213 827934
rect 26073 800400 26213 827600
rect 26073 800066 26213 800194
rect 26293 800146 27183 827854
rect 27263 827793 27383 827934
rect 27263 800400 27383 827600
rect 27263 800066 27383 800194
rect 27463 800146 28353 827854
rect 28433 827793 28573 827934
rect 28433 800400 28573 827600
rect 28433 800066 28573 800194
rect 0 793738 28573 800066
rect 28653 793818 28719 827854
rect 0 792072 28699 793738
rect 28779 792152 29375 1002182
rect 29455 1001990 40466 1002262
rect 29435 968946 29671 1001910
rect 29751 1001867 40466 1001990
rect 29455 954534 29651 968866
rect 29435 926746 29671 954454
rect 29455 912334 29651 926666
rect 29435 884546 29671 912254
rect 29455 870134 29651 884466
rect 29435 842346 29671 870054
rect 29455 827934 29651 842266
rect 29435 800146 29671 827854
rect 29455 795213 29651 800066
rect 29731 795293 30327 1001787
rect 30407 1001595 40466 1001867
rect 30387 842346 30453 1001515
rect 30533 1001477 40466 1001595
rect 40546 1001557 76454 1002487
rect 76534 1001477 90866 1002567
rect 90946 1001557 127854 1002487
rect 127934 1001477 142266 1002567
rect 142346 1001557 179254 1002487
rect 179334 1001477 193666 1002567
rect 193746 1001557 230543 1002487
rect 230623 1001477 245161 1002567
rect 245241 1001557 282143 1002487
rect 282223 1001477 296761 1002567
rect 296841 1001557 333654 1002487
rect 333734 1001477 348066 1002567
rect 348146 1001557 384054 1002487
rect 384134 1001477 398466 1002567
rect 398546 1001557 473054 1002487
rect 473134 1001477 487466 1002567
rect 487546 1001557 524454 1002487
rect 524534 1001477 538866 1002567
rect 538946 1001557 575854 1002487
rect 575934 1001477 590266 1002567
rect 590346 1001557 626254 1002487
rect 626334 1001477 640666 1002567
rect 640746 1001557 677905 1002487
rect 677985 1002315 717600 1002567
rect 677985 1002262 688801 1002315
rect 677985 1001595 688145 1002262
rect 677985 1001477 687067 1001595
rect 30533 1001357 40549 1001477
rect 76393 1001357 91007 1001477
rect 127793 1001357 142407 1001477
rect 179193 1001357 193807 1001477
rect 230448 1001357 246177 1001477
rect 282048 1001357 297777 1001477
rect 333593 1001357 348207 1001477
rect 383993 1001357 398607 1001477
rect 472993 1001357 487607 1001477
rect 524393 1001357 539007 1001477
rect 575793 1001357 590407 1001477
rect 626193 1001357 640807 1001477
rect 677600 1001357 687067 1001477
rect 30533 1000507 40469 1001357
rect 40549 1000587 76393 1001277
rect 76473 1000507 90927 1001357
rect 91007 1000587 127793 1001277
rect 127873 1000507 142327 1001357
rect 142407 1000587 179193 1001277
rect 179273 1000507 193727 1001357
rect 193807 1000587 230543 1001277
rect 230623 1000507 245161 1001357
rect 245241 1000587 282143 1001277
rect 282223 1000507 296761 1001357
rect 296841 1000587 333593 1001277
rect 333673 1000507 348127 1001357
rect 348207 1000587 381800 1001277
rect 382800 1000587 383993 1001277
rect 384073 1000507 398527 1001357
rect 398607 1000587 472993 1001277
rect 473073 1000507 487527 1001357
rect 487607 1000587 524393 1001277
rect 524473 1000507 538927 1001357
rect 539007 1000587 575793 1001277
rect 575873 1000507 590327 1001357
rect 590407 1000587 626193 1001277
rect 626273 1000507 640727 1001357
rect 640807 1000587 677894 1001277
rect 677974 1000507 687067 1001357
rect 30533 1000387 40549 1000507
rect 76393 1000387 91007 1000507
rect 127793 1000387 142407 1000507
rect 179193 1000387 193807 1000507
rect 230448 1000387 246177 1000507
rect 282048 1000387 297777 1000507
rect 333593 1000387 348207 1000507
rect 383993 1000387 398607 1000507
rect 472993 1000387 487607 1000507
rect 524393 1000387 539007 1000507
rect 575793 1000387 590407 1000507
rect 626193 1000387 640807 1000507
rect 677600 1000387 687067 1000507
rect 30533 999297 40466 1000387
rect 40546 999377 76454 1000307
rect 76534 999297 90866 1000387
rect 90946 999377 127854 1000307
rect 127934 999297 142266 1000387
rect 142346 999377 179254 1000307
rect 179334 999297 193666 1000387
rect 193746 999377 230543 1000307
rect 230623 999297 246097 1000387
rect 246177 999377 282143 1000307
rect 282223 999297 297697 1000387
rect 297777 999377 333654 1000307
rect 333734 999297 348066 1000387
rect 348146 999377 382800 1000307
rect 383800 999377 384054 1000307
rect 384134 999297 398466 1000387
rect 398546 999377 473054 1000307
rect 473134 999297 487466 1000387
rect 487546 999377 524454 1000307
rect 524534 999297 538866 1000387
rect 538946 999377 575854 1000307
rect 575934 999297 590266 1000387
rect 590346 999377 626254 1000307
rect 626334 999297 640666 1000387
rect 640746 999377 678357 1000307
rect 678437 999297 687067 1000387
rect 30533 999177 40549 999297
rect 76393 999177 91007 999297
rect 127793 999177 142407 999297
rect 179193 999177 193807 999297
rect 230448 999177 246177 999297
rect 282048 999177 297777 999297
rect 333593 999177 348207 999297
rect 383993 999177 398607 999297
rect 472993 999177 487607 999297
rect 524393 999177 539007 999297
rect 575793 999177 590407 999297
rect 626193 999177 640807 999297
rect 677600 999177 687067 999297
rect 30533 998437 40466 999177
rect 30533 998000 37213 998437
rect 30533 997975 33823 998000
rect 30533 997600 30673 997975
rect 31763 997957 33823 997975
rect 31763 997947 32853 997957
rect 30533 968866 30673 969007
rect 30753 968946 31683 997895
rect 31763 997600 31883 997947
rect 31763 968866 31883 969007
rect 31963 968946 32653 997867
rect 32733 997600 32853 997947
rect 32733 968866 32853 969007
rect 32933 968946 33623 997877
rect 33703 997600 33823 997957
rect 34913 997985 37213 998000
rect 33703 968866 33823 969007
rect 33903 968946 34833 997920
rect 34913 997600 35033 997985
rect 36123 997974 37213 997985
rect 34913 968866 35033 969007
rect 35113 968946 36043 997905
rect 36123 997600 36243 997974
rect 36323 969007 37013 997894
rect 37093 997600 37213 997974
rect 36123 968927 36243 969007
rect 37093 968927 37213 969007
rect 37293 968946 38223 998357
rect 38303 998150 40466 998437
rect 38303 997600 38423 998150
rect 36123 968866 37213 968927
rect 38303 968866 38423 969007
rect 38503 968946 39593 998070
rect 39673 997927 40466 998150
rect 40546 998007 76454 999097
rect 76534 998007 90866 999177
rect 90946 998007 127854 999097
rect 127934 998007 142266 999177
rect 142346 998007 179254 999097
rect 179334 998007 193666 999177
rect 193746 998007 230543 999097
rect 230623 998007 246097 999177
rect 246177 998007 282143 999097
rect 282223 998007 297697 999177
rect 297777 998007 333654 999097
rect 333734 998007 348066 999177
rect 348146 998007 384054 999097
rect 384134 998007 398466 999177
rect 398546 998007 473054 999097
rect 473134 998007 487466 999177
rect 487546 998007 524454 999097
rect 524534 998007 538866 999177
rect 538946 998007 575854 999097
rect 575934 998007 590266 999177
rect 590346 998007 626254 999097
rect 626334 998007 640666 999177
rect 640746 998007 678070 999097
rect 678150 997927 687067 999177
rect 39673 997600 40549 997927
rect 677600 997134 687067 997927
rect 677600 997051 677927 997134
rect 30533 954534 39593 968866
rect 678007 967457 679097 997054
rect 679177 997051 679297 997134
rect 680387 997131 681477 997134
rect 679177 967377 679297 967552
rect 679377 967457 680307 997054
rect 680387 997051 680507 997131
rect 681357 997051 681477 997131
rect 680387 967377 680507 967552
rect 680587 967457 681277 997051
rect 681357 967377 681477 967552
rect 681557 967457 682487 997054
rect 682567 997051 682687 997134
rect 682567 967377 682687 967552
rect 682767 967457 683697 997054
rect 683777 997051 683897 997134
rect 683777 967377 683897 967552
rect 683977 967457 684667 997054
rect 684747 997051 684867 997134
rect 684747 967377 684867 967552
rect 684947 967457 685637 997054
rect 685717 997051 685837 997134
rect 685717 967470 685837 967552
rect 685917 967550 686847 997054
rect 686927 997051 687067 997134
rect 686927 967470 687067 967552
rect 685717 967377 687067 967470
rect 30533 954393 30673 954534
rect 30533 926666 30673 927000
rect 30753 926746 31683 954454
rect 31763 954393 31883 954534
rect 31763 926666 31883 927000
rect 31963 926746 32653 954454
rect 32733 954393 32853 954534
rect 32733 926666 32853 927000
rect 32933 926746 33623 954454
rect 33703 954393 33823 954534
rect 33903 929187 34833 954454
rect 34913 954393 35033 954534
rect 36123 954473 37213 954534
rect 33703 926666 33823 927000
rect 33903 926987 34840 929187
rect 33903 926746 34833 926987
rect 34913 926666 35033 927000
rect 35113 926746 36043 954454
rect 36123 954393 36243 954473
rect 37093 954393 37213 954473
rect 36123 926727 36243 927000
rect 36323 926807 37013 954393
rect 37093 926727 37213 927000
rect 37293 926746 38223 954454
rect 38303 954393 38423 954534
rect 36123 926666 37213 926727
rect 38303 926666 38423 927000
rect 38503 926746 39593 954454
rect 678007 952839 687067 967377
rect 678007 951903 680507 952839
rect 679177 951823 679297 951903
rect 680387 951823 680507 951903
rect 30533 912334 39593 926666
rect 678007 922346 679097 951823
rect 679177 922266 679297 922600
rect 679377 922346 680307 951823
rect 680387 922327 680507 922600
rect 680587 922407 681277 952759
rect 681357 951823 681477 952839
rect 681357 922327 681477 922600
rect 681557 922346 682487 952759
rect 682567 951903 687067 952839
rect 682567 951823 682687 951903
rect 683777 951823 683897 951903
rect 684747 951823 684867 951903
rect 685717 951823 685837 951903
rect 686927 951823 687067 951903
rect 680387 922266 681477 922327
rect 682567 922266 682687 922600
rect 682767 922346 683697 951823
rect 683777 922266 683897 922600
rect 683977 922346 684667 951823
rect 684747 922266 684867 922600
rect 684947 922346 685637 951823
rect 685917 924795 686847 951823
rect 685717 922266 685837 922600
rect 685910 922586 686847 924795
rect 685917 922346 686847 922586
rect 686927 922266 687067 922600
rect 30533 912000 30673 912334
rect 30753 912014 31683 912254
rect 30753 909805 31690 912014
rect 31763 912000 31883 912334
rect 30533 884466 30673 884607
rect 30753 884546 31683 909805
rect 31763 884466 31883 884607
rect 31963 884546 32653 912254
rect 32733 912000 32853 912334
rect 32733 884466 32853 884607
rect 32933 884546 33623 912254
rect 33703 912000 33823 912334
rect 33703 884466 33823 884607
rect 33903 884546 34833 912254
rect 34913 912000 35033 912334
rect 36123 912273 37213 912334
rect 34913 884466 35033 884607
rect 35113 884546 36043 912254
rect 36123 912000 36243 912273
rect 36323 884607 37013 912193
rect 37093 912000 37213 912273
rect 36123 884527 36243 884607
rect 37093 884527 37213 884607
rect 37293 884546 38223 912254
rect 38303 912000 38423 912334
rect 36123 884466 37213 884527
rect 38303 884466 38423 884607
rect 38503 884546 39593 912254
rect 678007 907934 687067 922266
rect 30533 870134 39593 884466
rect 677707 878066 677927 878207
rect 678007 878146 679097 907854
rect 679177 907600 679297 907934
rect 680387 907873 681477 907934
rect 679177 878066 679297 878207
rect 679377 878146 680307 907854
rect 680387 907600 680507 907873
rect 680587 878207 681277 907793
rect 681357 907600 681477 907873
rect 680387 878127 680507 878207
rect 681357 878127 681477 878207
rect 681557 878146 682487 907854
rect 682567 907600 682687 907934
rect 682767 907613 683697 907854
rect 682760 905413 683697 907613
rect 683777 907600 683897 907934
rect 680387 878066 681477 878127
rect 682567 878066 682687 878207
rect 682767 878146 683697 905413
rect 683777 878066 683897 878207
rect 683977 878146 684667 907854
rect 684747 907600 684867 907934
rect 684747 878066 684867 878207
rect 684947 878146 685637 907854
rect 685717 907600 685837 907934
rect 685717 878066 685837 878207
rect 685917 878146 686847 907854
rect 686927 907600 687067 907934
rect 686927 878066 687067 878207
rect 677707 877798 687067 878066
rect 687147 877878 687213 1001515
rect 687293 1001191 688145 1001595
rect 687293 1001055 687849 1001191
rect 30533 869993 30673 870134
rect 30533 842266 30673 842407
rect 30753 842346 31683 870054
rect 31763 869993 31883 870134
rect 31763 842266 31883 842407
rect 31963 842346 32653 870054
rect 32733 869993 32853 870134
rect 32733 842266 32853 842407
rect 32933 842346 33623 870054
rect 33703 869993 33823 870134
rect 33703 842266 33823 842407
rect 33903 842346 34833 870054
rect 34913 869993 35033 870134
rect 36123 870073 37213 870134
rect 34913 842266 35033 842407
rect 35113 842346 36043 870054
rect 36123 869993 36243 870073
rect 37093 869993 37213 870073
rect 36323 842407 37013 869993
rect 36123 842327 36243 842407
rect 37093 842327 37213 842407
rect 37293 842346 38223 870054
rect 38303 869993 38423 870134
rect 36123 842266 37213 842327
rect 38303 842266 38423 842407
rect 38503 842346 39593 870054
rect 677707 869062 687193 877798
rect 677707 862734 687067 869062
rect 677707 862606 677927 862734
rect 30407 827934 39593 842266
rect 678007 833146 679097 862654
rect 679177 862606 679297 862734
rect 680387 862686 681477 862734
rect 679177 833066 679297 833207
rect 679377 833146 680307 862654
rect 680387 862606 680507 862686
rect 681357 862606 681477 862686
rect 680587 833207 681277 862606
rect 680387 833127 680507 833207
rect 681357 833127 681477 833207
rect 681557 833146 682487 862654
rect 682567 862606 682687 862734
rect 680387 833066 681477 833127
rect 682567 833066 682687 833207
rect 682767 833146 683697 862654
rect 683777 862606 683897 862734
rect 683777 833066 683897 833207
rect 683977 833146 684667 862654
rect 684747 862606 684867 862734
rect 684747 833066 684867 833207
rect 684947 833146 685637 862654
rect 685717 862606 685837 862734
rect 685717 833066 685837 833207
rect 685917 833146 686847 862654
rect 686927 862606 687067 862734
rect 686927 833066 687067 833207
rect 29455 794909 30307 795213
rect 29455 792072 29651 794909
rect 0 791768 29651 792072
rect 0 785002 28699 791768
rect 0 784734 28573 785002
rect 0 784400 4843 784654
rect 4923 784593 20920 784734
rect 0 757200 20920 784400
rect 0 756946 4843 757200
rect 4923 756866 20920 756994
rect 21000 756946 25993 784654
rect 26073 784593 26213 784734
rect 26073 757200 26213 784400
rect 26073 756866 26213 756994
rect 26293 756946 27183 784654
rect 27263 784593 27383 784734
rect 27263 757200 27383 784400
rect 27263 756866 27383 756994
rect 27463 756946 28353 784654
rect 28433 784593 28573 784734
rect 28433 757200 28573 784400
rect 28433 756866 28573 756994
rect 0 750538 28573 756866
rect 28653 750618 28719 784922
rect 0 748872 28699 750538
rect 28779 748952 29375 791688
rect 29455 784734 29651 791768
rect 29435 756946 29671 784654
rect 29455 752013 29651 756866
rect 29731 752093 30327 794829
rect 30387 793818 30453 827854
rect 30533 827793 30673 827934
rect 30533 800066 30673 800194
rect 30753 800146 31683 827854
rect 31763 827793 31883 827934
rect 31763 800066 31883 800194
rect 31963 800146 32653 827854
rect 32733 827793 32853 827934
rect 32733 800066 32853 800194
rect 32933 800146 33623 827854
rect 33703 827793 33823 827934
rect 33703 800066 33823 800194
rect 33903 800146 34833 827854
rect 34913 827793 35033 827934
rect 36123 827873 37213 827934
rect 34913 800066 35033 800194
rect 35113 800146 36043 827854
rect 36123 827793 36243 827873
rect 37093 827793 37213 827873
rect 36323 800194 37013 827793
rect 36123 800114 36243 800194
rect 37093 800114 37213 800194
rect 37293 800146 38223 827854
rect 38303 827793 38423 827934
rect 36123 800066 37213 800114
rect 38303 800066 38423 800194
rect 38503 800146 39593 827854
rect 678007 818734 687067 833066
rect 39673 800066 39893 800194
rect 30533 793738 39893 800066
rect 30407 785002 39893 793738
rect 29455 751709 30307 752013
rect 29455 748872 29651 751709
rect 0 748568 29651 748872
rect 0 741802 28699 748568
rect 0 741534 28573 741802
rect 0 741200 4843 741454
rect 4923 741393 20920 741534
rect 0 714000 20920 741200
rect 0 713746 4843 714000
rect 4923 713666 20920 713794
rect 21000 713746 25993 741454
rect 26073 741393 26213 741534
rect 26073 714000 26213 741200
rect 26073 713666 26213 713794
rect 26293 713746 27183 741454
rect 27263 741393 27383 741534
rect 27263 714000 27383 741200
rect 27263 713666 27383 713794
rect 27463 713746 28353 741454
rect 28433 741393 28573 741534
rect 28433 714000 28573 741200
rect 28433 713666 28573 713794
rect 0 707338 28573 713666
rect 28653 707418 28719 741722
rect 0 705672 28699 707338
rect 28779 705752 29375 748488
rect 29455 741534 29651 748568
rect 29435 713746 29671 741454
rect 29455 708813 29651 713666
rect 29731 708893 30327 751629
rect 30387 750618 30453 784922
rect 30533 784734 39893 785002
rect 30533 784593 30673 784734
rect 30533 756866 30673 756994
rect 30753 756946 31683 784654
rect 31763 784593 31883 784734
rect 31763 756866 31883 756994
rect 31963 756946 32653 784654
rect 32733 784593 32853 784734
rect 32733 756866 32853 756994
rect 32933 756946 33623 784654
rect 33703 784593 33823 784734
rect 33703 756866 33823 756994
rect 33903 756946 34833 784654
rect 34913 784593 35033 784734
rect 36123 784673 37213 784734
rect 34913 756866 35033 756994
rect 35113 756946 36043 784654
rect 36123 784593 36243 784673
rect 37093 784593 37213 784673
rect 36323 756994 37013 784593
rect 36123 756914 36243 756994
rect 37093 756914 37213 756994
rect 37293 756946 38223 784654
rect 38303 784593 38423 784734
rect 36123 756866 37213 756914
rect 38303 756866 38423 756994
rect 38503 756946 39593 784654
rect 39673 784593 39893 784734
rect 677707 788866 677927 789007
rect 678007 788946 679097 818654
rect 679177 818593 679297 818734
rect 680387 818673 681477 818734
rect 679177 788866 679297 789007
rect 679377 788946 680307 818654
rect 680387 818593 680507 818673
rect 681357 818593 681477 818673
rect 680587 789007 681277 818593
rect 680387 788927 680507 789007
rect 681357 788927 681477 789007
rect 681557 788946 682487 818654
rect 682567 818593 682687 818734
rect 680387 788866 681477 788927
rect 682567 788866 682687 789007
rect 682767 788946 683697 818654
rect 683777 818593 683897 818734
rect 683777 788866 683897 789007
rect 683977 788946 684667 818654
rect 684747 818593 684867 818734
rect 684747 788866 684867 789007
rect 684947 788946 685637 818654
rect 685717 818593 685837 818734
rect 685717 788866 685837 789007
rect 685917 788946 686847 818654
rect 686927 818593 687067 818734
rect 686927 788866 687067 789007
rect 677707 788598 687067 788866
rect 687147 788678 687213 868982
rect 687273 867971 687869 1000975
rect 687929 967552 688165 1001111
rect 687949 951903 688145 967472
rect 687929 922346 688165 951823
rect 687949 907934 688145 922266
rect 687929 878146 688165 907854
rect 687949 871032 688145 878066
rect 688225 871112 688821 1002182
rect 688881 877878 688947 1002235
rect 689027 997251 717600 1002315
rect 689027 997134 691527 997251
rect 689027 997051 689167 997134
rect 689027 977000 689167 996800
rect 689027 967377 689167 967552
rect 689247 967457 690137 997054
rect 690217 997051 690337 997134
rect 690217 977000 690337 996800
rect 690217 967377 690337 967552
rect 690417 967457 691307 997054
rect 691387 997051 691527 997134
rect 691387 977000 691527 996800
rect 691387 967377 691527 967552
rect 691607 967457 696600 997171
rect 696680 997134 717600 997251
rect 696680 997051 712677 997134
rect 712757 996800 717600 997054
rect 696680 977000 717600 996800
rect 696680 967377 712677 967552
rect 689027 967279 712677 967377
rect 712757 967359 717600 977000
rect 689027 951903 717600 967279
rect 689027 951823 689167 951903
rect 690217 951823 690337 951903
rect 691387 951823 691527 951903
rect 696680 951823 712677 951903
rect 689027 922266 689167 943200
rect 689247 922346 690137 951823
rect 690217 922266 690337 943200
rect 690417 922346 691307 951823
rect 691387 922266 691527 943200
rect 691607 922346 696600 951823
rect 712757 943200 717600 951823
rect 696680 922600 717600 943200
rect 696680 922266 712677 922600
rect 712757 922346 717600 922600
rect 689027 907934 717600 922266
rect 689027 878400 689167 907934
rect 689027 878066 689167 878207
rect 689247 878146 690137 907854
rect 690217 878400 690337 907934
rect 690217 878066 690337 878207
rect 690417 878146 691307 907854
rect 691387 878400 691527 907934
rect 691387 878066 691527 878207
rect 691607 878146 696600 907854
rect 696680 907600 712677 907934
rect 712757 907643 717600 907854
rect 712750 907600 717600 907643
rect 696680 878400 717600 907600
rect 696680 878066 712677 878207
rect 712757 878146 717600 878400
rect 689027 877798 717600 878066
rect 688901 871032 717600 877798
rect 687949 870728 717600 871032
rect 687949 867891 688145 870728
rect 687293 867587 688145 867891
rect 677707 779862 687193 788598
rect 677707 773534 687067 779862
rect 677707 773406 677927 773534
rect 39673 756866 39893 756994
rect 30533 750538 39893 756866
rect 30407 741802 39893 750538
rect 29455 708509 30307 708813
rect 29455 705672 29651 708509
rect 0 705368 29651 705672
rect 0 698602 28699 705368
rect 0 698334 28573 698602
rect 0 698000 4843 698254
rect 4923 698193 20920 698334
rect 0 670800 20920 698000
rect 0 670546 4843 670800
rect 4923 670466 20920 670594
rect 21000 670546 25993 698254
rect 26073 698193 26213 698334
rect 26073 670800 26213 698000
rect 26073 670466 26213 670594
rect 26293 670546 27183 698254
rect 27263 698193 27383 698334
rect 27263 670800 27383 698000
rect 27263 670466 27383 670594
rect 27463 670546 28353 698254
rect 28433 698193 28573 698334
rect 28433 670800 28573 698000
rect 28433 670466 28573 670594
rect 0 664138 28573 670466
rect 28653 664218 28719 698522
rect 0 662472 28699 664138
rect 28779 662552 29375 705288
rect 29455 698334 29651 705368
rect 29435 670546 29671 698254
rect 29455 665613 29651 670466
rect 29731 665693 30327 708429
rect 30387 707418 30453 741722
rect 30533 741534 39893 741802
rect 30533 741393 30673 741534
rect 30533 713666 30673 713794
rect 30753 713746 31683 741454
rect 31763 741393 31883 741534
rect 31763 713666 31883 713794
rect 31963 713746 32653 741454
rect 32733 741393 32853 741534
rect 32733 713666 32853 713794
rect 32933 713746 33623 741454
rect 33703 741393 33823 741534
rect 33703 713666 33823 713794
rect 33903 713746 34833 741454
rect 34913 741393 35033 741534
rect 36123 741473 37213 741534
rect 34913 713666 35033 713794
rect 35113 713746 36043 741454
rect 36123 741393 36243 741473
rect 37093 741393 37213 741473
rect 36323 713794 37013 741393
rect 36123 713714 36243 713794
rect 37093 713714 37213 713794
rect 37293 713746 38223 741454
rect 38303 741393 38423 741534
rect 36123 713666 37213 713714
rect 38303 713666 38423 713794
rect 38503 713746 39593 741454
rect 39673 741393 39893 741534
rect 677707 743866 677927 744007
rect 678007 743946 679097 773454
rect 679177 773406 679297 773534
rect 680387 773486 681477 773534
rect 679177 743866 679297 744007
rect 679377 743946 680307 773454
rect 680387 773406 680507 773486
rect 681357 773406 681477 773486
rect 680587 744007 681277 773406
rect 680387 743927 680507 744007
rect 681357 743927 681477 744007
rect 681557 743946 682487 773454
rect 682567 773406 682687 773534
rect 680387 743866 681477 743927
rect 682567 743866 682687 744007
rect 682767 743946 683697 773454
rect 683777 773406 683897 773534
rect 683777 743866 683897 744007
rect 683977 743946 684667 773454
rect 684747 773406 684867 773534
rect 684747 743866 684867 744007
rect 684947 743946 685637 773454
rect 685717 773406 685837 773534
rect 685717 743866 685837 744007
rect 685917 743946 686847 773454
rect 686927 773406 687067 773534
rect 686927 743866 687067 744007
rect 677707 743598 687067 743866
rect 687147 743678 687213 779782
rect 687273 778771 687869 867507
rect 687949 862734 688145 867587
rect 687929 833146 688165 862654
rect 687949 818734 688145 833066
rect 687929 788946 688165 818654
rect 687949 781832 688145 788866
rect 688225 781912 688821 870648
rect 688901 869062 717600 870728
rect 688881 788678 688947 868982
rect 689027 862734 717600 869062
rect 689027 862606 689167 862734
rect 689027 833400 689167 862400
rect 689027 833066 689167 833207
rect 689247 833146 690137 862654
rect 690217 862606 690337 862734
rect 690217 833400 690337 862400
rect 690217 833066 690337 833207
rect 690417 833146 691307 862654
rect 691387 862606 691527 862734
rect 691387 833400 691527 862400
rect 691387 833066 691527 833207
rect 691607 833146 696600 862654
rect 696680 862606 712677 862734
rect 712757 862400 717600 862654
rect 696680 833400 717600 862400
rect 696680 833066 712677 833207
rect 712757 833146 717600 833400
rect 689027 818734 717600 833066
rect 689027 818593 689167 818734
rect 689027 789200 689167 818400
rect 689027 788866 689167 789007
rect 689247 788946 690137 818654
rect 690217 818593 690337 818734
rect 690217 789200 690337 818400
rect 690217 788866 690337 789007
rect 690417 788946 691307 818654
rect 691387 818593 691527 818734
rect 691387 789200 691527 818400
rect 691387 788866 691527 789007
rect 691607 788946 696600 818654
rect 696680 818593 712677 818734
rect 712757 818400 717600 818654
rect 696680 789200 717600 818400
rect 696680 788866 712677 789007
rect 712757 788946 717600 789200
rect 689027 788598 717600 788866
rect 688901 781832 717600 788598
rect 687949 781528 717600 781832
rect 687949 778691 688145 781528
rect 687293 778387 688145 778691
rect 677707 734862 687193 743598
rect 677707 728534 687067 734862
rect 677707 728406 677927 728534
rect 39673 713666 39893 713794
rect 30533 707338 39893 713666
rect 30407 698602 39893 707338
rect 29455 665309 30307 665613
rect 29455 662472 29651 665309
rect 0 662168 29651 662472
rect 0 655402 28699 662168
rect 0 655134 28573 655402
rect 0 654800 4843 655054
rect 4923 654993 20920 655134
rect 0 627600 20920 654800
rect 0 627346 4843 627600
rect 4923 627266 20920 627394
rect 21000 627346 25993 655054
rect 26073 654993 26213 655134
rect 26073 627600 26213 654800
rect 26073 627266 26213 627394
rect 26293 627346 27183 655054
rect 27263 654993 27383 655134
rect 27263 627600 27383 654800
rect 27263 627266 27383 627394
rect 27463 627346 28353 655054
rect 28433 654993 28573 655134
rect 28433 627600 28573 654800
rect 28433 627266 28573 627394
rect 0 620938 28573 627266
rect 28653 621018 28719 655322
rect 0 619272 28699 620938
rect 28779 619352 29375 662088
rect 29455 655134 29651 662168
rect 29435 627346 29671 655054
rect 29455 622413 29651 627266
rect 29731 622493 30327 665229
rect 30387 664218 30453 698522
rect 30533 698334 39893 698602
rect 30533 698193 30673 698334
rect 30533 670466 30673 670594
rect 30753 670546 31683 698254
rect 31763 698193 31883 698334
rect 31763 670466 31883 670594
rect 31963 670546 32653 698254
rect 32733 698193 32853 698334
rect 32733 670466 32853 670594
rect 32933 670546 33623 698254
rect 33703 698193 33823 698334
rect 33703 670466 33823 670594
rect 33903 670546 34833 698254
rect 34913 698193 35033 698334
rect 36123 698273 37213 698334
rect 34913 670466 35033 670594
rect 35113 670546 36043 698254
rect 36123 698193 36243 698273
rect 37093 698193 37213 698273
rect 36323 670594 37013 698193
rect 36123 670514 36243 670594
rect 37093 670514 37213 670594
rect 37293 670546 38223 698254
rect 38303 698193 38423 698334
rect 36123 670466 37213 670514
rect 38303 670466 38423 670594
rect 38503 670546 39593 698254
rect 39673 698193 39893 698334
rect 677707 698866 677927 699007
rect 678007 698946 679097 728454
rect 679177 728406 679297 728534
rect 680387 728486 681477 728534
rect 679177 698866 679297 699007
rect 679377 698946 680307 728454
rect 680387 728406 680507 728486
rect 681357 728406 681477 728486
rect 680587 699007 681277 728406
rect 680387 698927 680507 699007
rect 681357 698927 681477 699007
rect 681557 698946 682487 728454
rect 682567 728406 682687 728534
rect 680387 698866 681477 698927
rect 682567 698866 682687 699007
rect 682767 698946 683697 728454
rect 683777 728406 683897 728534
rect 683777 698866 683897 699007
rect 683977 698946 684667 728454
rect 684747 728406 684867 728534
rect 684747 698866 684867 699007
rect 684947 698946 685637 728454
rect 685717 728406 685837 728534
rect 685717 698866 685837 699007
rect 685917 698946 686847 728454
rect 686927 728406 687067 728534
rect 686927 698866 687067 699007
rect 677707 698598 687067 698866
rect 687147 698678 687213 734782
rect 687273 733771 687869 778307
rect 687949 773534 688145 778387
rect 687929 743946 688165 773454
rect 687949 736832 688145 743866
rect 688225 736912 688821 781448
rect 688901 779862 717600 781528
rect 688881 743678 688947 779782
rect 689027 773534 717600 779862
rect 689027 773406 689167 773534
rect 689027 744200 689167 773200
rect 689027 743866 689167 744007
rect 689247 743946 690137 773454
rect 690217 773406 690337 773534
rect 690217 744200 690337 773200
rect 690217 743866 690337 744007
rect 690417 743946 691307 773454
rect 691387 773406 691527 773534
rect 691387 744200 691527 773200
rect 691387 743866 691527 744007
rect 691607 743946 696600 773454
rect 696680 773406 712677 773534
rect 712757 773200 717600 773454
rect 696680 744200 717600 773200
rect 696680 743866 712677 744007
rect 712757 743946 717600 744200
rect 689027 743598 717600 743866
rect 688901 736832 717600 743598
rect 687949 736528 717600 736832
rect 687949 733691 688145 736528
rect 687293 733387 688145 733691
rect 677707 689862 687193 698598
rect 677707 683534 687067 689862
rect 677707 683406 677927 683534
rect 39673 670466 39893 670594
rect 30533 664138 39893 670466
rect 30407 655402 39893 664138
rect 29455 622109 30307 622413
rect 29455 619272 29651 622109
rect 0 618968 29651 619272
rect 0 612202 28699 618968
rect 0 611934 28573 612202
rect 0 611600 4843 611854
rect 4923 611793 20920 611934
rect 0 584400 20920 611600
rect 0 584146 4843 584400
rect 4923 584066 20920 584194
rect 21000 584146 25993 611854
rect 26073 611793 26213 611934
rect 26073 584400 26213 611600
rect 26073 584066 26213 584194
rect 26293 584146 27183 611854
rect 27263 611793 27383 611934
rect 27263 584400 27383 611600
rect 27263 584066 27383 584194
rect 27463 584146 28353 611854
rect 28433 611793 28573 611934
rect 28433 584400 28573 611600
rect 28433 584066 28573 584194
rect 0 577738 28573 584066
rect 28653 577818 28719 612122
rect 0 576072 28699 577738
rect 28779 576152 29375 618888
rect 29455 611934 29651 618968
rect 29435 584146 29671 611854
rect 29455 579213 29651 584066
rect 29731 579293 30327 622029
rect 30387 621018 30453 655322
rect 30533 655134 39893 655402
rect 30533 654993 30673 655134
rect 30533 627266 30673 627394
rect 30753 627346 31683 655054
rect 31763 654993 31883 655134
rect 31763 627266 31883 627394
rect 31963 627346 32653 655054
rect 32733 654993 32853 655134
rect 32733 627266 32853 627394
rect 32933 627346 33623 655054
rect 33703 654993 33823 655134
rect 33703 627266 33823 627394
rect 33903 627346 34833 655054
rect 34913 654993 35033 655134
rect 36123 655073 37213 655134
rect 34913 627266 35033 627394
rect 35113 627346 36043 655054
rect 36123 654993 36243 655073
rect 37093 654993 37213 655073
rect 36323 627394 37013 654993
rect 36123 627314 36243 627394
rect 37093 627314 37213 627394
rect 37293 627346 38223 655054
rect 38303 654993 38423 655134
rect 36123 627266 37213 627314
rect 38303 627266 38423 627394
rect 38503 627346 39593 655054
rect 39673 654993 39893 655134
rect 677707 653666 677927 653807
rect 678007 653746 679097 683454
rect 679177 683406 679297 683534
rect 680387 683486 681477 683534
rect 679177 653666 679297 653807
rect 679377 653746 680307 683454
rect 680387 683406 680507 683486
rect 681357 683406 681477 683486
rect 680587 653807 681277 683406
rect 680387 653727 680507 653807
rect 681357 653727 681477 653807
rect 681557 653746 682487 683454
rect 682567 683406 682687 683534
rect 680387 653666 681477 653727
rect 682567 653666 682687 653807
rect 682767 653746 683697 683454
rect 683777 683406 683897 683534
rect 683777 653666 683897 653807
rect 683977 653746 684667 683454
rect 684747 683406 684867 683534
rect 684747 653666 684867 653807
rect 684947 653746 685637 683454
rect 685717 683406 685837 683534
rect 685717 653666 685837 653807
rect 685917 653746 686847 683454
rect 686927 683406 687067 683534
rect 686927 653666 687067 653807
rect 677707 653398 687067 653666
rect 687147 653478 687213 689782
rect 687273 688771 687869 733307
rect 687949 728534 688145 733387
rect 687929 698946 688165 728454
rect 687949 691832 688145 698866
rect 688225 691912 688821 736448
rect 688901 734862 717600 736528
rect 688881 698678 688947 734782
rect 689027 728534 717600 734862
rect 689027 728406 689167 728534
rect 689027 699200 689167 728200
rect 689027 698866 689167 699007
rect 689247 698946 690137 728454
rect 690217 728406 690337 728534
rect 690217 699200 690337 728200
rect 690217 698866 690337 699007
rect 690417 698946 691307 728454
rect 691387 728406 691527 728534
rect 691387 699200 691527 728200
rect 691387 698866 691527 699007
rect 691607 698946 696600 728454
rect 696680 728406 712677 728534
rect 712757 728200 717600 728454
rect 696680 699200 717600 728200
rect 696680 698866 712677 699007
rect 712757 698946 717600 699200
rect 689027 698598 717600 698866
rect 688901 691832 717600 698598
rect 687949 691528 717600 691832
rect 687949 688691 688145 691528
rect 687293 688387 688145 688691
rect 677707 644662 687193 653398
rect 677707 638334 687067 644662
rect 677707 638206 677927 638334
rect 39673 627266 39893 627394
rect 30533 620938 39893 627266
rect 30407 612202 39893 620938
rect 29455 578909 30307 579213
rect 29455 576072 29651 578909
rect 0 575768 29651 576072
rect 0 569002 28699 575768
rect 0 568734 28573 569002
rect 0 568400 4843 568654
rect 4923 568593 20920 568734
rect 0 541200 20920 568400
rect 0 540946 4843 541200
rect 4923 540866 20920 540994
rect 21000 540946 25993 568654
rect 26073 568593 26213 568734
rect 26073 541200 26213 568400
rect 26073 540866 26213 540994
rect 26293 540946 27183 568654
rect 27263 568593 27383 568734
rect 27263 541200 27383 568400
rect 27263 540866 27383 540994
rect 27463 540946 28353 568654
rect 28433 568593 28573 568734
rect 28433 541200 28573 568400
rect 28433 540866 28573 540994
rect 0 534538 28573 540866
rect 28653 534618 28719 568922
rect 0 532872 28699 534538
rect 28779 532952 29375 575688
rect 29455 568734 29651 575768
rect 29435 540946 29671 568654
rect 29455 536013 29651 540866
rect 29731 536093 30327 578829
rect 30387 577818 30453 612122
rect 30533 611934 39893 612202
rect 30533 611793 30673 611934
rect 30533 584066 30673 584194
rect 30753 584146 31683 611854
rect 31763 611793 31883 611934
rect 31763 584066 31883 584194
rect 31963 584146 32653 611854
rect 32733 611793 32853 611934
rect 32733 584066 32853 584194
rect 32933 584146 33623 611854
rect 33703 611793 33823 611934
rect 33703 584066 33823 584194
rect 33903 584146 34833 611854
rect 34913 611793 35033 611934
rect 36123 611873 37213 611934
rect 34913 584066 35033 584194
rect 35113 584146 36043 611854
rect 36123 611793 36243 611873
rect 37093 611793 37213 611873
rect 36323 584194 37013 611793
rect 36123 584114 36243 584194
rect 37093 584114 37213 584194
rect 37293 584146 38223 611854
rect 38303 611793 38423 611934
rect 36123 584066 37213 584114
rect 38303 584066 38423 584194
rect 38503 584146 39593 611854
rect 39673 611793 39893 611934
rect 677707 608666 677927 608807
rect 678007 608746 679097 638254
rect 679177 638206 679297 638334
rect 680387 638286 681477 638334
rect 679177 608666 679297 608807
rect 679377 608746 680307 638254
rect 680387 638206 680507 638286
rect 681357 638206 681477 638286
rect 680587 608807 681277 638206
rect 680387 608727 680507 608807
rect 681357 608727 681477 608807
rect 681557 608746 682487 638254
rect 682567 638206 682687 638334
rect 680387 608666 681477 608727
rect 682567 608666 682687 608807
rect 682767 608746 683697 638254
rect 683777 638206 683897 638334
rect 683777 608666 683897 608807
rect 683977 608746 684667 638254
rect 684747 638206 684867 638334
rect 684747 608666 684867 608807
rect 684947 608746 685637 638254
rect 685717 638206 685837 638334
rect 685717 608666 685837 608807
rect 685917 608746 686847 638254
rect 686927 638206 687067 638334
rect 686927 608666 687067 608807
rect 677707 608398 687067 608666
rect 687147 608478 687213 644582
rect 687273 643571 687869 688307
rect 687949 683534 688145 688387
rect 687929 653746 688165 683454
rect 687949 646632 688145 653666
rect 688225 646712 688821 691448
rect 688901 689862 717600 691528
rect 688881 653478 688947 689782
rect 689027 683534 717600 689862
rect 689027 683406 689167 683534
rect 689027 654000 689167 683200
rect 689027 653666 689167 653807
rect 689247 653746 690137 683454
rect 690217 683406 690337 683534
rect 690217 654000 690337 683200
rect 690217 653666 690337 653807
rect 690417 653746 691307 683454
rect 691387 683406 691527 683534
rect 691387 654000 691527 683200
rect 691387 653666 691527 653807
rect 691607 653746 696600 683454
rect 696680 683406 712677 683534
rect 712757 683200 717600 683454
rect 696680 654000 717600 683200
rect 696680 653666 712677 653807
rect 712757 653746 717600 654000
rect 689027 653398 717600 653666
rect 688901 646632 717600 653398
rect 687949 646328 717600 646632
rect 687949 643491 688145 646328
rect 687293 643187 688145 643491
rect 677707 599662 687193 608398
rect 677707 593334 687067 599662
rect 677707 593206 677927 593334
rect 39673 584066 39893 584194
rect 30533 577738 39893 584066
rect 30407 569002 39893 577738
rect 29455 535709 30307 536013
rect 29455 532872 29651 535709
rect 0 532568 29651 532872
rect 0 525802 28699 532568
rect 0 525534 28573 525802
rect 0 525200 4843 525454
rect 4923 525393 20920 525534
rect 0 498000 20920 525200
rect 0 497746 4843 498000
rect 4923 497666 20920 497807
rect 21000 497746 25993 525454
rect 26073 525393 26213 525534
rect 26073 498000 26213 525200
rect 26073 497666 26213 497807
rect 26293 497746 27183 525454
rect 27263 525393 27383 525534
rect 27263 498000 27383 525200
rect 27263 497666 27383 497807
rect 27463 497746 28353 525454
rect 28433 525393 28573 525534
rect 28433 498000 28573 525200
rect 28433 497666 28573 497807
rect 0 483334 28573 497666
rect 0 483000 4843 483254
rect 4923 483193 20920 483334
rect 0 456093 20920 483000
rect 0 455800 7 456093
rect 4843 455800 20920 456093
rect 4843 455757 4850 455800
rect 4923 455466 20920 455800
rect 21000 455546 25993 483254
rect 26073 483193 26213 483334
rect 26073 455466 26213 483000
rect 26293 455546 27183 483254
rect 27263 483193 27383 483334
rect 27263 455466 27383 483000
rect 27463 455546 28353 483254
rect 28433 483193 28573 483334
rect 28433 455466 28573 483000
rect 0 441134 28573 455466
rect 0 440800 4843 441054
rect 4923 440800 20920 441134
rect 0 413600 20920 440800
rect 0 413346 4843 413600
rect 4923 413266 20920 413394
rect 21000 413346 25993 441054
rect 26073 413600 26213 441134
rect 26073 413266 26213 413394
rect 26293 413346 27183 441054
rect 27263 413600 27383 441134
rect 27263 413266 27383 413394
rect 27463 413346 28353 441054
rect 28433 413600 28573 441134
rect 28433 413266 28573 413394
rect 0 406938 28573 413266
rect 0 405272 28699 406938
rect 28779 405352 29375 532488
rect 29455 525534 29651 532568
rect 29435 497746 29671 525454
rect 29455 483334 29651 497666
rect 29435 455546 29671 483254
rect 29455 441134 29651 455466
rect 29435 413346 29671 441054
rect 29455 408413 29651 413266
rect 29731 408493 30327 535629
rect 30387 534618 30453 568922
rect 30533 568734 39893 569002
rect 30533 568593 30673 568734
rect 30533 540866 30673 540994
rect 30753 540946 31683 568654
rect 31763 568593 31883 568734
rect 31763 540866 31883 540994
rect 31963 540946 32653 568654
rect 32733 568593 32853 568734
rect 32733 540866 32853 540994
rect 32933 540946 33623 568654
rect 33703 568593 33823 568734
rect 33703 540866 33823 540994
rect 33903 540946 34833 568654
rect 34913 568593 35033 568734
rect 36123 568673 37213 568734
rect 34913 540866 35033 540994
rect 35113 540946 36043 568654
rect 36123 568593 36243 568673
rect 37093 568593 37213 568673
rect 36323 540994 37013 568593
rect 36123 540914 36243 540994
rect 37093 540914 37213 540994
rect 37293 540946 38223 568654
rect 38303 568593 38423 568734
rect 36123 540866 37213 540914
rect 38303 540866 38423 540994
rect 38503 540946 39593 568654
rect 39673 568593 39893 568734
rect 677707 563466 677927 563607
rect 678007 563546 679097 593254
rect 679177 593206 679297 593334
rect 680387 593286 681477 593334
rect 679177 563466 679297 563607
rect 679377 563546 680307 593254
rect 680387 593206 680507 593286
rect 681357 593206 681477 593286
rect 680587 563607 681277 593206
rect 680387 563527 680507 563607
rect 681357 563527 681477 563607
rect 681557 563546 682487 593254
rect 682567 593206 682687 593334
rect 680387 563466 681477 563527
rect 682567 563466 682687 563607
rect 682767 563546 683697 593254
rect 683777 593206 683897 593334
rect 683777 563466 683897 563607
rect 683977 563546 684667 593254
rect 684747 593206 684867 593334
rect 684747 563466 684867 563607
rect 684947 563546 685637 593254
rect 685717 593206 685837 593334
rect 685717 563466 685837 563607
rect 685917 563546 686847 593254
rect 686927 593206 687067 593334
rect 686927 563466 687067 563607
rect 677707 563198 687067 563466
rect 687147 563278 687213 599582
rect 687273 598571 687869 643107
rect 687949 638334 688145 643187
rect 687929 608746 688165 638254
rect 687949 601632 688145 608666
rect 688225 601712 688821 646248
rect 688901 644662 717600 646328
rect 688881 608478 688947 644582
rect 689027 638334 717600 644662
rect 689027 638206 689167 638334
rect 689027 609000 689167 638000
rect 689027 608666 689167 608807
rect 689247 608746 690137 638254
rect 690217 638206 690337 638334
rect 690217 609000 690337 638000
rect 690217 608666 690337 608807
rect 690417 608746 691307 638254
rect 691387 638206 691527 638334
rect 691387 609000 691527 638000
rect 691387 608666 691527 608807
rect 691607 608746 696600 638254
rect 696680 638206 712677 638334
rect 712757 638000 717600 638254
rect 696680 609000 717600 638000
rect 696680 608666 712677 608807
rect 712757 608746 717600 609000
rect 689027 608398 717600 608666
rect 688901 601632 717600 608398
rect 687949 601328 717600 601632
rect 687949 598491 688145 601328
rect 687293 598187 688145 598491
rect 677707 554462 687193 563198
rect 677707 548134 687067 554462
rect 677707 548006 677927 548134
rect 39673 540866 39893 540994
rect 30533 534538 39893 540866
rect 30407 525802 39893 534538
rect 29455 408109 30307 408413
rect 29455 405272 29651 408109
rect 0 404968 29651 405272
rect 0 398202 28699 404968
rect 0 397934 28573 398202
rect 0 397600 4843 397854
rect 4923 397793 20920 397934
rect 0 370400 20920 397600
rect 0 370146 4843 370400
rect 4923 370066 20920 370194
rect 21000 370146 25993 397854
rect 26073 397793 26213 397934
rect 26073 370400 26213 397600
rect 26073 370066 26213 370194
rect 26293 370146 27183 397854
rect 27263 397793 27383 397934
rect 27263 370400 27383 397600
rect 27263 370066 27383 370194
rect 27463 370146 28353 397854
rect 28433 397793 28573 397934
rect 28433 370400 28573 397600
rect 28433 370066 28573 370194
rect 0 363738 28573 370066
rect 28653 363818 28719 398122
rect 0 362072 28699 363738
rect 28779 362152 29375 404888
rect 29455 397934 29651 404968
rect 29435 370146 29671 397854
rect 29455 365213 29651 370066
rect 29731 365293 30327 408029
rect 30387 407018 30453 525722
rect 30533 525534 39893 525802
rect 30533 525393 30673 525534
rect 30533 497666 30673 497807
rect 30753 497746 31683 525454
rect 31763 525393 31883 525534
rect 31763 497666 31883 497807
rect 31963 497746 32653 525454
rect 32733 525393 32853 525534
rect 32733 497666 32853 497807
rect 32933 497746 33623 525454
rect 33703 525393 33823 525534
rect 33703 497666 33823 497807
rect 33903 497746 34833 525454
rect 34913 525393 35033 525534
rect 36123 525473 37213 525534
rect 34913 497666 35033 497807
rect 35113 497746 36043 525454
rect 36123 525393 36243 525473
rect 37093 525393 37213 525473
rect 36323 497807 37013 525393
rect 36123 497727 36243 497807
rect 37093 497727 37213 497807
rect 37293 497746 38223 525454
rect 38303 525393 38423 525534
rect 36123 497666 37213 497727
rect 38303 497666 38423 497807
rect 38503 497746 39593 525454
rect 39673 525393 39893 525534
rect 678007 518546 679097 548054
rect 679177 548006 679297 548134
rect 680387 548086 681477 548134
rect 679177 518466 679297 518607
rect 679377 518546 680307 548054
rect 680387 548006 680507 548086
rect 681357 548006 681477 548086
rect 680587 518607 681277 548006
rect 680387 518527 680507 518607
rect 681357 518527 681477 518607
rect 681557 518546 682487 548054
rect 682567 548006 682687 548134
rect 680387 518466 681477 518527
rect 682567 518466 682687 518607
rect 682767 518546 683697 548054
rect 683777 548006 683897 548134
rect 683777 518466 683897 518607
rect 683977 518546 684667 548054
rect 684747 548006 684867 548134
rect 684747 518466 684867 518607
rect 684947 518546 685637 548054
rect 685717 548006 685837 548134
rect 685717 518466 685837 518607
rect 685917 518546 686847 548054
rect 686927 548006 687067 548134
rect 686927 518466 687067 518607
rect 678007 504134 687067 518466
rect 30533 483334 39593 497666
rect 30533 483193 30673 483334
rect 30533 455466 30673 455800
rect 30753 455546 31683 483254
rect 31763 483193 31883 483334
rect 31763 455466 31883 455800
rect 31963 455546 32653 483254
rect 32733 483193 32853 483334
rect 32733 455466 32853 455800
rect 33703 483193 33823 483334
rect 33903 457987 34833 483254
rect 34913 483193 35033 483334
rect 36123 483273 37213 483334
rect 33703 455466 33823 455800
rect 33903 455787 34840 457987
rect 33903 455546 34833 455787
rect 34913 455466 35033 455800
rect 35113 455546 36043 483254
rect 36123 483193 36243 483273
rect 37093 483193 37213 483273
rect 36123 455527 36243 455800
rect 37093 455527 37213 455800
rect 38303 483193 38423 483334
rect 36123 455466 37213 455527
rect 38303 455466 38423 455800
rect 678007 474546 679097 504054
rect 679177 503993 679297 504134
rect 680387 504073 681477 504134
rect 679177 474466 679297 474800
rect 679377 474546 680307 504054
rect 680387 503993 680507 504073
rect 681357 503993 681477 504073
rect 680387 474527 680507 474800
rect 680587 474607 681277 503993
rect 681357 474527 681477 474800
rect 681557 474546 682487 504054
rect 682567 503993 682687 504134
rect 680387 474466 681477 474527
rect 682567 474466 682687 474800
rect 682767 474546 683697 504054
rect 683777 503993 683897 504134
rect 683777 474466 683897 474800
rect 683977 474546 684667 504054
rect 684747 503993 684867 504134
rect 684747 474466 684867 474800
rect 684947 474546 685637 504054
rect 685717 503993 685837 504134
rect 685917 476995 686847 504054
rect 686927 503993 687067 504134
rect 685717 474466 685837 474800
rect 685910 474786 686847 476995
rect 685917 474546 686847 474786
rect 686927 474466 687067 474800
rect 678007 460134 687067 474466
rect 30533 441134 39593 455466
rect 30533 440800 30673 441134
rect 30753 440814 31683 441054
rect 30753 438605 31690 440814
rect 31763 440800 31883 441134
rect 30533 413266 30673 413394
rect 30753 413346 31683 438605
rect 31763 413266 31883 413394
rect 31963 413346 32653 441054
rect 32733 440800 32853 441134
rect 32733 413266 32853 413394
rect 32933 413346 33623 441054
rect 33703 440800 33823 441134
rect 33703 413266 33823 413394
rect 33903 413346 34833 441054
rect 34913 440800 35033 441134
rect 36123 441073 37213 441134
rect 34913 413266 35033 413394
rect 35113 413346 36043 441054
rect 36123 440800 36243 441073
rect 36323 413394 37013 440993
rect 37093 440800 37213 441073
rect 36123 413314 36243 413394
rect 37093 413314 37213 413394
rect 37293 413346 38223 441054
rect 38303 440800 38423 441134
rect 36123 413266 37213 413314
rect 38303 413266 38423 413394
rect 38503 413346 39593 441054
rect 678007 430346 679097 460054
rect 679177 459800 679297 460134
rect 680387 460073 681477 460134
rect 679177 430266 679297 430407
rect 680387 459800 680507 460073
rect 681357 459800 681477 460073
rect 680387 430327 680507 430407
rect 681357 430327 681477 430407
rect 681557 430346 682487 460054
rect 682567 459800 682687 460134
rect 682767 459813 683697 460054
rect 682760 457613 683697 459813
rect 683777 459800 683897 460134
rect 680387 430266 681477 430327
rect 682567 430266 682687 430407
rect 682767 430346 683697 457613
rect 683777 430266 683897 430407
rect 683977 430346 684667 460054
rect 684747 459800 684867 460134
rect 684747 430266 684867 430407
rect 684947 430346 685637 460054
rect 685717 459800 685837 460134
rect 685717 430266 685837 430407
rect 685917 430346 686847 460054
rect 686927 459800 687067 460134
rect 686927 430266 687067 430407
rect 687147 430346 687213 554382
rect 687273 553371 687869 598107
rect 687949 593334 688145 598187
rect 687929 563546 688165 593254
rect 687949 556432 688145 563466
rect 688225 556512 688821 601248
rect 688901 599662 717600 601328
rect 688881 563278 688947 599582
rect 689027 593334 717600 599662
rect 689027 593206 689167 593334
rect 689027 563800 689167 593000
rect 689027 563466 689167 563607
rect 689247 563546 690137 593254
rect 690217 593206 690337 593334
rect 690217 563800 690337 593000
rect 690217 563466 690337 563607
rect 690417 563546 691307 593254
rect 691387 593206 691527 593334
rect 691387 563800 691527 593000
rect 691387 563466 691527 563607
rect 691607 563546 696600 593254
rect 696680 593206 712677 593334
rect 712757 593000 717600 593254
rect 696680 563800 717600 593000
rect 696680 563466 712677 563607
rect 712757 563546 717600 563800
rect 689027 563198 717600 563466
rect 688901 556432 717600 563198
rect 687949 556128 717600 556432
rect 687949 553291 688145 556128
rect 687293 552987 688145 553291
rect 678007 415934 687193 430266
rect 39673 413266 39893 413394
rect 30533 406938 39893 413266
rect 30407 398202 39893 406938
rect 29455 364909 30307 365213
rect 29455 362072 29651 364909
rect 0 361768 29651 362072
rect 0 355002 28699 361768
rect 0 354734 28573 355002
rect 0 354400 4843 354654
rect 4923 354593 20920 354734
rect 0 327200 20920 354400
rect 0 326946 4843 327200
rect 4923 326866 20920 326994
rect 21000 326946 25993 354654
rect 26073 354593 26213 354734
rect 26073 327200 26213 354400
rect 26073 326866 26213 326994
rect 26293 326946 27183 354654
rect 27263 354593 27383 354734
rect 27263 327200 27383 354400
rect 27263 326866 27383 326994
rect 27463 326946 28353 354654
rect 28433 354593 28573 354734
rect 28433 327200 28573 354400
rect 28433 326866 28573 326994
rect 0 320538 28573 326866
rect 28653 320618 28719 354922
rect 0 318872 28699 320538
rect 28779 318952 29375 361688
rect 29455 354734 29651 361768
rect 29435 326946 29671 354654
rect 29455 322013 29651 326866
rect 29731 322093 30327 364829
rect 30387 363818 30453 398122
rect 30533 397934 39893 398202
rect 30533 397793 30673 397934
rect 30533 370066 30673 370194
rect 30753 370146 31683 397854
rect 31763 397793 31883 397934
rect 31763 370066 31883 370194
rect 31963 370146 32653 397854
rect 32733 397793 32853 397934
rect 32733 370066 32853 370194
rect 32933 370146 33623 397854
rect 33703 397793 33823 397934
rect 33703 370066 33823 370194
rect 33903 370146 34833 397854
rect 34913 397793 35033 397934
rect 36123 397873 37213 397934
rect 34913 370066 35033 370194
rect 35113 370146 36043 397854
rect 36123 397793 36243 397873
rect 37093 397793 37213 397873
rect 36323 370194 37013 397793
rect 36123 370114 36243 370194
rect 37093 370114 37213 370194
rect 37293 370146 38223 397854
rect 38303 397793 38423 397934
rect 36123 370066 37213 370114
rect 38303 370066 38423 370194
rect 38503 370146 39593 397854
rect 39673 397793 39893 397934
rect 677707 386266 677927 386407
rect 678007 386346 679097 415854
rect 679177 415793 679297 415934
rect 680387 415873 681477 415934
rect 679177 386266 679297 386407
rect 679377 386346 680307 415854
rect 680387 415793 680507 415873
rect 681357 415793 681477 415873
rect 680587 386407 681277 415793
rect 680387 386327 680507 386407
rect 681357 386327 681477 386407
rect 681557 386346 682487 415854
rect 682567 415793 682687 415934
rect 680387 386266 681477 386327
rect 682567 386266 682687 386407
rect 682767 386346 683697 415854
rect 683777 415793 683897 415934
rect 683777 386266 683897 386407
rect 683977 386346 684667 415854
rect 684747 415793 684867 415934
rect 684747 386266 684867 386407
rect 684947 386346 685637 415854
rect 685717 415793 685837 415934
rect 685717 386266 685837 386407
rect 685917 386346 686847 415854
rect 686927 415793 687067 415934
rect 686927 386266 687067 386407
rect 677707 385998 687067 386266
rect 687147 386078 687213 415854
rect 677707 377262 687193 385998
rect 677707 370934 687067 377262
rect 677707 370806 677927 370934
rect 39673 370066 39893 370194
rect 30533 363738 39893 370066
rect 30407 355002 39893 363738
rect 29455 321709 30307 322013
rect 29455 318872 29651 321709
rect 0 318568 29651 318872
rect 0 311802 28699 318568
rect 0 311534 28573 311802
rect 0 311200 4843 311454
rect 4923 311393 20920 311534
rect 0 284000 20920 311200
rect 0 283746 4843 284000
rect 4923 283666 20920 283794
rect 21000 283746 25993 311454
rect 26073 311393 26213 311534
rect 26073 284000 26213 311200
rect 26073 283666 26213 283794
rect 26293 283746 27183 311454
rect 27263 311393 27383 311534
rect 27263 284000 27383 311200
rect 27263 283666 27383 283794
rect 27463 283746 28353 311454
rect 28433 311393 28573 311534
rect 28433 284000 28573 311200
rect 28433 283666 28573 283794
rect 0 277338 28573 283666
rect 28653 277418 28719 311722
rect 0 275672 28699 277338
rect 28779 275752 29375 318488
rect 29455 311534 29651 318568
rect 29435 283746 29671 311454
rect 29455 278813 29651 283666
rect 29731 278893 30327 321629
rect 30387 320618 30453 354922
rect 30533 354734 39893 355002
rect 30533 354593 30673 354734
rect 30533 326866 30673 326994
rect 30753 326946 31683 354654
rect 31763 354593 31883 354734
rect 31763 326866 31883 326994
rect 31963 326946 32653 354654
rect 32733 354593 32853 354734
rect 32733 326866 32853 326994
rect 32933 326946 33623 354654
rect 33703 354593 33823 354734
rect 33703 326866 33823 326994
rect 33903 326946 34833 354654
rect 34913 354593 35033 354734
rect 36123 354673 37213 354734
rect 34913 326866 35033 326994
rect 35113 326946 36043 354654
rect 36123 354593 36243 354673
rect 37093 354593 37213 354673
rect 36323 326994 37013 354593
rect 36123 326914 36243 326994
rect 37093 326914 37213 326994
rect 37293 326946 38223 354654
rect 38303 354593 38423 354734
rect 36123 326866 37213 326914
rect 38303 326866 38423 326994
rect 38503 326946 39593 354654
rect 39673 354593 39893 354734
rect 677707 341066 677927 341207
rect 678007 341146 679097 370854
rect 679177 370806 679297 370934
rect 680387 370886 681477 370934
rect 679177 341066 679297 341207
rect 679377 341146 680307 370854
rect 680387 370806 680507 370886
rect 681357 370806 681477 370886
rect 680587 341207 681277 370806
rect 680387 341127 680507 341207
rect 681357 341127 681477 341207
rect 681557 341146 682487 370854
rect 682567 370806 682687 370934
rect 680387 341066 681477 341127
rect 682567 341066 682687 341207
rect 682767 341146 683697 370854
rect 683777 370806 683897 370934
rect 683777 341066 683897 341207
rect 683977 341146 684667 370854
rect 684747 370806 684867 370934
rect 684747 341066 684867 341207
rect 684947 341146 685637 370854
rect 685717 370806 685837 370934
rect 685717 341066 685837 341207
rect 685917 341146 686847 370854
rect 686927 370806 687067 370934
rect 686927 341066 687067 341207
rect 677707 340798 687067 341066
rect 687147 340878 687213 377182
rect 687273 376171 687869 552907
rect 687949 548134 688145 552987
rect 687929 518546 688165 548054
rect 687949 504134 688145 518466
rect 687929 474546 688165 504054
rect 687949 460134 688145 474466
rect 687929 430346 688165 460054
rect 687949 415934 688145 430266
rect 687929 386346 688165 415854
rect 687949 379232 688145 386266
rect 688225 379312 688821 556048
rect 688901 554462 717600 556128
rect 689027 548134 717600 554462
rect 689027 548006 689167 548134
rect 689027 518800 689167 547800
rect 689027 518466 689167 518607
rect 689247 518546 690137 548054
rect 690217 548006 690337 548134
rect 690217 518800 690337 547800
rect 690217 518466 690337 518607
rect 690417 518546 691307 548054
rect 691387 548006 691527 548134
rect 691387 518800 691527 547800
rect 691387 518466 691527 518607
rect 691607 518546 696600 548054
rect 696680 548006 712677 548134
rect 712757 547800 717600 548054
rect 696680 518800 717600 547800
rect 696680 518466 712677 518607
rect 712757 518546 717600 518800
rect 689027 504134 717600 518466
rect 689027 503993 689167 504134
rect 689027 474466 689167 503800
rect 689247 474546 690137 504054
rect 690217 503993 690337 504134
rect 690217 474466 690337 503800
rect 690417 474546 691307 504054
rect 691387 503993 691527 504134
rect 691387 474466 691527 503800
rect 691607 474546 696600 504054
rect 696680 503993 712677 504134
rect 712757 503800 717600 504054
rect 696680 474800 717600 503800
rect 696680 474466 712677 474800
rect 712757 474546 717600 474800
rect 689027 460134 717600 474466
rect 689027 430600 689167 460134
rect 689027 430266 689167 430407
rect 689247 430346 690137 460054
rect 690217 430600 690337 460134
rect 690217 430266 690337 430407
rect 690417 430346 691307 460054
rect 691387 430600 691527 460134
rect 691387 430266 691527 430407
rect 691607 430346 696600 460054
rect 696680 459800 712677 460134
rect 712757 459843 717600 460054
rect 712750 459800 717600 459843
rect 696680 430600 717600 459800
rect 696680 430266 712677 430407
rect 712757 430346 717600 430600
rect 688901 415934 717600 430266
rect 688881 386078 688947 415854
rect 689027 415793 689167 415934
rect 689027 386600 689167 415600
rect 689027 386266 689167 386407
rect 689247 386346 690137 415854
rect 690217 415793 690337 415934
rect 690217 386600 690337 415600
rect 690217 386266 690337 386407
rect 690417 386346 691307 415854
rect 691387 415793 691527 415934
rect 691387 386600 691527 415600
rect 691387 386266 691527 386407
rect 691607 386346 696600 415854
rect 696680 415793 712677 415934
rect 712757 415600 717600 415854
rect 696680 386600 717600 415600
rect 696680 386266 712677 386407
rect 712757 386346 717600 386600
rect 689027 385998 717600 386266
rect 688901 379232 717600 385998
rect 687949 378928 717600 379232
rect 687949 376091 688145 378928
rect 687293 375787 688145 376091
rect 677707 332062 687193 340798
rect 39673 326866 39893 326994
rect 30533 320538 39893 326866
rect 677707 325734 687067 332062
rect 677707 325606 677927 325734
rect 30407 311802 39893 320538
rect 29455 278509 30307 278813
rect 29455 275672 29651 278509
rect 0 275368 29651 275672
rect 0 268602 28699 275368
rect 0 268334 28573 268602
rect 0 268000 4843 268254
rect 4923 268193 20920 268334
rect 0 240800 20920 268000
rect 0 240546 4843 240800
rect 4923 240466 20920 240594
rect 21000 240546 25993 268254
rect 26073 268193 26213 268334
rect 26073 240800 26213 268000
rect 26073 240466 26213 240594
rect 26293 240546 27183 268254
rect 27263 268193 27383 268334
rect 27263 240800 27383 268000
rect 27263 240466 27383 240594
rect 27463 240546 28353 268254
rect 28433 268193 28573 268334
rect 28433 240800 28573 268000
rect 28433 240466 28573 240594
rect 0 234138 28573 240466
rect 28653 234218 28719 268522
rect 0 232472 28699 234138
rect 28779 232552 29375 275288
rect 29455 268334 29651 275368
rect 29435 240546 29671 268254
rect 29455 235613 29651 240466
rect 29731 235693 30327 278429
rect 30387 277418 30453 311722
rect 30533 311534 39893 311802
rect 30533 311393 30673 311534
rect 30533 283666 30673 283794
rect 30753 283746 31683 311454
rect 31763 311393 31883 311534
rect 31763 283666 31883 283794
rect 31963 283746 32653 311454
rect 32733 311393 32853 311534
rect 32733 283666 32853 283794
rect 32933 283746 33623 311454
rect 33703 311393 33823 311534
rect 33703 283666 33823 283794
rect 33903 283746 34833 311454
rect 34913 311393 35033 311534
rect 36123 311473 37213 311534
rect 34913 283666 35033 283794
rect 35113 283746 36043 311454
rect 36123 311393 36243 311473
rect 37093 311393 37213 311473
rect 36323 283794 37013 311393
rect 36123 283714 36243 283794
rect 37093 283714 37213 283794
rect 37293 283746 38223 311454
rect 38303 311393 38423 311534
rect 36123 283666 37213 283714
rect 38303 283666 38423 283794
rect 38503 283746 39593 311454
rect 39673 311393 39893 311534
rect 677707 296066 677927 296207
rect 678007 296146 679097 325654
rect 679177 325606 679297 325734
rect 680387 325686 681477 325734
rect 679177 296066 679297 296207
rect 679377 296146 680307 325654
rect 680387 325606 680507 325686
rect 681357 325606 681477 325686
rect 680587 296207 681277 325606
rect 680387 296127 680507 296207
rect 681357 296127 681477 296207
rect 681557 296146 682487 325654
rect 682567 325606 682687 325734
rect 680387 296066 681477 296127
rect 682567 296066 682687 296207
rect 682767 296146 683697 325654
rect 683777 325606 683897 325734
rect 683777 296066 683897 296207
rect 683977 296146 684667 325654
rect 684747 325606 684867 325734
rect 684747 296066 684867 296207
rect 684947 296146 685637 325654
rect 685717 325606 685837 325734
rect 685717 296066 685837 296207
rect 685917 296146 686847 325654
rect 686927 325606 687067 325734
rect 686927 296066 687067 296207
rect 677707 295798 687067 296066
rect 687147 295878 687213 331982
rect 687273 330971 687869 375707
rect 687949 370934 688145 375787
rect 687929 341146 688165 370854
rect 687949 334032 688145 341066
rect 688225 334112 688821 378848
rect 688901 377262 717600 378928
rect 688881 340878 688947 377182
rect 689027 370934 717600 377262
rect 689027 370806 689167 370934
rect 689027 341400 689167 370600
rect 689027 341066 689167 341207
rect 689247 341146 690137 370854
rect 690217 370806 690337 370934
rect 690217 341400 690337 370600
rect 690217 341066 690337 341207
rect 690417 341146 691307 370854
rect 691387 370806 691527 370934
rect 691387 341400 691527 370600
rect 691387 341066 691527 341207
rect 691607 341146 696600 370854
rect 696680 370806 712677 370934
rect 712757 370600 717600 370854
rect 696680 341400 717600 370600
rect 696680 341066 712677 341207
rect 712757 341146 717600 341400
rect 689027 340798 717600 341066
rect 688901 334032 717600 340798
rect 687949 333728 717600 334032
rect 687949 330891 688145 333728
rect 687293 330587 688145 330891
rect 677707 287062 687193 295798
rect 39673 283666 39893 283794
rect 30533 277338 39893 283666
rect 677707 280734 687067 287062
rect 677707 280606 677927 280734
rect 30407 268602 39893 277338
rect 29455 235309 30307 235613
rect 29455 232472 29651 235309
rect 0 232168 29651 232472
rect 0 225402 28699 232168
rect 0 225134 28573 225402
rect 0 224800 4843 225054
rect 4923 224993 20920 225134
rect 0 197600 20920 224800
rect 0 197346 4843 197600
rect 4923 197266 20920 197394
rect 21000 197346 25993 225054
rect 26073 224993 26213 225134
rect 26073 197600 26213 224800
rect 26073 197266 26213 197394
rect 26293 197346 27183 225054
rect 27263 224993 27383 225134
rect 27263 197600 27383 224800
rect 27263 197266 27383 197394
rect 27463 197346 28353 225054
rect 28433 224993 28573 225134
rect 28433 197600 28573 224800
rect 28433 197266 28573 197394
rect 0 190938 28573 197266
rect 28653 191018 28719 225322
rect 0 189272 28699 190938
rect 28779 189352 29375 232088
rect 29455 225134 29651 232168
rect 29435 197346 29671 225054
rect 29455 192413 29651 197266
rect 29731 192493 30327 235229
rect 30387 234218 30453 268522
rect 30533 268334 39893 268602
rect 30533 268193 30673 268334
rect 30533 240466 30673 240594
rect 30753 240546 31683 268254
rect 31763 268193 31883 268334
rect 31763 240466 31883 240594
rect 31963 240546 32653 268254
rect 32733 268193 32853 268334
rect 32733 240466 32853 240594
rect 32933 240546 33623 268254
rect 33703 268193 33823 268334
rect 33703 240466 33823 240594
rect 33903 240546 34833 268254
rect 34913 268193 35033 268334
rect 36123 268273 37213 268334
rect 34913 240466 35033 240594
rect 35113 240546 36043 268254
rect 36123 268193 36243 268273
rect 37093 268193 37213 268273
rect 36323 240594 37013 268193
rect 36123 240514 36243 240594
rect 37093 240514 37213 240594
rect 37293 240546 38223 268254
rect 38303 268193 38423 268334
rect 36123 240466 37213 240514
rect 38303 240466 38423 240594
rect 38503 240546 39593 268254
rect 39673 268193 39893 268334
rect 677707 251066 677927 251207
rect 678007 251146 679097 280654
rect 679177 280606 679297 280734
rect 680387 280686 681477 280734
rect 679177 251066 679297 251207
rect 679377 251146 680307 280654
rect 680387 280606 680507 280686
rect 681357 280606 681477 280686
rect 680587 251207 681277 280606
rect 680387 251127 680507 251207
rect 681357 251127 681477 251207
rect 681557 251146 682487 280654
rect 682567 280606 682687 280734
rect 680387 251066 681477 251127
rect 682567 251066 682687 251207
rect 682767 251146 683697 280654
rect 683777 280606 683897 280734
rect 683777 251066 683897 251207
rect 683977 251146 684667 280654
rect 684747 280606 684867 280734
rect 684747 251066 684867 251207
rect 684947 251146 685637 280654
rect 685717 280606 685837 280734
rect 685717 251066 685837 251207
rect 685917 251146 686847 280654
rect 686927 280606 687067 280734
rect 686927 251066 687067 251207
rect 677707 250798 687067 251066
rect 687147 250878 687213 286982
rect 687273 285971 687869 330507
rect 687949 325734 688145 330587
rect 687929 296146 688165 325654
rect 687949 289032 688145 296066
rect 688225 289112 688821 333648
rect 688901 332062 717600 333728
rect 688881 295878 688947 331982
rect 689027 325734 717600 332062
rect 689027 325606 689167 325734
rect 689027 296400 689167 325400
rect 689027 296066 689167 296207
rect 689247 296146 690137 325654
rect 690217 325606 690337 325734
rect 690217 296400 690337 325400
rect 690217 296066 690337 296207
rect 690417 296146 691307 325654
rect 691387 325606 691527 325734
rect 691387 296400 691527 325400
rect 691387 296066 691527 296207
rect 691607 296146 696600 325654
rect 696680 325606 712677 325734
rect 712757 325400 717600 325654
rect 696680 296400 717600 325400
rect 696680 296066 712677 296207
rect 712757 296146 717600 296400
rect 689027 295798 717600 296066
rect 688901 289032 717600 295798
rect 687949 288728 717600 289032
rect 687949 285891 688145 288728
rect 687293 285587 688145 285891
rect 677707 242062 687193 250798
rect 39673 240466 39893 240594
rect 30533 234138 39893 240466
rect 677707 235734 687067 242062
rect 677707 235606 677927 235734
rect 30407 225402 39893 234138
rect 29455 192109 30307 192413
rect 29455 189272 29651 192109
rect 0 188968 29651 189272
rect 0 182202 28699 188968
rect 0 181934 28573 182202
rect 0 181600 4843 181854
rect 4923 181793 20920 181934
rect 0 126200 20920 181600
rect 0 124946 4843 126200
rect 4923 124866 20920 125007
rect 21000 124946 25993 181854
rect 26073 181793 26213 181934
rect 26073 126200 26213 181600
rect 26073 124866 26213 125007
rect 26293 124946 27183 181854
rect 27263 181793 27383 181934
rect 27263 126200 27383 181600
rect 27263 124866 27383 125007
rect 27463 124946 28353 181854
rect 28433 181793 28573 181934
rect 28433 126200 28573 181600
rect 28653 126200 28719 182122
rect 28433 124866 28573 125007
rect 0 110534 28573 124866
rect 0 110200 4843 110454
rect 4923 110393 20920 110534
rect 0 83000 20920 110200
rect 0 82746 4843 83000
rect 4923 82666 20920 83000
rect 21000 82746 25993 110454
rect 26073 110393 26213 110534
rect 26073 82666 26213 110200
rect 26293 82746 27183 110454
rect 27263 110393 27383 110534
rect 27263 82666 27383 110200
rect 27463 82746 28353 110454
rect 28433 110393 28573 110534
rect 28433 82666 28573 110200
rect 0 68334 28573 82666
rect 0 68000 4843 68254
rect 4923 68193 20920 68334
rect 0 40800 20920 68000
rect 0 40546 4843 40800
rect 4923 40466 20920 40549
rect 0 40349 20920 40466
rect 21000 40429 25993 68254
rect 26073 68193 26213 68334
rect 26073 40800 26213 68000
rect 26073 40466 26213 40549
rect 26293 40546 27183 68254
rect 27263 68193 27383 68334
rect 27263 40800 27383 68000
rect 27263 40466 27383 40549
rect 27463 40546 28353 68254
rect 28433 68193 28573 68334
rect 28433 40800 28573 68000
rect 28433 40466 28573 40549
rect 26073 40349 28573 40466
rect 0 35285 28573 40349
rect 28653 35365 28719 125200
rect 28779 35418 29375 188888
rect 29455 181934 29651 188968
rect 29435 126200 29671 181854
rect 29435 124946 29671 125200
rect 29455 110534 29651 124866
rect 29435 82746 29671 110454
rect 29455 68334 29651 82666
rect 29435 36489 29671 68254
rect 29731 36625 30327 192029
rect 30387 191018 30453 225322
rect 30533 225134 39893 225402
rect 30533 224993 30673 225134
rect 30533 197266 30673 197394
rect 30753 197346 31683 225054
rect 31763 224993 31883 225134
rect 31763 197266 31883 197394
rect 31963 197346 32653 225054
rect 32733 224993 32853 225134
rect 32733 197266 32853 197394
rect 32933 197346 33623 225054
rect 33703 224993 33823 225134
rect 33703 197266 33823 197394
rect 33903 197346 34833 225054
rect 34913 224993 35033 225134
rect 36123 225073 37213 225134
rect 34913 197266 35033 197394
rect 35113 197346 36043 225054
rect 36123 224993 36243 225073
rect 37093 224993 37213 225073
rect 36323 197394 37013 224993
rect 36123 197314 36243 197394
rect 37093 197314 37213 197394
rect 37293 197346 38223 225054
rect 38303 224993 38423 225134
rect 36123 197266 37213 197314
rect 38303 197266 38423 197394
rect 38503 197346 39593 225054
rect 39673 224993 39893 225134
rect 677707 205866 677927 206007
rect 678007 205946 679097 235654
rect 679177 235606 679297 235734
rect 680387 235686 681477 235734
rect 679177 205866 679297 206007
rect 679377 205946 680307 235654
rect 680387 235606 680507 235686
rect 681357 235606 681477 235686
rect 680587 206007 681277 235606
rect 680387 205927 680507 206007
rect 681357 205927 681477 206007
rect 681557 205946 682487 235654
rect 682567 235606 682687 235734
rect 680387 205866 681477 205927
rect 682567 205866 682687 206007
rect 682767 205946 683697 235654
rect 683777 235606 683897 235734
rect 683777 205866 683897 206007
rect 683977 205946 684667 235654
rect 684747 235606 684867 235734
rect 684747 205866 684867 206007
rect 684947 205946 685637 235654
rect 685717 235606 685837 235734
rect 685717 205866 685837 206007
rect 685917 205946 686847 235654
rect 686927 235606 687067 235734
rect 686927 205866 687067 206007
rect 677707 205598 687067 205866
rect 687147 205678 687213 241982
rect 687273 240971 687869 285507
rect 687949 280734 688145 285587
rect 687929 251146 688165 280654
rect 687949 244032 688145 251066
rect 688225 244112 688821 288648
rect 688901 287062 717600 288728
rect 688881 250878 688947 286982
rect 689027 280734 717600 287062
rect 689027 280606 689167 280734
rect 689027 251400 689167 280400
rect 689027 251066 689167 251207
rect 689247 251146 690137 280654
rect 690217 280606 690337 280734
rect 690217 251400 690337 280400
rect 690217 251066 690337 251207
rect 690417 251146 691307 280654
rect 691387 280606 691527 280734
rect 691387 251400 691527 280400
rect 691387 251066 691527 251207
rect 691607 251146 696600 280654
rect 696680 280606 712677 280734
rect 712757 280400 717600 280654
rect 696680 251400 717600 280400
rect 696680 251066 712677 251207
rect 712757 251146 717600 251400
rect 689027 250798 717600 251066
rect 688901 244032 717600 250798
rect 687949 243728 717600 244032
rect 687949 240891 688145 243728
rect 687293 240587 688145 240891
rect 39673 197266 39893 197394
rect 30533 190938 39893 197266
rect 30407 182202 39893 190938
rect 677707 196862 687193 205598
rect 677707 190534 687067 196862
rect 677707 190406 677927 190534
rect 30387 126200 30453 182122
rect 30533 181934 39893 182202
rect 30533 181793 30673 181934
rect 30753 127200 31683 181854
rect 31763 181793 31883 181934
rect 31963 126200 32653 181854
rect 32733 181793 32853 181934
rect 29751 36409 30307 36545
rect 29455 36005 30307 36409
rect 30387 36085 30453 125200
rect 30533 124866 30673 125007
rect 30753 124946 31683 126200
rect 31763 124866 31883 125007
rect 31963 124946 32653 125200
rect 32733 124866 32853 125007
rect 32933 124946 33623 181854
rect 33703 181793 33823 181934
rect 33703 124866 33823 125007
rect 33903 124946 34833 181854
rect 34913 181793 35033 181934
rect 36123 181873 37213 181934
rect 34913 124866 35033 125007
rect 35113 124946 36043 181854
rect 36123 181793 36243 181873
rect 37093 181793 37213 181873
rect 36323 126200 37013 181793
rect 37293 127200 38223 181854
rect 38303 181793 38423 181934
rect 36323 125007 37013 125200
rect 36123 124927 36243 125007
rect 37093 124927 37213 125007
rect 37293 124946 38223 126200
rect 36123 124866 37213 124927
rect 38303 124866 38423 125007
rect 38503 124946 39593 181854
rect 39673 181793 39893 181934
rect 677707 160866 677927 161007
rect 678007 160946 679097 190454
rect 679177 190406 679297 190534
rect 680387 190486 681477 190534
rect 679177 160866 679297 161007
rect 679377 160946 680307 190454
rect 680387 190406 680507 190486
rect 681357 190406 681477 190486
rect 680587 161007 681277 190406
rect 680387 160927 680507 161007
rect 681357 160927 681477 161007
rect 681557 160946 682487 190454
rect 682567 190406 682687 190534
rect 680387 160866 681477 160927
rect 682567 160866 682687 161007
rect 682767 160946 683697 190454
rect 683777 190406 683897 190534
rect 683777 160866 683897 161007
rect 683977 160946 684667 190454
rect 684747 190406 684867 190534
rect 684747 160866 684867 161007
rect 684947 160946 685637 190454
rect 685717 190406 685837 190534
rect 685717 160866 685837 161007
rect 685917 160946 686847 190454
rect 686927 190406 687067 190534
rect 686927 160866 687067 161007
rect 677707 160598 687067 160866
rect 687147 160678 687213 196782
rect 687273 195771 687869 240507
rect 687949 235734 688145 240587
rect 687929 205946 688165 235654
rect 687949 198832 688145 205866
rect 688225 198912 688821 243648
rect 688901 242062 717600 243728
rect 688881 205678 688947 241982
rect 689027 235734 717600 242062
rect 689027 235606 689167 235734
rect 689027 206200 689167 235400
rect 689027 205866 689167 206007
rect 689247 205946 690137 235654
rect 690217 235606 690337 235734
rect 690217 206200 690337 235400
rect 690217 205866 690337 206007
rect 690417 205946 691307 235654
rect 691387 235606 691527 235734
rect 691387 206200 691527 235400
rect 691387 205866 691527 206007
rect 691607 205946 696600 235654
rect 696680 235606 712677 235734
rect 712757 235400 717600 235654
rect 696680 206200 717600 235400
rect 696680 205866 712677 206007
rect 712757 205946 717600 206200
rect 689027 205598 717600 205866
rect 688901 198832 717600 205598
rect 687949 198528 717600 198832
rect 687949 195691 688145 198528
rect 687293 195387 688145 195691
rect 677707 151862 687193 160598
rect 677707 145534 687067 151862
rect 677707 145406 677927 145534
rect 30533 110534 39593 124866
rect 677707 115666 677927 115807
rect 678007 115746 679097 145454
rect 679177 145406 679297 145534
rect 680387 145486 681477 145534
rect 679177 115666 679297 115807
rect 679377 115746 680307 145454
rect 680387 145406 680507 145486
rect 681357 145406 681477 145486
rect 680587 115807 681277 145406
rect 680387 115727 680507 115807
rect 681357 115727 681477 115807
rect 681557 115746 682487 145454
rect 682567 145406 682687 145534
rect 680387 115666 681477 115727
rect 682567 115666 682687 115807
rect 682767 115746 683697 145454
rect 683777 145406 683897 145534
rect 683777 115666 683897 115807
rect 683977 115746 684667 145454
rect 684747 145406 684867 145534
rect 684747 115666 684867 115807
rect 684947 115746 685637 145454
rect 685717 145406 685837 145534
rect 685717 115666 685837 115807
rect 685917 115746 686847 145454
rect 686927 145406 687067 145534
rect 686927 115666 687067 115807
rect 677707 115398 687067 115666
rect 687147 115478 687213 151782
rect 687273 150771 687869 195307
rect 687949 190534 688145 195387
rect 687929 160946 688165 190454
rect 687949 153832 688145 160866
rect 688225 153912 688821 198448
rect 688901 196862 717600 198528
rect 688881 160678 688947 196782
rect 689027 190534 717600 196862
rect 689027 190406 689167 190534
rect 689027 161200 689167 190200
rect 689027 160866 689167 161007
rect 689247 160946 690137 190454
rect 690217 190406 690337 190534
rect 690217 161200 690337 190200
rect 690217 160866 690337 161007
rect 690417 160946 691307 190454
rect 691387 190406 691527 190534
rect 691387 161200 691527 190200
rect 691387 160866 691527 161007
rect 691607 160946 696600 190454
rect 696680 190406 712677 190534
rect 712757 190200 717600 190454
rect 696680 161200 717600 190200
rect 696680 160866 712677 161007
rect 712757 160946 717600 161200
rect 689027 160598 717600 160866
rect 688901 153832 717600 160598
rect 687949 153528 717600 153832
rect 687949 150691 688145 153528
rect 687293 150387 688145 150691
rect 30533 110393 30673 110534
rect 30533 82666 30673 83000
rect 30753 82746 31683 110454
rect 31763 110393 31883 110534
rect 31763 82666 31883 83000
rect 31963 82746 32653 110454
rect 32733 110393 32853 110534
rect 32733 82666 32853 83000
rect 32933 82746 33623 110454
rect 33703 110393 33823 110534
rect 33703 82666 33823 83000
rect 33903 82746 34833 110454
rect 34913 110393 35033 110534
rect 36123 110473 37213 110534
rect 34913 82666 35033 83000
rect 35113 82746 36043 110454
rect 36123 110393 36243 110473
rect 37093 110393 37213 110473
rect 36123 82727 36243 83000
rect 36323 82807 37013 110393
rect 37093 82727 37213 83000
rect 37293 82746 38223 110454
rect 38303 110393 38423 110534
rect 36123 82666 37213 82727
rect 38303 82666 38423 83000
rect 38503 82746 39593 110454
rect 677707 106662 687193 115398
rect 677707 100334 687067 106662
rect 677707 100206 677927 100334
rect 30533 68334 39593 82666
rect 30533 68193 30673 68334
rect 30533 40466 30673 40549
rect 30753 40546 31683 68254
rect 31763 68193 31883 68334
rect 31763 40466 31883 40549
rect 31963 40546 32653 68254
rect 32733 68193 32853 68334
rect 32733 40466 32853 40549
rect 32933 40546 33623 68254
rect 33703 68193 33823 68334
rect 33703 40466 33823 40549
rect 33903 40546 34833 68254
rect 34913 68193 35033 68334
rect 36123 68273 37213 68334
rect 34913 40466 35033 40549
rect 35113 40546 36043 68254
rect 36123 68193 36243 68273
rect 37093 68193 37213 68273
rect 36323 40549 37013 68193
rect 36123 40469 36243 40549
rect 37093 40469 37213 40549
rect 37293 40546 38223 68254
rect 38303 68193 38423 68334
rect 36123 40466 37213 40469
rect 38303 40466 38423 40549
rect 38503 40546 39593 68254
rect 39673 40466 40000 40549
rect 30533 39673 40000 40466
rect 186606 39673 202207 39893
rect 295206 39673 310807 39893
rect 350006 39673 365607 39893
rect 404806 39673 420407 39893
rect 459606 39673 475207 39893
rect 514406 39673 530007 39893
rect 677051 39673 677927 40000
rect 30533 38423 39450 39673
rect 39530 38503 79054 39593
rect 79134 38423 93466 39593
rect 93546 38503 132854 39593
rect 132934 38423 147266 39593
rect 147346 38503 186654 39593
rect 186734 38423 202066 39673
rect 202146 38503 241454 39593
rect 241534 38423 255866 39593
rect 255946 38503 295254 39593
rect 295334 38423 310666 39673
rect 310746 38503 350054 39593
rect 350134 38423 365466 39673
rect 365546 38503 404854 39593
rect 404934 38423 420266 39673
rect 420346 38503 459654 39593
rect 459734 38423 475066 39673
rect 475146 38503 514454 39593
rect 514534 38423 529866 39673
rect 529946 38503 569254 39593
rect 569334 38423 583666 39593
rect 583746 38503 623054 39593
rect 623134 38423 637466 39593
rect 637546 38503 677054 39593
rect 677134 39450 677927 39673
rect 678007 39530 679097 100254
rect 679177 100206 679297 100334
rect 680387 100286 681477 100334
rect 679377 71000 680307 100254
rect 680387 100206 680507 100286
rect 681357 100206 681477 100286
rect 680587 70000 681277 100206
rect 679177 39450 679297 40000
rect 677134 39163 679297 39450
rect 679377 39243 680307 70000
rect 680387 39626 680507 40000
rect 680587 39706 681277 69000
rect 681357 39626 681477 40000
rect 681557 39695 682487 100254
rect 682567 100206 682687 100334
rect 680387 39615 681477 39626
rect 682567 39615 682687 40000
rect 682767 39680 683697 100254
rect 683777 100206 683897 100334
rect 680387 39600 682687 39615
rect 683777 39643 683897 40000
rect 683977 39723 684667 100254
rect 684747 100206 684867 100334
rect 684947 70000 685637 100254
rect 685717 100206 685837 100334
rect 685917 71000 686847 100254
rect 686927 100206 687067 100334
rect 687147 70000 687213 106582
rect 687273 105571 687869 150307
rect 687949 145534 688145 150387
rect 687929 115746 688165 145454
rect 687949 108632 688145 115666
rect 688225 108712 688821 153448
rect 688901 151862 717600 153528
rect 688881 115478 688947 151782
rect 689027 145534 717600 151862
rect 689027 145406 689167 145534
rect 689027 116000 689167 145200
rect 689027 115666 689167 115807
rect 689247 115746 690137 145454
rect 690217 145406 690337 145534
rect 690217 116000 690337 145200
rect 690217 115666 690337 115807
rect 690417 115746 691307 145454
rect 691387 145406 691527 145534
rect 691387 116000 691527 145200
rect 691387 115666 691527 115807
rect 691607 115746 696600 145454
rect 696680 145406 712677 145534
rect 712757 145200 717600 145454
rect 696680 116000 717600 145200
rect 696680 115666 712677 115807
rect 712757 115746 717600 116000
rect 689027 115398 717600 115666
rect 688901 108632 717600 115398
rect 687949 108328 717600 108632
rect 687949 105491 688145 108328
rect 687293 105187 688145 105491
rect 684747 39653 684867 40000
rect 684947 39733 685637 69000
rect 685717 39653 685837 40000
rect 685917 39705 686847 70000
rect 684747 39643 685837 39653
rect 683777 39625 685837 39643
rect 686927 39625 687067 40000
rect 683777 39600 687067 39625
rect 680387 39163 687067 39600
rect 677134 38423 687067 39163
rect 30533 38303 40000 38423
rect 78993 38303 93607 38423
rect 132793 38303 147407 38423
rect 186606 38303 202207 38423
rect 241200 38303 256007 38423
rect 295206 38303 310807 38423
rect 350006 38303 365607 38423
rect 404806 38303 420407 38423
rect 459606 38303 475207 38423
rect 514406 38303 530007 38423
rect 569193 38303 583807 38423
rect 622993 38303 637607 38423
rect 677051 38303 687067 38423
rect 30533 37213 39163 38303
rect 39243 37293 79054 38223
rect 79134 37213 93466 38303
rect 93546 37293 132854 38223
rect 132934 37213 147266 38303
rect 147346 37293 186654 38223
rect 186734 37213 202066 38303
rect 202146 37293 241454 38223
rect 241534 37213 255866 38303
rect 255946 37293 295254 38223
rect 295334 37213 310666 38303
rect 310746 37293 350054 38223
rect 350134 37213 365466 38303
rect 365546 37293 404854 38223
rect 404934 37213 420266 38303
rect 420346 37293 459654 38223
rect 459734 37213 475066 38303
rect 475146 37293 514454 38223
rect 514534 37213 529866 38303
rect 529946 37293 569254 38223
rect 569334 37213 583666 38303
rect 583746 37293 623054 38223
rect 623134 37213 637466 38303
rect 637546 37293 677054 38223
rect 677134 37213 687067 38303
rect 30533 37093 40000 37213
rect 78993 37093 93607 37213
rect 132793 37093 147407 37213
rect 186606 37093 202207 37213
rect 241200 37093 256007 37213
rect 295206 37093 310807 37213
rect 350006 37093 365607 37213
rect 404806 37093 420407 37213
rect 459606 37093 475207 37213
rect 514406 37093 530007 37213
rect 569193 37093 583807 37213
rect 622993 37093 637607 37213
rect 677051 37093 687067 37213
rect 30533 36243 39626 37093
rect 39706 36323 78993 37013
rect 79073 36243 93527 37093
rect 132873 36243 147327 37093
rect 147407 36323 186606 37013
rect 186686 36243 202127 37093
rect 202207 36323 241393 37013
rect 241473 36243 255927 37093
rect 256007 36323 295206 37013
rect 295286 36243 310727 37093
rect 310807 36323 350006 37013
rect 350086 36243 365527 37093
rect 365607 36323 404806 37013
rect 404886 36243 420327 37093
rect 420407 36323 459606 37013
rect 459686 36243 475127 37093
rect 475207 36323 514406 37013
rect 514486 36243 529927 37093
rect 530007 36323 569193 37013
rect 569273 36243 583727 37093
rect 583807 36323 622993 37013
rect 623073 36243 637527 37093
rect 637607 36323 677051 37013
rect 677131 36243 687067 37093
rect 30533 36123 40000 36243
rect 78993 36123 93607 36243
rect 132793 36123 147407 36243
rect 186606 36123 202207 36243
rect 241200 36123 256007 36243
rect 295206 36123 310807 36243
rect 350006 36123 365607 36243
rect 404806 36123 420407 36243
rect 459606 36123 475207 36243
rect 514406 36123 530007 36243
rect 569193 36123 583807 36243
rect 622993 36123 637607 36243
rect 677051 36123 687067 36243
rect 30533 36005 39615 36123
rect 29455 35338 39615 36005
rect 28799 35285 39615 35338
rect 0 35033 39615 35285
rect 39695 35113 79054 36043
rect 79134 35033 93466 36123
rect 93546 35113 132854 36043
rect 132934 35033 147266 36123
rect 147346 35113 186654 36043
rect 186734 35033 202066 36123
rect 202146 35113 241454 36043
rect 241534 35033 255866 36123
rect 255946 35113 295254 36043
rect 295334 35033 310666 36123
rect 310746 35113 350054 36043
rect 350134 35033 365466 36123
rect 365546 35113 404854 36043
rect 404934 35033 420266 36123
rect 420346 35113 459654 36043
rect 459734 35033 475066 36123
rect 475146 35113 514454 36043
rect 514534 35033 529866 36123
rect 529946 35113 569254 36043
rect 569334 35033 583666 36123
rect 583746 35113 623054 36043
rect 623134 35033 637466 36123
rect 637546 35113 677054 36043
rect 677134 36005 687067 36123
rect 687147 36085 687213 69000
rect 677134 35733 687193 36005
rect 687273 35813 687869 105107
rect 687949 100334 688145 105187
rect 687929 70000 688165 100254
rect 677134 35610 687849 35733
rect 687929 35690 688165 69000
rect 677134 35338 688145 35610
rect 688225 35418 688821 108248
rect 688901 106662 717600 108328
rect 688881 70000 688947 106582
rect 689027 100334 717600 106662
rect 689027 100206 689167 100334
rect 689027 70000 689167 100000
rect 688881 35365 688947 69000
rect 689027 39595 689167 69000
rect 689247 39675 690137 100254
rect 690217 100206 690337 100334
rect 690217 70000 690337 100000
rect 690217 39624 690337 69000
rect 690417 39704 691307 100254
rect 691387 100206 691527 100334
rect 691387 70000 691527 100000
rect 691387 39624 691527 69000
rect 690217 39595 691527 39624
rect 689027 39391 691527 39595
rect 691607 39471 696600 100254
rect 696680 100206 712677 100334
rect 712757 100000 717600 100254
rect 696680 70000 717600 100000
rect 712757 69000 717600 70000
rect 696680 40000 717600 69000
rect 696680 39633 712677 40000
rect 712757 39713 717600 40000
rect 696680 39391 717600 39633
rect 677134 35285 688801 35338
rect 689027 35285 717600 39391
rect 677134 35033 717600 35285
rect 0 34913 40000 35033
rect 78993 34913 93607 35033
rect 132793 34913 147407 35033
rect 186606 34913 202207 35033
rect 241200 34913 256007 35033
rect 295206 34913 310807 35033
rect 350006 34913 365607 35033
rect 404806 34913 420407 35033
rect 459606 34913 475207 35033
rect 514406 34913 530007 35033
rect 569193 34913 583807 35033
rect 622993 34913 637607 35033
rect 677051 34913 717600 35033
rect 0 33823 39600 34913
rect 39680 33903 79054 34833
rect 79134 33823 93466 34913
rect 93546 33903 132854 34833
rect 132934 33823 147266 34913
rect 147346 33903 186654 34833
rect 186734 33823 202066 34913
rect 202146 33903 241454 34833
rect 241534 33823 255866 34913
rect 255946 33903 295254 34833
rect 295334 33823 310666 34913
rect 310746 33903 350054 34833
rect 350134 33823 365466 34913
rect 365546 33903 404854 34833
rect 404934 33823 420266 34913
rect 420346 33903 459654 34833
rect 459734 33823 475066 34913
rect 475146 33903 514454 34833
rect 514534 33823 529866 34913
rect 529946 33903 569254 34833
rect 569334 33823 583666 34913
rect 583746 33903 623054 34833
rect 623134 33823 637466 34913
rect 637546 33903 677054 34833
rect 677134 33823 717600 34913
rect 0 33703 40000 33823
rect 78993 33703 93607 33823
rect 132793 33703 147407 33823
rect 186606 33703 202207 33823
rect 241200 33703 256007 33823
rect 295206 33703 310807 33823
rect 350006 33703 365607 33823
rect 404806 33703 420407 33823
rect 459606 33703 475207 33823
rect 514406 33703 530007 33823
rect 569193 33703 583807 33823
rect 622993 33703 637607 33823
rect 677051 33703 717600 33823
rect 0 32853 39643 33703
rect 39723 32933 79054 33623
rect 79134 32853 93466 33703
rect 93546 32933 132854 33623
rect 132934 32853 147266 33703
rect 147346 32933 186654 33623
rect 186734 32853 202066 33703
rect 202146 32933 241454 33623
rect 241534 32853 255866 33703
rect 255946 32933 295254 33623
rect 295334 32853 310666 33703
rect 310746 32933 350054 33623
rect 350134 32853 365466 33703
rect 365546 32933 404854 33623
rect 404934 32853 420266 33703
rect 420346 32933 459654 33623
rect 459734 32853 475066 33703
rect 475146 32933 514454 33623
rect 514534 32853 529866 33703
rect 529946 32933 569254 33623
rect 569334 32853 583666 33703
rect 583746 32933 623054 33623
rect 623134 32853 637466 33703
rect 637546 32933 677054 33623
rect 677134 32853 717600 33703
rect 0 32733 40000 32853
rect 78993 32733 93607 32853
rect 132793 32733 147407 32853
rect 186606 32733 202207 32853
rect 241200 32733 256007 32853
rect 295206 32733 310807 32853
rect 350006 32733 365607 32853
rect 404806 32733 420407 32853
rect 459606 32733 475207 32853
rect 514406 32733 530007 32853
rect 569193 32733 583807 32853
rect 622993 32733 637607 32853
rect 677051 32733 717600 32853
rect 0 31883 39653 32733
rect 39733 31963 79054 32653
rect 79134 31883 93466 32733
rect 93546 31963 132854 32653
rect 132934 31883 147266 32733
rect 147346 31963 186654 32653
rect 186734 31883 202066 32733
rect 202146 31963 241454 32653
rect 241534 31883 255866 32733
rect 255946 31963 295254 32653
rect 295334 31883 310666 32733
rect 310746 31963 350054 32653
rect 350134 31883 365466 32733
rect 365546 31963 404854 32653
rect 404934 31883 420266 32733
rect 420346 31963 459654 32653
rect 459734 31883 475066 32733
rect 475146 31963 514454 32653
rect 514534 31883 529866 32733
rect 529946 31963 569254 32653
rect 569334 31883 583666 32733
rect 583746 31963 623054 32653
rect 623134 31883 637466 32733
rect 637546 31963 677054 32653
rect 677134 31883 717600 32733
rect 0 31763 40000 31883
rect 78993 31763 93607 31883
rect 132793 31763 147407 31883
rect 186606 31763 202207 31883
rect 241200 31763 256007 31883
rect 295206 31763 310807 31883
rect 350006 31763 365607 31883
rect 404806 31763 420407 31883
rect 459606 31763 475207 31883
rect 514406 31763 530007 31883
rect 569193 31763 583807 31883
rect 622993 31763 637607 31883
rect 677051 31763 717600 31883
rect 0 30673 39625 31763
rect 39705 30753 79054 31683
rect 79134 30673 93466 31763
rect 132934 31754 147266 31763
rect 132949 30682 147266 31754
rect 147346 30753 186654 31683
rect 132934 30673 147266 30682
rect 186734 30673 202066 31763
rect 202146 30753 241454 31683
rect 241534 30673 255866 31763
rect 255946 30753 295254 31683
rect 295334 30673 310666 31763
rect 310746 30753 350054 31683
rect 350134 30673 365466 31763
rect 365546 30753 404854 31683
rect 404934 30673 420266 31763
rect 420346 30753 459654 31683
rect 459734 30673 475066 31763
rect 475146 30753 514454 31683
rect 514534 30673 529866 31763
rect 529946 30753 569254 31683
rect 569334 30673 583666 31763
rect 583746 30753 623054 31683
rect 623134 30673 637466 31763
rect 637546 30753 677054 31683
rect 677134 30673 717600 31763
rect 0 30533 40000 30673
rect 78993 30533 93607 30673
rect 132793 30533 147407 30673
rect 186606 30533 202207 30673
rect 241200 30533 256007 30673
rect 295206 30533 310807 30673
rect 350006 30533 365607 30673
rect 404806 30533 420407 30673
rect 459606 30533 475207 30673
rect 514406 30533 530007 30673
rect 569193 30533 583807 30673
rect 622993 30533 637607 30673
rect 677051 30533 717600 30673
rect 0 30407 36005 30533
rect 0 29751 35733 30407
rect 36085 30387 79054 30453
rect 79134 30407 93466 30533
rect 93546 30387 192982 30453
rect 193062 30407 201798 30533
rect 201878 30387 301582 30453
rect 301662 30407 310398 30533
rect 310478 30387 356382 30453
rect 356462 30407 365198 30533
rect 365278 30387 411182 30453
rect 411262 30407 419998 30533
rect 420078 30387 465982 30453
rect 466062 30407 474798 30533
rect 474878 30387 520782 30453
rect 520862 30407 529598 30533
rect 529678 30387 681515 30453
rect 0 29455 35610 29751
rect 35813 29731 191507 30327
rect 0 28799 35338 29455
rect 35690 29435 79054 29671
rect 79134 29455 93466 29651
rect 93546 29435 132854 29671
rect 132934 29455 147266 29651
rect 147346 29435 186654 29671
rect 191587 29651 191891 30307
rect 191971 29731 300107 30327
rect 186734 29455 202066 29651
rect 0 28573 35285 28799
rect 35418 28779 194648 29375
rect 35365 28653 79054 28719
rect 79134 28573 93466 28699
rect 194728 28699 195032 29455
rect 202146 29435 241454 29671
rect 241534 29455 255866 29651
rect 255946 29435 295254 29671
rect 300187 29651 300491 30307
rect 300571 29731 354907 30327
rect 295334 29455 310666 29651
rect 195112 28779 303248 29375
rect 193062 28573 201798 28699
rect 201878 28653 301582 28719
rect 303328 28699 303632 29455
rect 310746 29435 350054 29671
rect 354987 29651 355291 30307
rect 355371 29731 409707 30327
rect 350134 29455 365466 29651
rect 303712 28779 358048 29375
rect 301662 28573 310398 28699
rect 310478 28653 356382 28719
rect 358128 28699 358432 29455
rect 365546 29435 404854 29671
rect 409787 29651 410091 30307
rect 410171 29731 464507 30327
rect 404934 29455 420266 29651
rect 358512 28779 412848 29375
rect 356462 28573 365198 28699
rect 365278 28653 411182 28719
rect 412928 28699 413232 29455
rect 420346 29435 459654 29671
rect 464587 29651 464891 30307
rect 464971 29731 519307 30327
rect 459734 29455 475066 29651
rect 413312 28779 467648 29375
rect 411262 28573 419998 28699
rect 420078 28653 465982 28719
rect 467728 28699 468032 29455
rect 475146 29435 514454 29671
rect 519387 29651 519691 30307
rect 519771 29731 680975 30327
rect 681595 30307 717600 30533
rect 681055 29751 717600 30307
rect 514534 29455 529866 29651
rect 468112 28779 522448 29375
rect 466062 28573 474798 28699
rect 474878 28653 520782 28719
rect 522528 28699 522832 29455
rect 529946 29435 569254 29671
rect 569334 29455 583666 29651
rect 583746 29435 623054 29671
rect 623134 29455 637466 29651
rect 637546 29435 681111 29671
rect 681191 29455 717600 29751
rect 522912 28779 682182 29375
rect 682262 28799 717600 29455
rect 520862 28573 529598 28699
rect 529678 28653 682235 28719
rect 682315 28573 717600 28799
rect 0 28433 78800 28573
rect 78993 28433 93607 28573
rect 93800 28433 132600 28573
rect 132793 28433 147407 28573
rect 147600 28433 186400 28573
rect 186606 28433 202207 28573
rect 202400 28433 256007 28573
rect 256200 28433 295000 28573
rect 295206 28433 310807 28573
rect 311000 28433 349800 28573
rect 350006 28433 365607 28573
rect 365800 28433 404600 28573
rect 404806 28433 420407 28573
rect 420600 28433 459400 28573
rect 459606 28433 475207 28573
rect 475400 28433 514200 28573
rect 514406 28433 530007 28573
rect 530200 28433 569000 28573
rect 569193 28433 583807 28573
rect 584000 28433 622800 28573
rect 622993 28433 637607 28573
rect 637800 28433 676800 28573
rect 677051 28433 717600 28573
rect 0 27383 39595 28433
rect 39675 27463 79054 28353
rect 79134 27383 93466 28433
rect 93546 27463 132854 28353
rect 132934 27383 147266 28433
rect 147346 27463 186654 28353
rect 186734 27383 202066 28433
rect 202146 27463 241454 28353
rect 241534 27383 255866 28433
rect 255946 27463 295254 28353
rect 295334 27383 310666 28433
rect 310746 27463 350054 28353
rect 350134 27383 365466 28433
rect 365546 27463 404854 28353
rect 404934 27383 420266 28433
rect 420346 27463 459654 28353
rect 459734 27383 475066 28433
rect 475146 27463 514454 28353
rect 514534 27383 529866 28433
rect 529946 27463 569254 28353
rect 569334 27383 583666 28433
rect 583746 27463 623054 28353
rect 623134 27383 637466 28433
rect 637546 27463 677054 28353
rect 677134 27383 717600 28433
rect 0 27263 78800 27383
rect 78993 27263 93607 27383
rect 93800 27263 132600 27383
rect 132793 27263 147407 27383
rect 147600 27263 186400 27383
rect 186606 27263 202207 27383
rect 202400 27263 256007 27383
rect 256200 27263 295000 27383
rect 295206 27263 310807 27383
rect 311000 27263 349800 27383
rect 350006 27263 365607 27383
rect 365800 27263 404600 27383
rect 404806 27263 420407 27383
rect 420600 27263 459400 27383
rect 459606 27263 475207 27383
rect 475400 27263 514200 27383
rect 514406 27263 530007 27383
rect 530200 27263 569000 27383
rect 569193 27263 583807 27383
rect 584000 27263 622800 27383
rect 622993 27263 637607 27383
rect 637800 27263 676800 27383
rect 677051 27263 717600 27383
rect 0 26213 39624 27263
rect 39704 26293 79054 27183
rect 79134 26213 93466 27263
rect 93546 26293 132854 27183
rect 132934 26213 147266 27263
rect 147346 26293 186654 27183
rect 186734 26213 202066 27263
rect 202146 26293 241454 27183
rect 241534 26213 255866 27263
rect 255946 26293 295254 27183
rect 295334 26213 310666 27263
rect 310746 26293 350054 27183
rect 350134 26213 365466 27263
rect 365546 26293 404854 27183
rect 404934 26213 420266 27263
rect 420346 26293 459654 27183
rect 459734 26213 475066 27263
rect 475146 26293 514454 27183
rect 514534 26213 529866 27263
rect 529946 26293 569254 27183
rect 569334 26213 583666 27263
rect 583746 26293 623054 27183
rect 623134 26213 637466 27263
rect 637546 26293 677054 27183
rect 677134 26213 717600 27263
rect 0 26073 78800 26213
rect 78993 26073 93607 26213
rect 93800 26073 132600 26213
rect 132793 26073 147407 26213
rect 147600 26073 186400 26213
rect 186606 26073 202207 26213
rect 202400 26073 256007 26213
rect 256200 26073 295000 26213
rect 295206 26073 310807 26213
rect 311000 26073 349800 26213
rect 350006 26073 365607 26213
rect 365800 26073 404600 26213
rect 404806 26073 420407 26213
rect 420600 26073 459400 26213
rect 459606 26073 475207 26213
rect 475400 26073 514200 26213
rect 514406 26073 530007 26213
rect 530200 26073 569000 26213
rect 569193 26073 583807 26213
rect 584000 26073 622800 26213
rect 622993 26073 637607 26213
rect 637800 26073 676800 26213
rect 677051 26073 717600 26213
rect 0 20920 39391 26073
rect 39471 21000 79054 25993
rect 79134 20920 93466 26073
rect 93546 21000 132854 25993
rect 132934 20920 147266 26073
rect 147346 21000 186654 25993
rect 186734 20920 202066 26073
rect 202146 21000 241454 25993
rect 241534 20920 255866 26073
rect 255946 21000 295254 25993
rect 295334 20920 310666 26073
rect 310746 21000 350054 25993
rect 350134 20920 365466 26073
rect 365546 21000 404854 25993
rect 404934 20920 420266 26073
rect 420346 21000 459654 25993
rect 459734 20920 475066 26073
rect 475146 21000 514454 25993
rect 514534 20920 529866 26073
rect 529946 21000 569254 25993
rect 569334 20920 583666 26073
rect 583746 21000 623054 25993
rect 623134 20920 637466 26073
rect 637546 21000 677171 25993
rect 677251 20920 717600 26073
rect 0 4923 78800 20920
rect 78993 4923 93607 20920
rect 0 0 39633 4923
rect 40000 4843 78800 4923
rect 39713 0 79054 4843
rect 79134 0 93466 4923
rect 93800 4843 132600 20920
rect 132793 4923 147407 20920
rect 93546 0 132854 4843
rect 132934 0 147266 4923
rect 147600 4843 186400 20920
rect 186606 4923 202207 20920
rect 202400 4923 256007 20920
rect 147346 0 186654 4843
rect 186734 0 202066 4923
rect 202400 4843 241200 4923
rect 202146 0 241454 4843
rect 241534 0 255866 4923
rect 256200 4843 295000 20920
rect 295206 4923 310807 20920
rect 255946 0 295254 4843
rect 295334 0 310666 4923
rect 311000 4843 349800 20920
rect 350006 4923 365607 20920
rect 310746 0 350054 4843
rect 350134 0 365466 4923
rect 365800 4843 404600 20920
rect 404806 4923 420407 20920
rect 365546 0 404854 4843
rect 404934 0 420266 4923
rect 420600 4843 459400 20920
rect 459606 4923 475207 20920
rect 420346 0 459654 4843
rect 459734 0 475066 4923
rect 475400 4843 514200 20920
rect 514406 4923 530007 20920
rect 475146 0 514454 4843
rect 514534 0 529866 4923
rect 530200 4843 569000 20920
rect 569193 4923 583807 20920
rect 529946 0 569254 4843
rect 569334 0 583666 4923
rect 584000 4843 622800 20920
rect 622993 4923 637607 20920
rect 583746 0 623054 4843
rect 623134 0 637466 4923
rect 637800 4843 676800 20920
rect 677051 4923 717600 20920
rect 637546 0 677054 4843
rect 677134 0 717600 4923
<< metal5 >>
rect 77610 1018624 89778 1030789
rect 129010 1018624 141178 1030789
rect 180410 1018624 192578 1030789
rect 231810 1018624 243978 1030789
rect 283410 1018624 295578 1030789
rect 334810 1018624 346978 1030789
rect 385210 1018624 397378 1030789
rect 474210 1018624 486378 1030789
rect 525610 1018624 537778 1030789
rect 577010 1018624 589178 1030789
rect 627410 1018624 639578 1030789
rect 6811 955610 18976 967778
rect 698624 954022 710789 966190
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876180
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786620 19088 799160
rect 698512 774440 711002 786980
rect 6598 743420 19088 755960
rect 698512 729440 711002 741980
rect 6598 700220 19088 712760
rect 698512 684440 711002 696980
rect 6598 657020 19088 669560
rect 698512 639240 711002 651780
rect 6598 613820 19088 626360
rect 698512 594240 711002 606780
rect 6598 570620 19088 583160
rect 698512 549040 711002 561580
rect 6598 527420 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399820 19088 412360
rect 698512 371840 711002 384380
rect 6598 356620 19088 369160
rect 6598 313420 19088 325960
rect 698512 326640 711002 339180
rect 6598 270220 19088 282760
rect 698512 281640 711002 294180
rect 6598 227020 19088 239560
rect 698512 236640 711002 249180
rect 6598 183820 19088 196360
rect 698512 191440 711002 203980
rect 698512 146440 711002 158980
rect 6811 111610 18976 123778
rect 698512 101240 711002 113780
rect 6167 70054 19620 80934
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200180 19088
rect 243266 6167 254146 19620
rect 296240 6598 308780 19088
rect 351040 6598 363580 19088
rect 405840 6598 418380 19088
rect 460640 6598 473180 19088
rect 515440 6598 527980 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
<< obsm5 >>
rect 0 1032757 76454 1037600
rect 0 1016917 40800 1032757
rect 76774 1032437 90626 1037600
rect 90946 1032757 127854 1037600
rect 128174 1032437 142026 1037600
rect 142346 1032757 179254 1037600
rect 179574 1032437 193426 1037600
rect 193746 1032757 384054 1037600
rect 76200 1031109 91200 1032437
rect 76200 1018304 77290 1031109
rect 90098 1018304 91200 1031109
rect 76200 1016917 91200 1018304
rect 127600 1031109 142600 1032437
rect 127600 1018304 128690 1031109
rect 141498 1018304 142600 1031109
rect 127600 1016917 142600 1018304
rect 179000 1031109 194000 1032437
rect 179000 1018304 180090 1031109
rect 192898 1018304 194000 1031109
rect 179000 1016917 194000 1018304
rect 221000 1031109 254800 1032757
rect 221000 1018304 231490 1031109
rect 244298 1018304 254800 1031109
rect 221000 1016917 254800 1018304
rect 272600 1031109 306400 1032757
rect 272600 1018304 283090 1031109
rect 295898 1018304 306400 1031109
rect 272600 1016917 306400 1018304
rect 333400 1031109 348400 1032757
rect 384374 1032437 398226 1037600
rect 398546 1032757 473054 1037600
rect 473374 1032437 487226 1037600
rect 487546 1032757 524454 1037600
rect 524774 1032437 538626 1037600
rect 538946 1032757 626254 1037600
rect 333400 1018304 334490 1031109
rect 347298 1018304 348400 1031109
rect 333400 1016917 348400 1018304
rect 383800 1031109 398800 1032437
rect 383800 1018304 384890 1031109
rect 397698 1018304 398800 1031109
rect 383800 1016917 398800 1018304
rect 472800 1031109 487800 1032437
rect 472800 1018304 473890 1031109
rect 486698 1018304 487800 1031109
rect 472800 1016917 487800 1018304
rect 524200 1031109 539200 1032437
rect 524200 1018304 525290 1031109
rect 538098 1018304 539200 1031109
rect 524200 1016917 539200 1018304
rect 575600 1031109 590600 1032757
rect 626574 1032437 640426 1037600
rect 640746 1032757 717600 1037600
rect 575600 1018304 576690 1031109
rect 589498 1018304 590600 1031109
rect 575600 1016917 590600 1018304
rect 626000 1031109 641000 1032437
rect 626000 1018304 627090 1031109
rect 639898 1018304 641000 1031109
rect 626000 1016917 641000 1018304
rect 677600 1016917 717600 1032757
rect 0 1011287 40109 1016917
rect 40429 1011607 76454 1016597
rect 0 1009267 40226 1011287
rect 40546 1010437 76454 1011287
rect 40546 1009267 76454 1010117
rect 0 1006827 35049 1009267
rect 35369 1007147 76454 1008947
rect 0 1002551 40226 1006827
rect 40546 1005937 76454 1006827
rect 40546 1004968 76454 1005617
rect 76774 1004968 90626 1016917
rect 90946 1011607 127854 1016597
rect 90946 1010437 127854 1011287
rect 90946 1009267 127854 1010117
rect 90946 1007147 127854 1008947
rect 90946 1005937 127854 1006827
rect 90946 1004968 127854 1005617
rect 128174 1004968 142026 1016917
rect 142346 1011607 179254 1016597
rect 142346 1010437 179254 1011287
rect 142346 1009267 179254 1010117
rect 142346 1007147 179254 1008947
rect 142346 1005937 179254 1006827
rect 142346 1004968 179254 1005617
rect 179574 1004968 193426 1016917
rect 193746 1011607 230543 1016597
rect 193746 1010437 230543 1011287
rect 193746 1009267 230543 1010117
rect 230863 1008947 245857 1016917
rect 246177 1011607 282143 1016597
rect 246177 1010437 282143 1011287
rect 246177 1009267 282143 1010117
rect 282463 1008947 297457 1016917
rect 297777 1011607 333654 1016597
rect 297777 1010437 333654 1011287
rect 297777 1009267 333654 1010117
rect 193746 1007147 230448 1008947
rect 230768 1007147 245857 1008947
rect 246177 1007147 282048 1008947
rect 282368 1007147 297457 1008947
rect 297777 1007147 333654 1008947
rect 193746 1005937 230543 1006827
rect 193746 1004968 230543 1005617
rect 40800 1004967 230543 1004968
rect 40546 1003997 76454 1004647
rect 40546 1002787 76454 1003677
rect 0 998449 28333 1002551
rect 0 997600 20683 998449
rect 26313 998245 28333 998449
rect 26313 998216 27163 998245
rect 0 968946 4843 997600
rect 5163 968626 20683 969200
rect 21003 968946 25993 998129
rect 26313 968946 27163 997896
rect 27483 968946 28333 997925
rect 28653 968946 30453 1002231
rect 30773 1001257 40226 1002551
rect 40546 1001577 76454 1002467
rect 76774 1001257 90626 1004967
rect 90946 1003997 127854 1004647
rect 90946 1002787 127854 1003677
rect 90946 1001577 127854 1002467
rect 128174 1001257 142026 1004967
rect 142346 1003997 179254 1004647
rect 142346 1002787 179254 1003677
rect 142346 1001577 179254 1002467
rect 179574 1001257 193426 1004967
rect 193746 1003997 230543 1004647
rect 193746 1002787 230543 1003677
rect 193746 1001577 230543 1002467
rect 230863 1001577 245857 1007147
rect 246177 1005937 282143 1006827
rect 246177 1004967 282143 1005617
rect 246177 1003997 282143 1004647
rect 246177 1002787 282143 1003677
rect 246177 1001577 282143 1002467
rect 282463 1001577 297457 1007147
rect 297777 1005937 333654 1006827
rect 297777 1004968 333654 1005617
rect 333974 1004968 347826 1016917
rect 348146 1011607 384054 1016597
rect 348146 1010437 384054 1011287
rect 348146 1009267 384054 1010117
rect 348146 1007147 381800 1008947
rect 382800 1007147 384054 1008947
rect 348146 1005937 382800 1006827
rect 383800 1005937 384054 1006827
rect 348146 1004968 381800 1005617
rect 297777 1004967 381800 1004968
rect 382800 1004968 384054 1005617
rect 384374 1004968 398226 1016917
rect 398546 1011607 473054 1016597
rect 398546 1010437 473054 1011287
rect 398546 1009267 473054 1010117
rect 398546 1007147 473054 1008947
rect 398546 1005937 473054 1006827
rect 398546 1004968 473054 1005617
rect 473374 1004968 487226 1016917
rect 487546 1011607 524454 1016597
rect 487546 1010437 524454 1011287
rect 487546 1009267 524454 1010117
rect 487546 1007147 524454 1008947
rect 487546 1005937 524454 1006827
rect 487546 1004968 524454 1005617
rect 524774 1004968 538626 1016917
rect 538946 1011607 575854 1016597
rect 538946 1010437 575854 1011287
rect 538946 1009267 575854 1010117
rect 538946 1007147 575854 1008947
rect 538946 1005937 575854 1006827
rect 538946 1004968 575854 1005617
rect 576174 1004968 590026 1016917
rect 590346 1011607 626254 1016597
rect 590346 1010437 626254 1011287
rect 590346 1009267 626254 1010117
rect 590346 1007147 626254 1008947
rect 590346 1005937 626254 1006827
rect 590346 1004968 626254 1005617
rect 626574 1004968 640426 1016917
rect 640746 1011607 678129 1016597
rect 678449 1011287 717600 1016917
rect 640746 1010437 677896 1011287
rect 678216 1010437 717600 1011287
rect 640746 1009267 677925 1010117
rect 678245 1009267 717600 1010437
rect 640746 1007147 682231 1008947
rect 682551 1006827 717600 1009267
rect 640746 1005937 677895 1006827
rect 678215 1005617 717600 1006827
rect 640746 1004968 677867 1005617
rect 382800 1004967 677867 1004968
rect 678187 1004967 717600 1005617
rect 297777 1003997 333654 1004647
rect 297777 1002787 333654 1003677
rect 297777 1001577 333654 1002467
rect 30773 1000607 40229 1001257
rect 40549 1000607 76393 1001257
rect 76713 1000607 90687 1001257
rect 91007 1000607 127793 1001257
rect 128113 1000607 142087 1001257
rect 142407 1000607 179193 1001257
rect 179513 1000607 193487 1001257
rect 193807 1000607 230543 1001257
rect 30773 998677 40226 1000607
rect 40546 999397 76454 1000287
rect 30773 998240 36993 998677
rect 38523 998390 40226 998677
rect 30773 998215 33603 998240
rect 35133 998225 36993 998240
rect 31983 998197 33603 998215
rect 36343 998214 36993 998225
rect 31983 998187 32633 998197
rect 30773 968946 31663 997895
rect 31983 968946 32633 997867
rect 32953 968946 33603 997877
rect 33923 968946 34813 997920
rect 35133 968946 36023 997905
rect 36343 969007 36993 997894
rect 37313 968946 38203 998357
rect 38523 968946 39573 998070
rect 39893 997707 40226 998390
rect 40546 998027 76454 999077
rect 76774 998027 90626 1000607
rect 90946 999397 127854 1000287
rect 90946 998027 127854 999077
rect 128174 998027 142026 1000607
rect 142346 999397 179254 1000287
rect 142346 998027 179254 999077
rect 179574 998027 193426 1000607
rect 230863 1000287 244921 1001577
rect 245241 1000607 282143 1001257
rect 282463 1000287 296521 1001577
rect 333974 1001257 347826 1004967
rect 348146 1003997 384054 1004647
rect 348146 1002787 384054 1003677
rect 348146 1001577 384054 1002467
rect 384374 1001257 398226 1004967
rect 398546 1003997 473054 1004647
rect 398546 1002787 473054 1003677
rect 398546 1001577 473054 1002467
rect 473374 1001257 487226 1004967
rect 487546 1003997 524454 1004647
rect 487546 1002787 524454 1003677
rect 487546 1001577 524454 1002467
rect 524774 1001257 538626 1004967
rect 538946 1003997 575854 1004647
rect 538946 1002787 575854 1003677
rect 538946 1001577 575854 1002467
rect 576174 1001257 590026 1004967
rect 590346 1003997 626254 1004647
rect 590346 1002787 626254 1003677
rect 590346 1001577 626254 1002467
rect 626574 1001257 640426 1004967
rect 640746 1003997 677877 1004647
rect 678197 1003997 717600 1004967
rect 640746 1002787 677920 1003677
rect 678240 1002551 717600 1003997
rect 678240 1002467 686827 1002551
rect 640746 1001577 677905 1002467
rect 678225 1001257 686827 1002467
rect 296841 1000607 333593 1001257
rect 333913 1000607 347887 1001257
rect 348207 1000607 381800 1001257
rect 382800 1000607 383993 1001257
rect 384313 1000607 398287 1001257
rect 398607 1000607 472993 1001257
rect 473313 1000607 487287 1001257
rect 487607 1000607 524393 1001257
rect 524713 1000607 538687 1001257
rect 539007 1000607 575793 1001257
rect 576113 1000607 590087 1001257
rect 590407 1000607 626193 1001257
rect 626513 1000607 640487 1001257
rect 640807 1000607 677894 1001257
rect 678214 1000607 686827 1001257
rect 193746 999397 230543 1000287
rect 193746 998027 230543 999077
rect 230863 998027 245857 1000287
rect 246177 999397 282143 1000287
rect 246177 998027 282143 999077
rect 282463 998027 297457 1000287
rect 297777 999397 333654 1000287
rect 297777 998027 333654 999077
rect 333974 998027 347826 1000607
rect 348146 999397 382800 1000287
rect 383800 999397 384054 1000287
rect 348146 998027 384054 999077
rect 384374 998027 398226 1000607
rect 398546 999397 473054 1000287
rect 398546 998027 473054 999077
rect 473374 998027 487226 1000607
rect 487546 999397 524454 1000287
rect 487546 998027 524454 999077
rect 524774 998027 538626 1000607
rect 538946 999397 575854 1000287
rect 538946 998027 575854 999077
rect 576174 998027 590026 1000607
rect 590346 999397 626254 1000287
rect 590346 998027 626254 999077
rect 626574 998027 640426 1000607
rect 640746 999397 678357 1000287
rect 678677 999077 686827 1000607
rect 640746 998027 678070 999077
rect 678390 997707 686827 999077
rect 39893 997600 40800 997707
rect 677600 997374 686827 997707
rect 677600 996800 677707 997374
rect 680607 997371 681257 997374
rect 32632 968626 32633 968946
rect 36343 968626 36993 968687
rect 0 968098 39573 968626
rect 0 955290 6491 968098
rect 19296 955290 39573 968098
rect 678027 967457 679077 997054
rect 679397 967457 680287 997054
rect 680607 967457 681257 997051
rect 681577 967457 682467 997054
rect 682787 967457 683677 997054
rect 683997 967457 684647 997054
rect 684968 996800 685617 997054
rect 684967 967457 685617 996800
rect 685937 967457 686827 997054
rect 687147 967552 688947 1002231
rect 689267 997491 717600 1002551
rect 689267 997374 691287 997491
rect 689267 967457 690117 997054
rect 690437 967457 691287 997054
rect 691607 967457 696597 997171
rect 696917 996800 717600 997491
rect 712757 977000 717600 996800
rect 687147 967137 688947 967232
rect 696917 967137 717600 977000
rect 0 954774 39573 955290
rect 678027 966510 717600 967137
rect 0 927000 4843 954454
rect 5163 954200 20683 954774
rect 32632 954454 32633 954774
rect 36343 954713 36993 954774
rect 0 926426 20683 927000
rect 21003 926746 25993 954454
rect 26313 926746 27163 954454
rect 27483 926746 28333 954454
rect 28653 926746 30453 954454
rect 30773 926746 31663 954454
rect 31983 927000 32633 954454
rect 31983 926746 32632 927000
rect 32953 926746 33603 954454
rect 33923 926746 34813 954454
rect 35133 926746 36023 954454
rect 36343 926807 36993 954393
rect 37313 926746 38203 954454
rect 38523 926746 39573 954454
rect 678027 953702 698304 966510
rect 711109 953702 717600 966510
rect 678027 953079 717600 953702
rect 678027 952143 680287 953079
rect 36343 926426 36993 926487
rect 0 925254 39573 926426
rect 0 913734 5847 925254
rect 19940 913734 39573 925254
rect 678027 922346 679077 951823
rect 679397 922346 680287 951823
rect 680607 922407 681257 952759
rect 681577 952143 717600 953079
rect 681577 922346 682467 951823
rect 682787 922346 683677 951823
rect 683997 922346 684647 951823
rect 684967 922600 685617 951823
rect 684968 922346 685617 922600
rect 685937 922346 686827 951823
rect 687147 922346 688947 951823
rect 689267 922346 690117 951823
rect 690437 922346 691287 951823
rect 691607 922346 696597 951823
rect 696917 943200 717600 952143
rect 712757 922600 717600 943200
rect 680607 922026 681257 922087
rect 696917 922026 717600 922600
rect 0 912574 39573 913734
rect 678027 920866 717600 922026
rect 0 912000 20683 912574
rect 36343 912513 36993 912574
rect 0 884800 4843 912000
rect 0 884226 20683 884800
rect 21003 884546 25993 912254
rect 26313 884546 27163 912254
rect 27483 884546 28333 912254
rect 28653 884546 30453 912254
rect 30773 884546 31663 912254
rect 31983 912000 32632 912254
rect 31983 884546 32633 912000
rect 32953 884546 33603 912254
rect 33923 884546 34813 912254
rect 35133 884546 36023 912254
rect 36343 884607 36993 912193
rect 37313 884546 38203 912254
rect 38523 884546 39573 912254
rect 678027 909346 697660 920866
rect 711753 909346 717600 920866
rect 678027 908174 717600 909346
rect 680607 908113 681257 908174
rect 32632 884226 32633 884546
rect 36343 884226 36993 884287
rect 0 883698 39573 884226
rect 0 870890 6491 883698
rect 19296 870890 39573 883698
rect 678027 878146 679077 907854
rect 679397 878146 680287 907854
rect 680607 878207 681257 907793
rect 681577 878146 682467 907854
rect 682787 878146 683677 907854
rect 683997 878146 684647 907854
rect 684968 907600 685617 907854
rect 684967 878400 685617 907600
rect 684968 878146 685617 878400
rect 685937 878146 686827 907854
rect 687147 878146 688947 907854
rect 689267 878146 690117 907854
rect 690437 878146 691287 907854
rect 691607 878146 696597 907854
rect 696917 907600 717600 908174
rect 712757 878400 717600 907600
rect 680607 877826 681257 877887
rect 696917 877826 717600 878400
rect 0 870374 39573 870890
rect 678027 876500 717600 877826
rect 0 869800 20683 870374
rect 32632 870054 32633 870374
rect 36343 870313 36993 870374
rect 0 842600 4843 869800
rect 0 842026 20683 842600
rect 21003 842346 25993 870054
rect 26313 842346 27163 870054
rect 27483 842346 28333 870054
rect 28653 842346 30453 870054
rect 30773 842346 31663 870054
rect 31983 842346 32633 870054
rect 32953 842346 33603 870054
rect 33923 842346 34813 870054
rect 35133 842346 36023 870054
rect 36343 842407 36993 869993
rect 37313 842346 38203 870054
rect 38523 842346 39573 870054
rect 678027 863320 698192 876500
rect 711322 863320 717600 876500
rect 678027 862974 717600 863320
rect 680607 862926 681257 862974
rect 32632 842026 32633 842346
rect 36343 842026 36993 842087
rect 0 841498 39573 842026
rect 0 828690 6491 841498
rect 19296 828690 39573 841498
rect 678027 833146 679077 862654
rect 679397 833146 680287 862654
rect 680607 833207 681257 862606
rect 681577 833146 682467 862654
rect 682787 833146 683677 862654
rect 683997 833146 684647 862654
rect 684968 862400 685617 862654
rect 684967 833146 685617 862400
rect 685937 833146 686827 862654
rect 687147 833146 688947 862654
rect 689267 833146 690117 862654
rect 690437 833146 691287 862654
rect 691607 833146 696597 862654
rect 696917 862400 717600 862974
rect 712757 833400 717600 862400
rect 680607 832826 681257 832887
rect 684967 832826 684968 833146
rect 696917 832826 717600 833400
rect 0 828174 39573 828690
rect 678027 832310 717600 832826
rect 0 827600 20683 828174
rect 32632 827854 32633 828174
rect 36343 828113 36993 828174
rect 0 800400 4843 827600
rect 0 799826 20683 800400
rect 21003 800146 25993 827854
rect 26313 800146 27163 827854
rect 27483 800146 28333 827854
rect 28653 800146 30453 827854
rect 30773 800146 31663 827854
rect 31983 800400 32633 827854
rect 31983 800146 32632 800400
rect 32953 800146 33603 827854
rect 33923 800146 34813 827854
rect 35133 800146 36023 827854
rect 36343 800194 36993 827793
rect 37313 800146 38203 827854
rect 38523 800146 39573 827854
rect 678027 819502 698304 832310
rect 711109 819502 717600 832310
rect 678027 818974 717600 819502
rect 680607 818913 681257 818974
rect 684967 818654 684968 818974
rect 36343 799826 36993 799874
rect 0 799480 39573 799826
rect 0 786300 6278 799480
rect 19408 786300 39573 799480
rect 678027 788946 679077 818654
rect 679397 788946 680287 818654
rect 680607 789007 681257 818593
rect 681577 788946 682467 818654
rect 682787 788946 683677 818654
rect 683997 788946 684647 818654
rect 684967 789200 685617 818654
rect 684968 788946 685617 789200
rect 685937 788946 686827 818654
rect 687147 788946 688947 818654
rect 689267 788946 690117 818654
rect 690437 788946 691287 818654
rect 691607 788946 696597 818654
rect 696917 818400 717600 818974
rect 712757 789200 717600 818400
rect 680607 788626 681257 788687
rect 696917 788626 717600 789200
rect 0 784974 39573 786300
rect 678027 787300 717600 788626
rect 0 784400 20683 784974
rect 36343 784913 36993 784974
rect 0 757200 4843 784400
rect 0 756626 20683 757200
rect 21003 756946 25993 784654
rect 26313 756946 27163 784654
rect 27483 756946 28333 784654
rect 28653 756946 30453 784654
rect 30773 756946 31663 784654
rect 31983 784400 32632 784654
rect 31983 757200 32633 784400
rect 31983 756946 32632 757200
rect 32953 756946 33603 784654
rect 33923 756946 34813 784654
rect 35133 756946 36023 784654
rect 36343 756994 36993 784593
rect 37313 756946 38203 784654
rect 38523 756946 39573 784654
rect 678027 774120 698192 787300
rect 711322 774120 717600 787300
rect 678027 773774 717600 774120
rect 680607 773726 681257 773774
rect 36343 756626 36993 756674
rect 0 756280 39573 756626
rect 0 743100 6278 756280
rect 19408 743100 39573 756280
rect 678027 743946 679077 773454
rect 679397 743946 680287 773454
rect 680607 744007 681257 773406
rect 681577 743946 682467 773454
rect 682787 743946 683677 773454
rect 683997 743946 684647 773454
rect 684968 773200 685617 773454
rect 684967 744200 685617 773200
rect 684968 743946 685617 744200
rect 685937 743946 686827 773454
rect 687147 743946 688947 773454
rect 689267 743946 690117 773454
rect 690437 743946 691287 773454
rect 691607 743946 696597 773454
rect 696917 773200 717600 773774
rect 712757 744200 717600 773200
rect 680607 743626 681257 743687
rect 696917 743626 717600 744200
rect 0 741774 39573 743100
rect 678027 742300 717600 743626
rect 0 741200 20683 741774
rect 36343 741713 36993 741774
rect 0 714000 4843 741200
rect 0 713426 20683 714000
rect 21003 713746 25993 741454
rect 26313 713746 27163 741454
rect 27483 713746 28333 741454
rect 28653 713746 30453 741454
rect 30773 713746 31663 741454
rect 31983 741200 32632 741454
rect 31983 714000 32633 741200
rect 31983 713746 32632 714000
rect 32953 713746 33603 741454
rect 33923 713746 34813 741454
rect 35133 713746 36023 741454
rect 36343 713794 36993 741393
rect 37313 713746 38203 741454
rect 38523 713746 39573 741454
rect 678027 729120 698192 742300
rect 711322 729120 717600 742300
rect 678027 728774 717600 729120
rect 680607 728726 681257 728774
rect 36343 713426 36993 713474
rect 0 713080 39573 713426
rect 0 699900 6278 713080
rect 19408 699900 39573 713080
rect 0 698574 39573 699900
rect 678027 698946 679077 728454
rect 679397 698946 680287 728454
rect 680607 699007 681257 728406
rect 681577 698946 682467 728454
rect 682787 698946 683677 728454
rect 683997 698946 684647 728454
rect 684968 728200 685617 728454
rect 684967 699200 685617 728200
rect 684968 698946 685617 699200
rect 685937 698946 686827 728454
rect 687147 698946 688947 728454
rect 689267 698946 690117 728454
rect 690437 698946 691287 728454
rect 691607 698946 696597 728454
rect 696917 728200 717600 728774
rect 712757 699200 717600 728200
rect 680607 698626 681257 698687
rect 696917 698626 717600 699200
rect 0 698000 20683 698574
rect 36343 698513 36993 698574
rect 0 670800 4843 698000
rect 0 670226 20683 670800
rect 21003 670546 25993 698254
rect 26313 670546 27163 698254
rect 27483 670546 28333 698254
rect 28653 670546 30453 698254
rect 30773 670546 31663 698254
rect 31983 698000 32632 698254
rect 31983 670800 32633 698000
rect 31983 670546 32632 670800
rect 32953 670546 33603 698254
rect 33923 670546 34813 698254
rect 35133 670546 36023 698254
rect 36343 670594 36993 698193
rect 37313 670546 38203 698254
rect 38523 670546 39573 698254
rect 678027 697300 717600 698626
rect 678027 684120 698192 697300
rect 711322 684120 717600 697300
rect 678027 683774 717600 684120
rect 680607 683726 681257 683774
rect 36343 670226 36993 670274
rect 0 669880 39573 670226
rect 0 656700 6278 669880
rect 19408 656700 39573 669880
rect 0 655374 39573 656700
rect 0 654800 20683 655374
rect 36343 655313 36993 655374
rect 0 627600 4843 654800
rect 0 627026 20683 627600
rect 21003 627346 25993 655054
rect 26313 627346 27163 655054
rect 27483 627346 28333 655054
rect 28653 627346 30453 655054
rect 30773 627346 31663 655054
rect 31983 654800 32632 655054
rect 31983 627600 32633 654800
rect 31983 627346 32632 627600
rect 32953 627346 33603 655054
rect 33923 627346 34813 655054
rect 35133 627346 36023 655054
rect 36343 627394 36993 654993
rect 37313 627346 38203 655054
rect 38523 627346 39573 655054
rect 678027 653746 679077 683454
rect 679397 653746 680287 683454
rect 680607 653807 681257 683406
rect 681577 653746 682467 683454
rect 682787 653746 683677 683454
rect 683997 653746 684647 683454
rect 684968 683200 685617 683454
rect 684967 654000 685617 683200
rect 684968 653746 685617 654000
rect 685937 653746 686827 683454
rect 687147 653746 688947 683454
rect 689267 653746 690117 683454
rect 690437 653746 691287 683454
rect 691607 653746 696597 683454
rect 696917 683200 717600 683774
rect 712757 654000 717600 683200
rect 680607 653426 681257 653487
rect 696917 653426 717600 654000
rect 678027 652100 717600 653426
rect 678027 638920 698192 652100
rect 711322 638920 717600 652100
rect 678027 638574 717600 638920
rect 680607 638526 681257 638574
rect 36343 627026 36993 627074
rect 0 626680 39573 627026
rect 0 613500 6278 626680
rect 19408 613500 39573 626680
rect 0 612174 39573 613500
rect 0 611600 20683 612174
rect 36343 612113 36993 612174
rect 0 584400 4843 611600
rect 0 583826 20683 584400
rect 21003 584146 25993 611854
rect 26313 584146 27163 611854
rect 27483 584146 28333 611854
rect 28653 584146 30453 611854
rect 30773 584146 31663 611854
rect 31983 611600 32632 611854
rect 31983 584400 32633 611600
rect 31983 584146 32632 584400
rect 32953 584146 33603 611854
rect 33923 584146 34813 611854
rect 35133 584146 36023 611854
rect 36343 584194 36993 611793
rect 37313 584146 38203 611854
rect 38523 584146 39573 611854
rect 678027 608746 679077 638254
rect 679397 608746 680287 638254
rect 680607 608807 681257 638206
rect 681577 608746 682467 638254
rect 682787 608746 683677 638254
rect 683997 608746 684647 638254
rect 684968 638000 685617 638254
rect 684967 609000 685617 638000
rect 684968 608746 685617 609000
rect 685937 608746 686827 638254
rect 687147 608746 688947 638254
rect 689267 608746 690117 638254
rect 690437 608746 691287 638254
rect 691607 608746 696597 638254
rect 696917 638000 717600 638574
rect 712757 609000 717600 638000
rect 680607 608426 681257 608487
rect 696917 608426 717600 609000
rect 678027 607100 717600 608426
rect 678027 593920 698192 607100
rect 711322 593920 717600 607100
rect 678027 593574 717600 593920
rect 680607 593526 681257 593574
rect 36343 583826 36993 583874
rect 0 583480 39573 583826
rect 0 570300 6278 583480
rect 19408 570300 39573 583480
rect 0 568974 39573 570300
rect 0 568400 20683 568974
rect 36343 568913 36993 568974
rect 0 541200 4843 568400
rect 0 540626 20683 541200
rect 21003 540946 25993 568654
rect 26313 540946 27163 568654
rect 27483 540946 28333 568654
rect 28653 540946 30453 568654
rect 30773 540946 31663 568654
rect 31983 568400 32632 568654
rect 31983 541200 32633 568400
rect 31983 540946 32632 541200
rect 32953 540946 33603 568654
rect 33923 540946 34813 568654
rect 35133 540946 36023 568654
rect 36343 540994 36993 568593
rect 37313 540946 38203 568654
rect 38523 540946 39573 568654
rect 678027 563546 679077 593254
rect 679397 563546 680287 593254
rect 680607 563607 681257 593206
rect 681577 563546 682467 593254
rect 682787 563546 683677 593254
rect 683997 563546 684647 593254
rect 684968 593000 685617 593254
rect 684967 563800 685617 593000
rect 684968 563546 685617 563800
rect 685937 563546 686827 593254
rect 687147 563546 688947 593254
rect 689267 563546 690117 593254
rect 690437 563546 691287 593254
rect 691607 563546 696597 593254
rect 696917 593000 717600 593574
rect 712757 563800 717600 593000
rect 680607 563226 681257 563287
rect 696917 563226 717600 563800
rect 678027 561900 717600 563226
rect 678027 548720 698192 561900
rect 711322 548720 717600 561900
rect 678027 548374 717600 548720
rect 680607 548326 681257 548374
rect 36343 540626 36993 540674
rect 0 540280 39573 540626
rect 0 527100 6278 540280
rect 19408 527100 39573 540280
rect 0 525774 39573 527100
rect 0 525200 20683 525774
rect 36343 525713 36993 525774
rect 0 498000 4843 525200
rect 0 497426 20683 498000
rect 21003 497746 25993 525454
rect 26313 497746 27163 525454
rect 27483 497746 28333 525454
rect 28653 497746 30453 525454
rect 30773 497746 31663 525454
rect 31983 525200 32632 525454
rect 31983 497746 32633 525200
rect 32953 497746 33603 525454
rect 33923 497746 34813 525454
rect 35133 497746 36023 525454
rect 36343 497807 36993 525393
rect 37313 497746 38203 525454
rect 38523 497746 39573 525454
rect 678027 518546 679077 548054
rect 679397 518546 680287 548054
rect 680607 518607 681257 548006
rect 681577 518546 682467 548054
rect 682787 518546 683677 548054
rect 683997 518546 684647 548054
rect 684968 547800 685617 548054
rect 684967 518546 685617 547800
rect 685937 518546 686827 548054
rect 687147 518546 688947 548054
rect 689267 518546 690117 548054
rect 690437 518546 691287 548054
rect 691607 518546 696597 548054
rect 696917 547800 717600 548374
rect 712757 518800 717600 547800
rect 680607 518226 681257 518287
rect 684967 518226 684968 518546
rect 696917 518226 717600 518800
rect 678027 517710 717600 518226
rect 678027 504902 698304 517710
rect 711109 504902 717600 517710
rect 678027 504374 717600 504902
rect 680607 504313 681257 504374
rect 684967 504054 684968 504374
rect 32632 497426 32633 497746
rect 36343 497426 36993 497487
rect 0 496898 39573 497426
rect 0 484090 6491 496898
rect 19296 484090 39573 496898
rect 0 483574 39573 484090
rect 0 483000 20683 483574
rect 32632 483254 32633 483574
rect 36343 483513 36993 483574
rect 0 455800 4843 483000
rect 0 455226 20683 455800
rect 21003 455546 25993 483254
rect 26313 455546 27163 483254
rect 27483 455546 28333 483254
rect 28653 455546 30453 483254
rect 30773 455546 31663 483254
rect 31983 455800 32633 483254
rect 31983 455546 32632 455800
rect 32953 455546 33603 483254
rect 33923 455546 34813 483254
rect 35133 455546 36023 483254
rect 36343 455607 36993 483193
rect 37313 455546 38203 483254
rect 38523 455546 39573 483254
rect 678027 474546 679077 504054
rect 679397 474546 680287 504054
rect 680607 474607 681257 503993
rect 681577 474546 682467 504054
rect 682787 474546 683677 504054
rect 683997 474546 684647 504054
rect 684967 474800 685617 504054
rect 684968 474546 685617 474800
rect 685937 474546 686827 504054
rect 687147 474546 688947 504054
rect 689267 474546 690117 504054
rect 690437 474546 691287 504054
rect 691607 474546 696597 504054
rect 696917 503800 717600 504374
rect 712757 474800 717600 503800
rect 680607 474226 681257 474287
rect 696917 474226 717600 474800
rect 678027 473066 717600 474226
rect 678027 461546 697660 473066
rect 711753 461546 717600 473066
rect 678027 460374 717600 461546
rect 680607 460313 681257 460374
rect 36343 455226 36993 455287
rect 0 454054 39573 455226
rect 0 442534 5847 454054
rect 19940 442534 39573 454054
rect 0 441374 39573 442534
rect 0 440800 20683 441374
rect 36343 441313 36993 441374
rect 0 413600 4843 440800
rect 0 413026 20683 413600
rect 21003 413346 25993 441054
rect 26313 413346 27163 441054
rect 27483 413346 28333 441054
rect 28653 413346 30453 441054
rect 30773 413346 31663 441054
rect 31983 440800 32632 441054
rect 31983 413600 32633 440800
rect 31983 413346 32632 413600
rect 32953 413346 33603 441054
rect 33923 413346 34813 441054
rect 35133 413346 36023 441054
rect 36343 413394 36993 440993
rect 37313 413346 38203 441054
rect 38523 413346 39573 441054
rect 678027 430346 679077 460054
rect 679397 430346 680287 460054
rect 680607 430407 681257 459993
rect 681577 430346 682467 460054
rect 682787 430346 683677 460054
rect 683997 430346 684647 460054
rect 684968 459800 685617 460054
rect 684967 430346 685617 459800
rect 685937 430346 686827 460054
rect 687147 430346 688947 460054
rect 689267 430346 690117 460054
rect 690437 430346 691287 460054
rect 691607 430346 696597 460054
rect 696917 459800 717600 460374
rect 712757 430600 717600 459800
rect 680607 430026 681257 430087
rect 684967 430026 684968 430346
rect 696917 430026 717600 430600
rect 678027 429510 717600 430026
rect 678027 416702 698304 429510
rect 711109 416702 717600 429510
rect 678027 416174 717600 416702
rect 680607 416113 681257 416174
rect 684967 415854 684968 416174
rect 36343 413026 36993 413074
rect 0 412680 39573 413026
rect 0 399500 6278 412680
rect 19408 399500 39573 412680
rect 0 398174 39573 399500
rect 0 397600 20683 398174
rect 36343 398113 36993 398174
rect 0 370400 4843 397600
rect 0 369826 20683 370400
rect 21003 370146 25993 397854
rect 26313 370146 27163 397854
rect 27483 370146 28333 397854
rect 28653 370146 30453 397854
rect 30773 370146 31663 397854
rect 31983 397600 32632 397854
rect 31983 370400 32633 397600
rect 31983 370146 32632 370400
rect 32953 370146 33603 397854
rect 33923 370146 34813 397854
rect 35133 370146 36023 397854
rect 36343 370194 36993 397793
rect 37313 370146 38203 397854
rect 38523 370146 39573 397854
rect 678027 386346 679077 415854
rect 679397 386346 680287 415854
rect 680607 386407 681257 415793
rect 681577 386346 682467 415854
rect 682787 386346 683677 415854
rect 683997 386346 684647 415854
rect 684967 386600 685617 415854
rect 684968 386346 685617 386600
rect 685937 386346 686827 415854
rect 687147 386346 688947 415854
rect 689267 386346 690117 415854
rect 690437 386346 691287 415854
rect 691607 386346 696597 415854
rect 696917 415600 717600 416174
rect 712757 386600 717600 415600
rect 680607 386026 681257 386087
rect 696917 386026 717600 386600
rect 678027 384700 717600 386026
rect 678027 371520 698192 384700
rect 711322 371520 717600 384700
rect 678027 371174 717600 371520
rect 680607 371126 681257 371174
rect 36343 369826 36993 369874
rect 0 369480 39573 369826
rect 0 356300 6278 369480
rect 19408 356300 39573 369480
rect 0 354974 39573 356300
rect 0 354400 20683 354974
rect 36343 354913 36993 354974
rect 0 327200 4843 354400
rect 0 326626 20683 327200
rect 21003 326946 25993 354654
rect 26313 326946 27163 354654
rect 27483 326946 28333 354654
rect 28653 326946 30453 354654
rect 30773 326946 31663 354654
rect 31983 354400 32632 354654
rect 31983 327200 32633 354400
rect 31983 326946 32632 327200
rect 32953 326946 33603 354654
rect 33923 326946 34813 354654
rect 35133 326946 36023 354654
rect 36343 326994 36993 354593
rect 37313 326946 38203 354654
rect 38523 326946 39573 354654
rect 678027 341146 679077 370854
rect 679397 341146 680287 370854
rect 680607 341207 681257 370806
rect 681577 341146 682467 370854
rect 682787 341146 683677 370854
rect 683997 341146 684647 370854
rect 684968 370600 685617 370854
rect 684967 341400 685617 370600
rect 684968 341146 685617 341400
rect 685937 341146 686827 370854
rect 687147 341146 688947 370854
rect 689267 341146 690117 370854
rect 690437 341146 691287 370854
rect 691607 341146 696597 370854
rect 696917 370600 717600 371174
rect 712757 341400 717600 370600
rect 680607 340826 681257 340887
rect 696917 340826 717600 341400
rect 678027 339500 717600 340826
rect 36343 326626 36993 326674
rect 0 326280 39573 326626
rect 0 313100 6278 326280
rect 19408 313100 39573 326280
rect 678027 326320 698192 339500
rect 711322 326320 717600 339500
rect 678027 325974 717600 326320
rect 680607 325926 681257 325974
rect 0 311774 39573 313100
rect 0 311200 20683 311774
rect 36343 311713 36993 311774
rect 0 284000 4843 311200
rect 0 283426 20683 284000
rect 21003 283746 25993 311454
rect 26313 283746 27163 311454
rect 27483 283746 28333 311454
rect 28653 283746 30453 311454
rect 30773 283746 31663 311454
rect 31983 311200 32632 311454
rect 31983 284000 32633 311200
rect 31983 283746 32632 284000
rect 32953 283746 33603 311454
rect 33923 283746 34813 311454
rect 35133 283746 36023 311454
rect 36343 283794 36993 311393
rect 37313 283746 38203 311454
rect 38523 283746 39573 311454
rect 678027 296146 679077 325654
rect 679397 296146 680287 325654
rect 680607 296207 681257 325606
rect 681577 296146 682467 325654
rect 682787 296146 683677 325654
rect 683997 296146 684647 325654
rect 684968 325400 685617 325654
rect 684967 296400 685617 325400
rect 684968 296146 685617 296400
rect 685937 296146 686827 325654
rect 687147 296146 688947 325654
rect 689267 296146 690117 325654
rect 690437 296146 691287 325654
rect 691607 296146 696597 325654
rect 696917 325400 717600 325974
rect 712757 296400 717600 325400
rect 680607 295826 681257 295887
rect 696917 295826 717600 296400
rect 678027 294500 717600 295826
rect 36343 283426 36993 283474
rect 0 283080 39573 283426
rect 0 269900 6278 283080
rect 19408 269900 39573 283080
rect 678027 281320 698192 294500
rect 711322 281320 717600 294500
rect 678027 280974 717600 281320
rect 680607 280926 681257 280974
rect 0 268574 39573 269900
rect 0 268000 20683 268574
rect 36343 268513 36993 268574
rect 0 240800 4843 268000
rect 0 240226 20683 240800
rect 21003 240546 25993 268254
rect 26313 240546 27163 268254
rect 27483 240546 28333 268254
rect 28653 240546 30453 268254
rect 30773 240546 31663 268254
rect 31983 268000 32632 268254
rect 31983 240800 32633 268000
rect 31983 240546 32632 240800
rect 32953 240546 33603 268254
rect 33923 240546 34813 268254
rect 35133 240546 36023 268254
rect 36343 240594 36993 268193
rect 37313 240546 38203 268254
rect 38523 240546 39573 268254
rect 678027 251146 679077 280654
rect 679397 251146 680287 280654
rect 680607 251207 681257 280606
rect 681577 251146 682467 280654
rect 682787 251146 683677 280654
rect 683997 251146 684647 280654
rect 684968 280400 685617 280654
rect 684967 251400 685617 280400
rect 684968 251146 685617 251400
rect 685937 251146 686827 280654
rect 687147 251146 688947 280654
rect 689267 251146 690117 280654
rect 690437 251146 691287 280654
rect 691607 251146 696597 280654
rect 696917 280400 717600 280974
rect 712757 251400 717600 280400
rect 680607 250826 681257 250887
rect 696917 250826 717600 251400
rect 678027 249500 717600 250826
rect 36343 240226 36993 240274
rect 0 239880 39573 240226
rect 0 226700 6278 239880
rect 19408 226700 39573 239880
rect 678027 236320 698192 249500
rect 711322 236320 717600 249500
rect 678027 235974 717600 236320
rect 680607 235926 681257 235974
rect 0 225374 39573 226700
rect 0 224800 20683 225374
rect 36343 225313 36993 225374
rect 0 197600 4843 224800
rect 0 197026 20683 197600
rect 21003 197346 25993 225054
rect 26313 197346 27163 225054
rect 27483 197346 28333 225054
rect 28653 197346 30453 225054
rect 30773 197346 31663 225054
rect 31983 224800 32632 225054
rect 31983 197600 32633 224800
rect 31983 197346 32632 197600
rect 32953 197346 33603 225054
rect 33923 197346 34813 225054
rect 35133 197346 36023 225054
rect 36343 197394 36993 224993
rect 37313 197346 38203 225054
rect 38523 197346 39573 225054
rect 678027 205946 679077 235654
rect 679397 205946 680287 235654
rect 680607 206007 681257 235606
rect 681577 205946 682467 235654
rect 682787 205946 683677 235654
rect 683997 205946 684647 235654
rect 684968 235400 685617 235654
rect 684967 206200 685617 235400
rect 684968 205946 685617 206200
rect 685937 205946 686827 235654
rect 687147 205946 688947 235654
rect 689267 205946 690117 235654
rect 690437 205946 691287 235654
rect 691607 205946 696597 235654
rect 696917 235400 717600 235974
rect 712757 206200 717600 235400
rect 680607 205626 681257 205687
rect 696917 205626 717600 206200
rect 678027 204300 717600 205626
rect 36343 197026 36993 197074
rect 0 196680 39573 197026
rect 0 183500 6278 196680
rect 19408 183500 39573 196680
rect 678027 191120 698192 204300
rect 711322 191120 717600 204300
rect 678027 190774 717600 191120
rect 680607 190726 681257 190774
rect 0 182174 39573 183500
rect 0 181600 20683 182174
rect 36343 182113 36993 182174
rect 0 125200 4843 181600
rect 0 124626 20683 125200
rect 21003 124946 25993 181854
rect 26313 124946 27163 181854
rect 27483 124946 28333 181854
rect 28653 126200 30453 181854
rect 30773 127200 31663 181854
rect 31983 181600 32632 181854
rect 31983 126200 32633 181600
rect 28653 124946 30453 125200
rect 30773 124946 31663 126200
rect 31983 124946 32633 125200
rect 32953 124946 33603 181854
rect 33923 124946 34813 181854
rect 35133 124946 36023 181854
rect 36343 126200 36993 181793
rect 37313 127200 38203 181854
rect 36343 125007 36993 125200
rect 37313 124946 38203 126200
rect 38523 124946 39573 181854
rect 678027 160946 679077 190454
rect 679397 160946 680287 190454
rect 680607 161007 681257 190406
rect 681577 160946 682467 190454
rect 682787 160946 683677 190454
rect 683997 160946 684647 190454
rect 684968 190200 685617 190454
rect 684967 161200 685617 190200
rect 684968 160946 685617 161200
rect 685937 160946 686827 190454
rect 687147 160946 688947 190454
rect 689267 160946 690117 190454
rect 690437 160946 691287 190454
rect 691607 160946 696597 190454
rect 696917 190200 717600 190774
rect 712757 161200 717600 190200
rect 680607 160626 681257 160687
rect 696917 160626 717600 161200
rect 678027 159300 717600 160626
rect 678027 146120 698192 159300
rect 711322 146120 717600 159300
rect 678027 145774 717600 146120
rect 680607 145726 681257 145774
rect 32632 124626 32633 124946
rect 36343 124626 36993 124687
rect 0 124098 39573 124626
rect 0 111290 6491 124098
rect 19296 111290 39573 124098
rect 678027 115746 679077 145454
rect 679397 115746 680287 145454
rect 680607 115807 681257 145406
rect 681577 115746 682467 145454
rect 682787 115746 683677 145454
rect 683997 115746 684647 145454
rect 684968 145200 685617 145454
rect 684967 116000 685617 145200
rect 684968 115746 685617 116000
rect 685937 115746 686827 145454
rect 687147 115746 688947 145454
rect 689267 115746 690117 145454
rect 690437 115746 691287 145454
rect 691607 115746 696597 145454
rect 696917 145200 717600 145774
rect 712757 116000 717600 145200
rect 680607 115426 681257 115487
rect 696917 115426 717600 116000
rect 0 110774 39573 111290
rect 678027 114100 717600 115426
rect 0 110200 20683 110774
rect 32632 110454 32633 110774
rect 36343 110713 36993 110774
rect 0 83000 4843 110200
rect 0 82426 20683 83000
rect 21003 82746 25993 110454
rect 26313 82746 27163 110454
rect 27483 82746 28333 110454
rect 28653 82746 30453 110454
rect 30773 82746 31663 110454
rect 31983 82746 32633 110454
rect 32953 82746 33603 110454
rect 33923 82746 34813 110454
rect 35133 82746 36023 110454
rect 36343 82807 36993 110393
rect 37313 82746 38203 110454
rect 38523 82746 39573 110454
rect 678027 100920 698192 114100
rect 711322 100920 717600 114100
rect 678027 100574 717600 100920
rect 680607 100526 681257 100574
rect 32632 82426 32633 82746
rect 36343 82426 36993 82487
rect 0 81254 39573 82426
rect 0 69734 5847 81254
rect 19940 69734 39573 81254
rect 0 68574 39573 69734
rect 0 68000 20683 68574
rect 32632 68254 32633 68574
rect 36343 68513 36993 68574
rect 0 40800 4843 68000
rect 0 40109 20683 40800
rect 21003 40429 25993 68254
rect 26313 40546 27163 68254
rect 27483 40546 28333 68254
rect 26313 40109 28333 40226
rect 0 35049 28333 40109
rect 28653 35369 30453 68254
rect 30773 40546 31663 68254
rect 31983 40800 32633 68254
rect 31983 40546 32632 40800
rect 32953 40546 33603 68254
rect 33923 40546 34813 68254
rect 35133 40546 36023 68254
rect 36343 40549 36993 68193
rect 37313 40546 38203 68254
rect 38523 40546 39573 68254
rect 36343 40226 36993 40229
rect 39893 40226 40000 40800
rect 30773 39893 40000 40226
rect 676800 39893 677707 40000
rect 30773 38523 39210 39893
rect 39530 38523 79054 39573
rect 30773 36993 38923 38523
rect 47400 38203 71400 38523
rect 39243 37313 79054 38203
rect 79374 36993 93226 39573
rect 93546 38523 132854 39573
rect 101200 38203 125200 38523
rect 93546 37313 132854 38203
rect 133174 36993 147026 39573
rect 147346 38523 186654 39573
rect 155000 38203 179000 38523
rect 147346 37313 186654 38203
rect 186974 36993 201826 39573
rect 202146 38523 241454 39573
rect 209800 38203 233800 38523
rect 202146 37313 241454 38203
rect 241774 36993 255626 39573
rect 255946 38523 295254 39573
rect 263600 38203 287600 38523
rect 255946 37313 295254 38203
rect 295574 36993 310426 39573
rect 310746 38523 350054 39573
rect 318400 38203 342400 38523
rect 310746 37313 350054 38203
rect 350374 36993 365226 39573
rect 365546 38523 404854 39573
rect 373200 38203 397200 38523
rect 365546 37313 404854 38203
rect 405174 36993 420026 39573
rect 420346 38523 459654 39573
rect 428000 38203 452000 38523
rect 420346 37313 459654 38203
rect 459974 36993 474826 39573
rect 475146 38523 514454 39573
rect 482800 38203 506800 38523
rect 475146 37313 514454 38203
rect 514774 36993 529626 39573
rect 529946 38523 569254 39573
rect 537600 38203 561600 38523
rect 529946 37313 569254 38203
rect 569574 36993 583426 39573
rect 583746 38523 623054 39573
rect 591400 38203 615400 38523
rect 583746 37313 623054 38203
rect 623374 36993 637226 39573
rect 637546 38523 677054 39573
rect 677374 39210 677707 39893
rect 678027 39530 679077 100254
rect 679397 71000 680287 100254
rect 680607 70000 681257 100206
rect 679397 39243 680287 70000
rect 680607 39706 681257 69000
rect 681577 39695 682467 100254
rect 682787 39680 683677 100254
rect 683997 39723 684647 100254
rect 684968 100000 685617 100254
rect 684967 70000 685617 100000
rect 685937 71000 686827 100254
rect 687147 70000 688947 100254
rect 684967 39733 685617 69000
rect 685937 39705 686827 70000
rect 684967 39403 685617 39413
rect 680607 39375 681257 39386
rect 683997 39385 685617 39403
rect 680607 39360 682467 39375
rect 683997 39360 686827 39385
rect 677374 38923 679077 39210
rect 680607 38923 686827 39360
rect 645200 38203 669200 38523
rect 637546 37313 677054 38203
rect 677374 36993 686827 38923
rect 30773 36343 39386 36993
rect 39706 36343 78993 36993
rect 79313 36343 93287 36993
rect 93607 36343 132793 36993
rect 133113 36343 147087 36993
rect 147407 36343 186606 36993
rect 186926 36343 201887 36993
rect 202207 36343 241393 36993
rect 241713 36343 255687 36993
rect 256007 36343 295206 36993
rect 295526 36343 310487 36993
rect 310807 36343 350006 36993
rect 350326 36343 365287 36993
rect 365607 36343 404806 36993
rect 405126 36343 420087 36993
rect 420407 36343 459606 36993
rect 459926 36343 474887 36993
rect 475207 36343 514406 36993
rect 514726 36343 529687 36993
rect 530007 36343 569193 36993
rect 569513 36343 583487 36993
rect 583807 36343 622993 36993
rect 623313 36343 637287 36993
rect 637607 36343 677051 36993
rect 677371 36343 686827 36993
rect 30773 35133 39375 36343
rect 39695 35133 79054 36023
rect 30773 35049 39360 35133
rect 0 33603 39360 35049
rect 39680 33923 79054 34813
rect 0 32633 39403 33603
rect 39723 32953 79054 33603
rect 79374 32633 93226 36343
rect 93546 35133 132854 36023
rect 93546 33923 132854 34813
rect 93546 32953 132854 33603
rect 0 31983 39413 32633
rect 39733 32632 132600 32633
rect 39733 31983 79054 32632
rect 0 30773 39385 31983
rect 39705 30773 79054 31663
rect 0 28333 35049 30773
rect 35369 28653 79054 30453
rect 0 27163 39355 28333
rect 39675 27483 79054 28333
rect 0 26313 39384 27163
rect 39704 26313 79054 27163
rect 0 20683 39151 26313
rect 39471 21003 79054 25993
rect 79374 20683 93226 32632
rect 93546 31983 132854 32632
rect 93546 30773 132854 31663
rect 93546 28653 132854 30453
rect 93546 27483 132854 28333
rect 93546 26313 132854 27163
rect 93546 21003 132854 25993
rect 133174 20683 147026 36343
rect 147346 35133 186654 36023
rect 147346 33923 186654 34813
rect 147346 32953 186654 33603
rect 147600 32632 186400 32633
rect 147346 31983 186654 32632
rect 147346 30773 186654 31663
rect 147346 28653 186654 30453
rect 147346 27483 186654 28333
rect 147346 26313 186654 27163
rect 147346 21003 186654 25993
rect 186974 20683 201826 36343
rect 202146 35133 241454 36023
rect 202146 33923 241454 34813
rect 202146 32953 241454 33603
rect 241774 32633 255626 36343
rect 255946 35133 295254 36023
rect 255946 33923 295254 34813
rect 255946 32953 295254 33603
rect 202400 32632 295000 32633
rect 202146 31983 241454 32632
rect 202146 30773 241454 31663
rect 202146 28653 241454 30453
rect 202146 27483 241454 28333
rect 202146 26313 241454 27163
rect 202146 21003 241454 25993
rect 241774 20683 255626 32632
rect 255946 31983 295254 32632
rect 255946 30773 295254 31663
rect 255946 28653 295254 30453
rect 255946 27483 295254 28333
rect 255946 26313 295254 27163
rect 255946 21003 295254 25993
rect 295574 20683 310426 36343
rect 310746 35133 350054 36023
rect 310746 33923 350054 34813
rect 310746 32953 350054 33603
rect 311000 32632 349800 32633
rect 310746 31983 350054 32632
rect 310746 30773 350054 31663
rect 310746 28653 350054 30453
rect 310746 27483 350054 28333
rect 310746 26313 350054 27163
rect 310746 21003 350054 25993
rect 350374 20683 365226 36343
rect 365546 35133 404854 36023
rect 365546 33923 404854 34813
rect 365546 32953 404854 33603
rect 365800 32632 404600 32633
rect 365546 31983 404854 32632
rect 365546 30773 404854 31663
rect 365546 28653 404854 30453
rect 365546 27483 404854 28333
rect 365546 26313 404854 27163
rect 365546 21003 404854 25993
rect 405174 20683 420026 36343
rect 420346 35133 459654 36023
rect 420346 33923 459654 34813
rect 420346 32953 459654 33603
rect 420600 32632 459400 32633
rect 420346 31983 459654 32632
rect 420346 30773 459654 31663
rect 420346 28653 459654 30453
rect 420346 27483 459654 28333
rect 420346 26313 459654 27163
rect 420346 21003 459654 25993
rect 459974 20683 474826 36343
rect 475146 35133 514454 36023
rect 475146 33923 514454 34813
rect 475146 32953 514454 33603
rect 475400 32632 514200 32633
rect 475146 31983 514454 32632
rect 475146 30773 514454 31663
rect 475146 28653 514454 30453
rect 475146 27483 514454 28333
rect 475146 26313 514454 27163
rect 475146 21003 514454 25993
rect 514774 20683 529626 36343
rect 529946 35133 569254 36023
rect 529946 33923 569254 34813
rect 529946 32953 569254 33603
rect 569574 32633 583426 36343
rect 583746 35133 623054 36023
rect 583746 33923 623054 34813
rect 583746 32953 623054 33603
rect 623374 32633 637226 36343
rect 637546 35133 677054 36023
rect 677374 35049 686827 36343
rect 687147 35369 688947 69000
rect 689267 39675 690117 100254
rect 690437 39704 691287 100254
rect 691607 39471 696597 100254
rect 696917 100000 717600 100574
rect 712757 40000 717600 100000
rect 690437 39355 691287 39384
rect 689267 39151 691287 39355
rect 696917 39151 717600 40000
rect 689267 35049 717600 39151
rect 637546 33923 677054 34813
rect 637546 32953 677054 33603
rect 530200 32632 676800 32633
rect 529946 31983 569254 32632
rect 529946 30773 569254 31663
rect 529946 28653 569254 30453
rect 529946 27483 569254 28333
rect 529946 26313 569254 27163
rect 529946 21003 569254 25993
rect 569574 20683 583426 32632
rect 583746 31983 623054 32632
rect 583746 30773 623054 31663
rect 583746 28653 623054 30453
rect 583746 27483 623054 28333
rect 583746 26313 623054 27163
rect 583746 21003 623054 25993
rect 623374 20683 637226 32632
rect 637546 31983 677054 32632
rect 637546 30773 677054 31663
rect 677374 30773 717600 35049
rect 637546 28653 682231 30453
rect 682551 28333 717600 30773
rect 637546 27483 677054 28333
rect 637546 26313 677054 27163
rect 677374 26313 717600 28333
rect 637546 21003 677171 25993
rect 677491 20683 717600 26313
rect 0 4843 40000 20683
rect 78800 19296 93800 20683
rect 78800 6491 79902 19296
rect 92710 6491 93800 19296
rect 78800 4843 93800 6491
rect 132600 18629 147600 20683
rect 132600 6823 136393 18629
rect 144470 6823 147600 18629
rect 132600 5163 147600 6823
rect 186400 19408 202400 20683
rect 186400 6278 187320 19408
rect 200500 6278 202400 19408
rect 0 0 132854 4843
rect 133174 0 147026 5163
rect 186400 4843 202400 6278
rect 241200 19940 256200 20683
rect 241200 5847 242946 19940
rect 254466 5847 256200 19940
rect 241200 4843 256200 5847
rect 295000 19408 311000 20683
rect 295000 6278 295920 19408
rect 309100 6278 311000 19408
rect 295000 4843 311000 6278
rect 349800 19408 365800 20683
rect 349800 6278 350720 19408
rect 363900 6278 365800 19408
rect 349800 4843 365800 6278
rect 404600 19408 420600 20683
rect 404600 6278 405520 19408
rect 418700 6278 420600 19408
rect 404600 4843 420600 6278
rect 459400 19408 475400 20683
rect 459400 6278 460320 19408
rect 473500 6278 475400 19408
rect 459400 4843 475400 6278
rect 514200 19408 530200 20683
rect 514200 6278 515120 19408
rect 528300 6278 530200 19408
rect 514200 4843 530200 6278
rect 569000 19296 584000 20683
rect 569000 6491 570102 19296
rect 582910 6491 584000 19296
rect 569000 4843 584000 6491
rect 622800 19296 637800 20683
rect 622800 6491 623902 19296
rect 636710 6491 637800 19296
rect 622800 4843 637800 6491
rect 676800 4843 717600 20683
rect 147346 0 717600 4843
<< labels >>
rlabel metal5 s 187640 6598 200180 19088 6 clock
port 1 nsew signal input
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 2 nsew signal output
rlabel metal2 s 194043 41713 194099 42193 6 por
port 3 nsew signal input
rlabel metal5 s 351040 6598 363580 19088 6 flash_clk
port 4 nsew signal output
rlabel metal2 s 361767 41713 361823 42193 6 flash_clk_core
port 5 nsew signal input
rlabel metal2 s 357443 41713 357499 42193 6 flash_clk_ieb_core
port 6 nsew signal input
rlabel metal2 s 364895 41713 364951 42193 6 flash_clk_oeb_core
port 7 nsew signal input
rlabel metal5 s 296240 6598 308780 19088 6 flash_csb
port 8 nsew signal output
rlabel metal2 s 306967 41713 307023 42193 6 flash_csb_core
port 9 nsew signal input
rlabel metal2 s 302643 41713 302699 42193 6 flash_csb_ieb_core
port 10 nsew signal input
rlabel metal2 s 310095 41713 310151 42193 6 flash_csb_oeb_core
port 11 nsew signal input
rlabel metal5 s 405840 6598 418380 19088 6 flash_io0
port 12 nsew signal bidirectional
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 13 nsew signal output
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 14 nsew signal input
rlabel metal2 s 415371 41713 415427 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415216 41754 415268 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415216 41806 415427 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412364 41754 412416 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41713 412299 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41806 412416 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409328 41754 409380 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41713 409263 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41806 409380 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415228 41818 415427 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41818 412404 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41818 409368 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415371 41834 415427 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41834 412299 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41834 409263 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 415216 41760 415268 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 412364 41760 412416 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 409328 41760 409380 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 415210 41760 415274 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 412358 41760 412422 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41760 409386 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41772 415274 41800 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 415210 41800 415274 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 412358 41800 412422 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41800 409386 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal3 s 419717 44371 419783 44374 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 411069 44371 411135 44374 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 411069 44374 419783 44434 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 419717 44434 419783 44437 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 411069 44434 411135 44437 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel via2 s 419722 44376 419778 44432 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel via2 s 411074 44376 411130 44432 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419695 41713 419751 41820 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411047 41713 411103 41820 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419695 41820 419764 42193 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411047 41820 411116 42193 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419736 42193 419764 44367 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411088 42193 411116 44367 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419722 44367 419778 44441 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411074 44367 411130 44441 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal5 s 460640 6598 473180 19088 6 flash_io1
port 17 nsew signal bidirectional
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 18 nsew signal output
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 19 nsew signal input
rlabel metal2 s 470171 41713 470227 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470048 41754 470100 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470048 41806 470227 41818 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467196 41754 467248 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41713 467099 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41806 467248 41818 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464160 41754 464212 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41713 464063 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41806 464212 41818 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470060 41818 470227 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41818 467236 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41818 464200 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470171 41834 470227 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41834 467099 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41834 464063 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 470048 41760 470100 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 467196 41760 467248 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 464160 41760 464212 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 470042 41760 470106 41772 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 467190 41760 467254 41772 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41760 464218 41772 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41772 470106 41800 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 470042 41800 470106 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 467190 41800 467254 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41800 464218 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal3 s 474457 44371 474523 44374 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44371 465875 44374 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44374 474523 44434 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 474457 44434 474523 44437 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44434 465875 44437 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel via2 s 474462 44376 474518 44432 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel via2 s 465814 44376 465870 44432 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474495 41713 474551 41806 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465847 41713 465903 41806 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474476 41806 474551 42193 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465828 41806 465903 42193 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474476 42193 474504 44367 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465828 42193 465856 44367 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474462 44367 474518 44441 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465814 44367 465870 44441 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal5 s 515440 6598 527980 19088 6 gpio
port 22 nsew signal bidirectional
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 23 nsew signal output
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 24 nsew signal input
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 25 nsew signal input
rlabel metal3 s 524965 44235 525031 44238 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44235 518867 44238 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44238 525031 44298 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 524965 44298 525031 44301 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44298 518867 44301 6 gpio_mode1_core
port 26 nsew signal input
rlabel via2 s 524970 44240 525026 44296 6 gpio_mode1_core
port 26 nsew signal input
rlabel via2 s 518806 44240 518862 44296 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524971 41713 525027 42193 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518807 41713 518863 42193 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524984 42193 525012 44231 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518820 42193 518848 44231 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524970 44231 525026 44305 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518806 44231 518862 44305 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 27 nsew signal input
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 28 nsew signal input
rlabel metal5 s 6167 70054 19620 80934 6 vccd_pad
port 29 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda_pad
port 30 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio_pad
port 31 nsew signal bidirectional
rlabel metal5 s 6811 871210 18976 883378 6 vddio_pad2
port 32 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa_pad
port 33 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19620 6 vssd_pad
port 34 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio_pad
port 35 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_pad2
port 36 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113780 6 mprj_io[0]
port 37 nsew signal bidirectional
rlabel metal2 s 675407 105803 675887 105859 6 mprj_io_analog_en[0]
port 38 nsew signal input
rlabel metal2 s 675407 107091 675887 107147 6 mprj_io_analog_pol[0]
port 39 nsew signal input
rlabel metal2 s 675407 110127 675887 110183 6 mprj_io_analog_sel[0]
port 40 nsew signal input
rlabel metal2 s 675407 106447 675887 106503 6 mprj_io_dm[0]
port 41 nsew signal input
rlabel metal2 s 675407 104607 675887 104663 6 mprj_io_dm[1]
port 42 nsew signal input
rlabel metal2 s 675407 110771 675887 110827 6 mprj_io_dm[2]
port 43 nsew signal input
rlabel metal2 s 675407 111415 675887 111471 6 mprj_io_holdover[0]
port 44 nsew signal input
rlabel metal2 s 675407 114451 675887 114507 6 mprj_io_ib_mode_sel[0]
port 45 nsew signal input
rlabel metal2 s 675407 107643 675887 107699 6 mprj_io_inp_dis[0]
port 46 nsew signal input
rlabel metal2 s 675407 115095 675887 115151 6 mprj_io_oeb[0]
port 47 nsew signal input
rlabel metal2 s 675407 111967 675887 112023 6 mprj_io_out[0]
port 48 nsew signal input
rlabel metal2 s 675407 102767 675887 102823 6 mprj_io_slow_sel[0]
port 49 nsew signal input
rlabel metal2 s 675407 113807 675887 113863 6 mprj_io_vtrip_sel[0]
port 50 nsew signal input
rlabel metal2 s 675407 100927 675887 100983 6 mprj_io_in[0]
port 51 nsew signal output
rlabel metal2 s 675407 115647 675887 115703 6 mprj_io_in_3v3[0]
port 52 nsew signal output
rlabel metal2 s 675407 686611 675887 686667 6 mprj_gpio_analog[3]
port 53 nsew signal bidirectional
rlabel metal2 s 675407 688451 675887 688507 6 mprj_gpio_noesd[3]
port 54 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696980 6 mprj_io[10]
port 55 nsew signal bidirectional
rlabel metal2 s 675407 689003 675887 689059 6 mprj_io_analog_en[10]
port 56 nsew signal input
rlabel metal2 s 675407 690291 675887 690347 6 mprj_io_analog_pol[10]
port 57 nsew signal input
rlabel metal2 s 675407 693327 675887 693383 6 mprj_io_analog_sel[10]
port 58 nsew signal input
rlabel metal2 s 675407 689647 675887 689703 6 mprj_io_dm[30]
port 59 nsew signal input
rlabel metal2 s 675407 687807 675887 687863 6 mprj_io_dm[31]
port 60 nsew signal input
rlabel metal2 s 675407 693971 675887 694027 6 mprj_io_dm[32]
port 61 nsew signal input
rlabel metal2 s 675407 694615 675887 694671 6 mprj_io_holdover[10]
port 62 nsew signal input
rlabel metal2 s 675407 697651 675887 697707 6 mprj_io_ib_mode_sel[10]
port 63 nsew signal input
rlabel metal2 s 675407 690843 675887 690899 6 mprj_io_inp_dis[10]
port 64 nsew signal input
rlabel metal2 s 675407 698295 675887 698351 6 mprj_io_oeb[10]
port 65 nsew signal input
rlabel metal2 s 675407 695167 675887 695223 6 mprj_io_out[10]
port 66 nsew signal input
rlabel metal2 s 675407 685967 675887 686023 6 mprj_io_slow_sel[10]
port 67 nsew signal input
rlabel metal2 s 675407 697007 675887 697063 6 mprj_io_vtrip_sel[10]
port 68 nsew signal input
rlabel metal2 s 675407 684127 675887 684183 6 mprj_io_in[10]
port 69 nsew signal output
rlabel metal2 s 675407 698847 675887 698903 6 mprj_io_in_3v3[10]
port 70 nsew signal output
rlabel metal2 s 675407 731611 675887 731667 6 mprj_gpio_analog[4]
port 71 nsew signal bidirectional
rlabel metal2 s 675407 733451 675887 733507 6 mprj_gpio_noesd[4]
port 72 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741980 6 mprj_io[11]
port 73 nsew signal bidirectional
rlabel metal2 s 675407 734003 675887 734059 6 mprj_io_analog_en[11]
port 74 nsew signal input
rlabel metal2 s 675407 735291 675887 735347 6 mprj_io_analog_pol[11]
port 75 nsew signal input
rlabel metal2 s 675407 738327 675887 738383 6 mprj_io_analog_sel[11]
port 76 nsew signal input
rlabel metal2 s 675407 734647 675887 734703 6 mprj_io_dm[33]
port 77 nsew signal input
rlabel metal2 s 675407 732807 675887 732863 6 mprj_io_dm[34]
port 78 nsew signal input
rlabel metal2 s 675407 738971 675887 739027 6 mprj_io_dm[35]
port 79 nsew signal input
rlabel metal2 s 675407 739615 675887 739671 6 mprj_io_holdover[11]
port 80 nsew signal input
rlabel metal2 s 675407 742651 675887 742707 6 mprj_io_ib_mode_sel[11]
port 81 nsew signal input
rlabel metal2 s 675407 735843 675887 735899 6 mprj_io_inp_dis[11]
port 82 nsew signal input
rlabel metal2 s 675407 743295 675887 743351 6 mprj_io_oeb[11]
port 83 nsew signal input
rlabel metal2 s 675407 740167 675887 740223 6 mprj_io_out[11]
port 84 nsew signal input
rlabel metal2 s 675407 730967 675887 731023 6 mprj_io_slow_sel[11]
port 85 nsew signal input
rlabel metal2 s 675407 742007 675887 742063 6 mprj_io_vtrip_sel[11]
port 86 nsew signal input
rlabel metal2 s 675407 729127 675887 729183 6 mprj_io_in[11]
port 87 nsew signal output
rlabel metal2 s 675407 743847 675887 743903 6 mprj_io_in_3v3[11]
port 88 nsew signal output
rlabel metal2 s 675407 776611 675887 776667 6 mprj_gpio_analog[5]
port 89 nsew signal bidirectional
rlabel metal2 s 675407 778451 675887 778507 6 mprj_gpio_noesd[5]
port 90 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786980 6 mprj_io[12]
port 91 nsew signal bidirectional
rlabel metal2 s 675407 779003 675887 779059 6 mprj_io_analog_en[12]
port 92 nsew signal input
rlabel metal2 s 675407 780291 675887 780347 6 mprj_io_analog_pol[12]
port 93 nsew signal input
rlabel metal2 s 675407 783327 675887 783383 6 mprj_io_analog_sel[12]
port 94 nsew signal input
rlabel metal2 s 675407 779647 675887 779703 6 mprj_io_dm[36]
port 95 nsew signal input
rlabel metal2 s 675407 777807 675887 777863 6 mprj_io_dm[37]
port 96 nsew signal input
rlabel metal2 s 675407 783971 675887 784027 6 mprj_io_dm[38]
port 97 nsew signal input
rlabel metal2 s 675407 784615 675887 784671 6 mprj_io_holdover[12]
port 98 nsew signal input
rlabel metal2 s 675407 787651 675887 787707 6 mprj_io_ib_mode_sel[12]
port 99 nsew signal input
rlabel metal2 s 675407 780843 675887 780899 6 mprj_io_inp_dis[12]
port 100 nsew signal input
rlabel metal2 s 675407 788295 675887 788351 6 mprj_io_oeb[12]
port 101 nsew signal input
rlabel metal2 s 675407 785167 675887 785223 6 mprj_io_out[12]
port 102 nsew signal input
rlabel metal2 s 675407 775967 675887 776023 6 mprj_io_slow_sel[12]
port 103 nsew signal input
rlabel metal2 s 675407 787007 675887 787063 6 mprj_io_vtrip_sel[12]
port 104 nsew signal input
rlabel metal2 s 675407 774127 675887 774183 6 mprj_io_in[12]
port 105 nsew signal output
rlabel metal2 s 675407 788847 675887 788903 6 mprj_io_in_3v3[12]
port 106 nsew signal output
rlabel metal2 s 675407 865811 675887 865867 6 mprj_gpio_analog[6]
port 107 nsew signal bidirectional
rlabel metal2 s 675407 867651 675887 867707 6 mprj_gpio_noesd[6]
port 108 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876180 6 mprj_io[13]
port 109 nsew signal bidirectional
rlabel metal2 s 675407 868203 675887 868259 6 mprj_io_analog_en[13]
port 110 nsew signal input
rlabel metal2 s 675407 869491 675887 869547 6 mprj_io_analog_pol[13]
port 111 nsew signal input
rlabel metal2 s 675407 872527 675887 872583 6 mprj_io_analog_sel[13]
port 112 nsew signal input
rlabel metal2 s 675407 868847 675887 868903 6 mprj_io_dm[39]
port 113 nsew signal input
rlabel metal2 s 675407 867007 675887 867063 6 mprj_io_dm[40]
port 114 nsew signal input
rlabel metal2 s 675407 873171 675887 873227 6 mprj_io_dm[41]
port 115 nsew signal input
rlabel metal2 s 675407 873815 675887 873871 6 mprj_io_holdover[13]
port 116 nsew signal input
rlabel metal2 s 675407 876851 675887 876907 6 mprj_io_ib_mode_sel[13]
port 117 nsew signal input
rlabel metal2 s 675407 870043 675887 870099 6 mprj_io_inp_dis[13]
port 118 nsew signal input
rlabel metal2 s 675407 877495 675887 877551 6 mprj_io_oeb[13]
port 119 nsew signal input
rlabel metal2 s 675407 874367 675887 874423 6 mprj_io_out[13]
port 120 nsew signal input
rlabel metal2 s 675407 865167 675887 865223 6 mprj_io_slow_sel[13]
port 121 nsew signal input
rlabel metal2 s 675407 876207 675887 876263 6 mprj_io_vtrip_sel[13]
port 122 nsew signal input
rlabel metal2 s 675407 863327 675887 863383 6 mprj_io_in[13]
port 123 nsew signal output
rlabel metal2 s 675407 878047 675887 878103 6 mprj_io_in_3v3[13]
port 124 nsew signal output
rlabel metal5 s 698512 146440 711002 158980 6 mprj_io[1]
port 125 nsew signal bidirectional
rlabel metal2 s 675407 151003 675887 151059 6 mprj_io_analog_en[1]
port 126 nsew signal input
rlabel metal2 s 675407 152291 675887 152347 6 mprj_io_analog_pol[1]
port 127 nsew signal input
rlabel metal2 s 675407 155327 675887 155383 6 mprj_io_analog_sel[1]
port 128 nsew signal input
rlabel metal2 s 675407 151647 675887 151703 6 mprj_io_dm[3]
port 129 nsew signal input
rlabel metal2 s 675407 149807 675887 149863 6 mprj_io_dm[4]
port 130 nsew signal input
rlabel metal2 s 675407 155971 675887 156027 6 mprj_io_dm[5]
port 131 nsew signal input
rlabel metal2 s 675407 156615 675887 156671 6 mprj_io_holdover[1]
port 132 nsew signal input
rlabel metal2 s 675407 159651 675887 159707 6 mprj_io_ib_mode_sel[1]
port 133 nsew signal input
rlabel metal2 s 675407 152843 675887 152899 6 mprj_io_inp_dis[1]
port 134 nsew signal input
rlabel metal2 s 675407 160295 675887 160351 6 mprj_io_oeb[1]
port 135 nsew signal input
rlabel metal2 s 675407 157167 675887 157223 6 mprj_io_out[1]
port 136 nsew signal input
rlabel metal2 s 675407 147967 675887 148023 6 mprj_io_slow_sel[1]
port 137 nsew signal input
rlabel metal2 s 675407 159007 675887 159063 6 mprj_io_vtrip_sel[1]
port 138 nsew signal input
rlabel metal2 s 675407 146127 675887 146183 6 mprj_io_in[1]
port 139 nsew signal output
rlabel metal2 s 675407 160847 675887 160903 6 mprj_io_in_3v3[1]
port 140 nsew signal output
rlabel metal5 s 698512 191440 711002 203980 6 mprj_io[2]
port 141 nsew signal bidirectional
rlabel metal2 s 675407 196003 675887 196059 6 mprj_io_analog_en[2]
port 142 nsew signal input
rlabel metal2 s 675407 197291 675887 197347 6 mprj_io_analog_pol[2]
port 143 nsew signal input
rlabel metal2 s 675407 200327 675887 200383 6 mprj_io_analog_sel[2]
port 144 nsew signal input
rlabel metal2 s 675407 196647 675887 196703 6 mprj_io_dm[6]
port 145 nsew signal input
rlabel metal2 s 675407 194807 675887 194863 6 mprj_io_dm[7]
port 146 nsew signal input
rlabel metal2 s 675407 200971 675887 201027 6 mprj_io_dm[8]
port 147 nsew signal input
rlabel metal2 s 675407 201615 675887 201671 6 mprj_io_holdover[2]
port 148 nsew signal input
rlabel metal2 s 675407 204651 675887 204707 6 mprj_io_ib_mode_sel[2]
port 149 nsew signal input
rlabel metal2 s 675407 197843 675887 197899 6 mprj_io_inp_dis[2]
port 150 nsew signal input
rlabel metal2 s 675407 205295 675887 205351 6 mprj_io_oeb[2]
port 151 nsew signal input
rlabel metal2 s 675407 202167 675887 202223 6 mprj_io_out[2]
port 152 nsew signal input
rlabel metal2 s 675407 192967 675887 193023 6 mprj_io_slow_sel[2]
port 153 nsew signal input
rlabel metal2 s 675407 204007 675887 204063 6 mprj_io_vtrip_sel[2]
port 154 nsew signal input
rlabel metal2 s 675407 191127 675887 191183 6 mprj_io_in[2]
port 155 nsew signal output
rlabel metal2 s 675407 205847 675887 205903 6 mprj_io_in_3v3[2]
port 156 nsew signal output
rlabel metal5 s 698512 236640 711002 249180 6 mprj_io[3]
port 157 nsew signal bidirectional
rlabel metal2 s 675407 241203 675887 241259 6 mprj_io_analog_en[3]
port 158 nsew signal input
rlabel metal2 s 675407 242491 675887 242547 6 mprj_io_analog_pol[3]
port 159 nsew signal input
rlabel metal2 s 675407 245527 675887 245583 6 mprj_io_analog_sel[3]
port 160 nsew signal input
rlabel metal2 s 675407 240007 675887 240063 6 mprj_io_dm[10]
port 161 nsew signal input
rlabel metal2 s 675407 246171 675887 246227 6 mprj_io_dm[11]
port 162 nsew signal input
rlabel metal2 s 675407 241847 675887 241903 6 mprj_io_dm[9]
port 163 nsew signal input
rlabel metal2 s 675407 246815 675887 246871 6 mprj_io_holdover[3]
port 164 nsew signal input
rlabel metal2 s 675407 249851 675887 249907 6 mprj_io_ib_mode_sel[3]
port 165 nsew signal input
rlabel metal2 s 675407 243043 675887 243099 6 mprj_io_inp_dis[3]
port 166 nsew signal input
rlabel metal2 s 675407 250495 675887 250551 6 mprj_io_oeb[3]
port 167 nsew signal input
rlabel metal2 s 675407 247367 675887 247423 6 mprj_io_out[3]
port 168 nsew signal input
rlabel metal2 s 675407 238167 675887 238223 6 mprj_io_slow_sel[3]
port 169 nsew signal input
rlabel metal2 s 675407 249207 675887 249263 6 mprj_io_vtrip_sel[3]
port 170 nsew signal input
rlabel metal2 s 675407 236327 675887 236383 6 mprj_io_in[3]
port 171 nsew signal output
rlabel metal2 s 675407 251047 675887 251103 6 mprj_io_in_3v3[3]
port 172 nsew signal output
rlabel metal5 s 698512 281640 711002 294180 6 mprj_io[4]
port 173 nsew signal bidirectional
rlabel metal2 s 675407 286203 675887 286259 6 mprj_io_analog_en[4]
port 174 nsew signal input
rlabel metal2 s 675407 287491 675887 287547 6 mprj_io_analog_pol[4]
port 175 nsew signal input
rlabel metal2 s 675407 290527 675887 290583 6 mprj_io_analog_sel[4]
port 176 nsew signal input
rlabel metal2 s 675407 286847 675887 286903 6 mprj_io_dm[12]
port 177 nsew signal input
rlabel metal2 s 675407 285007 675887 285063 6 mprj_io_dm[13]
port 178 nsew signal input
rlabel metal2 s 675407 291171 675887 291227 6 mprj_io_dm[14]
port 179 nsew signal input
rlabel metal2 s 675407 291815 675887 291871 6 mprj_io_holdover[4]
port 180 nsew signal input
rlabel metal2 s 675407 294851 675887 294907 6 mprj_io_ib_mode_sel[4]
port 181 nsew signal input
rlabel metal2 s 675407 288043 675887 288099 6 mprj_io_inp_dis[4]
port 182 nsew signal input
rlabel metal2 s 675407 295495 675887 295551 6 mprj_io_oeb[4]
port 183 nsew signal input
rlabel metal2 s 675407 292367 675887 292423 6 mprj_io_out[4]
port 184 nsew signal input
rlabel metal2 s 675407 283167 675887 283223 6 mprj_io_slow_sel[4]
port 185 nsew signal input
rlabel metal2 s 675407 294207 675887 294263 6 mprj_io_vtrip_sel[4]
port 186 nsew signal input
rlabel metal2 s 675407 281327 675887 281383 6 mprj_io_in[4]
port 187 nsew signal output
rlabel metal2 s 675407 296047 675887 296103 6 mprj_io_in_3v3[4]
port 188 nsew signal output
rlabel metal5 s 698512 326640 711002 339180 6 mprj_io[5]
port 189 nsew signal bidirectional
rlabel metal2 s 675407 331203 675887 331259 6 mprj_io_analog_en[5]
port 190 nsew signal input
rlabel metal2 s 675407 332491 675887 332547 6 mprj_io_analog_pol[5]
port 191 nsew signal input
rlabel metal2 s 675407 335527 675887 335583 6 mprj_io_analog_sel[5]
port 192 nsew signal input
rlabel metal2 s 675407 331847 675887 331903 6 mprj_io_dm[15]
port 193 nsew signal input
rlabel metal2 s 675407 330007 675887 330063 6 mprj_io_dm[16]
port 194 nsew signal input
rlabel metal2 s 675407 336171 675887 336227 6 mprj_io_dm[17]
port 195 nsew signal input
rlabel metal2 s 675407 336815 675887 336871 6 mprj_io_holdover[5]
port 196 nsew signal input
rlabel metal2 s 675407 339851 675887 339907 6 mprj_io_ib_mode_sel[5]
port 197 nsew signal input
rlabel metal2 s 675407 333043 675887 333099 6 mprj_io_inp_dis[5]
port 198 nsew signal input
rlabel metal2 s 675407 340495 675887 340551 6 mprj_io_oeb[5]
port 199 nsew signal input
rlabel metal2 s 675407 337367 675887 337423 6 mprj_io_out[5]
port 200 nsew signal input
rlabel metal2 s 675407 328167 675887 328223 6 mprj_io_slow_sel[5]
port 201 nsew signal input
rlabel metal2 s 675407 339207 675887 339263 6 mprj_io_vtrip_sel[5]
port 202 nsew signal input
rlabel metal2 s 675407 326327 675887 326383 6 mprj_io_in[5]
port 203 nsew signal output
rlabel metal2 s 675407 341047 675887 341103 6 mprj_io_in_3v3[5]
port 204 nsew signal output
rlabel metal5 s 698512 371840 711002 384380 6 mprj_io[6]
port 205 nsew signal bidirectional
rlabel metal2 s 675407 376403 675887 376459 6 mprj_io_analog_en[6]
port 206 nsew signal input
rlabel metal2 s 675407 377691 675887 377747 6 mprj_io_analog_pol[6]
port 207 nsew signal input
rlabel metal2 s 675407 380727 675887 380783 6 mprj_io_analog_sel[6]
port 208 nsew signal input
rlabel metal2 s 675407 377047 675887 377103 6 mprj_io_dm[18]
port 209 nsew signal input
rlabel metal2 s 675407 375207 675887 375263 6 mprj_io_dm[19]
port 210 nsew signal input
rlabel metal2 s 675407 381371 675887 381427 6 mprj_io_dm[20]
port 211 nsew signal input
rlabel metal2 s 675407 382015 675887 382071 6 mprj_io_holdover[6]
port 212 nsew signal input
rlabel metal2 s 675407 385051 675887 385107 6 mprj_io_ib_mode_sel[6]
port 213 nsew signal input
rlabel metal2 s 675407 378243 675887 378299 6 mprj_io_inp_dis[6]
port 214 nsew signal input
rlabel metal2 s 675407 385695 675887 385751 6 mprj_io_oeb[6]
port 215 nsew signal input
rlabel metal2 s 675407 382567 675887 382623 6 mprj_io_out[6]
port 216 nsew signal input
rlabel metal2 s 675407 373367 675887 373423 6 mprj_io_slow_sel[6]
port 217 nsew signal input
rlabel metal2 s 675407 384407 675887 384463 6 mprj_io_vtrip_sel[6]
port 218 nsew signal input
rlabel metal2 s 675407 371527 675887 371583 6 mprj_io_in[6]
port 219 nsew signal output
rlabel metal2 s 675407 386247 675887 386303 6 mprj_io_in_3v3[6]
port 220 nsew signal output
rlabel metal2 s 675407 551211 675887 551267 6 mprj_gpio_analog[0]
port 221 nsew signal bidirectional
rlabel metal2 s 675407 553051 675887 553107 6 mprj_gpio_noesd[0]
port 222 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561580 6 mprj_io[7]
port 223 nsew signal bidirectional
rlabel metal2 s 675407 553603 675887 553659 6 mprj_io_analog_en[7]
port 224 nsew signal input
rlabel metal2 s 675407 554891 675887 554947 6 mprj_io_analog_pol[7]
port 225 nsew signal input
rlabel metal2 s 675407 557927 675887 557983 6 mprj_io_analog_sel[7]
port 226 nsew signal input
rlabel metal2 s 675407 554247 675887 554303 6 mprj_io_dm[21]
port 227 nsew signal input
rlabel metal2 s 675407 552407 675887 552463 6 mprj_io_dm[22]
port 228 nsew signal input
rlabel metal2 s 675407 558571 675887 558627 6 mprj_io_dm[23]
port 229 nsew signal input
rlabel metal2 s 675407 559215 675887 559271 6 mprj_io_holdover[7]
port 230 nsew signal input
rlabel metal2 s 675407 562251 675887 562307 6 mprj_io_ib_mode_sel[7]
port 231 nsew signal input
rlabel metal2 s 675407 555443 675887 555499 6 mprj_io_inp_dis[7]
port 232 nsew signal input
rlabel metal2 s 675407 562895 675887 562951 6 mprj_io_oeb[7]
port 233 nsew signal input
rlabel metal2 s 675407 559767 675887 559823 6 mprj_io_out[7]
port 234 nsew signal input
rlabel metal2 s 675407 550567 675887 550623 6 mprj_io_slow_sel[7]
port 235 nsew signal input
rlabel metal2 s 675407 561607 675887 561663 6 mprj_io_vtrip_sel[7]
port 236 nsew signal input
rlabel metal2 s 675407 548727 675887 548783 6 mprj_io_in[7]
port 237 nsew signal output
rlabel metal2 s 675407 563447 675887 563503 6 mprj_io_in_3v3[7]
port 238 nsew signal output
rlabel metal2 s 675407 596411 675887 596467 6 mprj_gpio_analog[1]
port 239 nsew signal bidirectional
rlabel metal2 s 675407 598251 675887 598307 6 mprj_gpio_noesd[1]
port 240 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606780 6 mprj_io[8]
port 241 nsew signal bidirectional
rlabel metal2 s 675407 598803 675887 598859 6 mprj_io_analog_en[8]
port 242 nsew signal input
rlabel metal2 s 675407 600091 675887 600147 6 mprj_io_analog_pol[8]
port 243 nsew signal input
rlabel metal2 s 675407 603127 675887 603183 6 mprj_io_analog_sel[8]
port 244 nsew signal input
rlabel metal2 s 675407 599447 675887 599503 6 mprj_io_dm[24]
port 245 nsew signal input
rlabel metal2 s 675407 597607 675887 597663 6 mprj_io_dm[25]
port 246 nsew signal input
rlabel metal2 s 675407 603771 675887 603827 6 mprj_io_dm[26]
port 247 nsew signal input
rlabel metal2 s 675407 604415 675887 604471 6 mprj_io_holdover[8]
port 248 nsew signal input
rlabel metal2 s 675407 607451 675887 607507 6 mprj_io_ib_mode_sel[8]
port 249 nsew signal input
rlabel metal2 s 675407 600643 675887 600699 6 mprj_io_inp_dis[8]
port 250 nsew signal input
rlabel metal2 s 675407 608095 675887 608151 6 mprj_io_oeb[8]
port 251 nsew signal input
rlabel metal2 s 675407 604967 675887 605023 6 mprj_io_out[8]
port 252 nsew signal input
rlabel metal2 s 675407 595767 675887 595823 6 mprj_io_slow_sel[8]
port 253 nsew signal input
rlabel metal2 s 675407 606807 675887 606863 6 mprj_io_vtrip_sel[8]
port 254 nsew signal input
rlabel metal2 s 675407 593927 675887 593983 6 mprj_io_in[8]
port 255 nsew signal output
rlabel metal2 s 675407 608647 675887 608703 6 mprj_io_in_3v3[8]
port 256 nsew signal output
rlabel metal2 s 675407 641411 675887 641467 6 mprj_gpio_analog[2]
port 257 nsew signal bidirectional
rlabel metal2 s 675407 643251 675887 643307 6 mprj_gpio_noesd[2]
port 258 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651780 6 mprj_io[9]
port 259 nsew signal bidirectional
rlabel metal2 s 675407 643803 675887 643859 6 mprj_io_analog_en[9]
port 260 nsew signal input
rlabel metal2 s 675407 645091 675887 645147 6 mprj_io_analog_pol[9]
port 261 nsew signal input
rlabel metal2 s 675407 648127 675887 648183 6 mprj_io_analog_sel[9]
port 262 nsew signal input
rlabel metal2 s 675407 644447 675887 644503 6 mprj_io_dm[27]
port 263 nsew signal input
rlabel metal2 s 675407 642607 675887 642663 6 mprj_io_dm[28]
port 264 nsew signal input
rlabel metal2 s 675407 648771 675887 648827 6 mprj_io_dm[29]
port 265 nsew signal input
rlabel metal2 s 675407 649415 675887 649471 6 mprj_io_holdover[9]
port 266 nsew signal input
rlabel metal2 s 675407 652451 675887 652507 6 mprj_io_ib_mode_sel[9]
port 267 nsew signal input
rlabel metal2 s 675407 645643 675887 645699 6 mprj_io_inp_dis[9]
port 268 nsew signal input
rlabel metal2 s 675407 653095 675887 653151 6 mprj_io_oeb[9]
port 269 nsew signal input
rlabel metal2 s 675407 649967 675887 650023 6 mprj_io_out[9]
port 270 nsew signal input
rlabel metal2 s 675407 640767 675887 640823 6 mprj_io_slow_sel[9]
port 271 nsew signal input
rlabel metal2 s 675407 651807 675887 651863 6 mprj_io_vtrip_sel[9]
port 272 nsew signal input
rlabel metal2 s 675407 638927 675887 638983 6 mprj_io_in[9]
port 273 nsew signal output
rlabel metal2 s 675407 653647 675887 653703 6 mprj_io_in_3v3[9]
port 274 nsew signal output
rlabel metal2 s 41713 796933 42193 796989 6 mprj_gpio_analog[7]
port 275 nsew signal bidirectional
rlabel metal2 s 41713 795093 42193 795149 6 mprj_gpio_noesd[7]
port 276 nsew signal bidirectional
rlabel metal5 s 6598 786620 19088 799160 6 mprj_io[25]
port 277 nsew signal bidirectional
rlabel metal2 s 41713 794541 42193 794597 6 mprj_io_analog_en[14]
port 278 nsew signal input
rlabel metal2 s 41713 793253 42193 793309 6 mprj_io_analog_pol[14]
port 279 nsew signal input
rlabel metal2 s 41713 790217 42193 790273 6 mprj_io_analog_sel[14]
port 280 nsew signal input
rlabel metal2 s 41713 793897 42193 793953 6 mprj_io_dm[42]
port 281 nsew signal input
rlabel metal2 s 41713 795737 42193 795793 6 mprj_io_dm[43]
port 282 nsew signal input
rlabel metal2 s 41713 789573 42193 789629 6 mprj_io_dm[44]
port 283 nsew signal input
rlabel metal2 s 41713 788929 42193 788985 6 mprj_io_holdover[14]
port 284 nsew signal input
rlabel metal2 s 41713 785893 42193 785949 6 mprj_io_ib_mode_sel[14]
port 285 nsew signal input
rlabel metal2 s 41713 792701 42193 792757 6 mprj_io_inp_dis[14]
port 286 nsew signal input
rlabel metal2 s 41713 785249 42193 785305 6 mprj_io_oeb[14]
port 287 nsew signal input
rlabel metal2 s 41713 788377 42193 788433 6 mprj_io_out[14]
port 288 nsew signal input
rlabel metal2 s 41713 797577 42193 797633 6 mprj_io_slow_sel[14]
port 289 nsew signal input
rlabel metal2 s 41713 786537 42193 786593 6 mprj_io_vtrip_sel[14]
port 290 nsew signal input
rlabel metal2 s 41713 799417 42193 799473 6 mprj_io_in[14]
port 291 nsew signal output
rlabel metal2 s 41713 784697 42193 784753 6 mprj_io_in_3v3[14]
port 292 nsew signal output
rlabel metal2 s 41713 280533 42193 280589 6 mprj_gpio_analog[17]
port 293 nsew signal bidirectional
rlabel metal2 s 41713 278693 42193 278749 6 mprj_gpio_noesd[17]
port 294 nsew signal bidirectional
rlabel metal5 s 6598 270220 19088 282760 6 mprj_io[35]
port 295 nsew signal bidirectional
rlabel metal2 s 41713 278141 42193 278197 6 mprj_io_analog_en[24]
port 296 nsew signal input
rlabel metal2 s 41713 276853 42193 276909 6 mprj_io_analog_pol[24]
port 297 nsew signal input
rlabel metal2 s 41713 273817 42193 273873 6 mprj_io_analog_sel[24]
port 298 nsew signal input
rlabel metal2 s 41713 277497 42193 277553 6 mprj_io_dm[72]
port 299 nsew signal input
rlabel metal2 s 41713 279337 42193 279393 6 mprj_io_dm[73]
port 300 nsew signal input
rlabel metal2 s 41713 273173 42193 273229 6 mprj_io_dm[74]
port 301 nsew signal input
rlabel metal2 s 41713 272529 42193 272585 6 mprj_io_holdover[24]
port 302 nsew signal input
rlabel metal2 s 41713 269493 42193 269549 6 mprj_io_ib_mode_sel[24]
port 303 nsew signal input
rlabel metal2 s 41713 276301 42193 276357 6 mprj_io_inp_dis[24]
port 304 nsew signal input
rlabel metal2 s 41713 268849 42193 268905 6 mprj_io_oeb[24]
port 305 nsew signal input
rlabel metal2 s 41713 271977 42193 272033 6 mprj_io_out[24]
port 306 nsew signal input
rlabel metal2 s 41713 281177 42193 281233 6 mprj_io_slow_sel[24]
port 307 nsew signal input
rlabel metal2 s 41713 270137 42193 270193 6 mprj_io_vtrip_sel[24]
port 308 nsew signal input
rlabel metal2 s 41713 283017 42193 283073 6 mprj_io_in[24]
port 309 nsew signal output
rlabel metal2 s 41713 268297 42193 268353 6 mprj_io_in_3v3[24]
port 310 nsew signal output
rlabel metal5 s 6598 227020 19088 239560 6 mprj_io[36]
port 311 nsew signal bidirectional
rlabel metal2 s 41713 234941 42193 234997 6 mprj_io_analog_en[25]
port 312 nsew signal input
rlabel metal2 s 41713 233653 42193 233709 6 mprj_io_analog_pol[25]
port 313 nsew signal input
rlabel metal2 s 41713 230617 42193 230673 6 mprj_io_analog_sel[25]
port 314 nsew signal input
rlabel metal2 s 41713 234297 42193 234353 6 mprj_io_dm[75]
port 315 nsew signal input
rlabel metal2 s 41713 236137 42193 236193 6 mprj_io_dm[76]
port 316 nsew signal input
rlabel metal2 s 41713 229973 42193 230029 6 mprj_io_dm[77]
port 317 nsew signal input
rlabel metal2 s 41713 229329 42193 229385 6 mprj_io_holdover[25]
port 318 nsew signal input
rlabel metal2 s 41713 226293 42193 226349 6 mprj_io_ib_mode_sel[25]
port 319 nsew signal input
rlabel metal2 s 41713 233101 42193 233157 6 mprj_io_inp_dis[25]
port 320 nsew signal input
rlabel metal2 s 41713 225649 42193 225705 6 mprj_io_oeb[25]
port 321 nsew signal input
rlabel metal2 s 41713 228777 42193 228833 6 mprj_io_out[25]
port 322 nsew signal input
rlabel metal2 s 41713 237977 42193 238033 6 mprj_io_slow_sel[25]
port 323 nsew signal input
rlabel metal2 s 41713 226937 42193 226993 6 mprj_io_vtrip_sel[25]
port 324 nsew signal input
rlabel metal2 s 41713 239817 42193 239873 6 mprj_io_in[25]
port 325 nsew signal output
rlabel metal2 s 41713 225097 42193 225153 6 mprj_io_in_3v3[25]
port 326 nsew signal output
rlabel metal5 s 6598 183820 19088 196360 6 mprj_io[37]
port 327 nsew signal bidirectional
rlabel metal2 s 41713 191741 42193 191797 6 mprj_io_analog_en[26]
port 328 nsew signal input
rlabel metal2 s 41713 190453 42193 190509 6 mprj_io_analog_pol[26]
port 329 nsew signal input
rlabel metal2 s 41713 187417 42193 187473 6 mprj_io_analog_sel[26]
port 330 nsew signal input
rlabel metal2 s 41713 191097 42193 191153 6 mprj_io_dm[78]
port 331 nsew signal input
rlabel metal2 s 41713 192937 42193 192993 6 mprj_io_dm[79]
port 332 nsew signal input
rlabel metal2 s 41713 186773 42193 186829 6 mprj_io_dm[80]
port 333 nsew signal input
rlabel metal2 s 41713 186129 42193 186185 6 mprj_io_holdover[26]
port 334 nsew signal input
rlabel metal2 s 41713 183093 42193 183149 6 mprj_io_ib_mode_sel[26]
port 335 nsew signal input
rlabel metal2 s 41713 189901 42193 189957 6 mprj_io_inp_dis[26]
port 336 nsew signal input
rlabel metal2 s 41713 182449 42193 182505 6 mprj_io_oeb[26]
port 337 nsew signal input
rlabel metal2 s 41713 185577 42193 185633 6 mprj_io_out[26]
port 338 nsew signal input
rlabel metal2 s 41713 194777 42193 194833 6 mprj_io_slow_sel[26]
port 339 nsew signal input
rlabel metal2 s 41713 183737 42193 183793 6 mprj_io_vtrip_sel[26]
port 340 nsew signal input
rlabel metal2 s 41713 196617 42193 196673 6 mprj_io_in[26]
port 341 nsew signal output
rlabel metal2 s 41713 181897 42193 181953 6 mprj_io_in_3v3[26]
port 342 nsew signal output
rlabel metal2 s 41713 753733 42193 753789 6 mprj_gpio_analog[8]
port 343 nsew signal bidirectional
rlabel metal2 s 41713 751893 42193 751949 6 mprj_gpio_noesd[8]
port 344 nsew signal bidirectional
rlabel metal5 s 6598 743420 19088 755960 6 mprj_io[26]
port 345 nsew signal bidirectional
rlabel metal2 s 41713 751341 42193 751397 6 mprj_io_analog_en[15]
port 346 nsew signal input
rlabel metal2 s 41713 750053 42193 750109 6 mprj_io_analog_pol[15]
port 347 nsew signal input
rlabel metal2 s 41713 747017 42193 747073 6 mprj_io_analog_sel[15]
port 348 nsew signal input
rlabel metal2 s 41713 750697 42193 750753 6 mprj_io_dm[45]
port 349 nsew signal input
rlabel metal2 s 41713 752537 42193 752593 6 mprj_io_dm[46]
port 350 nsew signal input
rlabel metal2 s 41713 746373 42193 746429 6 mprj_io_dm[47]
port 351 nsew signal input
rlabel metal2 s 41713 745729 42193 745785 6 mprj_io_holdover[15]
port 352 nsew signal input
rlabel metal2 s 41713 742693 42193 742749 6 mprj_io_ib_mode_sel[15]
port 353 nsew signal input
rlabel metal2 s 41713 749501 42193 749557 6 mprj_io_inp_dis[15]
port 354 nsew signal input
rlabel metal2 s 41713 742049 42193 742105 6 mprj_io_oeb[15]
port 355 nsew signal input
rlabel metal2 s 41713 745177 42193 745233 6 mprj_io_out[15]
port 356 nsew signal input
rlabel metal2 s 41713 754377 42193 754433 6 mprj_io_slow_sel[15]
port 357 nsew signal input
rlabel metal2 s 41713 743337 42193 743393 6 mprj_io_vtrip_sel[15]
port 358 nsew signal input
rlabel metal2 s 41713 756217 42193 756273 6 mprj_io_in[15]
port 359 nsew signal output
rlabel metal2 s 41713 741497 42193 741553 6 mprj_io_in_3v3[15]
port 360 nsew signal output
rlabel metal2 s 41713 710533 42193 710589 6 mprj_gpio_analog[9]
port 361 nsew signal bidirectional
rlabel metal2 s 41713 708693 42193 708749 6 mprj_gpio_noesd[9]
port 362 nsew signal bidirectional
rlabel metal5 s 6598 700220 19088 712760 6 mprj_io[27]
port 363 nsew signal bidirectional
rlabel metal2 s 41713 708141 42193 708197 6 mprj_io_analog_en[16]
port 364 nsew signal input
rlabel metal2 s 41713 706853 42193 706909 6 mprj_io_analog_pol[16]
port 365 nsew signal input
rlabel metal2 s 41713 703817 42193 703873 6 mprj_io_analog_sel[16]
port 366 nsew signal input
rlabel metal2 s 41713 707497 42193 707553 6 mprj_io_dm[48]
port 367 nsew signal input
rlabel metal2 s 41713 709337 42193 709393 6 mprj_io_dm[49]
port 368 nsew signal input
rlabel metal2 s 41713 703173 42193 703229 6 mprj_io_dm[50]
port 369 nsew signal input
rlabel metal2 s 41713 702529 42193 702585 6 mprj_io_holdover[16]
port 370 nsew signal input
rlabel metal2 s 41713 699493 42193 699549 6 mprj_io_ib_mode_sel[16]
port 371 nsew signal input
rlabel metal2 s 41713 706301 42193 706357 6 mprj_io_inp_dis[16]
port 372 nsew signal input
rlabel metal2 s 41713 698849 42193 698905 6 mprj_io_oeb[16]
port 373 nsew signal input
rlabel metal2 s 41713 701977 42193 702033 6 mprj_io_out[16]
port 374 nsew signal input
rlabel metal2 s 41713 711177 42193 711233 6 mprj_io_slow_sel[16]
port 375 nsew signal input
rlabel metal2 s 41713 700137 42193 700193 6 mprj_io_vtrip_sel[16]
port 376 nsew signal input
rlabel metal2 s 41713 713017 42193 713073 6 mprj_io_in[16]
port 377 nsew signal output
rlabel metal2 s 41713 698297 42193 698353 6 mprj_io_in_3v3[16]
port 378 nsew signal output
rlabel metal2 s 41713 667333 42193 667389 6 mprj_gpio_analog[10]
port 379 nsew signal bidirectional
rlabel metal2 s 41713 665493 42193 665549 6 mprj_gpio_noesd[10]
port 380 nsew signal bidirectional
rlabel metal5 s 6598 657020 19088 669560 6 mprj_io[28]
port 381 nsew signal bidirectional
rlabel metal2 s 41713 664941 42193 664997 6 mprj_io_analog_en[17]
port 382 nsew signal input
rlabel metal2 s 41713 663653 42193 663709 6 mprj_io_analog_pol[17]
port 383 nsew signal input
rlabel metal2 s 41713 660617 42193 660673 6 mprj_io_analog_sel[17]
port 384 nsew signal input
rlabel metal2 s 41713 664297 42193 664353 6 mprj_io_dm[51]
port 385 nsew signal input
rlabel metal2 s 41713 666137 42193 666193 6 mprj_io_dm[52]
port 386 nsew signal input
rlabel metal2 s 41713 659973 42193 660029 6 mprj_io_dm[53]
port 387 nsew signal input
rlabel metal2 s 41713 659329 42193 659385 6 mprj_io_holdover[17]
port 388 nsew signal input
rlabel metal2 s 41713 656293 42193 656349 6 mprj_io_ib_mode_sel[17]
port 389 nsew signal input
rlabel metal2 s 41713 663101 42193 663157 6 mprj_io_inp_dis[17]
port 390 nsew signal input
rlabel metal2 s 41713 655649 42193 655705 6 mprj_io_oeb[17]
port 391 nsew signal input
rlabel metal2 s 41713 658777 42193 658833 6 mprj_io_out[17]
port 392 nsew signal input
rlabel metal2 s 41713 667977 42193 668033 6 mprj_io_slow_sel[17]
port 393 nsew signal input
rlabel metal2 s 41713 656937 42193 656993 6 mprj_io_vtrip_sel[17]
port 394 nsew signal input
rlabel metal2 s 41713 669817 42193 669873 6 mprj_io_in[17]
port 395 nsew signal output
rlabel metal2 s 41713 655097 42193 655153 6 mprj_io_in_3v3[17]
port 396 nsew signal output
rlabel metal2 s 41713 624133 42193 624189 6 mprj_gpio_analog[11]
port 397 nsew signal bidirectional
rlabel metal2 s 41713 622293 42193 622349 6 mprj_gpio_noesd[11]
port 398 nsew signal bidirectional
rlabel metal5 s 6598 613820 19088 626360 6 mprj_io[29]
port 399 nsew signal bidirectional
rlabel metal2 s 41713 621741 42193 621797 6 mprj_io_analog_en[18]
port 400 nsew signal input
rlabel metal2 s 41713 620453 42193 620509 6 mprj_io_analog_pol[18]
port 401 nsew signal input
rlabel metal2 s 41713 617417 42193 617473 6 mprj_io_analog_sel[18]
port 402 nsew signal input
rlabel metal2 s 41713 621097 42193 621153 6 mprj_io_dm[54]
port 403 nsew signal input
rlabel metal2 s 41713 622937 42193 622993 6 mprj_io_dm[55]
port 404 nsew signal input
rlabel metal2 s 41713 616773 42193 616829 6 mprj_io_dm[56]
port 405 nsew signal input
rlabel metal2 s 41713 616129 42193 616185 6 mprj_io_holdover[18]
port 406 nsew signal input
rlabel metal2 s 41713 613093 42193 613149 6 mprj_io_ib_mode_sel[18]
port 407 nsew signal input
rlabel metal2 s 41713 619901 42193 619957 6 mprj_io_inp_dis[18]
port 408 nsew signal input
rlabel metal2 s 41713 612449 42193 612505 6 mprj_io_oeb[18]
port 409 nsew signal input
rlabel metal2 s 41713 615577 42193 615633 6 mprj_io_out[18]
port 410 nsew signal input
rlabel metal2 s 41713 624777 42193 624833 6 mprj_io_slow_sel[18]
port 411 nsew signal input
rlabel metal2 s 41713 613737 42193 613793 6 mprj_io_vtrip_sel[18]
port 412 nsew signal input
rlabel metal2 s 41713 626617 42193 626673 6 mprj_io_in[18]
port 413 nsew signal output
rlabel metal2 s 41713 611897 42193 611953 6 mprj_io_in_3v3[18]
port 414 nsew signal output
rlabel metal2 s 41713 580933 42193 580989 6 mprj_gpio_analog[12]
port 415 nsew signal bidirectional
rlabel metal2 s 41713 579093 42193 579149 6 mprj_gpio_noesd[12]
port 416 nsew signal bidirectional
rlabel metal5 s 6598 570620 19088 583160 6 mprj_io[30]
port 417 nsew signal bidirectional
rlabel metal2 s 41713 578541 42193 578597 6 mprj_io_analog_en[19]
port 418 nsew signal input
rlabel metal2 s 41713 577253 42193 577309 6 mprj_io_analog_pol[19]
port 419 nsew signal input
rlabel metal2 s 41713 574217 42193 574273 6 mprj_io_analog_sel[19]
port 420 nsew signal input
rlabel metal2 s 41713 577897 42193 577953 6 mprj_io_dm[57]
port 421 nsew signal input
rlabel metal2 s 41713 579737 42193 579793 6 mprj_io_dm[58]
port 422 nsew signal input
rlabel metal2 s 41713 573573 42193 573629 6 mprj_io_dm[59]
port 423 nsew signal input
rlabel metal2 s 41713 572929 42193 572985 6 mprj_io_holdover[19]
port 424 nsew signal input
rlabel metal2 s 41713 569893 42193 569949 6 mprj_io_ib_mode_sel[19]
port 425 nsew signal input
rlabel metal2 s 41713 576701 42193 576757 6 mprj_io_inp_dis[19]
port 426 nsew signal input
rlabel metal2 s 41713 569249 42193 569305 6 mprj_io_oeb[19]
port 427 nsew signal input
rlabel metal2 s 41713 572377 42193 572433 6 mprj_io_out[19]
port 428 nsew signal input
rlabel metal2 s 41713 581577 42193 581633 6 mprj_io_slow_sel[19]
port 429 nsew signal input
rlabel metal2 s 41713 570537 42193 570593 6 mprj_io_vtrip_sel[19]
port 430 nsew signal input
rlabel metal2 s 41713 583417 42193 583473 6 mprj_io_in[19]
port 431 nsew signal output
rlabel metal2 s 41713 568697 42193 568753 6 mprj_io_in_3v3[19]
port 432 nsew signal output
rlabel metal2 s 41713 537733 42193 537789 6 mprj_gpio_analog[13]
port 433 nsew signal bidirectional
rlabel metal2 s 41713 535893 42193 535949 6 mprj_gpio_noesd[13]
port 434 nsew signal bidirectional
rlabel metal5 s 6598 527420 19088 539960 6 mprj_io[31]
port 435 nsew signal bidirectional
rlabel metal2 s 41713 535341 42193 535397 6 mprj_io_analog_en[20]
port 436 nsew signal input
rlabel metal2 s 41713 534053 42193 534109 6 mprj_io_analog_pol[20]
port 437 nsew signal input
rlabel metal2 s 41713 531017 42193 531073 6 mprj_io_analog_sel[20]
port 438 nsew signal input
rlabel metal2 s 41713 534697 42193 534753 6 mprj_io_dm[60]
port 439 nsew signal input
rlabel metal2 s 41713 536537 42193 536593 6 mprj_io_dm[61]
port 440 nsew signal input
rlabel metal2 s 41713 530373 42193 530429 6 mprj_io_dm[62]
port 441 nsew signal input
rlabel metal2 s 41713 529729 42193 529785 6 mprj_io_holdover[20]
port 442 nsew signal input
rlabel metal2 s 41713 526693 42193 526749 6 mprj_io_ib_mode_sel[20]
port 443 nsew signal input
rlabel metal2 s 41713 533501 42193 533557 6 mprj_io_inp_dis[20]
port 444 nsew signal input
rlabel metal2 s 41713 526049 42193 526105 6 mprj_io_oeb[20]
port 445 nsew signal input
rlabel metal2 s 41713 529177 42193 529233 6 mprj_io_out[20]
port 446 nsew signal input
rlabel metal2 s 41713 538377 42193 538433 6 mprj_io_slow_sel[20]
port 447 nsew signal input
rlabel metal2 s 41713 527337 42193 527393 6 mprj_io_vtrip_sel[20]
port 448 nsew signal input
rlabel metal2 s 41713 540217 42193 540273 6 mprj_io_in[20]
port 449 nsew signal output
rlabel metal2 s 41713 525497 42193 525553 6 mprj_io_in_3v3[20]
port 450 nsew signal output
rlabel metal2 s 41713 410133 42193 410189 6 mprj_gpio_analog[14]
port 451 nsew signal bidirectional
rlabel metal2 s 41713 408293 42193 408349 6 mprj_gpio_noesd[14]
port 452 nsew signal bidirectional
rlabel metal5 s 6598 399820 19088 412360 6 mprj_io[32]
port 453 nsew signal bidirectional
rlabel metal2 s 41713 407741 42193 407797 6 mprj_io_analog_en[21]
port 454 nsew signal input
rlabel metal2 s 41713 406453 42193 406509 6 mprj_io_analog_pol[21]
port 455 nsew signal input
rlabel metal2 s 41713 403417 42193 403473 6 mprj_io_analog_sel[21]
port 456 nsew signal input
rlabel metal2 s 41713 407097 42193 407153 6 mprj_io_dm[63]
port 457 nsew signal input
rlabel metal2 s 41713 408937 42193 408993 6 mprj_io_dm[64]
port 458 nsew signal input
rlabel metal2 s 41713 402773 42193 402829 6 mprj_io_dm[65]
port 459 nsew signal input
rlabel metal2 s 41713 402129 42193 402185 6 mprj_io_holdover[21]
port 460 nsew signal input
rlabel metal2 s 41713 399093 42193 399149 6 mprj_io_ib_mode_sel[21]
port 461 nsew signal input
rlabel metal2 s 41713 405901 42193 405957 6 mprj_io_inp_dis[21]
port 462 nsew signal input
rlabel metal2 s 41713 398449 42193 398505 6 mprj_io_oeb[21]
port 463 nsew signal input
rlabel metal2 s 41713 401577 42193 401633 6 mprj_io_out[21]
port 464 nsew signal input
rlabel metal2 s 41713 410777 42193 410833 6 mprj_io_slow_sel[21]
port 465 nsew signal input
rlabel metal2 s 41713 399737 42193 399793 6 mprj_io_vtrip_sel[21]
port 466 nsew signal input
rlabel metal2 s 41713 412617 42193 412673 6 mprj_io_in[21]
port 467 nsew signal output
rlabel metal2 s 41713 397897 42193 397953 6 mprj_io_in_3v3[21]
port 468 nsew signal output
rlabel metal2 s 41713 366933 42193 366989 6 mprj_gpio_analog[15]
port 469 nsew signal bidirectional
rlabel metal2 s 41713 365093 42193 365149 6 mprj_gpio_noesd[15]
port 470 nsew signal bidirectional
rlabel metal5 s 6598 356620 19088 369160 6 mprj_io[33]
port 471 nsew signal bidirectional
rlabel metal2 s 41713 364541 42193 364597 6 mprj_io_analog_en[22]
port 472 nsew signal input
rlabel metal2 s 41713 363253 42193 363309 6 mprj_io_analog_pol[22]
port 473 nsew signal input
rlabel metal2 s 41713 360217 42193 360273 6 mprj_io_analog_sel[22]
port 474 nsew signal input
rlabel metal2 s 41713 363897 42193 363953 6 mprj_io_dm[66]
port 475 nsew signal input
rlabel metal2 s 41713 365737 42193 365793 6 mprj_io_dm[67]
port 476 nsew signal input
rlabel metal2 s 41713 359573 42193 359629 6 mprj_io_dm[68]
port 477 nsew signal input
rlabel metal2 s 41713 358929 42193 358985 6 mprj_io_holdover[22]
port 478 nsew signal input
rlabel metal2 s 41713 355893 42193 355949 6 mprj_io_ib_mode_sel[22]
port 479 nsew signal input
rlabel metal2 s 41713 362701 42193 362757 6 mprj_io_inp_dis[22]
port 480 nsew signal input
rlabel metal2 s 41713 355249 42193 355305 6 mprj_io_oeb[22]
port 481 nsew signal input
rlabel metal2 s 41713 358377 42193 358433 6 mprj_io_out[22]
port 482 nsew signal input
rlabel metal2 s 41713 367577 42193 367633 6 mprj_io_slow_sel[22]
port 483 nsew signal input
rlabel metal2 s 41713 356537 42193 356593 6 mprj_io_vtrip_sel[22]
port 484 nsew signal input
rlabel metal2 s 41713 369417 42193 369473 6 mprj_io_in[22]
port 485 nsew signal output
rlabel metal2 s 41713 354697 42193 354753 6 mprj_io_in_3v3[22]
port 486 nsew signal output
rlabel metal2 s 41713 323733 42193 323789 6 mprj_gpio_analog[16]
port 487 nsew signal bidirectional
rlabel metal2 s 41713 321893 42193 321949 6 mprj_gpio_noesd[16]
port 488 nsew signal bidirectional
rlabel metal5 s 6598 313420 19088 325960 6 mprj_io[34]
port 489 nsew signal bidirectional
rlabel metal2 s 41713 321341 42193 321397 6 mprj_io_analog_en[23]
port 490 nsew signal input
rlabel metal2 s 41713 320053 42193 320109 6 mprj_io_analog_pol[23]
port 491 nsew signal input
rlabel metal2 s 41713 317017 42193 317073 6 mprj_io_analog_sel[23]
port 492 nsew signal input
rlabel metal2 s 41713 320697 42193 320753 6 mprj_io_dm[69]
port 493 nsew signal input
rlabel metal2 s 41713 322537 42193 322593 6 mprj_io_dm[70]
port 494 nsew signal input
rlabel metal2 s 41713 316373 42193 316429 6 mprj_io_dm[71]
port 495 nsew signal input
rlabel metal2 s 41713 315729 42193 315785 6 mprj_io_holdover[23]
port 496 nsew signal input
rlabel metal2 s 41713 312693 42193 312749 6 mprj_io_ib_mode_sel[23]
port 497 nsew signal input
rlabel metal2 s 41713 319501 42193 319557 6 mprj_io_inp_dis[23]
port 498 nsew signal input
rlabel metal2 s 41713 312049 42193 312105 6 mprj_io_oeb[23]
port 499 nsew signal input
rlabel metal2 s 41713 315177 42193 315233 6 mprj_io_out[23]
port 500 nsew signal input
rlabel metal2 s 41713 324377 42193 324433 6 mprj_io_slow_sel[23]
port 501 nsew signal input
rlabel metal2 s 41713 313337 42193 313393 6 mprj_io_vtrip_sel[23]
port 502 nsew signal input
rlabel metal2 s 41713 326217 42193 326273 6 mprj_io_in[23]
port 503 nsew signal output
rlabel metal2 s 41713 311497 42193 311553 6 mprj_io_in_3v3[23]
port 504 nsew signal output
rlabel metal3 s 52453 46819 52519 46822 6 porb_h
port 505 nsew signal input
rlabel metal3 s 44774 46822 52519 46882 6 porb_h
port 505 nsew signal input
rlabel metal3 s 52453 46882 52519 46885 6 porb_h
port 505 nsew signal input
rlabel metal3 s 44774 46882 44834 46958 6 porb_h
port 505 nsew signal input
rlabel metal3 s 42333 46955 42399 46958 6 porb_h
port 505 nsew signal input
rlabel metal3 s 42333 46958 44834 47018 6 porb_h
port 505 nsew signal input
rlabel metal3 s 42333 47018 42399 47021 6 porb_h
port 505 nsew signal input
rlabel via2 s 52458 46824 52514 46880 6 porb_h
port 505 nsew signal input
rlabel via2 s 42338 46960 42394 47016 6 porb_h
port 505 nsew signal input
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 505 nsew signal input
rlabel metal2 s 145103 40000 145131 40174 6 porb_h
port 505 nsew signal input
rlabel metal2 s 145103 40174 145144 40202 6 porb_h
port 505 nsew signal input
rlabel metal2 s 527455 41713 527511 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 523131 41713 523187 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 472655 41713 472711 41806 6 porb_h
port 505 nsew signal input
rlabel metal2 s 468331 41713 468387 41806 6 porb_h
port 505 nsew signal input
rlabel metal2 s 472636 41806 472711 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 468312 41806 468387 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 417855 41713 417911 41820 6 porb_h
port 505 nsew signal input
rlabel metal2 s 413531 41713 413587 41820 6 porb_h
port 505 nsew signal input
rlabel metal2 s 527468 42193 527496 44134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 523144 42193 523172 44134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 527456 44134 527508 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 523132 44134 523184 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 527468 44198 527496 46854 6 porb_h
port 505 nsew signal input
rlabel metal2 s 472636 42193 472664 44338 6 porb_h
port 505 nsew signal input
rlabel metal2 s 468312 42193 468340 44338 6 porb_h
port 505 nsew signal input
rlabel metal2 s 417855 41820 417924 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 413531 41820 413600 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 363055 41713 363111 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 358731 41713 358787 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 308255 41713 308311 41806 6 porb_h
port 505 nsew signal input
rlabel metal2 s 303931 41713 303987 41806 6 porb_h
port 505 nsew signal input
rlabel metal2 s 308232 41806 308311 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 303908 41806 303987 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 199655 41713 199711 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 195331 41713 195387 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 417896 42193 417924 44202 6 porb_h
port 505 nsew signal input
rlabel metal2 s 413572 42193 413600 44202 6 porb_h
port 505 nsew signal input
rlabel metal2 s 417884 44202 417936 44266 6 porb_h
port 505 nsew signal input
rlabel metal2 s 413560 44202 413612 44266 6 porb_h
port 505 nsew signal input
rlabel metal2 s 363064 42193 363092 44270 6 porb_h
port 505 nsew signal input
rlabel metal2 s 358740 42193 358768 44270 6 porb_h
port 505 nsew signal input
rlabel metal2 s 308232 42193 308260 44202 6 porb_h
port 505 nsew signal input
rlabel metal2 s 303908 42193 303936 44202 6 porb_h
port 505 nsew signal input
rlabel metal2 s 199672 42193 199700 44134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 195348 42193 195376 44134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 145116 40202 145144 44134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 199660 44134 199712 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 195336 44134 195388 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 145104 44134 145156 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 143540 44134 143592 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 308220 44202 308272 44266 6 porb_h
port 505 nsew signal input
rlabel metal2 s 303896 44202 303948 44266 6 porb_h
port 505 nsew signal input
rlabel metal2 s 363052 44270 363104 44334 6 porb_h
port 505 nsew signal input
rlabel metal2 s 358728 44270 358780 44334 6 porb_h
port 505 nsew signal input
rlabel metal2 s 472624 44338 472676 44402 6 porb_h
port 505 nsew signal input
rlabel metal2 s 468300 44338 468352 44402 6 porb_h
port 505 nsew signal input
rlabel metal2 s 143552 44198 143580 46854 6 porb_h
port 505 nsew signal input
rlabel metal2 s 527456 46854 527508 46918 6 porb_h
port 505 nsew signal input
rlabel metal2 s 143540 46854 143592 46918 6 porb_h
port 505 nsew signal input
rlabel metal2 s 52458 46815 52514 46889 6 porb_h
port 505 nsew signal input
rlabel metal2 s 52460 46889 52512 46918 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 46922 673696 46986 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673656 46986 673684 108394 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42338 46951 42394 47025 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 108394 675444 108458 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 108394 673696 108458 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 108458 675432 108931 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 108931 675887 108945 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 108945 675887 108973 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 108973 675887 108987 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 113255 675887 113269 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 108973 675340 113269 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 113269 675887 113297 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 113297 675887 113311 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 113311 675432 113698 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 113698 675444 113762 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 113698 673696 113762 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 154059 675340 154090 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673656 113762 673684 154090 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 154131 675887 154142 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 154090 675352 154142 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 154142 675887 154154 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 154090 673696 154154 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 154154 675887 154170 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 154170 675887 154187 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 158455 675887 158494 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 154170 675340 158494 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 158494 675887 158511 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 158511 675432 158522 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 158522 675432 158578 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 158578 675444 158642 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 158578 673788 158642 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 158642 673776 199038 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 47025 42380 184303 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 184289 42193 184303 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 184303 42380 184331 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 184331 42288 188006 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 184331 42193 184345 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 188006 42472 188034 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42444 188034 42472 189110 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 188613 42193 188669 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 188669 41828 189110 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42432 189110 42484 189174 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41788 189110 41840 189174 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42444 189174 42472 197526 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 197526 42472 197554 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 199038 675444 199102 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 199038 673788 199102 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 199102 675432 199131 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 199131 675887 199158 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 199158 675887 199186 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 199186 675887 199187 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 203455 675887 203469 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 199186 675340 203458 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 203458 675352 203469 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 203469 675887 203497 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 203497 675887 203511 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 203497 675352 203522 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673828 203458 673880 203522 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 203522 675340 203580 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673840 203522 673868 243782 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 197554 42380 227582 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 227489 42193 227545 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 227545 41828 227582 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 227582 42380 227610 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 227610 42288 231827 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 231813 42193 231827 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 231827 42380 231855 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 243782 675444 243846 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673828 243782 673880 243846 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 243846 675432 244331 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 244331 675887 244345 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 244345 675887 244373 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 244373 675887 244387 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 248655 675887 248662 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 244373 675340 248662 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 248662 675887 248690 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 248690 675887 248711 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 248711 675432 249086 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 249086 675444 249150 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 249086 673696 249150 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673656 249150 673684 288798 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 231855 42380 264946 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 231855 42193 231869 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 264946 42380 264974 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 264974 42288 270830 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 270689 42193 270745 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 270745 41920 270830 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 270830 42288 270858 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 270858 42288 275182 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 275013 42193 275069 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41722 275069 41828 275074 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 275074 41828 275182 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 275182 42380 275210 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 288798 675444 288862 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 288798 673696 288862 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 288862 675432 289326 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 289326 675432 289331 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 289331 675887 289354 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 289354 675887 289387 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 293655 675887 293678 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 289354 675340 293678 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 293678 675887 293706 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 293706 675887 293711 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 293706 675340 294646 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 294646 675352 294710 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673828 294646 673880 294710 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673840 294710 673868 334222 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 275210 42380 303586 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 303586 42380 303614 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 303614 42288 313806 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 313806 42288 313834 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 313834 42288 318227 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 313834 41828 313889 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 313889 42193 313945 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 318213 42193 318227 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 318227 42380 318255 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 318255 42380 332574 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 318255 42193 318269 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 332574 42380 332602 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 334222 675444 334286 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673828 334222 673880 334286 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 334286 675432 334331 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 334331 675887 334342 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 334342 675887 334370 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 334370 675887 334387 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 334370 675340 338150 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 338150 675432 338178 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 338178 675432 338655 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 338655 675887 338711 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 338711 675432 338778 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 338778 675444 338842 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 338778 673696 338842 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673656 338842 673684 379034 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 332602 42288 356646 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41984 356646 42288 356674 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 356674 42288 361406 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41984 356674 42012 357089 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 357089 42193 357145 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41722 361406 42288 361413 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 361413 42288 361434 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 379034 675444 379098 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 379034 673696 379098 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 379098 675432 379531 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 379531 675887 379545 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 379545 675887 379573 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 379573 675887 379587 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 383855 675887 383860 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 383860 675887 383911 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 383911 675432 383982 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 379573 675340 383982 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 383982 675432 384010 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 384010 675432 384270 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 384270 675444 384334 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 384270 673696 384334 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673656 384334 673684 556582 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 361434 42288 400302 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 361434 42193 361469 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 400289 42193 400302 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 400302 42288 400330 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 400330 42288 405198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 400330 42193 400345 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 404613 42193 404669 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41722 404669 41828 404682 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 404682 41828 405198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 405198 42380 405226 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 405226 42380 419506 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 419506 42380 419534 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 419534 42288 527870 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41708 527870 42288 527898 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 527898 42288 532086 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41708 527898 42193 527917 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 527917 42193 527945 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 532086 42380 532114 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 556582 675444 556646 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 556582 675260 556646 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 556582 673696 556646 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 556646 675432 556731 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 556731 675887 556759 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 556759 675887 556787 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 556646 675248 561054 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 561054 675418 561055 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 561055 675887 561070 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 561070 675887 561082 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 561082 675887 561111 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 561082 675260 561134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 561070 673788 561134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 561134 675248 561165 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 561134 673776 601802 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 532114 42380 571254 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 532114 41920 532213 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 532213 42193 532269 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 571089 42193 571145 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41722 571145 41828 571146 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 571146 41828 571254 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 571254 42380 571282 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 571282 42288 575427 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 575413 42193 575427 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 575427 42380 575455 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 601802 675444 601866 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 601802 675260 601866 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 601802 673788 601866 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 601866 675432 601931 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 601931 675887 601959 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 601959 675887 601987 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 601866 675248 605746 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 605746 675444 605810 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 605746 675260 605810 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 605746 673788 605810 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 605810 675432 606255 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 606255 675887 606283 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 606283 675887 606311 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 605810 673776 646410 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 575455 42380 612706 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 575455 42193 575469 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 612706 42380 612734 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 612734 42288 614303 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 614289 42193 614303 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 614303 42288 614331 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 614331 42288 618718 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 614331 42193 614345 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 618613 42193 618669 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 618669 41828 618718 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 618718 42380 618746 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 646410 675444 646474 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 646410 673788 646474 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 646474 675432 646931 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 646931 675887 646959 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 646959 675887 646987 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 646474 673776 651102 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 651102 675444 651166 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 651102 673788 651166 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 651166 675432 651255 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 651255 675887 651283 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 651283 675887 651311 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 651166 673776 692038 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 618746 42380 651346 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 651346 42380 651374 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 651374 42288 657614 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41722 657478 41920 657489 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 657489 42193 657545 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 657545 41920 657614 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 657614 42288 657642 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 657642 42288 661966 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 661813 42193 661869 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 661869 41828 661966 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 661966 42380 661994 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 661994 42380 689986 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 689986 42380 690014 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 692038 675444 692102 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 692038 675260 692102 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 692038 673788 692102 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 692102 675432 692131 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 692131 675887 692172 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 692172 675887 692187 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 692102 675248 695914 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 695914 675444 695978 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 695914 675260 695978 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 695914 673788 695978 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 695978 675432 696455 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 696455 675887 696483 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 696483 675887 696511 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 695978 673776 736986 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 690014 42288 700590 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 700590 42288 700618 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 700618 42288 704942 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 700618 41920 700689 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 700689 42193 700745 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41722 700745 41920 700754 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 704942 42380 704970 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 704970 42380 728626 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 704970 41920 705013 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 705013 42193 705069 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 728626 42380 728654 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 736986 675444 737050 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 736986 675260 737050 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 736986 673788 737050 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 737050 675432 737131 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 737131 675887 737159 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 737159 675887 737187 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 737050 675248 740930 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 740930 675444 740994 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 740930 675260 740994 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 740930 673788 740994 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 740994 675432 741455 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 741455 675887 741483 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 741483 675887 741511 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 740994 673776 781594 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 728654 42288 743702 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 743702 42288 743730 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 743730 42288 747946 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 743730 41828 743889 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 743889 42193 743945 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 747946 42472 747974 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 781594 675444 781658 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 781594 675260 781658 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 781594 673788 781658 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 781658 675432 782131 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 782131 675887 782159 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 782159 675887 782187 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 781658 675248 785946 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 785946 675444 786010 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 785946 675260 786010 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 785946 673788 786010 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 786010 675432 786455 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 786455 675887 786483 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 786483 675887 786511 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 786010 673776 870810 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42444 747974 42472 787238 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 747974 41920 748213 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 748213 42193 748269 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41722 787086 41920 787089 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 787089 42193 787145 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 787145 41920 787222 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 787222 42288 787238 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42432 787238 42484 787302 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 787238 42300 787250 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42248 787250 42300 787302 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 787302 42288 791438 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 791413 42193 791438 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 791438 42288 791466 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 791466 42193 791469 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 870810 675444 870874 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 870810 673788 870874 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 870874 675432 871331 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 871331 675887 871345 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 871345 675887 871373 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 871373 675887 871387 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 875655 675887 875669 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 871373 675340 875669 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 875669 675887 875697 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 875697 675887 875711 6 porb_h
port 505 nsew signal input
rlabel via1 s 527456 44140 527508 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 523132 44140 523184 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 417884 44208 417936 44260 6 porb_h
port 505 nsew signal input
rlabel via1 s 413560 44208 413612 44260 6 porb_h
port 505 nsew signal input
rlabel via1 s 472624 44344 472676 44396 6 porb_h
port 505 nsew signal input
rlabel via1 s 468300 44344 468352 44396 6 porb_h
port 505 nsew signal input
rlabel via1 s 363052 44276 363104 44328 6 porb_h
port 505 nsew signal input
rlabel via1 s 358728 44276 358780 44328 6 porb_h
port 505 nsew signal input
rlabel via1 s 308220 44208 308272 44260 6 porb_h
port 505 nsew signal input
rlabel via1 s 303896 44208 303948 44260 6 porb_h
port 505 nsew signal input
rlabel via1 s 199660 44140 199712 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 195336 44140 195388 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 145104 44140 145156 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 143540 44140 143592 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 527456 46860 527508 46912 6 porb_h
port 505 nsew signal input
rlabel via1 s 143540 46860 143592 46912 6 porb_h
port 505 nsew signal input
rlabel via1 s 52460 46860 52512 46912 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 46928 673696 46980 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 108400 675444 108452 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 108400 673696 108452 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 113704 675444 113756 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 113704 673696 113756 6 porb_h
port 505 nsew signal input
rlabel via1 s 675300 154096 675352 154148 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 154096 673696 154148 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 158584 675444 158636 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 158584 673788 158636 6 porb_h
port 505 nsew signal input
rlabel via1 s 42432 189116 42484 189168 6 porb_h
port 505 nsew signal input
rlabel via1 s 41788 189116 41840 189168 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 199044 675444 199096 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 199044 673788 199096 6 porb_h
port 505 nsew signal input
rlabel via1 s 675300 203464 675352 203516 6 porb_h
port 505 nsew signal input
rlabel via1 s 673828 203464 673880 203516 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 243788 675444 243840 6 porb_h
port 505 nsew signal input
rlabel via1 s 673828 243788 673880 243840 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 249092 675444 249144 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 249092 673696 249144 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 288804 675444 288856 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 288804 673696 288856 6 porb_h
port 505 nsew signal input
rlabel via1 s 675300 294652 675352 294704 6 porb_h
port 505 nsew signal input
rlabel via1 s 673828 294652 673880 294704 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 334228 675444 334280 6 porb_h
port 505 nsew signal input
rlabel via1 s 673828 334228 673880 334280 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 338784 675444 338836 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 338784 673696 338836 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 379040 675444 379092 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 379040 673696 379092 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 384276 675444 384328 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 384276 673696 384328 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 556588 675444 556640 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 556588 675260 556640 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 556588 673696 556640 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 561076 675260 561128 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 561076 673788 561128 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 601808 675444 601860 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 601808 675260 601860 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 601808 673788 601860 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 605752 675444 605804 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 605752 675260 605804 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 605752 673788 605804 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 646416 675444 646468 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 646416 673788 646468 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 651108 675444 651160 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 651108 673788 651160 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 692044 675444 692096 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 692044 675260 692096 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 692044 673788 692096 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 695920 675444 695972 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 695920 675260 695972 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 695920 673788 695972 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 736992 675444 737044 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 736992 675260 737044 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 736992 673788 737044 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 740936 675444 740988 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 740936 675260 740988 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 740936 673788 740988 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 781600 675444 781652 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 781600 675260 781652 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 781600 673788 781652 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 785952 675444 786004 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 785952 675260 786004 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 785952 673788 786004 6 porb_h
port 505 nsew signal input
rlabel via1 s 42432 787244 42484 787296 6 porb_h
port 505 nsew signal input
rlabel via1 s 42248 787244 42300 787296 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 870816 675444 870868 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 870816 673788 870868 6 porb_h
port 505 nsew signal input
rlabel metal1 s 527450 44140 527514 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 523126 44140 523190 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 199654 44140 199718 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 195330 44140 195394 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 145098 44140 145162 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 143534 44140 143598 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 523126 44152 527514 44180 6 porb_h
port 505 nsew signal input
rlabel metal1 s 527450 44180 527514 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 523126 44180 523190 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 143534 44152 207014 44180 6 porb_h
port 505 nsew signal input
rlabel metal1 s 523144 44192 523172 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 417878 44208 417942 44220 6 porb_h
port 505 nsew signal input
rlabel metal1 s 413554 44208 413618 44220 6 porb_h
port 505 nsew signal input
rlabel metal1 s 308214 44208 308278 44220 6 porb_h
port 505 nsew signal input
rlabel metal1 s 303890 44208 303954 44220 6 porb_h
port 505 nsew signal input
rlabel metal1 s 206986 44180 207014 44220 6 porb_h
port 505 nsew signal input
rlabel metal1 s 199654 44180 199718 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 195330 44180 195394 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 145098 44180 145162 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 143534 44180 143598 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 363340 44220 417942 44248 6 porb_h
port 505 nsew signal input
rlabel metal1 s 417878 44248 417942 44260 6 porb_h
port 505 nsew signal input
rlabel metal1 s 413554 44248 413618 44260 6 porb_h
port 505 nsew signal input
rlabel metal1 s 477466 44288 523172 44316 6 porb_h
port 505 nsew signal input
rlabel metal1 s 477466 44316 477494 44356 6 porb_h
port 505 nsew signal input
rlabel metal1 s 472618 44344 472682 44356 6 porb_h
port 505 nsew signal input
rlabel metal1 s 468294 44344 468358 44356 6 porb_h
port 505 nsew signal input
rlabel metal1 s 417896 44260 417924 44356 6 porb_h
port 505 nsew signal input
rlabel metal1 s 363340 44248 363368 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 206986 44220 349936 44248 6 porb_h
port 505 nsew signal input
rlabel metal1 s 363046 44276 363110 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 358722 44276 358786 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 349908 44248 349936 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 308214 44248 308278 44260 6 porb_h
port 505 nsew signal input
rlabel metal1 s 303890 44248 303954 44260 6 porb_h
port 505 nsew signal input
rlabel metal1 s 349908 44288 363368 44316 6 porb_h
port 505 nsew signal input
rlabel metal1 s 363046 44316 363110 44328 6 porb_h
port 505 nsew signal input
rlabel metal1 s 358722 44316 358786 44328 6 porb_h
port 505 nsew signal input
rlabel metal1 s 417896 44356 477494 44384 6 porb_h
port 505 nsew signal input
rlabel metal1 s 472618 44384 472682 44396 6 porb_h
port 505 nsew signal input
rlabel metal1 s 468294 44384 468358 44396 6 porb_h
port 505 nsew signal input
rlabel metal1 s 527450 46860 527514 46912 6 porb_h
port 505 nsew signal input
rlabel metal1 s 143534 46860 143598 46872 6 porb_h
port 505 nsew signal input
rlabel metal1 s 52454 46860 52518 46872 6 porb_h
port 505 nsew signal input
rlabel metal1 s 52454 46872 143598 46900 6 porb_h
port 505 nsew signal input
rlabel metal1 s 143534 46900 143598 46912 6 porb_h
port 505 nsew signal input
rlabel metal1 s 52454 46900 52518 46912 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 46928 673702 46940 6 porb_h
port 505 nsew signal input
rlabel metal1 s 527468 46912 527496 46940 6 porb_h
port 505 nsew signal input
rlabel metal1 s 527468 46940 673702 46968 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 46968 673702 46980 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 108400 675450 108412 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 108400 673702 108412 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 108412 675450 108440 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 108440 675450 108452 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 108440 673702 108452 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 113704 675450 113716 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 113704 673702 113716 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 113716 675450 113744 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 113744 675450 113756 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 113744 673702 113756 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 154096 675358 154108 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 154096 673702 154108 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 154108 675358 154136 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 154136 675358 154148 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 154136 673702 154148 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 158584 675450 158596 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 158584 673794 158596 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 158596 675450 158624 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 158624 675450 158636 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 158624 673794 158636 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42426 189116 42490 189128 6 porb_h
port 505 nsew signal input
rlabel metal1 s 41782 189116 41846 189128 6 porb_h
port 505 nsew signal input
rlabel metal1 s 41782 189128 42490 189156 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42426 189156 42490 189168 6 porb_h
port 505 nsew signal input
rlabel metal1 s 41782 189156 41846 189168 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 199044 675450 199056 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 199044 673794 199056 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 199056 675450 199084 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 199084 675450 199096 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 199084 673794 199096 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 203464 675358 203476 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 203464 673886 203476 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 203476 675358 203504 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 203504 675358 203516 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 203504 673886 203516 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 243788 675450 243800 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 243788 673886 243800 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 243800 675450 243828 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 243828 675450 243840 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 243828 673886 243840 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 249092 675450 249104 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 249092 673702 249104 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 249104 675450 249132 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 249132 675450 249144 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 249132 673702 249144 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 288804 675450 288816 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 288804 673702 288816 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 288816 675450 288844 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 288844 675450 288856 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 288844 673702 288856 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 294652 675358 294664 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 294652 673886 294664 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 294664 675358 294692 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 294692 675358 294704 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 294692 673886 294704 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 334228 675450 334240 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 334228 673886 334240 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 334240 675450 334268 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 334268 675450 334280 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 334268 673886 334280 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 338784 675450 338796 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 338784 673702 338796 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 338796 675450 338824 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 338824 675450 338836 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 338824 673702 338836 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 379040 675450 379052 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 379040 673702 379052 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 379052 675450 379080 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 379080 675450 379092 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 379080 673702 379092 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 384276 675450 384288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 384276 673702 384288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 384288 675450 384316 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 384316 675450 384328 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 384316 673702 384328 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 556588 675450 556600 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 556588 675266 556600 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 556588 673702 556600 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 556600 675450 556628 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 556628 675450 556640 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 556628 675266 556640 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 556628 673702 556640 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 561076 675266 561088 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 561076 673794 561088 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 561088 675266 561116 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 561116 675266 561128 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 561116 673794 561128 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 601808 675450 601820 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 601808 675266 601820 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 601808 673794 601820 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 601820 675450 601848 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 601848 675450 601860 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 601848 675266 601860 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 601848 673794 601860 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 605752 675450 605764 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 605752 675266 605764 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 605752 673794 605764 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 605764 675450 605792 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 605792 675450 605804 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 605792 675266 605804 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 605792 673794 605804 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 646416 675450 646428 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 646416 673794 646428 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 646428 675450 646456 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 646456 675450 646468 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 646456 673794 646468 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 651108 675450 651120 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 651108 673794 651120 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 651120 675450 651148 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 651148 675450 651160 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 651148 673794 651160 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 692044 675450 692056 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 692044 675266 692056 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 692044 673794 692056 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 692056 675450 692084 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 692084 675450 692096 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 692084 675266 692096 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 692084 673794 692096 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 695920 675450 695932 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 695920 675266 695932 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 695920 673794 695932 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 695932 675450 695960 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 695960 675450 695972 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 695960 675266 695972 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 695960 673794 695972 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 736992 675450 737004 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 736992 675266 737004 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 736992 673794 737004 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 737004 675450 737032 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 737032 675450 737044 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 737032 675266 737044 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 737032 673794 737044 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 740936 675450 740948 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 740936 675266 740948 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 740936 673794 740948 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 740948 675450 740976 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 740976 675450 740988 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 740976 675266 740988 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 740976 673794 740988 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 781600 675450 781612 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 781600 675266 781612 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 781600 673794 781612 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 781612 675450 781640 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 781640 675450 781652 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 781640 675266 781652 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 781640 673794 781652 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 785952 675450 785964 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 785952 675266 785964 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 785952 673794 785964 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 785964 675450 785992 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 785992 675450 786004 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 785992 675266 786004 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 785992 673794 786004 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42426 787244 42490 787256 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42242 787244 42306 787256 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42242 787256 42490 787284 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42426 787284 42490 787296 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42242 787284 42306 787296 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 870816 675450 870828 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 870816 673794 870828 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 870828 675450 870856 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 870856 675450 870868 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 870856 673794 870868 6 porb_h
port 505 nsew signal input
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 506 nsew signal input
rlabel metal3 s 141820 37046 141966 37818 6 resetb_core_h
port 507 nsew signal output
rlabel metal3 s 141667 37818 141966 37911 6 resetb_core_h
port 507 nsew signal output
rlabel metal3 s 141873 37911 141966 37971 6 resetb_core_h
port 507 nsew signal output
rlabel metal3 s 141667 37911 141820 37971 6 resetb_core_h
port 507 nsew signal output
rlabel metal3 s 141667 37971 141873 38031 6 resetb_core_h
port 507 nsew signal output
rlabel metal3 s 141667 38031 141813 40000 6 resetb_core_h
port 507 nsew signal output
rlabel metal4 s 93607 36323 132793 37013 6 vdda
port 508 nsew signal bidirectional
rlabel metal4 s 93546 28653 192982 28719 6 vssa
port 509 nsew signal bidirectional
rlabel metal4 s 93546 30753 132854 30762 6 vssd
port 510 nsew signal bidirectional
rlabel metal4 s 93546 30762 132869 31674 6 vssd
port 510 nsew signal bidirectional
rlabel metal4 s 93546 31674 132854 31683 6 vssd
port 510 nsew signal bidirectional
rlabel metal3 s 630944 997600 635944 1014070 6 mprj_analog[1]
port 511 nsew signal bidirectional
rlabel metal5 s 627410 1018624 639578 1030789 6 mprj_io[15]
port 512 nsew signal bidirectional
rlabel metal3 s 529144 997600 534144 1014070 6 mprj_analog[2]
port 513 nsew signal bidirectional
rlabel metal5 s 525610 1018624 537778 1030789 6 mprj_io[16]
port 514 nsew signal bidirectional
rlabel metal3 s 477744 997600 482744 1014070 6 mprj_analog[3]
port 515 nsew signal bidirectional
rlabel metal5 s 474210 1018624 486378 1030789 6 mprj_io[17]
port 516 nsew signal bidirectional
rlabel metal3 s 388744 997600 393744 1014070 6 mprj_analog[4]
port 517 nsew signal bidirectional
rlabel metal5 s 385210 1018624 397378 1030789 6 mprj_io[18]
port 518 nsew signal bidirectional
rlabel metal3 s 677600 943200 680737 957522 6 mprj_analog[0]
port 519 nsew signal bidirectional
rlabel metal2 s 677600 952742 682732 957522 6 mprj_clamp_high[0]
port 520 nsew signal input
rlabel metal2 s 677600 962721 678011 967501 6 mprj_clamp_low[0]
port 521 nsew signal input
rlabel metal5 s 698624 954022 710789 966190 6 mprj_io[14]
port 522 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1_pad
port 523 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1_pad
port 524 nsew signal bidirectional
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_pad2
port 525 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1_pad
port 526 nsew signal bidirectional
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_pad2
port 527 nsew signal bidirectional
rlabel metal4 s 679377 430346 680307 460054 6 vccd1
port 528 nsew signal bidirectional
rlabel metal4 s 680587 430407 681277 459993 6 vdda1
port 529 nsew signal bidirectional
rlabel metal4 s 688881 430346 688947 554382 6 vssa1
port 530 nsew signal bidirectional
rlabel metal3 s 678000 469900 685920 474700 6 vssd1
port 531 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1_pad
port 532 nsew signal bidirectional
rlabel metal3 s 183944 997600 188944 1014070 6 mprj_analog[7]
port 533 nsew signal bidirectional
rlabel metal5 s 180410 1018624 192578 1030789 6 mprj_io[21]
port 534 nsew signal bidirectional
rlabel metal3 s 132544 997600 137544 1014070 6 mprj_analog[8]
port 535 nsew signal bidirectional
rlabel metal5 s 129010 1018624 141178 1030789 6 mprj_io[22]
port 536 nsew signal bidirectional
rlabel metal3 s 81144 997600 86144 1014070 6 mprj_analog[9]
port 537 nsew signal bidirectional
rlabel metal5 s 77610 1018624 89778 1030789 6 mprj_io[23]
port 538 nsew signal bidirectional
rlabel metal3 s 23530 959144 40000 964144 6 mprj_analog[10]
port 539 nsew signal bidirectional
rlabel metal5 s 6811 955610 18976 967778 6 mprj_io[24]
port 540 nsew signal bidirectional
rlabel metal3 s 292078 997600 306400 1000737 6 mprj_analog[5]
port 541 nsew signal bidirectional
rlabel metal2 s 292078 997600 296858 1002732 6 mprj_clamp_high[1]
port 542 nsew signal input
rlabel metal2 s 282099 997600 286879 998011 6 mprj_clamp_low[1]
port 543 nsew signal input
rlabel metal5 s 283410 1018624 295578 1030789 6 mprj_io[19]
port 544 nsew signal bidirectional
rlabel metal3 s 240478 997600 254800 1000737 6 mprj_analog[6]
port 545 nsew signal bidirectional
rlabel metal2 s 240478 997600 245258 1002732 6 mprj_clamp_high[2]
port 546 nsew signal input
rlabel metal2 s 230499 997600 235279 998011 6 mprj_clamp_low[2]
port 547 nsew signal input
rlabel metal5 s 231810 1018624 243978 1030789 6 mprj_io[20]
port 548 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2_pad
port 549 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2_pad
port 550 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2_pad
port 551 nsew signal bidirectional
rlabel metal4 s 38503 455546 39593 483254 6 vccd
port 552 nsew signal bidirectional
rlabel metal4 s 37293 455546 38223 483254 6 vccd2
port 553 nsew signal bidirectional
rlabel metal4 s 36323 455607 37013 483193 6 vdda2
port 554 nsew signal bidirectional
rlabel metal4 s 32933 455546 33623 483254 6 vddio
port 555 nsew signal bidirectional
rlabel metal4 s 28653 407018 28719 525722 6 vssa2
port 556 nsew signal bidirectional
rlabel metal3 s 31680 440900 39600 445700 6 vssd2
port 557 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2_pad
port 558 nsew signal bidirectional
rlabel metal4 s 0 455546 4843 455800 6 vssio
port 559 nsew signal bidirectional
rlabel metal4 s 7 455800 4843 456093 6 vssio
port 559 nsew signal bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 717600 1037600
string LEFview TRUE
string GDS_FILE /project/openlane/chip_io_alt/runs/chip_io_alt/results/magic/chip_io_alt.gds
string GDS_END 36735404
string GDS_START 36371924
<< end >>

