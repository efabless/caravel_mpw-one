VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM
  CLASS BLOCK ;
  FOREIGN DFFRAM ;
  ORIGIN 0.000 0.000 ;
  SIZE 745.115 BY 525.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.400 19.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.400 56.400 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.400 93.800 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.400 131.200 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 2.400 168.600 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 2.400 206.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 2.400 243.400 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 2.400 281.480 ;
    END
  END A[7]
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 2.400 318.880 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 522.600 11.870 525.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 245.730 522.600 246.010 525.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.190 522.600 269.470 525.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 292.650 522.600 292.930 525.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.110 522.600 316.390 525.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 339.570 522.600 339.850 525.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.030 522.600 363.310 525.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.490 522.600 386.770 525.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 409.490 522.600 409.770 525.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.950 522.600 433.230 525.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 456.410 522.600 456.690 525.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 522.600 34.870 525.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.870 522.600 480.150 525.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 503.330 522.600 503.610 525.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 526.790 522.600 527.070 525.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 550.250 522.600 550.530 525.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 573.710 522.600 573.990 525.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.170 522.600 597.450 525.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.630 522.600 620.910 525.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.090 522.600 644.370 525.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 667.550 522.600 667.830 525.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 691.010 522.600 691.290 525.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 522.600 58.330 525.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.470 522.600 714.750 525.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 737.930 522.600 738.210 525.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 522.600 81.790 525.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 522.600 105.250 525.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.430 522.600 128.710 525.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.890 522.600 152.170 525.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 175.350 522.600 175.630 525.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 198.810 522.600 199.090 525.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.270 522.600 222.550 525.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 2.400 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 2.400 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 2.400 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 2.400 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 2.400 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 2.400 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 2.400 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 2.400 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 2.400 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 2.400 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 2.400 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 2.400 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 2.400 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 2.400 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.710 0.000 573.990 2.400 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 597.170 0.000 597.450 2.400 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 2.400 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 2.400 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 2.400 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 2.400 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.400 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 2.400 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 737.930 0.000 738.210 2.400 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 2.400 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 2.400 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 2.400 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 2.400 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 2.400 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 2.400 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 2.400 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.280 2.400 505.880 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 2.400 356.280 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 2.400 393.680 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 2.400 431.080 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 2.400 468.480 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 514.320 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 514.320 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 745.055 514.165 ;
      LAYER met1 ;
        RECT 5.520 9.900 745.115 514.320 ;
      LAYER met2 ;
        RECT 6.990 522.320 11.310 522.600 ;
        RECT 12.150 522.320 34.310 522.600 ;
        RECT 35.150 522.320 57.770 522.600 ;
        RECT 58.610 522.320 81.230 522.600 ;
        RECT 82.070 522.320 104.690 522.600 ;
        RECT 105.530 522.320 128.150 522.600 ;
        RECT 128.990 522.320 151.610 522.600 ;
        RECT 152.450 522.320 175.070 522.600 ;
        RECT 175.910 522.320 198.530 522.600 ;
        RECT 199.370 522.320 221.990 522.600 ;
        RECT 222.830 522.320 245.450 522.600 ;
        RECT 246.290 522.320 268.910 522.600 ;
        RECT 269.750 522.320 292.370 522.600 ;
        RECT 293.210 522.320 315.830 522.600 ;
        RECT 316.670 522.320 339.290 522.600 ;
        RECT 340.130 522.320 362.750 522.600 ;
        RECT 363.590 522.320 386.210 522.600 ;
        RECT 387.050 522.320 409.210 522.600 ;
        RECT 410.050 522.320 432.670 522.600 ;
        RECT 433.510 522.320 456.130 522.600 ;
        RECT 456.970 522.320 479.590 522.600 ;
        RECT 480.430 522.320 503.050 522.600 ;
        RECT 503.890 522.320 526.510 522.600 ;
        RECT 527.350 522.320 549.970 522.600 ;
        RECT 550.810 522.320 573.430 522.600 ;
        RECT 574.270 522.320 596.890 522.600 ;
        RECT 597.730 522.320 620.350 522.600 ;
        RECT 621.190 522.320 643.810 522.600 ;
        RECT 644.650 522.320 667.270 522.600 ;
        RECT 668.110 522.320 690.730 522.600 ;
        RECT 691.570 522.320 714.190 522.600 ;
        RECT 715.030 522.320 737.650 522.600 ;
        RECT 738.490 522.320 742.800 522.600 ;
        RECT 6.990 2.680 742.800 522.320 ;
        RECT 6.990 2.400 11.310 2.680 ;
        RECT 12.150 2.400 34.310 2.680 ;
        RECT 35.150 2.400 57.770 2.680 ;
        RECT 58.610 2.400 81.230 2.680 ;
        RECT 82.070 2.400 104.690 2.680 ;
        RECT 105.530 2.400 128.150 2.680 ;
        RECT 128.990 2.400 151.610 2.680 ;
        RECT 152.450 2.400 175.070 2.680 ;
        RECT 175.910 2.400 198.530 2.680 ;
        RECT 199.370 2.400 221.990 2.680 ;
        RECT 222.830 2.400 245.450 2.680 ;
        RECT 246.290 2.400 268.910 2.680 ;
        RECT 269.750 2.400 292.370 2.680 ;
        RECT 293.210 2.400 315.830 2.680 ;
        RECT 316.670 2.400 339.290 2.680 ;
        RECT 340.130 2.400 362.750 2.680 ;
        RECT 363.590 2.400 386.210 2.680 ;
        RECT 387.050 2.400 409.210 2.680 ;
        RECT 410.050 2.400 432.670 2.680 ;
        RECT 433.510 2.400 456.130 2.680 ;
        RECT 456.970 2.400 479.590 2.680 ;
        RECT 480.430 2.400 503.050 2.680 ;
        RECT 503.890 2.400 526.510 2.680 ;
        RECT 527.350 2.400 549.970 2.680 ;
        RECT 550.810 2.400 573.430 2.680 ;
        RECT 574.270 2.400 596.890 2.680 ;
        RECT 597.730 2.400 620.350 2.680 ;
        RECT 621.190 2.400 643.810 2.680 ;
        RECT 644.650 2.400 667.270 2.680 ;
        RECT 668.110 2.400 690.730 2.680 ;
        RECT 691.570 2.400 714.190 2.680 ;
        RECT 715.030 2.400 737.650 2.680 ;
        RECT 738.490 2.400 742.800 2.680 ;
      LAYER met3 ;
        RECT 2.400 506.280 735.935 514.245 ;
        RECT 2.800 504.880 735.935 506.280 ;
        RECT 2.400 468.880 735.935 504.880 ;
        RECT 2.800 467.480 735.935 468.880 ;
        RECT 2.400 431.480 735.935 467.480 ;
        RECT 2.800 430.080 735.935 431.480 ;
        RECT 2.400 394.080 735.935 430.080 ;
        RECT 2.800 392.680 735.935 394.080 ;
        RECT 2.400 356.680 735.935 392.680 ;
        RECT 2.800 355.280 735.935 356.680 ;
        RECT 2.400 319.280 735.935 355.280 ;
        RECT 2.800 317.880 735.935 319.280 ;
        RECT 2.400 281.880 735.935 317.880 ;
        RECT 2.800 280.480 735.935 281.880 ;
        RECT 2.400 243.800 735.935 280.480 ;
        RECT 2.800 242.400 735.935 243.800 ;
        RECT 2.400 206.400 735.935 242.400 ;
        RECT 2.800 205.000 735.935 206.400 ;
        RECT 2.400 169.000 735.935 205.000 ;
        RECT 2.800 167.600 735.935 169.000 ;
        RECT 2.400 131.600 735.935 167.600 ;
        RECT 2.800 130.200 735.935 131.600 ;
        RECT 2.400 94.200 735.935 130.200 ;
        RECT 2.800 92.800 735.935 94.200 ;
        RECT 2.400 56.800 735.935 92.800 ;
        RECT 2.800 55.400 735.935 56.800 ;
        RECT 2.400 19.400 735.935 55.400 ;
        RECT 2.800 18.000 735.935 19.400 ;
        RECT 2.400 10.715 735.935 18.000 ;
      LAYER met4 ;
        RECT 96.895 10.640 97.440 514.320 ;
        RECT 99.840 10.640 713.840 514.320 ;
  END
END DFFRAM
END LIBRARY

