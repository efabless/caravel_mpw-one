magic
tech sky130A
magscale 1 2
timestamp 1622487809
<< obsli1 >>
rect 1104 1309 428967 171683
<< obsm1 >>
rect 290 1300 429626 171964
<< metal2 >>
rect 294 171200 350 172000
rect 938 171200 994 172000
rect 1582 171200 1638 172000
rect 2226 171200 2282 172000
rect 2870 171200 2926 172000
rect 3514 171200 3570 172000
rect 4158 171200 4214 172000
rect 4802 171200 4858 172000
rect 5446 171200 5502 172000
rect 6090 171200 6146 172000
rect 6734 171200 6790 172000
rect 7378 171200 7434 172000
rect 8022 171200 8078 172000
rect 8666 171200 8722 172000
rect 9310 171200 9366 172000
rect 9954 171200 10010 172000
rect 10598 171200 10654 172000
rect 11334 171200 11390 172000
rect 11978 171200 12034 172000
rect 12622 171200 12678 172000
rect 13266 171200 13322 172000
rect 13910 171200 13966 172000
rect 14554 171200 14610 172000
rect 15198 171200 15254 172000
rect 15842 171200 15898 172000
rect 16486 171200 16542 172000
rect 17130 171200 17186 172000
rect 17774 171200 17830 172000
rect 18418 171200 18474 172000
rect 19062 171200 19118 172000
rect 19706 171200 19762 172000
rect 20350 171200 20406 172000
rect 20994 171200 21050 172000
rect 21638 171200 21694 172000
rect 22374 171200 22430 172000
rect 23018 171200 23074 172000
rect 23662 171200 23718 172000
rect 24306 171200 24362 172000
rect 24950 171200 25006 172000
rect 25594 171200 25650 172000
rect 26238 171200 26294 172000
rect 26882 171200 26938 172000
rect 27526 171200 27582 172000
rect 28170 171200 28226 172000
rect 28814 171200 28870 172000
rect 29458 171200 29514 172000
rect 30102 171200 30158 172000
rect 30746 171200 30802 172000
rect 31390 171200 31446 172000
rect 32034 171200 32090 172000
rect 32770 171200 32826 172000
rect 33414 171200 33470 172000
rect 34058 171200 34114 172000
rect 34702 171200 34758 172000
rect 35346 171200 35402 172000
rect 35990 171200 36046 172000
rect 36634 171200 36690 172000
rect 37278 171200 37334 172000
rect 37922 171200 37978 172000
rect 38566 171200 38622 172000
rect 39210 171200 39266 172000
rect 39854 171200 39910 172000
rect 40498 171200 40554 172000
rect 41142 171200 41198 172000
rect 41786 171200 41842 172000
rect 42430 171200 42486 172000
rect 43074 171200 43130 172000
rect 43810 171200 43866 172000
rect 44454 171200 44510 172000
rect 45098 171200 45154 172000
rect 45742 171200 45798 172000
rect 46386 171200 46442 172000
rect 47030 171200 47086 172000
rect 47674 171200 47730 172000
rect 48318 171200 48374 172000
rect 48962 171200 49018 172000
rect 49606 171200 49662 172000
rect 50250 171200 50306 172000
rect 50894 171200 50950 172000
rect 51538 171200 51594 172000
rect 52182 171200 52238 172000
rect 52826 171200 52882 172000
rect 53470 171200 53526 172000
rect 54206 171200 54262 172000
rect 54850 171200 54906 172000
rect 55494 171200 55550 172000
rect 56138 171200 56194 172000
rect 56782 171200 56838 172000
rect 57426 171200 57482 172000
rect 58070 171200 58126 172000
rect 58714 171200 58770 172000
rect 59358 171200 59414 172000
rect 60002 171200 60058 172000
rect 60646 171200 60702 172000
rect 61290 171200 61346 172000
rect 61934 171200 61990 172000
rect 62578 171200 62634 172000
rect 63222 171200 63278 172000
rect 63866 171200 63922 172000
rect 64510 171200 64566 172000
rect 65246 171200 65302 172000
rect 65890 171200 65946 172000
rect 66534 171200 66590 172000
rect 67178 171200 67234 172000
rect 67822 171200 67878 172000
rect 68466 171200 68522 172000
rect 69110 171200 69166 172000
rect 69754 171200 69810 172000
rect 70398 171200 70454 172000
rect 71042 171200 71098 172000
rect 71686 171200 71742 172000
rect 72330 171200 72386 172000
rect 72974 171200 73030 172000
rect 73618 171200 73674 172000
rect 74262 171200 74318 172000
rect 74906 171200 74962 172000
rect 75642 171200 75698 172000
rect 76286 171200 76342 172000
rect 76930 171200 76986 172000
rect 77574 171200 77630 172000
rect 78218 171200 78274 172000
rect 78862 171200 78918 172000
rect 79506 171200 79562 172000
rect 80150 171200 80206 172000
rect 80794 171200 80850 172000
rect 81438 171200 81494 172000
rect 82082 171200 82138 172000
rect 82726 171200 82782 172000
rect 83370 171200 83426 172000
rect 84014 171200 84070 172000
rect 84658 171200 84714 172000
rect 85302 171200 85358 172000
rect 85946 171200 86002 172000
rect 86682 171200 86738 172000
rect 87326 171200 87382 172000
rect 87970 171200 88026 172000
rect 88614 171200 88670 172000
rect 89258 171200 89314 172000
rect 89902 171200 89958 172000
rect 90546 171200 90602 172000
rect 91190 171200 91246 172000
rect 91834 171200 91890 172000
rect 92478 171200 92534 172000
rect 93122 171200 93178 172000
rect 93766 171200 93822 172000
rect 94410 171200 94466 172000
rect 95054 171200 95110 172000
rect 95698 171200 95754 172000
rect 96342 171200 96398 172000
rect 97078 171200 97134 172000
rect 97722 171200 97778 172000
rect 98366 171200 98422 172000
rect 99010 171200 99066 172000
rect 99654 171200 99710 172000
rect 100298 171200 100354 172000
rect 100942 171200 100998 172000
rect 101586 171200 101642 172000
rect 102230 171200 102286 172000
rect 102874 171200 102930 172000
rect 103518 171200 103574 172000
rect 104162 171200 104218 172000
rect 104806 171200 104862 172000
rect 105450 171200 105506 172000
rect 106094 171200 106150 172000
rect 106738 171200 106794 172000
rect 107382 171200 107438 172000
rect 108118 171200 108174 172000
rect 108762 171200 108818 172000
rect 109406 171200 109462 172000
rect 110050 171200 110106 172000
rect 110694 171200 110750 172000
rect 111338 171200 111394 172000
rect 111982 171200 112038 172000
rect 112626 171200 112682 172000
rect 113270 171200 113326 172000
rect 113914 171200 113970 172000
rect 114558 171200 114614 172000
rect 115202 171200 115258 172000
rect 115846 171200 115902 172000
rect 116490 171200 116546 172000
rect 117134 171200 117190 172000
rect 117778 171200 117834 172000
rect 118422 171200 118478 172000
rect 119158 171200 119214 172000
rect 119802 171200 119858 172000
rect 120446 171200 120502 172000
rect 121090 171200 121146 172000
rect 121734 171200 121790 172000
rect 122378 171200 122434 172000
rect 123022 171200 123078 172000
rect 123666 171200 123722 172000
rect 124310 171200 124366 172000
rect 124954 171200 125010 172000
rect 125598 171200 125654 172000
rect 126242 171200 126298 172000
rect 126886 171200 126942 172000
rect 127530 171200 127586 172000
rect 128174 171200 128230 172000
rect 128818 171200 128874 172000
rect 129554 171200 129610 172000
rect 130198 171200 130254 172000
rect 130842 171200 130898 172000
rect 131486 171200 131542 172000
rect 132130 171200 132186 172000
rect 132774 171200 132830 172000
rect 133418 171200 133474 172000
rect 134062 171200 134118 172000
rect 134706 171200 134762 172000
rect 135350 171200 135406 172000
rect 135994 171200 136050 172000
rect 136638 171200 136694 172000
rect 137282 171200 137338 172000
rect 137926 171200 137982 172000
rect 138570 171200 138626 172000
rect 139214 171200 139270 172000
rect 139858 171200 139914 172000
rect 140594 171200 140650 172000
rect 141238 171200 141294 172000
rect 141882 171200 141938 172000
rect 142526 171200 142582 172000
rect 143170 171200 143226 172000
rect 143814 171200 143870 172000
rect 144458 171200 144514 172000
rect 145102 171200 145158 172000
rect 145746 171200 145802 172000
rect 146390 171200 146446 172000
rect 147034 171200 147090 172000
rect 147678 171200 147734 172000
rect 148322 171200 148378 172000
rect 148966 171200 149022 172000
rect 149610 171200 149666 172000
rect 150254 171200 150310 172000
rect 150990 171200 151046 172000
rect 151634 171200 151690 172000
rect 152278 171200 152334 172000
rect 152922 171200 152978 172000
rect 153566 171200 153622 172000
rect 154210 171200 154266 172000
rect 154854 171200 154910 172000
rect 155498 171200 155554 172000
rect 156142 171200 156198 172000
rect 156786 171200 156842 172000
rect 157430 171200 157486 172000
rect 158074 171200 158130 172000
rect 158718 171200 158774 172000
rect 159362 171200 159418 172000
rect 160006 171200 160062 172000
rect 160650 171200 160706 172000
rect 161294 171200 161350 172000
rect 162030 171200 162086 172000
rect 162674 171200 162730 172000
rect 163318 171200 163374 172000
rect 163962 171200 164018 172000
rect 164606 171200 164662 172000
rect 165250 171200 165306 172000
rect 165894 171200 165950 172000
rect 166538 171200 166594 172000
rect 167182 171200 167238 172000
rect 167826 171200 167882 172000
rect 168470 171200 168526 172000
rect 169114 171200 169170 172000
rect 169758 171200 169814 172000
rect 170402 171200 170458 172000
rect 171046 171200 171102 172000
rect 171690 171200 171746 172000
rect 172426 171200 172482 172000
rect 173070 171200 173126 172000
rect 173714 171200 173770 172000
rect 174358 171200 174414 172000
rect 175002 171200 175058 172000
rect 175646 171200 175702 172000
rect 176290 171200 176346 172000
rect 176934 171200 176990 172000
rect 177578 171200 177634 172000
rect 178222 171200 178278 172000
rect 178866 171200 178922 172000
rect 179510 171200 179566 172000
rect 180154 171200 180210 172000
rect 180798 171200 180854 172000
rect 181442 171200 181498 172000
rect 182086 171200 182142 172000
rect 182730 171200 182786 172000
rect 183466 171200 183522 172000
rect 184110 171200 184166 172000
rect 184754 171200 184810 172000
rect 185398 171200 185454 172000
rect 186042 171200 186098 172000
rect 186686 171200 186742 172000
rect 187330 171200 187386 172000
rect 187974 171200 188030 172000
rect 188618 171200 188674 172000
rect 189262 171200 189318 172000
rect 189906 171200 189962 172000
rect 190550 171200 190606 172000
rect 191194 171200 191250 172000
rect 191838 171200 191894 172000
rect 192482 171200 192538 172000
rect 193126 171200 193182 172000
rect 193862 171200 193918 172000
rect 194506 171200 194562 172000
rect 195150 171200 195206 172000
rect 195794 171200 195850 172000
rect 196438 171200 196494 172000
rect 197082 171200 197138 172000
rect 197726 171200 197782 172000
rect 198370 171200 198426 172000
rect 199014 171200 199070 172000
rect 199658 171200 199714 172000
rect 200302 171200 200358 172000
rect 200946 171200 201002 172000
rect 201590 171200 201646 172000
rect 202234 171200 202290 172000
rect 202878 171200 202934 172000
rect 203522 171200 203578 172000
rect 204166 171200 204222 172000
rect 204902 171200 204958 172000
rect 205546 171200 205602 172000
rect 206190 171200 206246 172000
rect 206834 171200 206890 172000
rect 207478 171200 207534 172000
rect 208122 171200 208178 172000
rect 208766 171200 208822 172000
rect 209410 171200 209466 172000
rect 210054 171200 210110 172000
rect 210698 171200 210754 172000
rect 211342 171200 211398 172000
rect 211986 171200 212042 172000
rect 212630 171200 212686 172000
rect 213274 171200 213330 172000
rect 213918 171200 213974 172000
rect 214562 171200 214618 172000
rect 215298 171200 215354 172000
rect 215942 171200 215998 172000
rect 216586 171200 216642 172000
rect 217230 171200 217286 172000
rect 217874 171200 217930 172000
rect 218518 171200 218574 172000
rect 219162 171200 219218 172000
rect 219806 171200 219862 172000
rect 220450 171200 220506 172000
rect 221094 171200 221150 172000
rect 221738 171200 221794 172000
rect 222382 171200 222438 172000
rect 223026 171200 223082 172000
rect 223670 171200 223726 172000
rect 224314 171200 224370 172000
rect 224958 171200 225014 172000
rect 225602 171200 225658 172000
rect 226338 171200 226394 172000
rect 226982 171200 227038 172000
rect 227626 171200 227682 172000
rect 228270 171200 228326 172000
rect 228914 171200 228970 172000
rect 229558 171200 229614 172000
rect 230202 171200 230258 172000
rect 230846 171200 230902 172000
rect 231490 171200 231546 172000
rect 232134 171200 232190 172000
rect 232778 171200 232834 172000
rect 233422 171200 233478 172000
rect 234066 171200 234122 172000
rect 234710 171200 234766 172000
rect 235354 171200 235410 172000
rect 235998 171200 236054 172000
rect 236642 171200 236698 172000
rect 237378 171200 237434 172000
rect 238022 171200 238078 172000
rect 238666 171200 238722 172000
rect 239310 171200 239366 172000
rect 239954 171200 240010 172000
rect 240598 171200 240654 172000
rect 241242 171200 241298 172000
rect 241886 171200 241942 172000
rect 242530 171200 242586 172000
rect 243174 171200 243230 172000
rect 243818 171200 243874 172000
rect 244462 171200 244518 172000
rect 245106 171200 245162 172000
rect 245750 171200 245806 172000
rect 246394 171200 246450 172000
rect 247038 171200 247094 172000
rect 247774 171200 247830 172000
rect 248418 171200 248474 172000
rect 249062 171200 249118 172000
rect 249706 171200 249762 172000
rect 250350 171200 250406 172000
rect 250994 171200 251050 172000
rect 251638 171200 251694 172000
rect 252282 171200 252338 172000
rect 252926 171200 252982 172000
rect 253570 171200 253626 172000
rect 254214 171200 254270 172000
rect 254858 171200 254914 172000
rect 255502 171200 255558 172000
rect 256146 171200 256202 172000
rect 256790 171200 256846 172000
rect 257434 171200 257490 172000
rect 258078 171200 258134 172000
rect 258814 171200 258870 172000
rect 259458 171200 259514 172000
rect 260102 171200 260158 172000
rect 260746 171200 260802 172000
rect 261390 171200 261446 172000
rect 262034 171200 262090 172000
rect 262678 171200 262734 172000
rect 263322 171200 263378 172000
rect 263966 171200 264022 172000
rect 264610 171200 264666 172000
rect 265254 171200 265310 172000
rect 265898 171200 265954 172000
rect 266542 171200 266598 172000
rect 267186 171200 267242 172000
rect 267830 171200 267886 172000
rect 268474 171200 268530 172000
rect 269210 171200 269266 172000
rect 269854 171200 269910 172000
rect 270498 171200 270554 172000
rect 271142 171200 271198 172000
rect 271786 171200 271842 172000
rect 272430 171200 272486 172000
rect 273074 171200 273130 172000
rect 273718 171200 273774 172000
rect 274362 171200 274418 172000
rect 275006 171200 275062 172000
rect 275650 171200 275706 172000
rect 276294 171200 276350 172000
rect 276938 171200 276994 172000
rect 277582 171200 277638 172000
rect 278226 171200 278282 172000
rect 278870 171200 278926 172000
rect 279514 171200 279570 172000
rect 280250 171200 280306 172000
rect 280894 171200 280950 172000
rect 281538 171200 281594 172000
rect 282182 171200 282238 172000
rect 282826 171200 282882 172000
rect 283470 171200 283526 172000
rect 284114 171200 284170 172000
rect 284758 171200 284814 172000
rect 285402 171200 285458 172000
rect 286046 171200 286102 172000
rect 286690 171200 286746 172000
rect 287334 171200 287390 172000
rect 287978 171200 288034 172000
rect 288622 171200 288678 172000
rect 289266 171200 289322 172000
rect 289910 171200 289966 172000
rect 290646 171200 290702 172000
rect 291290 171200 291346 172000
rect 291934 171200 291990 172000
rect 292578 171200 292634 172000
rect 293222 171200 293278 172000
rect 293866 171200 293922 172000
rect 294510 171200 294566 172000
rect 295154 171200 295210 172000
rect 295798 171200 295854 172000
rect 296442 171200 296498 172000
rect 297086 171200 297142 172000
rect 297730 171200 297786 172000
rect 298374 171200 298430 172000
rect 299018 171200 299074 172000
rect 299662 171200 299718 172000
rect 300306 171200 300362 172000
rect 300950 171200 301006 172000
rect 301686 171200 301742 172000
rect 302330 171200 302386 172000
rect 302974 171200 303030 172000
rect 303618 171200 303674 172000
rect 304262 171200 304318 172000
rect 304906 171200 304962 172000
rect 305550 171200 305606 172000
rect 306194 171200 306250 172000
rect 306838 171200 306894 172000
rect 307482 171200 307538 172000
rect 308126 171200 308182 172000
rect 308770 171200 308826 172000
rect 309414 171200 309470 172000
rect 310058 171200 310114 172000
rect 310702 171200 310758 172000
rect 311346 171200 311402 172000
rect 312082 171200 312138 172000
rect 312726 171200 312782 172000
rect 313370 171200 313426 172000
rect 314014 171200 314070 172000
rect 314658 171200 314714 172000
rect 315302 171200 315358 172000
rect 315946 171200 316002 172000
rect 316590 171200 316646 172000
rect 317234 171200 317290 172000
rect 317878 171200 317934 172000
rect 318522 171200 318578 172000
rect 319166 171200 319222 172000
rect 319810 171200 319866 172000
rect 320454 171200 320510 172000
rect 321098 171200 321154 172000
rect 321742 171200 321798 172000
rect 322386 171200 322442 172000
rect 323122 171200 323178 172000
rect 323766 171200 323822 172000
rect 324410 171200 324466 172000
rect 325054 171200 325110 172000
rect 325698 171200 325754 172000
rect 326342 171200 326398 172000
rect 326986 171200 327042 172000
rect 327630 171200 327686 172000
rect 328274 171200 328330 172000
rect 328918 171200 328974 172000
rect 329562 171200 329618 172000
rect 330206 171200 330262 172000
rect 330850 171200 330906 172000
rect 331494 171200 331550 172000
rect 332138 171200 332194 172000
rect 332782 171200 332838 172000
rect 333426 171200 333482 172000
rect 334162 171200 334218 172000
rect 334806 171200 334862 172000
rect 335450 171200 335506 172000
rect 336094 171200 336150 172000
rect 336738 171200 336794 172000
rect 337382 171200 337438 172000
rect 338026 171200 338082 172000
rect 338670 171200 338726 172000
rect 339314 171200 339370 172000
rect 339958 171200 340014 172000
rect 340602 171200 340658 172000
rect 341246 171200 341302 172000
rect 341890 171200 341946 172000
rect 342534 171200 342590 172000
rect 343178 171200 343234 172000
rect 343822 171200 343878 172000
rect 344558 171200 344614 172000
rect 345202 171200 345258 172000
rect 345846 171200 345902 172000
rect 346490 171200 346546 172000
rect 347134 171200 347190 172000
rect 347778 171200 347834 172000
rect 348422 171200 348478 172000
rect 349066 171200 349122 172000
rect 349710 171200 349766 172000
rect 350354 171200 350410 172000
rect 350998 171200 351054 172000
rect 351642 171200 351698 172000
rect 352286 171200 352342 172000
rect 352930 171200 352986 172000
rect 353574 171200 353630 172000
rect 354218 171200 354274 172000
rect 354862 171200 354918 172000
rect 355598 171200 355654 172000
rect 356242 171200 356298 172000
rect 356886 171200 356942 172000
rect 357530 171200 357586 172000
rect 358174 171200 358230 172000
rect 358818 171200 358874 172000
rect 359462 171200 359518 172000
rect 360106 171200 360162 172000
rect 360750 171200 360806 172000
rect 361394 171200 361450 172000
rect 362038 171200 362094 172000
rect 362682 171200 362738 172000
rect 363326 171200 363382 172000
rect 363970 171200 364026 172000
rect 364614 171200 364670 172000
rect 365258 171200 365314 172000
rect 365994 171200 366050 172000
rect 366638 171200 366694 172000
rect 367282 171200 367338 172000
rect 367926 171200 367982 172000
rect 368570 171200 368626 172000
rect 369214 171200 369270 172000
rect 369858 171200 369914 172000
rect 370502 171200 370558 172000
rect 371146 171200 371202 172000
rect 371790 171200 371846 172000
rect 372434 171200 372490 172000
rect 373078 171200 373134 172000
rect 373722 171200 373778 172000
rect 374366 171200 374422 172000
rect 375010 171200 375066 172000
rect 375654 171200 375710 172000
rect 376298 171200 376354 172000
rect 377034 171200 377090 172000
rect 377678 171200 377734 172000
rect 378322 171200 378378 172000
rect 378966 171200 379022 172000
rect 379610 171200 379666 172000
rect 380254 171200 380310 172000
rect 380898 171200 380954 172000
rect 381542 171200 381598 172000
rect 382186 171200 382242 172000
rect 382830 171200 382886 172000
rect 383474 171200 383530 172000
rect 384118 171200 384174 172000
rect 384762 171200 384818 172000
rect 385406 171200 385462 172000
rect 386050 171200 386106 172000
rect 386694 171200 386750 172000
rect 387430 171200 387486 172000
rect 388074 171200 388130 172000
rect 388718 171200 388774 172000
rect 389362 171200 389418 172000
rect 390006 171200 390062 172000
rect 390650 171200 390706 172000
rect 391294 171200 391350 172000
rect 391938 171200 391994 172000
rect 392582 171200 392638 172000
rect 393226 171200 393282 172000
rect 393870 171200 393926 172000
rect 394514 171200 394570 172000
rect 395158 171200 395214 172000
rect 395802 171200 395858 172000
rect 396446 171200 396502 172000
rect 397090 171200 397146 172000
rect 397734 171200 397790 172000
rect 398470 171200 398526 172000
rect 399114 171200 399170 172000
rect 399758 171200 399814 172000
rect 400402 171200 400458 172000
rect 401046 171200 401102 172000
rect 401690 171200 401746 172000
rect 402334 171200 402390 172000
rect 402978 171200 403034 172000
rect 403622 171200 403678 172000
rect 404266 171200 404322 172000
rect 404910 171200 404966 172000
rect 405554 171200 405610 172000
rect 406198 171200 406254 172000
rect 406842 171200 406898 172000
rect 407486 171200 407542 172000
rect 408130 171200 408186 172000
rect 408866 171200 408922 172000
rect 409510 171200 409566 172000
rect 410154 171200 410210 172000
rect 410798 171200 410854 172000
rect 411442 171200 411498 172000
rect 412086 171200 412142 172000
rect 412730 171200 412786 172000
rect 413374 171200 413430 172000
rect 414018 171200 414074 172000
rect 414662 171200 414718 172000
rect 415306 171200 415362 172000
rect 415950 171200 416006 172000
rect 416594 171200 416650 172000
rect 417238 171200 417294 172000
rect 417882 171200 417938 172000
rect 418526 171200 418582 172000
rect 419170 171200 419226 172000
rect 419906 171200 419962 172000
rect 420550 171200 420606 172000
rect 421194 171200 421250 172000
rect 421838 171200 421894 172000
rect 422482 171200 422538 172000
rect 423126 171200 423182 172000
rect 423770 171200 423826 172000
rect 424414 171200 424470 172000
rect 425058 171200 425114 172000
rect 425702 171200 425758 172000
rect 426346 171200 426402 172000
rect 426990 171200 427046 172000
rect 427634 171200 427690 172000
rect 428278 171200 428334 172000
rect 428922 171200 428978 172000
rect 429566 171200 429622 172000
rect 9770 0 9826 800
rect 29274 0 29330 800
rect 48778 0 48834 800
rect 68374 0 68430 800
rect 87878 0 87934 800
rect 107474 0 107530 800
rect 126978 0 127034 800
rect 146574 0 146630 800
rect 166078 0 166134 800
rect 185674 0 185730 800
rect 205178 0 205234 800
rect 224774 0 224830 800
rect 244278 0 244334 800
rect 263782 0 263838 800
rect 283378 0 283434 800
rect 302882 0 302938 800
rect 322478 0 322534 800
rect 341982 0 342038 800
rect 361578 0 361634 800
rect 381082 0 381138 800
rect 400678 0 400734 800
rect 420182 0 420238 800
<< obsm2 >>
rect 406 171144 882 171970
rect 1050 171144 1526 171970
rect 1694 171144 2170 171970
rect 2338 171144 2814 171970
rect 2982 171144 3458 171970
rect 3626 171144 4102 171970
rect 4270 171144 4746 171970
rect 4914 171144 5390 171970
rect 5558 171144 6034 171970
rect 6202 171144 6678 171970
rect 6846 171144 7322 171970
rect 7490 171144 7966 171970
rect 8134 171144 8610 171970
rect 8778 171144 9254 171970
rect 9422 171144 9898 171970
rect 10066 171144 10542 171970
rect 10710 171144 11278 171970
rect 11446 171144 11922 171970
rect 12090 171144 12566 171970
rect 12734 171144 13210 171970
rect 13378 171144 13854 171970
rect 14022 171144 14498 171970
rect 14666 171144 15142 171970
rect 15310 171144 15786 171970
rect 15954 171144 16430 171970
rect 16598 171144 17074 171970
rect 17242 171144 17718 171970
rect 17886 171144 18362 171970
rect 18530 171144 19006 171970
rect 19174 171144 19650 171970
rect 19818 171144 20294 171970
rect 20462 171144 20938 171970
rect 21106 171144 21582 171970
rect 21750 171144 22318 171970
rect 22486 171144 22962 171970
rect 23130 171144 23606 171970
rect 23774 171144 24250 171970
rect 24418 171144 24894 171970
rect 25062 171144 25538 171970
rect 25706 171144 26182 171970
rect 26350 171144 26826 171970
rect 26994 171144 27470 171970
rect 27638 171144 28114 171970
rect 28282 171144 28758 171970
rect 28926 171144 29402 171970
rect 29570 171144 30046 171970
rect 30214 171144 30690 171970
rect 30858 171144 31334 171970
rect 31502 171144 31978 171970
rect 32146 171144 32714 171970
rect 32882 171144 33358 171970
rect 33526 171144 34002 171970
rect 34170 171144 34646 171970
rect 34814 171144 35290 171970
rect 35458 171144 35934 171970
rect 36102 171144 36578 171970
rect 36746 171144 37222 171970
rect 37390 171144 37866 171970
rect 38034 171144 38510 171970
rect 38678 171144 39154 171970
rect 39322 171144 39798 171970
rect 39966 171144 40442 171970
rect 40610 171144 41086 171970
rect 41254 171144 41730 171970
rect 41898 171144 42374 171970
rect 42542 171144 43018 171970
rect 43186 171144 43754 171970
rect 43922 171144 44398 171970
rect 44566 171144 45042 171970
rect 45210 171144 45686 171970
rect 45854 171144 46330 171970
rect 46498 171144 46974 171970
rect 47142 171144 47618 171970
rect 47786 171144 48262 171970
rect 48430 171144 48906 171970
rect 49074 171144 49550 171970
rect 49718 171144 50194 171970
rect 50362 171144 50838 171970
rect 51006 171144 51482 171970
rect 51650 171144 52126 171970
rect 52294 171144 52770 171970
rect 52938 171144 53414 171970
rect 53582 171144 54150 171970
rect 54318 171144 54794 171970
rect 54962 171144 55438 171970
rect 55606 171144 56082 171970
rect 56250 171144 56726 171970
rect 56894 171144 57370 171970
rect 57538 171144 58014 171970
rect 58182 171144 58658 171970
rect 58826 171144 59302 171970
rect 59470 171144 59946 171970
rect 60114 171144 60590 171970
rect 60758 171144 61234 171970
rect 61402 171144 61878 171970
rect 62046 171144 62522 171970
rect 62690 171144 63166 171970
rect 63334 171144 63810 171970
rect 63978 171144 64454 171970
rect 64622 171144 65190 171970
rect 65358 171144 65834 171970
rect 66002 171144 66478 171970
rect 66646 171144 67122 171970
rect 67290 171144 67766 171970
rect 67934 171144 68410 171970
rect 68578 171144 69054 171970
rect 69222 171144 69698 171970
rect 69866 171144 70342 171970
rect 70510 171144 70986 171970
rect 71154 171144 71630 171970
rect 71798 171144 72274 171970
rect 72442 171144 72918 171970
rect 73086 171144 73562 171970
rect 73730 171144 74206 171970
rect 74374 171144 74850 171970
rect 75018 171144 75586 171970
rect 75754 171144 76230 171970
rect 76398 171144 76874 171970
rect 77042 171144 77518 171970
rect 77686 171144 78162 171970
rect 78330 171144 78806 171970
rect 78974 171144 79450 171970
rect 79618 171144 80094 171970
rect 80262 171144 80738 171970
rect 80906 171144 81382 171970
rect 81550 171144 82026 171970
rect 82194 171144 82670 171970
rect 82838 171144 83314 171970
rect 83482 171144 83958 171970
rect 84126 171144 84602 171970
rect 84770 171144 85246 171970
rect 85414 171144 85890 171970
rect 86058 171144 86626 171970
rect 86794 171144 87270 171970
rect 87438 171144 87914 171970
rect 88082 171144 88558 171970
rect 88726 171144 89202 171970
rect 89370 171144 89846 171970
rect 90014 171144 90490 171970
rect 90658 171144 91134 171970
rect 91302 171144 91778 171970
rect 91946 171144 92422 171970
rect 92590 171144 93066 171970
rect 93234 171144 93710 171970
rect 93878 171144 94354 171970
rect 94522 171144 94998 171970
rect 95166 171144 95642 171970
rect 95810 171144 96286 171970
rect 96454 171144 97022 171970
rect 97190 171144 97666 171970
rect 97834 171144 98310 171970
rect 98478 171144 98954 171970
rect 99122 171144 99598 171970
rect 99766 171144 100242 171970
rect 100410 171144 100886 171970
rect 101054 171144 101530 171970
rect 101698 171144 102174 171970
rect 102342 171144 102818 171970
rect 102986 171144 103462 171970
rect 103630 171144 104106 171970
rect 104274 171144 104750 171970
rect 104918 171144 105394 171970
rect 105562 171144 106038 171970
rect 106206 171144 106682 171970
rect 106850 171144 107326 171970
rect 107494 171144 108062 171970
rect 108230 171144 108706 171970
rect 108874 171144 109350 171970
rect 109518 171144 109994 171970
rect 110162 171144 110638 171970
rect 110806 171144 111282 171970
rect 111450 171144 111926 171970
rect 112094 171144 112570 171970
rect 112738 171144 113214 171970
rect 113382 171144 113858 171970
rect 114026 171144 114502 171970
rect 114670 171144 115146 171970
rect 115314 171144 115790 171970
rect 115958 171144 116434 171970
rect 116602 171144 117078 171970
rect 117246 171144 117722 171970
rect 117890 171144 118366 171970
rect 118534 171144 119102 171970
rect 119270 171144 119746 171970
rect 119914 171144 120390 171970
rect 120558 171144 121034 171970
rect 121202 171144 121678 171970
rect 121846 171144 122322 171970
rect 122490 171144 122966 171970
rect 123134 171144 123610 171970
rect 123778 171144 124254 171970
rect 124422 171144 124898 171970
rect 125066 171144 125542 171970
rect 125710 171144 126186 171970
rect 126354 171144 126830 171970
rect 126998 171144 127474 171970
rect 127642 171144 128118 171970
rect 128286 171144 128762 171970
rect 128930 171144 129498 171970
rect 129666 171144 130142 171970
rect 130310 171144 130786 171970
rect 130954 171144 131430 171970
rect 131598 171144 132074 171970
rect 132242 171144 132718 171970
rect 132886 171144 133362 171970
rect 133530 171144 134006 171970
rect 134174 171144 134650 171970
rect 134818 171144 135294 171970
rect 135462 171144 135938 171970
rect 136106 171144 136582 171970
rect 136750 171144 137226 171970
rect 137394 171144 137870 171970
rect 138038 171144 138514 171970
rect 138682 171144 139158 171970
rect 139326 171144 139802 171970
rect 139970 171144 140538 171970
rect 140706 171144 141182 171970
rect 141350 171144 141826 171970
rect 141994 171144 142470 171970
rect 142638 171144 143114 171970
rect 143282 171144 143758 171970
rect 143926 171144 144402 171970
rect 144570 171144 145046 171970
rect 145214 171144 145690 171970
rect 145858 171144 146334 171970
rect 146502 171144 146978 171970
rect 147146 171144 147622 171970
rect 147790 171144 148266 171970
rect 148434 171144 148910 171970
rect 149078 171144 149554 171970
rect 149722 171144 150198 171970
rect 150366 171144 150934 171970
rect 151102 171144 151578 171970
rect 151746 171144 152222 171970
rect 152390 171144 152866 171970
rect 153034 171144 153510 171970
rect 153678 171144 154154 171970
rect 154322 171144 154798 171970
rect 154966 171144 155442 171970
rect 155610 171144 156086 171970
rect 156254 171144 156730 171970
rect 156898 171144 157374 171970
rect 157542 171144 158018 171970
rect 158186 171144 158662 171970
rect 158830 171144 159306 171970
rect 159474 171144 159950 171970
rect 160118 171144 160594 171970
rect 160762 171144 161238 171970
rect 161406 171144 161974 171970
rect 162142 171144 162618 171970
rect 162786 171144 163262 171970
rect 163430 171144 163906 171970
rect 164074 171144 164550 171970
rect 164718 171144 165194 171970
rect 165362 171144 165838 171970
rect 166006 171144 166482 171970
rect 166650 171144 167126 171970
rect 167294 171144 167770 171970
rect 167938 171144 168414 171970
rect 168582 171144 169058 171970
rect 169226 171144 169702 171970
rect 169870 171144 170346 171970
rect 170514 171144 170990 171970
rect 171158 171144 171634 171970
rect 171802 171144 172370 171970
rect 172538 171144 173014 171970
rect 173182 171144 173658 171970
rect 173826 171144 174302 171970
rect 174470 171144 174946 171970
rect 175114 171144 175590 171970
rect 175758 171144 176234 171970
rect 176402 171144 176878 171970
rect 177046 171144 177522 171970
rect 177690 171144 178166 171970
rect 178334 171144 178810 171970
rect 178978 171144 179454 171970
rect 179622 171144 180098 171970
rect 180266 171144 180742 171970
rect 180910 171144 181386 171970
rect 181554 171144 182030 171970
rect 182198 171144 182674 171970
rect 182842 171144 183410 171970
rect 183578 171144 184054 171970
rect 184222 171144 184698 171970
rect 184866 171144 185342 171970
rect 185510 171144 185986 171970
rect 186154 171144 186630 171970
rect 186798 171144 187274 171970
rect 187442 171144 187918 171970
rect 188086 171144 188562 171970
rect 188730 171144 189206 171970
rect 189374 171144 189850 171970
rect 190018 171144 190494 171970
rect 190662 171144 191138 171970
rect 191306 171144 191782 171970
rect 191950 171144 192426 171970
rect 192594 171144 193070 171970
rect 193238 171144 193806 171970
rect 193974 171144 194450 171970
rect 194618 171144 195094 171970
rect 195262 171144 195738 171970
rect 195906 171144 196382 171970
rect 196550 171144 197026 171970
rect 197194 171144 197670 171970
rect 197838 171144 198314 171970
rect 198482 171144 198958 171970
rect 199126 171144 199602 171970
rect 199770 171144 200246 171970
rect 200414 171144 200890 171970
rect 201058 171144 201534 171970
rect 201702 171144 202178 171970
rect 202346 171144 202822 171970
rect 202990 171144 203466 171970
rect 203634 171144 204110 171970
rect 204278 171144 204846 171970
rect 205014 171144 205490 171970
rect 205658 171144 206134 171970
rect 206302 171144 206778 171970
rect 206946 171144 207422 171970
rect 207590 171144 208066 171970
rect 208234 171144 208710 171970
rect 208878 171144 209354 171970
rect 209522 171144 209998 171970
rect 210166 171144 210642 171970
rect 210810 171144 211286 171970
rect 211454 171144 211930 171970
rect 212098 171144 212574 171970
rect 212742 171144 213218 171970
rect 213386 171144 213862 171970
rect 214030 171144 214506 171970
rect 214674 171144 215242 171970
rect 215410 171144 215886 171970
rect 216054 171144 216530 171970
rect 216698 171144 217174 171970
rect 217342 171144 217818 171970
rect 217986 171144 218462 171970
rect 218630 171144 219106 171970
rect 219274 171144 219750 171970
rect 219918 171144 220394 171970
rect 220562 171144 221038 171970
rect 221206 171144 221682 171970
rect 221850 171144 222326 171970
rect 222494 171144 222970 171970
rect 223138 171144 223614 171970
rect 223782 171144 224258 171970
rect 224426 171144 224902 171970
rect 225070 171144 225546 171970
rect 225714 171144 226282 171970
rect 226450 171144 226926 171970
rect 227094 171144 227570 171970
rect 227738 171144 228214 171970
rect 228382 171144 228858 171970
rect 229026 171144 229502 171970
rect 229670 171144 230146 171970
rect 230314 171144 230790 171970
rect 230958 171144 231434 171970
rect 231602 171144 232078 171970
rect 232246 171144 232722 171970
rect 232890 171144 233366 171970
rect 233534 171144 234010 171970
rect 234178 171144 234654 171970
rect 234822 171144 235298 171970
rect 235466 171144 235942 171970
rect 236110 171144 236586 171970
rect 236754 171144 237322 171970
rect 237490 171144 237966 171970
rect 238134 171144 238610 171970
rect 238778 171144 239254 171970
rect 239422 171144 239898 171970
rect 240066 171144 240542 171970
rect 240710 171144 241186 171970
rect 241354 171144 241830 171970
rect 241998 171144 242474 171970
rect 242642 171144 243118 171970
rect 243286 171144 243762 171970
rect 243930 171144 244406 171970
rect 244574 171144 245050 171970
rect 245218 171144 245694 171970
rect 245862 171144 246338 171970
rect 246506 171144 246982 171970
rect 247150 171144 247718 171970
rect 247886 171144 248362 171970
rect 248530 171144 249006 171970
rect 249174 171144 249650 171970
rect 249818 171144 250294 171970
rect 250462 171144 250938 171970
rect 251106 171144 251582 171970
rect 251750 171144 252226 171970
rect 252394 171144 252870 171970
rect 253038 171144 253514 171970
rect 253682 171144 254158 171970
rect 254326 171144 254802 171970
rect 254970 171144 255446 171970
rect 255614 171144 256090 171970
rect 256258 171144 256734 171970
rect 256902 171144 257378 171970
rect 257546 171144 258022 171970
rect 258190 171144 258758 171970
rect 258926 171144 259402 171970
rect 259570 171144 260046 171970
rect 260214 171144 260690 171970
rect 260858 171144 261334 171970
rect 261502 171144 261978 171970
rect 262146 171144 262622 171970
rect 262790 171144 263266 171970
rect 263434 171144 263910 171970
rect 264078 171144 264554 171970
rect 264722 171144 265198 171970
rect 265366 171144 265842 171970
rect 266010 171144 266486 171970
rect 266654 171144 267130 171970
rect 267298 171144 267774 171970
rect 267942 171144 268418 171970
rect 268586 171144 269154 171970
rect 269322 171144 269798 171970
rect 269966 171144 270442 171970
rect 270610 171144 271086 171970
rect 271254 171144 271730 171970
rect 271898 171144 272374 171970
rect 272542 171144 273018 171970
rect 273186 171144 273662 171970
rect 273830 171144 274306 171970
rect 274474 171144 274950 171970
rect 275118 171144 275594 171970
rect 275762 171144 276238 171970
rect 276406 171144 276882 171970
rect 277050 171144 277526 171970
rect 277694 171144 278170 171970
rect 278338 171144 278814 171970
rect 278982 171144 279458 171970
rect 279626 171144 280194 171970
rect 280362 171144 280838 171970
rect 281006 171144 281482 171970
rect 281650 171144 282126 171970
rect 282294 171144 282770 171970
rect 282938 171144 283414 171970
rect 283582 171144 284058 171970
rect 284226 171144 284702 171970
rect 284870 171144 285346 171970
rect 285514 171144 285990 171970
rect 286158 171144 286634 171970
rect 286802 171144 287278 171970
rect 287446 171144 287922 171970
rect 288090 171144 288566 171970
rect 288734 171144 289210 171970
rect 289378 171144 289854 171970
rect 290022 171144 290590 171970
rect 290758 171144 291234 171970
rect 291402 171144 291878 171970
rect 292046 171144 292522 171970
rect 292690 171144 293166 171970
rect 293334 171144 293810 171970
rect 293978 171144 294454 171970
rect 294622 171144 295098 171970
rect 295266 171144 295742 171970
rect 295910 171144 296386 171970
rect 296554 171144 297030 171970
rect 297198 171144 297674 171970
rect 297842 171144 298318 171970
rect 298486 171144 298962 171970
rect 299130 171144 299606 171970
rect 299774 171144 300250 171970
rect 300418 171144 300894 171970
rect 301062 171144 301630 171970
rect 301798 171144 302274 171970
rect 302442 171144 302918 171970
rect 303086 171144 303562 171970
rect 303730 171144 304206 171970
rect 304374 171144 304850 171970
rect 305018 171144 305494 171970
rect 305662 171144 306138 171970
rect 306306 171144 306782 171970
rect 306950 171144 307426 171970
rect 307594 171144 308070 171970
rect 308238 171144 308714 171970
rect 308882 171144 309358 171970
rect 309526 171144 310002 171970
rect 310170 171144 310646 171970
rect 310814 171144 311290 171970
rect 311458 171144 312026 171970
rect 312194 171144 312670 171970
rect 312838 171144 313314 171970
rect 313482 171144 313958 171970
rect 314126 171144 314602 171970
rect 314770 171144 315246 171970
rect 315414 171144 315890 171970
rect 316058 171144 316534 171970
rect 316702 171144 317178 171970
rect 317346 171144 317822 171970
rect 317990 171144 318466 171970
rect 318634 171144 319110 171970
rect 319278 171144 319754 171970
rect 319922 171144 320398 171970
rect 320566 171144 321042 171970
rect 321210 171144 321686 171970
rect 321854 171144 322330 171970
rect 322498 171144 323066 171970
rect 323234 171144 323710 171970
rect 323878 171144 324354 171970
rect 324522 171144 324998 171970
rect 325166 171144 325642 171970
rect 325810 171144 326286 171970
rect 326454 171144 326930 171970
rect 327098 171144 327574 171970
rect 327742 171144 328218 171970
rect 328386 171144 328862 171970
rect 329030 171144 329506 171970
rect 329674 171144 330150 171970
rect 330318 171144 330794 171970
rect 330962 171144 331438 171970
rect 331606 171144 332082 171970
rect 332250 171144 332726 171970
rect 332894 171144 333370 171970
rect 333538 171144 334106 171970
rect 334274 171144 334750 171970
rect 334918 171144 335394 171970
rect 335562 171144 336038 171970
rect 336206 171144 336682 171970
rect 336850 171144 337326 171970
rect 337494 171144 337970 171970
rect 338138 171144 338614 171970
rect 338782 171144 339258 171970
rect 339426 171144 339902 171970
rect 340070 171144 340546 171970
rect 340714 171144 341190 171970
rect 341358 171144 341834 171970
rect 342002 171144 342478 171970
rect 342646 171144 343122 171970
rect 343290 171144 343766 171970
rect 343934 171144 344502 171970
rect 344670 171144 345146 171970
rect 345314 171144 345790 171970
rect 345958 171144 346434 171970
rect 346602 171144 347078 171970
rect 347246 171144 347722 171970
rect 347890 171144 348366 171970
rect 348534 171144 349010 171970
rect 349178 171144 349654 171970
rect 349822 171144 350298 171970
rect 350466 171144 350942 171970
rect 351110 171144 351586 171970
rect 351754 171144 352230 171970
rect 352398 171144 352874 171970
rect 353042 171144 353518 171970
rect 353686 171144 354162 171970
rect 354330 171144 354806 171970
rect 354974 171144 355542 171970
rect 355710 171144 356186 171970
rect 356354 171144 356830 171970
rect 356998 171144 357474 171970
rect 357642 171144 358118 171970
rect 358286 171144 358762 171970
rect 358930 171144 359406 171970
rect 359574 171144 360050 171970
rect 360218 171144 360694 171970
rect 360862 171144 361338 171970
rect 361506 171144 361982 171970
rect 362150 171144 362626 171970
rect 362794 171144 363270 171970
rect 363438 171144 363914 171970
rect 364082 171144 364558 171970
rect 364726 171144 365202 171970
rect 365370 171144 365938 171970
rect 366106 171144 366582 171970
rect 366750 171144 367226 171970
rect 367394 171144 367870 171970
rect 368038 171144 368514 171970
rect 368682 171144 369158 171970
rect 369326 171144 369802 171970
rect 369970 171144 370446 171970
rect 370614 171144 371090 171970
rect 371258 171144 371734 171970
rect 371902 171144 372378 171970
rect 372546 171144 373022 171970
rect 373190 171144 373666 171970
rect 373834 171144 374310 171970
rect 374478 171144 374954 171970
rect 375122 171144 375598 171970
rect 375766 171144 376242 171970
rect 376410 171144 376978 171970
rect 377146 171144 377622 171970
rect 377790 171144 378266 171970
rect 378434 171144 378910 171970
rect 379078 171144 379554 171970
rect 379722 171144 380198 171970
rect 380366 171144 380842 171970
rect 381010 171144 381486 171970
rect 381654 171144 382130 171970
rect 382298 171144 382774 171970
rect 382942 171144 383418 171970
rect 383586 171144 384062 171970
rect 384230 171144 384706 171970
rect 384874 171144 385350 171970
rect 385518 171144 385994 171970
rect 386162 171144 386638 171970
rect 386806 171144 387374 171970
rect 387542 171144 388018 171970
rect 388186 171144 388662 171970
rect 388830 171144 389306 171970
rect 389474 171144 389950 171970
rect 390118 171144 390594 171970
rect 390762 171144 391238 171970
rect 391406 171144 391882 171970
rect 392050 171144 392526 171970
rect 392694 171144 393170 171970
rect 393338 171144 393814 171970
rect 393982 171144 394458 171970
rect 394626 171144 395102 171970
rect 395270 171144 395746 171970
rect 395914 171144 396390 171970
rect 396558 171144 397034 171970
rect 397202 171144 397678 171970
rect 397846 171144 398414 171970
rect 398582 171144 399058 171970
rect 399226 171144 399702 171970
rect 399870 171144 400346 171970
rect 400514 171144 400990 171970
rect 401158 171144 401634 171970
rect 401802 171144 402278 171970
rect 402446 171144 402922 171970
rect 403090 171144 403566 171970
rect 403734 171144 404210 171970
rect 404378 171144 404854 171970
rect 405022 171144 405498 171970
rect 405666 171144 406142 171970
rect 406310 171144 406786 171970
rect 406954 171144 407430 171970
rect 407598 171144 408074 171970
rect 408242 171144 408810 171970
rect 408978 171144 409454 171970
rect 409622 171144 410098 171970
rect 410266 171144 410742 171970
rect 410910 171144 411386 171970
rect 411554 171144 412030 171970
rect 412198 171144 412674 171970
rect 412842 171144 413318 171970
rect 413486 171144 413962 171970
rect 414130 171144 414606 171970
rect 414774 171144 415250 171970
rect 415418 171144 415894 171970
rect 416062 171144 416538 171970
rect 416706 171144 417182 171970
rect 417350 171144 417826 171970
rect 417994 171144 418470 171970
rect 418638 171144 419114 171970
rect 419282 171144 419850 171970
rect 420018 171144 420494 171970
rect 420662 171144 421138 171970
rect 421306 171144 421782 171970
rect 421950 171144 422426 171970
rect 422594 171144 423070 171970
rect 423238 171144 423714 171970
rect 423882 171144 424358 171970
rect 424526 171144 425002 171970
rect 425170 171144 425646 171970
rect 425814 171144 426290 171970
rect 426458 171144 426934 171970
rect 427102 171144 427578 171970
rect 427746 171144 428222 171970
rect 428390 171144 428866 171970
rect 429034 171144 429510 171970
rect 296 856 429620 171144
rect 296 439 9714 856
rect 9882 439 29218 856
rect 29386 439 48722 856
rect 48890 439 68318 856
rect 68486 439 87822 856
rect 87990 439 107418 856
rect 107586 439 126922 856
rect 127090 439 146518 856
rect 146686 439 166022 856
rect 166190 439 185618 856
rect 185786 439 205122 856
rect 205290 439 224718 856
rect 224886 439 244222 856
rect 244390 439 263726 856
rect 263894 439 283322 856
rect 283490 439 302826 856
rect 302994 439 322422 856
rect 322590 439 341926 856
rect 342094 439 361522 856
rect 361690 439 381026 856
rect 381194 439 400622 856
rect 400790 439 420126 856
rect 420294 439 429620 856
<< metal3 >>
rect 0 171368 800 171488
rect 429200 170960 430000 171080
rect 0 170280 800 170400
rect 0 169192 800 169312
rect 429200 169056 430000 169176
rect 0 168104 800 168224
rect 0 167016 800 167136
rect 429200 167152 430000 167272
rect 0 165928 800 166048
rect 429200 165248 430000 165368
rect 0 164840 800 164960
rect 0 163752 800 163872
rect 429200 163208 430000 163328
rect 0 162664 800 162784
rect 0 161576 800 161696
rect 429200 161304 430000 161424
rect 0 160624 800 160744
rect 0 159536 800 159656
rect 429200 159400 430000 159520
rect 0 158448 800 158568
rect 0 157360 800 157480
rect 429200 157496 430000 157616
rect 0 156272 800 156392
rect 429200 155592 430000 155712
rect 0 155184 800 155304
rect 0 154096 800 154216
rect 429200 153552 430000 153672
rect 0 153008 800 153128
rect 0 151920 800 152040
rect 429200 151648 430000 151768
rect 0 150832 800 150952
rect 0 149744 800 149864
rect 429200 149744 430000 149864
rect 0 148792 800 148912
rect 0 147704 800 147824
rect 429200 147840 430000 147960
rect 0 146616 800 146736
rect 429200 145936 430000 146056
rect 0 145528 800 145648
rect 0 144440 800 144560
rect 429200 143896 430000 144016
rect 0 143352 800 143472
rect 0 142264 800 142384
rect 429200 141992 430000 142112
rect 0 141176 800 141296
rect 0 140088 800 140208
rect 429200 140088 430000 140208
rect 0 139000 800 139120
rect 0 138048 800 138168
rect 429200 138184 430000 138304
rect 0 136960 800 137080
rect 429200 136144 430000 136264
rect 0 135872 800 135992
rect 0 134784 800 134904
rect 429200 134240 430000 134360
rect 0 133696 800 133816
rect 0 132608 800 132728
rect 429200 132336 430000 132456
rect 0 131520 800 131640
rect 0 130432 800 130552
rect 429200 130432 430000 130552
rect 0 129344 800 129464
rect 429200 128528 430000 128648
rect 0 128256 800 128376
rect 0 127168 800 127288
rect 429200 126488 430000 126608
rect 0 126216 800 126336
rect 0 125128 800 125248
rect 429200 124584 430000 124704
rect 0 124040 800 124160
rect 0 122952 800 123072
rect 429200 122680 430000 122800
rect 0 121864 800 121984
rect 0 120776 800 120896
rect 429200 120776 430000 120896
rect 0 119688 800 119808
rect 429200 118872 430000 118992
rect 0 118600 800 118720
rect 0 117512 800 117632
rect 429200 116832 430000 116952
rect 0 116424 800 116544
rect 0 115336 800 115456
rect 429200 114928 430000 115048
rect 0 114384 800 114504
rect 0 113296 800 113416
rect 429200 113024 430000 113144
rect 0 112208 800 112328
rect 0 111120 800 111240
rect 429200 111120 430000 111240
rect 0 110032 800 110152
rect 0 108944 800 109064
rect 429200 109080 430000 109200
rect 0 107856 800 107976
rect 429200 107176 430000 107296
rect 0 106768 800 106888
rect 0 105680 800 105800
rect 429200 105272 430000 105392
rect 0 104592 800 104712
rect 0 103640 800 103760
rect 429200 103368 430000 103488
rect 0 102552 800 102672
rect 0 101464 800 101584
rect 429200 101464 430000 101584
rect 0 100376 800 100496
rect 0 99288 800 99408
rect 429200 99424 430000 99544
rect 0 98200 800 98320
rect 429200 97520 430000 97640
rect 0 97112 800 97232
rect 0 96024 800 96144
rect 429200 95616 430000 95736
rect 0 94936 800 95056
rect 0 93848 800 93968
rect 429200 93712 430000 93832
rect 0 92760 800 92880
rect 0 91808 800 91928
rect 429200 91808 430000 91928
rect 0 90720 800 90840
rect 0 89632 800 89752
rect 429200 89768 430000 89888
rect 0 88544 800 88664
rect 429200 87864 430000 87984
rect 0 87456 800 87576
rect 0 86368 800 86488
rect 429200 85960 430000 86080
rect 0 85280 800 85400
rect 0 84192 800 84312
rect 429200 84056 430000 84176
rect 0 83104 800 83224
rect 0 82016 800 82136
rect 429200 82016 430000 82136
rect 0 80928 800 81048
rect 0 79976 800 80096
rect 429200 80112 430000 80232
rect 0 78888 800 79008
rect 429200 78208 430000 78328
rect 0 77800 800 77920
rect 0 76712 800 76832
rect 429200 76304 430000 76424
rect 0 75624 800 75744
rect 0 74536 800 74656
rect 429200 74400 430000 74520
rect 0 73448 800 73568
rect 0 72360 800 72480
rect 429200 72360 430000 72480
rect 0 71272 800 71392
rect 429200 70456 430000 70576
rect 0 70184 800 70304
rect 0 69232 800 69352
rect 429200 68552 430000 68672
rect 0 68144 800 68264
rect 0 67056 800 67176
rect 429200 66648 430000 66768
rect 0 65968 800 66088
rect 0 64880 800 65000
rect 429200 64744 430000 64864
rect 0 63792 800 63912
rect 0 62704 800 62824
rect 429200 62704 430000 62824
rect 0 61616 800 61736
rect 429200 60800 430000 60920
rect 0 60528 800 60648
rect 0 59440 800 59560
rect 429200 58896 430000 59016
rect 0 58352 800 58472
rect 0 57400 800 57520
rect 429200 56992 430000 57112
rect 0 56312 800 56432
rect 0 55224 800 55344
rect 429200 54952 430000 55072
rect 0 54136 800 54256
rect 0 53048 800 53168
rect 429200 53048 430000 53168
rect 0 51960 800 52080
rect 429200 51144 430000 51264
rect 0 50872 800 50992
rect 0 49784 800 49904
rect 429200 49240 430000 49360
rect 0 48696 800 48816
rect 0 47608 800 47728
rect 429200 47336 430000 47456
rect 0 46520 800 46640
rect 0 45568 800 45688
rect 429200 45296 430000 45416
rect 0 44480 800 44600
rect 0 43392 800 43512
rect 429200 43392 430000 43512
rect 0 42304 800 42424
rect 429200 41488 430000 41608
rect 0 41216 800 41336
rect 0 40128 800 40248
rect 429200 39584 430000 39704
rect 0 39040 800 39160
rect 0 37952 800 38072
rect 429200 37680 430000 37800
rect 0 36864 800 36984
rect 0 35776 800 35896
rect 429200 35640 430000 35760
rect 0 34824 800 34944
rect 0 33736 800 33856
rect 429200 33736 430000 33856
rect 0 32648 800 32768
rect 429200 31832 430000 31952
rect 0 31560 800 31680
rect 0 30472 800 30592
rect 429200 29928 430000 30048
rect 0 29384 800 29504
rect 0 28296 800 28416
rect 429200 27888 430000 28008
rect 0 27208 800 27328
rect 0 26120 800 26240
rect 429200 25984 430000 26104
rect 0 25032 800 25152
rect 0 23944 800 24064
rect 429200 24080 430000 24200
rect 0 22992 800 23112
rect 429200 22176 430000 22296
rect 0 21904 800 22024
rect 0 20816 800 20936
rect 429200 20272 430000 20392
rect 0 19728 800 19848
rect 0 18640 800 18760
rect 429200 18232 430000 18352
rect 0 17552 800 17672
rect 0 16464 800 16584
rect 429200 16328 430000 16448
rect 0 15376 800 15496
rect 0 14288 800 14408
rect 429200 14424 430000 14544
rect 0 13200 800 13320
rect 429200 12520 430000 12640
rect 0 12112 800 12232
rect 0 11160 800 11280
rect 429200 10616 430000 10736
rect 0 10072 800 10192
rect 0 8984 800 9104
rect 429200 8576 430000 8696
rect 0 7896 800 8016
rect 0 6808 800 6928
rect 429200 6672 430000 6792
rect 0 5720 800 5840
rect 0 4632 800 4752
rect 429200 4768 430000 4888
rect 0 3544 800 3664
rect 429200 2864 430000 2984
rect 0 2456 800 2576
rect 0 1368 800 1488
rect 429200 960 430000 1080
rect 0 416 800 536
<< obsm3 >>
rect 880 171288 429200 171461
rect 800 171160 429200 171288
rect 800 170880 429120 171160
rect 800 170480 429200 170880
rect 880 170200 429200 170480
rect 800 169392 429200 170200
rect 880 169256 429200 169392
rect 880 169112 429120 169256
rect 800 168976 429120 169112
rect 800 168304 429200 168976
rect 880 168024 429200 168304
rect 800 167352 429200 168024
rect 800 167216 429120 167352
rect 880 167072 429120 167216
rect 880 166936 429200 167072
rect 800 166128 429200 166936
rect 880 165848 429200 166128
rect 800 165448 429200 165848
rect 800 165168 429120 165448
rect 800 165040 429200 165168
rect 880 164760 429200 165040
rect 800 163952 429200 164760
rect 880 163672 429200 163952
rect 800 163408 429200 163672
rect 800 163128 429120 163408
rect 800 162864 429200 163128
rect 880 162584 429200 162864
rect 800 161776 429200 162584
rect 880 161504 429200 161776
rect 880 161496 429120 161504
rect 800 161224 429120 161496
rect 800 160824 429200 161224
rect 880 160544 429200 160824
rect 800 159736 429200 160544
rect 880 159600 429200 159736
rect 880 159456 429120 159600
rect 800 159320 429120 159456
rect 800 158648 429200 159320
rect 880 158368 429200 158648
rect 800 157696 429200 158368
rect 800 157560 429120 157696
rect 880 157416 429120 157560
rect 880 157280 429200 157416
rect 800 156472 429200 157280
rect 880 156192 429200 156472
rect 800 155792 429200 156192
rect 800 155512 429120 155792
rect 800 155384 429200 155512
rect 880 155104 429200 155384
rect 800 154296 429200 155104
rect 880 154016 429200 154296
rect 800 153752 429200 154016
rect 800 153472 429120 153752
rect 800 153208 429200 153472
rect 880 152928 429200 153208
rect 800 152120 429200 152928
rect 880 151848 429200 152120
rect 880 151840 429120 151848
rect 800 151568 429120 151840
rect 800 151032 429200 151568
rect 880 150752 429200 151032
rect 800 149944 429200 150752
rect 880 149664 429120 149944
rect 800 148992 429200 149664
rect 880 148712 429200 148992
rect 800 148040 429200 148712
rect 800 147904 429120 148040
rect 880 147760 429120 147904
rect 880 147624 429200 147760
rect 800 146816 429200 147624
rect 880 146536 429200 146816
rect 800 146136 429200 146536
rect 800 145856 429120 146136
rect 800 145728 429200 145856
rect 880 145448 429200 145728
rect 800 144640 429200 145448
rect 880 144360 429200 144640
rect 800 144096 429200 144360
rect 800 143816 429120 144096
rect 800 143552 429200 143816
rect 880 143272 429200 143552
rect 800 142464 429200 143272
rect 880 142192 429200 142464
rect 880 142184 429120 142192
rect 800 141912 429120 142184
rect 800 141376 429200 141912
rect 880 141096 429200 141376
rect 800 140288 429200 141096
rect 880 140008 429120 140288
rect 800 139200 429200 140008
rect 880 138920 429200 139200
rect 800 138384 429200 138920
rect 800 138248 429120 138384
rect 880 138104 429120 138248
rect 880 137968 429200 138104
rect 800 137160 429200 137968
rect 880 136880 429200 137160
rect 800 136344 429200 136880
rect 800 136072 429120 136344
rect 880 136064 429120 136072
rect 880 135792 429200 136064
rect 800 134984 429200 135792
rect 880 134704 429200 134984
rect 800 134440 429200 134704
rect 800 134160 429120 134440
rect 800 133896 429200 134160
rect 880 133616 429200 133896
rect 800 132808 429200 133616
rect 880 132536 429200 132808
rect 880 132528 429120 132536
rect 800 132256 429120 132528
rect 800 131720 429200 132256
rect 880 131440 429200 131720
rect 800 130632 429200 131440
rect 880 130352 429120 130632
rect 800 129544 429200 130352
rect 880 129264 429200 129544
rect 800 128728 429200 129264
rect 800 128456 429120 128728
rect 880 128448 429120 128456
rect 880 128176 429200 128448
rect 800 127368 429200 128176
rect 880 127088 429200 127368
rect 800 126688 429200 127088
rect 800 126416 429120 126688
rect 880 126408 429120 126416
rect 880 126136 429200 126408
rect 800 125328 429200 126136
rect 880 125048 429200 125328
rect 800 124784 429200 125048
rect 800 124504 429120 124784
rect 800 124240 429200 124504
rect 880 123960 429200 124240
rect 800 123152 429200 123960
rect 880 122880 429200 123152
rect 880 122872 429120 122880
rect 800 122600 429120 122872
rect 800 122064 429200 122600
rect 880 121784 429200 122064
rect 800 120976 429200 121784
rect 880 120696 429120 120976
rect 800 119888 429200 120696
rect 880 119608 429200 119888
rect 800 119072 429200 119608
rect 800 118800 429120 119072
rect 880 118792 429120 118800
rect 880 118520 429200 118792
rect 800 117712 429200 118520
rect 880 117432 429200 117712
rect 800 117032 429200 117432
rect 800 116752 429120 117032
rect 800 116624 429200 116752
rect 880 116344 429200 116624
rect 800 115536 429200 116344
rect 880 115256 429200 115536
rect 800 115128 429200 115256
rect 800 114848 429120 115128
rect 800 114584 429200 114848
rect 880 114304 429200 114584
rect 800 113496 429200 114304
rect 880 113224 429200 113496
rect 880 113216 429120 113224
rect 800 112944 429120 113216
rect 800 112408 429200 112944
rect 880 112128 429200 112408
rect 800 111320 429200 112128
rect 880 111040 429120 111320
rect 800 110232 429200 111040
rect 880 109952 429200 110232
rect 800 109280 429200 109952
rect 800 109144 429120 109280
rect 880 109000 429120 109144
rect 880 108864 429200 109000
rect 800 108056 429200 108864
rect 880 107776 429200 108056
rect 800 107376 429200 107776
rect 800 107096 429120 107376
rect 800 106968 429200 107096
rect 880 106688 429200 106968
rect 800 105880 429200 106688
rect 880 105600 429200 105880
rect 800 105472 429200 105600
rect 800 105192 429120 105472
rect 800 104792 429200 105192
rect 880 104512 429200 104792
rect 800 103840 429200 104512
rect 880 103568 429200 103840
rect 880 103560 429120 103568
rect 800 103288 429120 103560
rect 800 102752 429200 103288
rect 880 102472 429200 102752
rect 800 101664 429200 102472
rect 880 101384 429120 101664
rect 800 100576 429200 101384
rect 880 100296 429200 100576
rect 800 99624 429200 100296
rect 800 99488 429120 99624
rect 880 99344 429120 99488
rect 880 99208 429200 99344
rect 800 98400 429200 99208
rect 880 98120 429200 98400
rect 800 97720 429200 98120
rect 800 97440 429120 97720
rect 800 97312 429200 97440
rect 880 97032 429200 97312
rect 800 96224 429200 97032
rect 880 95944 429200 96224
rect 800 95816 429200 95944
rect 800 95536 429120 95816
rect 800 95136 429200 95536
rect 880 94856 429200 95136
rect 800 94048 429200 94856
rect 880 93912 429200 94048
rect 880 93768 429120 93912
rect 800 93632 429120 93768
rect 800 92960 429200 93632
rect 880 92680 429200 92960
rect 800 92008 429200 92680
rect 880 91728 429120 92008
rect 800 90920 429200 91728
rect 880 90640 429200 90920
rect 800 89968 429200 90640
rect 800 89832 429120 89968
rect 880 89688 429120 89832
rect 880 89552 429200 89688
rect 800 88744 429200 89552
rect 880 88464 429200 88744
rect 800 88064 429200 88464
rect 800 87784 429120 88064
rect 800 87656 429200 87784
rect 880 87376 429200 87656
rect 800 86568 429200 87376
rect 880 86288 429200 86568
rect 800 86160 429200 86288
rect 800 85880 429120 86160
rect 800 85480 429200 85880
rect 880 85200 429200 85480
rect 800 84392 429200 85200
rect 880 84256 429200 84392
rect 880 84112 429120 84256
rect 800 83976 429120 84112
rect 800 83304 429200 83976
rect 880 83024 429200 83304
rect 800 82216 429200 83024
rect 880 81936 429120 82216
rect 800 81128 429200 81936
rect 880 80848 429200 81128
rect 800 80312 429200 80848
rect 800 80176 429120 80312
rect 880 80032 429120 80176
rect 880 79896 429200 80032
rect 800 79088 429200 79896
rect 880 78808 429200 79088
rect 800 78408 429200 78808
rect 800 78128 429120 78408
rect 800 78000 429200 78128
rect 880 77720 429200 78000
rect 800 76912 429200 77720
rect 880 76632 429200 76912
rect 800 76504 429200 76632
rect 800 76224 429120 76504
rect 800 75824 429200 76224
rect 880 75544 429200 75824
rect 800 74736 429200 75544
rect 880 74600 429200 74736
rect 880 74456 429120 74600
rect 800 74320 429120 74456
rect 800 73648 429200 74320
rect 880 73368 429200 73648
rect 800 72560 429200 73368
rect 880 72280 429120 72560
rect 800 71472 429200 72280
rect 880 71192 429200 71472
rect 800 70656 429200 71192
rect 800 70384 429120 70656
rect 880 70376 429120 70384
rect 880 70104 429200 70376
rect 800 69432 429200 70104
rect 880 69152 429200 69432
rect 800 68752 429200 69152
rect 800 68472 429120 68752
rect 800 68344 429200 68472
rect 880 68064 429200 68344
rect 800 67256 429200 68064
rect 880 66976 429200 67256
rect 800 66848 429200 66976
rect 800 66568 429120 66848
rect 800 66168 429200 66568
rect 880 65888 429200 66168
rect 800 65080 429200 65888
rect 880 64944 429200 65080
rect 880 64800 429120 64944
rect 800 64664 429120 64800
rect 800 63992 429200 64664
rect 880 63712 429200 63992
rect 800 62904 429200 63712
rect 880 62624 429120 62904
rect 800 61816 429200 62624
rect 880 61536 429200 61816
rect 800 61000 429200 61536
rect 800 60728 429120 61000
rect 880 60720 429120 60728
rect 880 60448 429200 60720
rect 800 59640 429200 60448
rect 880 59360 429200 59640
rect 800 59096 429200 59360
rect 800 58816 429120 59096
rect 800 58552 429200 58816
rect 880 58272 429200 58552
rect 800 57600 429200 58272
rect 880 57320 429200 57600
rect 800 57192 429200 57320
rect 800 56912 429120 57192
rect 800 56512 429200 56912
rect 880 56232 429200 56512
rect 800 55424 429200 56232
rect 880 55152 429200 55424
rect 880 55144 429120 55152
rect 800 54872 429120 55144
rect 800 54336 429200 54872
rect 880 54056 429200 54336
rect 800 53248 429200 54056
rect 880 52968 429120 53248
rect 800 52160 429200 52968
rect 880 51880 429200 52160
rect 800 51344 429200 51880
rect 800 51072 429120 51344
rect 880 51064 429120 51072
rect 880 50792 429200 51064
rect 800 49984 429200 50792
rect 880 49704 429200 49984
rect 800 49440 429200 49704
rect 800 49160 429120 49440
rect 800 48896 429200 49160
rect 880 48616 429200 48896
rect 800 47808 429200 48616
rect 880 47536 429200 47808
rect 880 47528 429120 47536
rect 800 47256 429120 47528
rect 800 46720 429200 47256
rect 880 46440 429200 46720
rect 800 45768 429200 46440
rect 880 45496 429200 45768
rect 880 45488 429120 45496
rect 800 45216 429120 45488
rect 800 44680 429200 45216
rect 880 44400 429200 44680
rect 800 43592 429200 44400
rect 880 43312 429120 43592
rect 800 42504 429200 43312
rect 880 42224 429200 42504
rect 800 41688 429200 42224
rect 800 41416 429120 41688
rect 880 41408 429120 41416
rect 880 41136 429200 41408
rect 800 40328 429200 41136
rect 880 40048 429200 40328
rect 800 39784 429200 40048
rect 800 39504 429120 39784
rect 800 39240 429200 39504
rect 880 38960 429200 39240
rect 800 38152 429200 38960
rect 880 37880 429200 38152
rect 880 37872 429120 37880
rect 800 37600 429120 37872
rect 800 37064 429200 37600
rect 880 36784 429200 37064
rect 800 35976 429200 36784
rect 880 35840 429200 35976
rect 880 35696 429120 35840
rect 800 35560 429120 35696
rect 800 35024 429200 35560
rect 880 34744 429200 35024
rect 800 33936 429200 34744
rect 880 33656 429120 33936
rect 800 32848 429200 33656
rect 880 32568 429200 32848
rect 800 32032 429200 32568
rect 800 31760 429120 32032
rect 880 31752 429120 31760
rect 880 31480 429200 31752
rect 800 30672 429200 31480
rect 880 30392 429200 30672
rect 800 30128 429200 30392
rect 800 29848 429120 30128
rect 800 29584 429200 29848
rect 880 29304 429200 29584
rect 800 28496 429200 29304
rect 880 28216 429200 28496
rect 800 28088 429200 28216
rect 800 27808 429120 28088
rect 800 27408 429200 27808
rect 880 27128 429200 27408
rect 800 26320 429200 27128
rect 880 26184 429200 26320
rect 880 26040 429120 26184
rect 800 25904 429120 26040
rect 800 25232 429200 25904
rect 880 24952 429200 25232
rect 800 24280 429200 24952
rect 800 24144 429120 24280
rect 880 24000 429120 24144
rect 880 23864 429200 24000
rect 800 23192 429200 23864
rect 880 22912 429200 23192
rect 800 22376 429200 22912
rect 800 22104 429120 22376
rect 880 22096 429120 22104
rect 880 21824 429200 22096
rect 800 21016 429200 21824
rect 880 20736 429200 21016
rect 800 20472 429200 20736
rect 800 20192 429120 20472
rect 800 19928 429200 20192
rect 880 19648 429200 19928
rect 800 18840 429200 19648
rect 880 18560 429200 18840
rect 800 18432 429200 18560
rect 800 18152 429120 18432
rect 800 17752 429200 18152
rect 880 17472 429200 17752
rect 800 16664 429200 17472
rect 880 16528 429200 16664
rect 880 16384 429120 16528
rect 800 16248 429120 16384
rect 800 15576 429200 16248
rect 880 15296 429200 15576
rect 800 14624 429200 15296
rect 800 14488 429120 14624
rect 880 14344 429120 14488
rect 880 14208 429200 14344
rect 800 13400 429200 14208
rect 880 13120 429200 13400
rect 800 12720 429200 13120
rect 800 12440 429120 12720
rect 800 12312 429200 12440
rect 880 12032 429200 12312
rect 800 11360 429200 12032
rect 880 11080 429200 11360
rect 800 10816 429200 11080
rect 800 10536 429120 10816
rect 800 10272 429200 10536
rect 880 9992 429200 10272
rect 800 9184 429200 9992
rect 880 8904 429200 9184
rect 800 8776 429200 8904
rect 800 8496 429120 8776
rect 800 8096 429200 8496
rect 880 7816 429200 8096
rect 800 7008 429200 7816
rect 880 6872 429200 7008
rect 880 6728 429120 6872
rect 800 6592 429120 6728
rect 800 5920 429200 6592
rect 880 5640 429200 5920
rect 800 4968 429200 5640
rect 800 4832 429120 4968
rect 880 4688 429120 4832
rect 880 4552 429200 4688
rect 800 3744 429200 4552
rect 880 3464 429200 3744
rect 800 3064 429200 3464
rect 800 2784 429120 3064
rect 800 2656 429200 2784
rect 880 2376 429200 2656
rect 800 1568 429200 2376
rect 880 1288 429200 1568
rect 800 1160 429200 1288
rect 800 880 429120 1160
rect 800 616 429200 880
rect 880 443 429200 616
<< metal4 >>
rect 4208 2128 4528 169776
rect 9208 2128 9528 169776
rect 14208 2128 14528 169776
rect 19208 2128 19528 169776
rect 24208 128152 24528 169776
rect 29208 128152 29528 169776
rect 34208 128152 34528 169776
rect 39208 128152 39528 169776
rect 44208 128152 44528 169776
rect 49208 128152 49528 169776
rect 54208 128152 54528 169776
rect 59208 128152 59528 169776
rect 64208 128152 64528 169776
rect 69208 128152 69528 169776
rect 74208 128152 74528 169776
rect 79208 128152 79528 169776
rect 84208 128152 84528 169776
rect 89208 128152 89528 169776
rect 94208 128152 94528 169776
rect 99208 128152 99528 169776
rect 104208 128152 104528 169776
rect 109208 128152 109528 169776
rect 114208 128152 114528 169776
rect 119208 128152 119528 169776
rect 124208 128152 124528 169776
rect 129208 128152 129528 169776
rect 134208 128152 134528 169776
rect 139208 128152 139528 169776
rect 144208 128152 144528 169776
rect 149208 128152 149528 169776
rect 154208 128152 154528 169776
rect 159208 128152 159528 169776
rect 164208 128152 164528 169776
rect 169208 128152 169528 169776
rect 174208 128152 174528 169776
rect 24208 2128 24528 21248
rect 29208 2128 29528 21248
rect 34208 2128 34528 21248
rect 39208 2128 39528 21248
rect 44208 2128 44528 21248
rect 49208 2128 49528 21248
rect 54208 2128 54528 21248
rect 59208 2128 59528 21248
rect 64208 2128 64528 21248
rect 69208 2128 69528 21248
rect 74208 2128 74528 21248
rect 79208 2128 79528 21248
rect 84208 2128 84528 21248
rect 89208 2128 89528 21248
rect 94208 2128 94528 21248
rect 99208 2128 99528 21248
rect 104208 2128 104528 21248
rect 109208 2128 109528 21248
rect 114208 2128 114528 21248
rect 119208 2128 119528 21248
rect 124208 2128 124528 21248
rect 129208 2128 129528 21248
rect 134208 2128 134528 21248
rect 139208 2128 139528 21248
rect 144208 2128 144528 21248
rect 149208 2128 149528 21248
rect 154208 2128 154528 21248
rect 159208 2128 159528 21248
rect 164208 2128 164528 21248
rect 169208 2128 169528 21248
rect 174208 2128 174528 21248
rect 179208 2128 179528 169776
rect 184208 2128 184528 169776
rect 189208 2128 189528 169776
rect 194208 2128 194528 169776
rect 199208 2128 199528 169776
rect 204208 2128 204528 169776
rect 209208 2128 209528 169776
rect 214208 2128 214528 169776
rect 219208 2128 219528 169776
rect 224208 2128 224528 169776
rect 229208 2128 229528 169776
rect 234208 2128 234528 169776
rect 239208 2128 239528 169776
rect 244208 2128 244528 169776
rect 249208 2128 249528 169776
rect 254208 2128 254528 169776
rect 259208 2128 259528 169776
rect 264208 2128 264528 169776
rect 269208 2128 269528 169776
rect 274208 2128 274528 169776
rect 279208 2128 279528 169776
rect 284208 2128 284528 169776
rect 289208 2128 289528 169776
rect 294208 2128 294528 169776
rect 299208 2128 299528 169776
rect 304208 2128 304528 169776
rect 309208 2128 309528 169776
rect 314208 2128 314528 169776
rect 319208 2128 319528 169776
rect 324208 2128 324528 169776
rect 329208 2128 329528 169776
rect 334208 2128 334528 169776
rect 339208 2128 339528 169776
rect 344208 2128 344528 169776
rect 349208 2128 349528 169776
rect 354208 2128 354528 169776
rect 359208 2128 359528 169776
rect 364208 2128 364528 169776
rect 369208 2128 369528 169776
rect 374208 2128 374528 169776
rect 379208 2128 379528 169776
rect 384208 2128 384528 169776
rect 389208 164296 389528 169776
rect 394208 164296 394528 169776
rect 399208 164296 399528 169776
rect 389208 2128 389528 145392
rect 394208 2128 394528 145392
rect 399208 2128 399528 145392
rect 404208 2128 404528 169776
rect 409208 2128 409528 169776
rect 414208 2128 414528 169776
rect 419208 2128 419528 169776
rect 424208 2128 424528 169776
<< obsm4 >>
rect 1715 169856 426453 171189
rect 1715 2347 4128 169856
rect 4608 2347 9128 169856
rect 9608 2347 14128 169856
rect 14608 2347 19128 169856
rect 19608 128072 24128 169856
rect 24608 128072 29128 169856
rect 29608 128072 34128 169856
rect 34608 128072 39128 169856
rect 39608 128072 44128 169856
rect 44608 128072 49128 169856
rect 49608 128072 54128 169856
rect 54608 128072 59128 169856
rect 59608 128072 64128 169856
rect 64608 128072 69128 169856
rect 69608 128072 74128 169856
rect 74608 128072 79128 169856
rect 79608 128072 84128 169856
rect 84608 128072 89128 169856
rect 89608 128072 94128 169856
rect 94608 128072 99128 169856
rect 99608 128072 104128 169856
rect 104608 128072 109128 169856
rect 109608 128072 114128 169856
rect 114608 128072 119128 169856
rect 119608 128072 124128 169856
rect 124608 128072 129128 169856
rect 129608 128072 134128 169856
rect 134608 128072 139128 169856
rect 139608 128072 144128 169856
rect 144608 128072 149128 169856
rect 149608 128072 154128 169856
rect 154608 128072 159128 169856
rect 159608 128072 164128 169856
rect 164608 128072 169128 169856
rect 169608 128072 174128 169856
rect 174608 128072 179128 169856
rect 19608 21328 179128 128072
rect 19608 2347 24128 21328
rect 24608 2347 29128 21328
rect 29608 2347 34128 21328
rect 34608 2347 39128 21328
rect 39608 2347 44128 21328
rect 44608 2347 49128 21328
rect 49608 2347 54128 21328
rect 54608 2347 59128 21328
rect 59608 2347 64128 21328
rect 64608 2347 69128 21328
rect 69608 2347 74128 21328
rect 74608 2347 79128 21328
rect 79608 2347 84128 21328
rect 84608 2347 89128 21328
rect 89608 2347 94128 21328
rect 94608 2347 99128 21328
rect 99608 2347 104128 21328
rect 104608 2347 109128 21328
rect 109608 2347 114128 21328
rect 114608 2347 119128 21328
rect 119608 2347 124128 21328
rect 124608 2347 129128 21328
rect 129608 2347 134128 21328
rect 134608 2347 139128 21328
rect 139608 2347 144128 21328
rect 144608 2347 149128 21328
rect 149608 2347 154128 21328
rect 154608 2347 159128 21328
rect 159608 2347 164128 21328
rect 164608 2347 169128 21328
rect 169608 2347 174128 21328
rect 174608 2347 179128 21328
rect 179608 2347 184128 169856
rect 184608 2347 189128 169856
rect 189608 2347 194128 169856
rect 194608 2347 199128 169856
rect 199608 2347 204128 169856
rect 204608 2347 209128 169856
rect 209608 2347 214128 169856
rect 214608 2347 219128 169856
rect 219608 2347 224128 169856
rect 224608 2347 229128 169856
rect 229608 2347 234128 169856
rect 234608 2347 239128 169856
rect 239608 2347 244128 169856
rect 244608 2347 249128 169856
rect 249608 2347 254128 169856
rect 254608 2347 259128 169856
rect 259608 2347 264128 169856
rect 264608 2347 269128 169856
rect 269608 2347 274128 169856
rect 274608 2347 279128 169856
rect 279608 2347 284128 169856
rect 284608 2347 289128 169856
rect 289608 2347 294128 169856
rect 294608 2347 299128 169856
rect 299608 2347 304128 169856
rect 304608 2347 309128 169856
rect 309608 2347 314128 169856
rect 314608 2347 319128 169856
rect 319608 2347 324128 169856
rect 324608 2347 329128 169856
rect 329608 2347 334128 169856
rect 334608 2347 339128 169856
rect 339608 2347 344128 169856
rect 344608 2347 349128 169856
rect 349608 2347 354128 169856
rect 354608 2347 359128 169856
rect 359608 2347 364128 169856
rect 364608 2347 369128 169856
rect 369608 2347 374128 169856
rect 374608 2347 379128 169856
rect 379608 2347 384128 169856
rect 384608 164216 389128 169856
rect 389608 164216 394128 169856
rect 394608 164216 399128 169856
rect 399608 164216 404128 169856
rect 384608 145472 404128 164216
rect 384608 2347 389128 145472
rect 389608 2347 394128 145472
rect 394608 2347 399128 145472
rect 399608 2347 404128 145472
rect 404608 2347 409128 169856
rect 409608 2347 414128 169856
rect 414608 2347 419128 169856
rect 419608 2347 424128 169856
rect 424608 2347 426453 169856
<< metal5 >>
rect 1104 161298 428812 161618
rect 1104 148298 428812 148618
rect 1104 135298 428812 135618
rect 1104 122298 428812 122618
rect 1104 109298 428812 109618
rect 1104 96298 428812 96618
rect 1104 83298 428812 83618
rect 1104 70298 428812 70618
rect 1104 57298 428812 57618
rect 1104 44298 428812 44618
rect 1104 31298 428812 31618
rect 1104 18298 428812 18618
rect 1104 5298 428812 5618
<< labels >>
rlabel metal2 s 29274 0 29330 800 6 clock
port 1 nsew signal input
rlabel metal2 s 294 171200 350 172000 6 core_clk
port 2 nsew signal output
rlabel metal2 s 938 171200 994 172000 6 core_rstn
port 3 nsew signal output
rlabel metal2 s 224774 0 224830 800 6 flash_clk
port 4 nsew signal output
rlabel metal2 s 244278 0 244334 800 6 flash_clk_ieb
port 5 nsew signal output
rlabel metal2 s 263782 0 263838 800 6 flash_clk_oeb
port 6 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 flash_csb
port 7 nsew signal output
rlabel metal2 s 185674 0 185730 800 6 flash_csb_ieb
port 8 nsew signal output
rlabel metal2 s 205178 0 205234 800 6 flash_csb_oeb
port 9 nsew signal output
rlabel metal2 s 283378 0 283434 800 6 flash_io0_di
port 10 nsew signal input
rlabel metal2 s 302882 0 302938 800 6 flash_io0_do
port 11 nsew signal output
rlabel metal2 s 322478 0 322534 800 6 flash_io0_ieb
port 12 nsew signal output
rlabel metal2 s 341982 0 342038 800 6 flash_io0_oeb
port 13 nsew signal output
rlabel metal2 s 361578 0 361634 800 6 flash_io1_di
port 14 nsew signal input
rlabel metal2 s 381082 0 381138 800 6 flash_io1_do
port 15 nsew signal output
rlabel metal2 s 400678 0 400734 800 6 flash_io1_ieb
port 16 nsew signal output
rlabel metal2 s 420182 0 420238 800 6 flash_io1_oeb
port 17 nsew signal output
rlabel metal3 s 0 169192 800 169312 6 flash_io2_do
port 18 nsew signal output
rlabel metal3 s 429200 169056 430000 169176 6 flash_io2_oeb
port 19 nsew signal output
rlabel metal3 s 429200 170960 430000 171080 6 flash_io3_do
port 20 nsew signal output
rlabel metal3 s 0 170280 800 170400 6 flash_io3_oeb
port 21 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 gpio_inenb_pad
port 23 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 gpio_mode0_pad
port 24 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 gpio_mode1_pad
port 25 nsew signal output
rlabel metal2 s 126978 0 127034 800 6 gpio_out_pad
port 26 nsew signal output
rlabel metal2 s 146574 0 146630 800 6 gpio_outenb_pad
port 27 nsew signal output
rlabel metal3 s 429200 64744 430000 64864 6 jtag_out
port 28 nsew signal output
rlabel metal3 s 429200 66648 430000 66768 6 jtag_outenb
port 29 nsew signal output
rlabel metal2 s 87970 171200 88026 172000 6 la_iena[0]
port 30 nsew signal output
rlabel metal2 s 152922 171200 152978 172000 6 la_iena[100]
port 31 nsew signal output
rlabel metal2 s 153566 171200 153622 172000 6 la_iena[101]
port 32 nsew signal output
rlabel metal2 s 154210 171200 154266 172000 6 la_iena[102]
port 33 nsew signal output
rlabel metal2 s 154854 171200 154910 172000 6 la_iena[103]
port 34 nsew signal output
rlabel metal2 s 155498 171200 155554 172000 6 la_iena[104]
port 35 nsew signal output
rlabel metal2 s 156142 171200 156198 172000 6 la_iena[105]
port 36 nsew signal output
rlabel metal2 s 156786 171200 156842 172000 6 la_iena[106]
port 37 nsew signal output
rlabel metal2 s 157430 171200 157486 172000 6 la_iena[107]
port 38 nsew signal output
rlabel metal2 s 158074 171200 158130 172000 6 la_iena[108]
port 39 nsew signal output
rlabel metal2 s 158718 171200 158774 172000 6 la_iena[109]
port 40 nsew signal output
rlabel metal2 s 94410 171200 94466 172000 6 la_iena[10]
port 41 nsew signal output
rlabel metal2 s 159362 171200 159418 172000 6 la_iena[110]
port 42 nsew signal output
rlabel metal2 s 160006 171200 160062 172000 6 la_iena[111]
port 43 nsew signal output
rlabel metal2 s 160650 171200 160706 172000 6 la_iena[112]
port 44 nsew signal output
rlabel metal2 s 161294 171200 161350 172000 6 la_iena[113]
port 45 nsew signal output
rlabel metal2 s 162030 171200 162086 172000 6 la_iena[114]
port 46 nsew signal output
rlabel metal2 s 162674 171200 162730 172000 6 la_iena[115]
port 47 nsew signal output
rlabel metal2 s 163318 171200 163374 172000 6 la_iena[116]
port 48 nsew signal output
rlabel metal2 s 163962 171200 164018 172000 6 la_iena[117]
port 49 nsew signal output
rlabel metal2 s 164606 171200 164662 172000 6 la_iena[118]
port 50 nsew signal output
rlabel metal2 s 165250 171200 165306 172000 6 la_iena[119]
port 51 nsew signal output
rlabel metal2 s 95054 171200 95110 172000 6 la_iena[11]
port 52 nsew signal output
rlabel metal2 s 165894 171200 165950 172000 6 la_iena[120]
port 53 nsew signal output
rlabel metal2 s 166538 171200 166594 172000 6 la_iena[121]
port 54 nsew signal output
rlabel metal2 s 167182 171200 167238 172000 6 la_iena[122]
port 55 nsew signal output
rlabel metal2 s 167826 171200 167882 172000 6 la_iena[123]
port 56 nsew signal output
rlabel metal2 s 168470 171200 168526 172000 6 la_iena[124]
port 57 nsew signal output
rlabel metal2 s 169114 171200 169170 172000 6 la_iena[125]
port 58 nsew signal output
rlabel metal2 s 169758 171200 169814 172000 6 la_iena[126]
port 59 nsew signal output
rlabel metal2 s 170402 171200 170458 172000 6 la_iena[127]
port 60 nsew signal output
rlabel metal2 s 95698 171200 95754 172000 6 la_iena[12]
port 61 nsew signal output
rlabel metal2 s 96342 171200 96398 172000 6 la_iena[13]
port 62 nsew signal output
rlabel metal2 s 97078 171200 97134 172000 6 la_iena[14]
port 63 nsew signal output
rlabel metal2 s 97722 171200 97778 172000 6 la_iena[15]
port 64 nsew signal output
rlabel metal2 s 98366 171200 98422 172000 6 la_iena[16]
port 65 nsew signal output
rlabel metal2 s 99010 171200 99066 172000 6 la_iena[17]
port 66 nsew signal output
rlabel metal2 s 99654 171200 99710 172000 6 la_iena[18]
port 67 nsew signal output
rlabel metal2 s 100298 171200 100354 172000 6 la_iena[19]
port 68 nsew signal output
rlabel metal2 s 88614 171200 88670 172000 6 la_iena[1]
port 69 nsew signal output
rlabel metal2 s 100942 171200 100998 172000 6 la_iena[20]
port 70 nsew signal output
rlabel metal2 s 101586 171200 101642 172000 6 la_iena[21]
port 71 nsew signal output
rlabel metal2 s 102230 171200 102286 172000 6 la_iena[22]
port 72 nsew signal output
rlabel metal2 s 102874 171200 102930 172000 6 la_iena[23]
port 73 nsew signal output
rlabel metal2 s 103518 171200 103574 172000 6 la_iena[24]
port 74 nsew signal output
rlabel metal2 s 104162 171200 104218 172000 6 la_iena[25]
port 75 nsew signal output
rlabel metal2 s 104806 171200 104862 172000 6 la_iena[26]
port 76 nsew signal output
rlabel metal2 s 105450 171200 105506 172000 6 la_iena[27]
port 77 nsew signal output
rlabel metal2 s 106094 171200 106150 172000 6 la_iena[28]
port 78 nsew signal output
rlabel metal2 s 106738 171200 106794 172000 6 la_iena[29]
port 79 nsew signal output
rlabel metal2 s 89258 171200 89314 172000 6 la_iena[2]
port 80 nsew signal output
rlabel metal2 s 107382 171200 107438 172000 6 la_iena[30]
port 81 nsew signal output
rlabel metal2 s 108118 171200 108174 172000 6 la_iena[31]
port 82 nsew signal output
rlabel metal2 s 108762 171200 108818 172000 6 la_iena[32]
port 83 nsew signal output
rlabel metal2 s 109406 171200 109462 172000 6 la_iena[33]
port 84 nsew signal output
rlabel metal2 s 110050 171200 110106 172000 6 la_iena[34]
port 85 nsew signal output
rlabel metal2 s 110694 171200 110750 172000 6 la_iena[35]
port 86 nsew signal output
rlabel metal2 s 111338 171200 111394 172000 6 la_iena[36]
port 87 nsew signal output
rlabel metal2 s 111982 171200 112038 172000 6 la_iena[37]
port 88 nsew signal output
rlabel metal2 s 112626 171200 112682 172000 6 la_iena[38]
port 89 nsew signal output
rlabel metal2 s 113270 171200 113326 172000 6 la_iena[39]
port 90 nsew signal output
rlabel metal2 s 89902 171200 89958 172000 6 la_iena[3]
port 91 nsew signal output
rlabel metal2 s 113914 171200 113970 172000 6 la_iena[40]
port 92 nsew signal output
rlabel metal2 s 114558 171200 114614 172000 6 la_iena[41]
port 93 nsew signal output
rlabel metal2 s 115202 171200 115258 172000 6 la_iena[42]
port 94 nsew signal output
rlabel metal2 s 115846 171200 115902 172000 6 la_iena[43]
port 95 nsew signal output
rlabel metal2 s 116490 171200 116546 172000 6 la_iena[44]
port 96 nsew signal output
rlabel metal2 s 117134 171200 117190 172000 6 la_iena[45]
port 97 nsew signal output
rlabel metal2 s 117778 171200 117834 172000 6 la_iena[46]
port 98 nsew signal output
rlabel metal2 s 118422 171200 118478 172000 6 la_iena[47]
port 99 nsew signal output
rlabel metal2 s 119158 171200 119214 172000 6 la_iena[48]
port 100 nsew signal output
rlabel metal2 s 119802 171200 119858 172000 6 la_iena[49]
port 101 nsew signal output
rlabel metal2 s 90546 171200 90602 172000 6 la_iena[4]
port 102 nsew signal output
rlabel metal2 s 120446 171200 120502 172000 6 la_iena[50]
port 103 nsew signal output
rlabel metal2 s 121090 171200 121146 172000 6 la_iena[51]
port 104 nsew signal output
rlabel metal2 s 121734 171200 121790 172000 6 la_iena[52]
port 105 nsew signal output
rlabel metal2 s 122378 171200 122434 172000 6 la_iena[53]
port 106 nsew signal output
rlabel metal2 s 123022 171200 123078 172000 6 la_iena[54]
port 107 nsew signal output
rlabel metal2 s 123666 171200 123722 172000 6 la_iena[55]
port 108 nsew signal output
rlabel metal2 s 124310 171200 124366 172000 6 la_iena[56]
port 109 nsew signal output
rlabel metal2 s 124954 171200 125010 172000 6 la_iena[57]
port 110 nsew signal output
rlabel metal2 s 125598 171200 125654 172000 6 la_iena[58]
port 111 nsew signal output
rlabel metal2 s 126242 171200 126298 172000 6 la_iena[59]
port 112 nsew signal output
rlabel metal2 s 91190 171200 91246 172000 6 la_iena[5]
port 113 nsew signal output
rlabel metal2 s 126886 171200 126942 172000 6 la_iena[60]
port 114 nsew signal output
rlabel metal2 s 127530 171200 127586 172000 6 la_iena[61]
port 115 nsew signal output
rlabel metal2 s 128174 171200 128230 172000 6 la_iena[62]
port 116 nsew signal output
rlabel metal2 s 128818 171200 128874 172000 6 la_iena[63]
port 117 nsew signal output
rlabel metal2 s 129554 171200 129610 172000 6 la_iena[64]
port 118 nsew signal output
rlabel metal2 s 130198 171200 130254 172000 6 la_iena[65]
port 119 nsew signal output
rlabel metal2 s 130842 171200 130898 172000 6 la_iena[66]
port 120 nsew signal output
rlabel metal2 s 131486 171200 131542 172000 6 la_iena[67]
port 121 nsew signal output
rlabel metal2 s 132130 171200 132186 172000 6 la_iena[68]
port 122 nsew signal output
rlabel metal2 s 132774 171200 132830 172000 6 la_iena[69]
port 123 nsew signal output
rlabel metal2 s 91834 171200 91890 172000 6 la_iena[6]
port 124 nsew signal output
rlabel metal2 s 133418 171200 133474 172000 6 la_iena[70]
port 125 nsew signal output
rlabel metal2 s 134062 171200 134118 172000 6 la_iena[71]
port 126 nsew signal output
rlabel metal2 s 134706 171200 134762 172000 6 la_iena[72]
port 127 nsew signal output
rlabel metal2 s 135350 171200 135406 172000 6 la_iena[73]
port 128 nsew signal output
rlabel metal2 s 135994 171200 136050 172000 6 la_iena[74]
port 129 nsew signal output
rlabel metal2 s 136638 171200 136694 172000 6 la_iena[75]
port 130 nsew signal output
rlabel metal2 s 137282 171200 137338 172000 6 la_iena[76]
port 131 nsew signal output
rlabel metal2 s 137926 171200 137982 172000 6 la_iena[77]
port 132 nsew signal output
rlabel metal2 s 138570 171200 138626 172000 6 la_iena[78]
port 133 nsew signal output
rlabel metal2 s 139214 171200 139270 172000 6 la_iena[79]
port 134 nsew signal output
rlabel metal2 s 92478 171200 92534 172000 6 la_iena[7]
port 135 nsew signal output
rlabel metal2 s 139858 171200 139914 172000 6 la_iena[80]
port 136 nsew signal output
rlabel metal2 s 140594 171200 140650 172000 6 la_iena[81]
port 137 nsew signal output
rlabel metal2 s 141238 171200 141294 172000 6 la_iena[82]
port 138 nsew signal output
rlabel metal2 s 141882 171200 141938 172000 6 la_iena[83]
port 139 nsew signal output
rlabel metal2 s 142526 171200 142582 172000 6 la_iena[84]
port 140 nsew signal output
rlabel metal2 s 143170 171200 143226 172000 6 la_iena[85]
port 141 nsew signal output
rlabel metal2 s 143814 171200 143870 172000 6 la_iena[86]
port 142 nsew signal output
rlabel metal2 s 144458 171200 144514 172000 6 la_iena[87]
port 143 nsew signal output
rlabel metal2 s 145102 171200 145158 172000 6 la_iena[88]
port 144 nsew signal output
rlabel metal2 s 145746 171200 145802 172000 6 la_iena[89]
port 145 nsew signal output
rlabel metal2 s 93122 171200 93178 172000 6 la_iena[8]
port 146 nsew signal output
rlabel metal2 s 146390 171200 146446 172000 6 la_iena[90]
port 147 nsew signal output
rlabel metal2 s 147034 171200 147090 172000 6 la_iena[91]
port 148 nsew signal output
rlabel metal2 s 147678 171200 147734 172000 6 la_iena[92]
port 149 nsew signal output
rlabel metal2 s 148322 171200 148378 172000 6 la_iena[93]
port 150 nsew signal output
rlabel metal2 s 148966 171200 149022 172000 6 la_iena[94]
port 151 nsew signal output
rlabel metal2 s 149610 171200 149666 172000 6 la_iena[95]
port 152 nsew signal output
rlabel metal2 s 150254 171200 150310 172000 6 la_iena[96]
port 153 nsew signal output
rlabel metal2 s 150990 171200 151046 172000 6 la_iena[97]
port 154 nsew signal output
rlabel metal2 s 151634 171200 151690 172000 6 la_iena[98]
port 155 nsew signal output
rlabel metal2 s 152278 171200 152334 172000 6 la_iena[99]
port 156 nsew signal output
rlabel metal2 s 93766 171200 93822 172000 6 la_iena[9]
port 157 nsew signal output
rlabel metal2 s 171046 171200 171102 172000 6 la_input[0]
port 158 nsew signal input
rlabel metal2 s 235998 171200 236054 172000 6 la_input[100]
port 159 nsew signal input
rlabel metal2 s 236642 171200 236698 172000 6 la_input[101]
port 160 nsew signal input
rlabel metal2 s 237378 171200 237434 172000 6 la_input[102]
port 161 nsew signal input
rlabel metal2 s 238022 171200 238078 172000 6 la_input[103]
port 162 nsew signal input
rlabel metal2 s 238666 171200 238722 172000 6 la_input[104]
port 163 nsew signal input
rlabel metal2 s 239310 171200 239366 172000 6 la_input[105]
port 164 nsew signal input
rlabel metal2 s 239954 171200 240010 172000 6 la_input[106]
port 165 nsew signal input
rlabel metal2 s 240598 171200 240654 172000 6 la_input[107]
port 166 nsew signal input
rlabel metal2 s 241242 171200 241298 172000 6 la_input[108]
port 167 nsew signal input
rlabel metal2 s 241886 171200 241942 172000 6 la_input[109]
port 168 nsew signal input
rlabel metal2 s 177578 171200 177634 172000 6 la_input[10]
port 169 nsew signal input
rlabel metal2 s 242530 171200 242586 172000 6 la_input[110]
port 170 nsew signal input
rlabel metal2 s 243174 171200 243230 172000 6 la_input[111]
port 171 nsew signal input
rlabel metal2 s 243818 171200 243874 172000 6 la_input[112]
port 172 nsew signal input
rlabel metal2 s 244462 171200 244518 172000 6 la_input[113]
port 173 nsew signal input
rlabel metal2 s 245106 171200 245162 172000 6 la_input[114]
port 174 nsew signal input
rlabel metal2 s 245750 171200 245806 172000 6 la_input[115]
port 175 nsew signal input
rlabel metal2 s 246394 171200 246450 172000 6 la_input[116]
port 176 nsew signal input
rlabel metal2 s 247038 171200 247094 172000 6 la_input[117]
port 177 nsew signal input
rlabel metal2 s 247774 171200 247830 172000 6 la_input[118]
port 178 nsew signal input
rlabel metal2 s 248418 171200 248474 172000 6 la_input[119]
port 179 nsew signal input
rlabel metal2 s 178222 171200 178278 172000 6 la_input[11]
port 180 nsew signal input
rlabel metal2 s 249062 171200 249118 172000 6 la_input[120]
port 181 nsew signal input
rlabel metal2 s 249706 171200 249762 172000 6 la_input[121]
port 182 nsew signal input
rlabel metal2 s 250350 171200 250406 172000 6 la_input[122]
port 183 nsew signal input
rlabel metal2 s 250994 171200 251050 172000 6 la_input[123]
port 184 nsew signal input
rlabel metal2 s 251638 171200 251694 172000 6 la_input[124]
port 185 nsew signal input
rlabel metal2 s 252282 171200 252338 172000 6 la_input[125]
port 186 nsew signal input
rlabel metal2 s 252926 171200 252982 172000 6 la_input[126]
port 187 nsew signal input
rlabel metal2 s 253570 171200 253626 172000 6 la_input[127]
port 188 nsew signal input
rlabel metal2 s 178866 171200 178922 172000 6 la_input[12]
port 189 nsew signal input
rlabel metal2 s 179510 171200 179566 172000 6 la_input[13]
port 190 nsew signal input
rlabel metal2 s 180154 171200 180210 172000 6 la_input[14]
port 191 nsew signal input
rlabel metal2 s 180798 171200 180854 172000 6 la_input[15]
port 192 nsew signal input
rlabel metal2 s 181442 171200 181498 172000 6 la_input[16]
port 193 nsew signal input
rlabel metal2 s 182086 171200 182142 172000 6 la_input[17]
port 194 nsew signal input
rlabel metal2 s 182730 171200 182786 172000 6 la_input[18]
port 195 nsew signal input
rlabel metal2 s 183466 171200 183522 172000 6 la_input[19]
port 196 nsew signal input
rlabel metal2 s 171690 171200 171746 172000 6 la_input[1]
port 197 nsew signal input
rlabel metal2 s 184110 171200 184166 172000 6 la_input[20]
port 198 nsew signal input
rlabel metal2 s 184754 171200 184810 172000 6 la_input[21]
port 199 nsew signal input
rlabel metal2 s 185398 171200 185454 172000 6 la_input[22]
port 200 nsew signal input
rlabel metal2 s 186042 171200 186098 172000 6 la_input[23]
port 201 nsew signal input
rlabel metal2 s 186686 171200 186742 172000 6 la_input[24]
port 202 nsew signal input
rlabel metal2 s 187330 171200 187386 172000 6 la_input[25]
port 203 nsew signal input
rlabel metal2 s 187974 171200 188030 172000 6 la_input[26]
port 204 nsew signal input
rlabel metal2 s 188618 171200 188674 172000 6 la_input[27]
port 205 nsew signal input
rlabel metal2 s 189262 171200 189318 172000 6 la_input[28]
port 206 nsew signal input
rlabel metal2 s 189906 171200 189962 172000 6 la_input[29]
port 207 nsew signal input
rlabel metal2 s 172426 171200 172482 172000 6 la_input[2]
port 208 nsew signal input
rlabel metal2 s 190550 171200 190606 172000 6 la_input[30]
port 209 nsew signal input
rlabel metal2 s 191194 171200 191250 172000 6 la_input[31]
port 210 nsew signal input
rlabel metal2 s 191838 171200 191894 172000 6 la_input[32]
port 211 nsew signal input
rlabel metal2 s 192482 171200 192538 172000 6 la_input[33]
port 212 nsew signal input
rlabel metal2 s 193126 171200 193182 172000 6 la_input[34]
port 213 nsew signal input
rlabel metal2 s 193862 171200 193918 172000 6 la_input[35]
port 214 nsew signal input
rlabel metal2 s 194506 171200 194562 172000 6 la_input[36]
port 215 nsew signal input
rlabel metal2 s 195150 171200 195206 172000 6 la_input[37]
port 216 nsew signal input
rlabel metal2 s 195794 171200 195850 172000 6 la_input[38]
port 217 nsew signal input
rlabel metal2 s 196438 171200 196494 172000 6 la_input[39]
port 218 nsew signal input
rlabel metal2 s 173070 171200 173126 172000 6 la_input[3]
port 219 nsew signal input
rlabel metal2 s 197082 171200 197138 172000 6 la_input[40]
port 220 nsew signal input
rlabel metal2 s 197726 171200 197782 172000 6 la_input[41]
port 221 nsew signal input
rlabel metal2 s 198370 171200 198426 172000 6 la_input[42]
port 222 nsew signal input
rlabel metal2 s 199014 171200 199070 172000 6 la_input[43]
port 223 nsew signal input
rlabel metal2 s 199658 171200 199714 172000 6 la_input[44]
port 224 nsew signal input
rlabel metal2 s 200302 171200 200358 172000 6 la_input[45]
port 225 nsew signal input
rlabel metal2 s 200946 171200 201002 172000 6 la_input[46]
port 226 nsew signal input
rlabel metal2 s 201590 171200 201646 172000 6 la_input[47]
port 227 nsew signal input
rlabel metal2 s 202234 171200 202290 172000 6 la_input[48]
port 228 nsew signal input
rlabel metal2 s 202878 171200 202934 172000 6 la_input[49]
port 229 nsew signal input
rlabel metal2 s 173714 171200 173770 172000 6 la_input[4]
port 230 nsew signal input
rlabel metal2 s 203522 171200 203578 172000 6 la_input[50]
port 231 nsew signal input
rlabel metal2 s 204166 171200 204222 172000 6 la_input[51]
port 232 nsew signal input
rlabel metal2 s 204902 171200 204958 172000 6 la_input[52]
port 233 nsew signal input
rlabel metal2 s 205546 171200 205602 172000 6 la_input[53]
port 234 nsew signal input
rlabel metal2 s 206190 171200 206246 172000 6 la_input[54]
port 235 nsew signal input
rlabel metal2 s 206834 171200 206890 172000 6 la_input[55]
port 236 nsew signal input
rlabel metal2 s 207478 171200 207534 172000 6 la_input[56]
port 237 nsew signal input
rlabel metal2 s 208122 171200 208178 172000 6 la_input[57]
port 238 nsew signal input
rlabel metal2 s 208766 171200 208822 172000 6 la_input[58]
port 239 nsew signal input
rlabel metal2 s 209410 171200 209466 172000 6 la_input[59]
port 240 nsew signal input
rlabel metal2 s 174358 171200 174414 172000 6 la_input[5]
port 241 nsew signal input
rlabel metal2 s 210054 171200 210110 172000 6 la_input[60]
port 242 nsew signal input
rlabel metal2 s 210698 171200 210754 172000 6 la_input[61]
port 243 nsew signal input
rlabel metal2 s 211342 171200 211398 172000 6 la_input[62]
port 244 nsew signal input
rlabel metal2 s 211986 171200 212042 172000 6 la_input[63]
port 245 nsew signal input
rlabel metal2 s 212630 171200 212686 172000 6 la_input[64]
port 246 nsew signal input
rlabel metal2 s 213274 171200 213330 172000 6 la_input[65]
port 247 nsew signal input
rlabel metal2 s 213918 171200 213974 172000 6 la_input[66]
port 248 nsew signal input
rlabel metal2 s 214562 171200 214618 172000 6 la_input[67]
port 249 nsew signal input
rlabel metal2 s 215298 171200 215354 172000 6 la_input[68]
port 250 nsew signal input
rlabel metal2 s 215942 171200 215998 172000 6 la_input[69]
port 251 nsew signal input
rlabel metal2 s 175002 171200 175058 172000 6 la_input[6]
port 252 nsew signal input
rlabel metal2 s 216586 171200 216642 172000 6 la_input[70]
port 253 nsew signal input
rlabel metal2 s 217230 171200 217286 172000 6 la_input[71]
port 254 nsew signal input
rlabel metal2 s 217874 171200 217930 172000 6 la_input[72]
port 255 nsew signal input
rlabel metal2 s 218518 171200 218574 172000 6 la_input[73]
port 256 nsew signal input
rlabel metal2 s 219162 171200 219218 172000 6 la_input[74]
port 257 nsew signal input
rlabel metal2 s 219806 171200 219862 172000 6 la_input[75]
port 258 nsew signal input
rlabel metal2 s 220450 171200 220506 172000 6 la_input[76]
port 259 nsew signal input
rlabel metal2 s 221094 171200 221150 172000 6 la_input[77]
port 260 nsew signal input
rlabel metal2 s 221738 171200 221794 172000 6 la_input[78]
port 261 nsew signal input
rlabel metal2 s 222382 171200 222438 172000 6 la_input[79]
port 262 nsew signal input
rlabel metal2 s 175646 171200 175702 172000 6 la_input[7]
port 263 nsew signal input
rlabel metal2 s 223026 171200 223082 172000 6 la_input[80]
port 264 nsew signal input
rlabel metal2 s 223670 171200 223726 172000 6 la_input[81]
port 265 nsew signal input
rlabel metal2 s 224314 171200 224370 172000 6 la_input[82]
port 266 nsew signal input
rlabel metal2 s 224958 171200 225014 172000 6 la_input[83]
port 267 nsew signal input
rlabel metal2 s 225602 171200 225658 172000 6 la_input[84]
port 268 nsew signal input
rlabel metal2 s 226338 171200 226394 172000 6 la_input[85]
port 269 nsew signal input
rlabel metal2 s 226982 171200 227038 172000 6 la_input[86]
port 270 nsew signal input
rlabel metal2 s 227626 171200 227682 172000 6 la_input[87]
port 271 nsew signal input
rlabel metal2 s 228270 171200 228326 172000 6 la_input[88]
port 272 nsew signal input
rlabel metal2 s 228914 171200 228970 172000 6 la_input[89]
port 273 nsew signal input
rlabel metal2 s 176290 171200 176346 172000 6 la_input[8]
port 274 nsew signal input
rlabel metal2 s 229558 171200 229614 172000 6 la_input[90]
port 275 nsew signal input
rlabel metal2 s 230202 171200 230258 172000 6 la_input[91]
port 276 nsew signal input
rlabel metal2 s 230846 171200 230902 172000 6 la_input[92]
port 277 nsew signal input
rlabel metal2 s 231490 171200 231546 172000 6 la_input[93]
port 278 nsew signal input
rlabel metal2 s 232134 171200 232190 172000 6 la_input[94]
port 279 nsew signal input
rlabel metal2 s 232778 171200 232834 172000 6 la_input[95]
port 280 nsew signal input
rlabel metal2 s 233422 171200 233478 172000 6 la_input[96]
port 281 nsew signal input
rlabel metal2 s 234066 171200 234122 172000 6 la_input[97]
port 282 nsew signal input
rlabel metal2 s 234710 171200 234766 172000 6 la_input[98]
port 283 nsew signal input
rlabel metal2 s 235354 171200 235410 172000 6 la_input[99]
port 284 nsew signal input
rlabel metal2 s 176934 171200 176990 172000 6 la_input[9]
port 285 nsew signal input
rlabel metal2 s 254214 171200 254270 172000 6 la_oenb[0]
port 286 nsew signal output
rlabel metal2 s 319166 171200 319222 172000 6 la_oenb[100]
port 287 nsew signal output
rlabel metal2 s 319810 171200 319866 172000 6 la_oenb[101]
port 288 nsew signal output
rlabel metal2 s 320454 171200 320510 172000 6 la_oenb[102]
port 289 nsew signal output
rlabel metal2 s 321098 171200 321154 172000 6 la_oenb[103]
port 290 nsew signal output
rlabel metal2 s 321742 171200 321798 172000 6 la_oenb[104]
port 291 nsew signal output
rlabel metal2 s 322386 171200 322442 172000 6 la_oenb[105]
port 292 nsew signal output
rlabel metal2 s 323122 171200 323178 172000 6 la_oenb[106]
port 293 nsew signal output
rlabel metal2 s 323766 171200 323822 172000 6 la_oenb[107]
port 294 nsew signal output
rlabel metal2 s 324410 171200 324466 172000 6 la_oenb[108]
port 295 nsew signal output
rlabel metal2 s 325054 171200 325110 172000 6 la_oenb[109]
port 296 nsew signal output
rlabel metal2 s 260746 171200 260802 172000 6 la_oenb[10]
port 297 nsew signal output
rlabel metal2 s 325698 171200 325754 172000 6 la_oenb[110]
port 298 nsew signal output
rlabel metal2 s 326342 171200 326398 172000 6 la_oenb[111]
port 299 nsew signal output
rlabel metal2 s 326986 171200 327042 172000 6 la_oenb[112]
port 300 nsew signal output
rlabel metal2 s 327630 171200 327686 172000 6 la_oenb[113]
port 301 nsew signal output
rlabel metal2 s 328274 171200 328330 172000 6 la_oenb[114]
port 302 nsew signal output
rlabel metal2 s 328918 171200 328974 172000 6 la_oenb[115]
port 303 nsew signal output
rlabel metal2 s 329562 171200 329618 172000 6 la_oenb[116]
port 304 nsew signal output
rlabel metal2 s 330206 171200 330262 172000 6 la_oenb[117]
port 305 nsew signal output
rlabel metal2 s 330850 171200 330906 172000 6 la_oenb[118]
port 306 nsew signal output
rlabel metal2 s 331494 171200 331550 172000 6 la_oenb[119]
port 307 nsew signal output
rlabel metal2 s 261390 171200 261446 172000 6 la_oenb[11]
port 308 nsew signal output
rlabel metal2 s 332138 171200 332194 172000 6 la_oenb[120]
port 309 nsew signal output
rlabel metal2 s 332782 171200 332838 172000 6 la_oenb[121]
port 310 nsew signal output
rlabel metal2 s 333426 171200 333482 172000 6 la_oenb[122]
port 311 nsew signal output
rlabel metal2 s 334162 171200 334218 172000 6 la_oenb[123]
port 312 nsew signal output
rlabel metal2 s 334806 171200 334862 172000 6 la_oenb[124]
port 313 nsew signal output
rlabel metal2 s 335450 171200 335506 172000 6 la_oenb[125]
port 314 nsew signal output
rlabel metal2 s 336094 171200 336150 172000 6 la_oenb[126]
port 315 nsew signal output
rlabel metal2 s 336738 171200 336794 172000 6 la_oenb[127]
port 316 nsew signal output
rlabel metal2 s 262034 171200 262090 172000 6 la_oenb[12]
port 317 nsew signal output
rlabel metal2 s 262678 171200 262734 172000 6 la_oenb[13]
port 318 nsew signal output
rlabel metal2 s 263322 171200 263378 172000 6 la_oenb[14]
port 319 nsew signal output
rlabel metal2 s 263966 171200 264022 172000 6 la_oenb[15]
port 320 nsew signal output
rlabel metal2 s 264610 171200 264666 172000 6 la_oenb[16]
port 321 nsew signal output
rlabel metal2 s 265254 171200 265310 172000 6 la_oenb[17]
port 322 nsew signal output
rlabel metal2 s 265898 171200 265954 172000 6 la_oenb[18]
port 323 nsew signal output
rlabel metal2 s 266542 171200 266598 172000 6 la_oenb[19]
port 324 nsew signal output
rlabel metal2 s 254858 171200 254914 172000 6 la_oenb[1]
port 325 nsew signal output
rlabel metal2 s 267186 171200 267242 172000 6 la_oenb[20]
port 326 nsew signal output
rlabel metal2 s 267830 171200 267886 172000 6 la_oenb[21]
port 327 nsew signal output
rlabel metal2 s 268474 171200 268530 172000 6 la_oenb[22]
port 328 nsew signal output
rlabel metal2 s 269210 171200 269266 172000 6 la_oenb[23]
port 329 nsew signal output
rlabel metal2 s 269854 171200 269910 172000 6 la_oenb[24]
port 330 nsew signal output
rlabel metal2 s 270498 171200 270554 172000 6 la_oenb[25]
port 331 nsew signal output
rlabel metal2 s 271142 171200 271198 172000 6 la_oenb[26]
port 332 nsew signal output
rlabel metal2 s 271786 171200 271842 172000 6 la_oenb[27]
port 333 nsew signal output
rlabel metal2 s 272430 171200 272486 172000 6 la_oenb[28]
port 334 nsew signal output
rlabel metal2 s 273074 171200 273130 172000 6 la_oenb[29]
port 335 nsew signal output
rlabel metal2 s 255502 171200 255558 172000 6 la_oenb[2]
port 336 nsew signal output
rlabel metal2 s 273718 171200 273774 172000 6 la_oenb[30]
port 337 nsew signal output
rlabel metal2 s 274362 171200 274418 172000 6 la_oenb[31]
port 338 nsew signal output
rlabel metal2 s 275006 171200 275062 172000 6 la_oenb[32]
port 339 nsew signal output
rlabel metal2 s 275650 171200 275706 172000 6 la_oenb[33]
port 340 nsew signal output
rlabel metal2 s 276294 171200 276350 172000 6 la_oenb[34]
port 341 nsew signal output
rlabel metal2 s 276938 171200 276994 172000 6 la_oenb[35]
port 342 nsew signal output
rlabel metal2 s 277582 171200 277638 172000 6 la_oenb[36]
port 343 nsew signal output
rlabel metal2 s 278226 171200 278282 172000 6 la_oenb[37]
port 344 nsew signal output
rlabel metal2 s 278870 171200 278926 172000 6 la_oenb[38]
port 345 nsew signal output
rlabel metal2 s 279514 171200 279570 172000 6 la_oenb[39]
port 346 nsew signal output
rlabel metal2 s 256146 171200 256202 172000 6 la_oenb[3]
port 347 nsew signal output
rlabel metal2 s 280250 171200 280306 172000 6 la_oenb[40]
port 348 nsew signal output
rlabel metal2 s 280894 171200 280950 172000 6 la_oenb[41]
port 349 nsew signal output
rlabel metal2 s 281538 171200 281594 172000 6 la_oenb[42]
port 350 nsew signal output
rlabel metal2 s 282182 171200 282238 172000 6 la_oenb[43]
port 351 nsew signal output
rlabel metal2 s 282826 171200 282882 172000 6 la_oenb[44]
port 352 nsew signal output
rlabel metal2 s 283470 171200 283526 172000 6 la_oenb[45]
port 353 nsew signal output
rlabel metal2 s 284114 171200 284170 172000 6 la_oenb[46]
port 354 nsew signal output
rlabel metal2 s 284758 171200 284814 172000 6 la_oenb[47]
port 355 nsew signal output
rlabel metal2 s 285402 171200 285458 172000 6 la_oenb[48]
port 356 nsew signal output
rlabel metal2 s 286046 171200 286102 172000 6 la_oenb[49]
port 357 nsew signal output
rlabel metal2 s 256790 171200 256846 172000 6 la_oenb[4]
port 358 nsew signal output
rlabel metal2 s 286690 171200 286746 172000 6 la_oenb[50]
port 359 nsew signal output
rlabel metal2 s 287334 171200 287390 172000 6 la_oenb[51]
port 360 nsew signal output
rlabel metal2 s 287978 171200 288034 172000 6 la_oenb[52]
port 361 nsew signal output
rlabel metal2 s 288622 171200 288678 172000 6 la_oenb[53]
port 362 nsew signal output
rlabel metal2 s 289266 171200 289322 172000 6 la_oenb[54]
port 363 nsew signal output
rlabel metal2 s 289910 171200 289966 172000 6 la_oenb[55]
port 364 nsew signal output
rlabel metal2 s 290646 171200 290702 172000 6 la_oenb[56]
port 365 nsew signal output
rlabel metal2 s 291290 171200 291346 172000 6 la_oenb[57]
port 366 nsew signal output
rlabel metal2 s 291934 171200 291990 172000 6 la_oenb[58]
port 367 nsew signal output
rlabel metal2 s 292578 171200 292634 172000 6 la_oenb[59]
port 368 nsew signal output
rlabel metal2 s 257434 171200 257490 172000 6 la_oenb[5]
port 369 nsew signal output
rlabel metal2 s 293222 171200 293278 172000 6 la_oenb[60]
port 370 nsew signal output
rlabel metal2 s 293866 171200 293922 172000 6 la_oenb[61]
port 371 nsew signal output
rlabel metal2 s 294510 171200 294566 172000 6 la_oenb[62]
port 372 nsew signal output
rlabel metal2 s 295154 171200 295210 172000 6 la_oenb[63]
port 373 nsew signal output
rlabel metal2 s 295798 171200 295854 172000 6 la_oenb[64]
port 374 nsew signal output
rlabel metal2 s 296442 171200 296498 172000 6 la_oenb[65]
port 375 nsew signal output
rlabel metal2 s 297086 171200 297142 172000 6 la_oenb[66]
port 376 nsew signal output
rlabel metal2 s 297730 171200 297786 172000 6 la_oenb[67]
port 377 nsew signal output
rlabel metal2 s 298374 171200 298430 172000 6 la_oenb[68]
port 378 nsew signal output
rlabel metal2 s 299018 171200 299074 172000 6 la_oenb[69]
port 379 nsew signal output
rlabel metal2 s 258078 171200 258134 172000 6 la_oenb[6]
port 380 nsew signal output
rlabel metal2 s 299662 171200 299718 172000 6 la_oenb[70]
port 381 nsew signal output
rlabel metal2 s 300306 171200 300362 172000 6 la_oenb[71]
port 382 nsew signal output
rlabel metal2 s 300950 171200 301006 172000 6 la_oenb[72]
port 383 nsew signal output
rlabel metal2 s 301686 171200 301742 172000 6 la_oenb[73]
port 384 nsew signal output
rlabel metal2 s 302330 171200 302386 172000 6 la_oenb[74]
port 385 nsew signal output
rlabel metal2 s 302974 171200 303030 172000 6 la_oenb[75]
port 386 nsew signal output
rlabel metal2 s 303618 171200 303674 172000 6 la_oenb[76]
port 387 nsew signal output
rlabel metal2 s 304262 171200 304318 172000 6 la_oenb[77]
port 388 nsew signal output
rlabel metal2 s 304906 171200 304962 172000 6 la_oenb[78]
port 389 nsew signal output
rlabel metal2 s 305550 171200 305606 172000 6 la_oenb[79]
port 390 nsew signal output
rlabel metal2 s 258814 171200 258870 172000 6 la_oenb[7]
port 391 nsew signal output
rlabel metal2 s 306194 171200 306250 172000 6 la_oenb[80]
port 392 nsew signal output
rlabel metal2 s 306838 171200 306894 172000 6 la_oenb[81]
port 393 nsew signal output
rlabel metal2 s 307482 171200 307538 172000 6 la_oenb[82]
port 394 nsew signal output
rlabel metal2 s 308126 171200 308182 172000 6 la_oenb[83]
port 395 nsew signal output
rlabel metal2 s 308770 171200 308826 172000 6 la_oenb[84]
port 396 nsew signal output
rlabel metal2 s 309414 171200 309470 172000 6 la_oenb[85]
port 397 nsew signal output
rlabel metal2 s 310058 171200 310114 172000 6 la_oenb[86]
port 398 nsew signal output
rlabel metal2 s 310702 171200 310758 172000 6 la_oenb[87]
port 399 nsew signal output
rlabel metal2 s 311346 171200 311402 172000 6 la_oenb[88]
port 400 nsew signal output
rlabel metal2 s 312082 171200 312138 172000 6 la_oenb[89]
port 401 nsew signal output
rlabel metal2 s 259458 171200 259514 172000 6 la_oenb[8]
port 402 nsew signal output
rlabel metal2 s 312726 171200 312782 172000 6 la_oenb[90]
port 403 nsew signal output
rlabel metal2 s 313370 171200 313426 172000 6 la_oenb[91]
port 404 nsew signal output
rlabel metal2 s 314014 171200 314070 172000 6 la_oenb[92]
port 405 nsew signal output
rlabel metal2 s 314658 171200 314714 172000 6 la_oenb[93]
port 406 nsew signal output
rlabel metal2 s 315302 171200 315358 172000 6 la_oenb[94]
port 407 nsew signal output
rlabel metal2 s 315946 171200 316002 172000 6 la_oenb[95]
port 408 nsew signal output
rlabel metal2 s 316590 171200 316646 172000 6 la_oenb[96]
port 409 nsew signal output
rlabel metal2 s 317234 171200 317290 172000 6 la_oenb[97]
port 410 nsew signal output
rlabel metal2 s 317878 171200 317934 172000 6 la_oenb[98]
port 411 nsew signal output
rlabel metal2 s 318522 171200 318578 172000 6 la_oenb[99]
port 412 nsew signal output
rlabel metal2 s 260102 171200 260158 172000 6 la_oenb[9]
port 413 nsew signal output
rlabel metal2 s 337382 171200 337438 172000 6 la_output[0]
port 414 nsew signal output
rlabel metal2 s 402334 171200 402390 172000 6 la_output[100]
port 415 nsew signal output
rlabel metal2 s 402978 171200 403034 172000 6 la_output[101]
port 416 nsew signal output
rlabel metal2 s 403622 171200 403678 172000 6 la_output[102]
port 417 nsew signal output
rlabel metal2 s 404266 171200 404322 172000 6 la_output[103]
port 418 nsew signal output
rlabel metal2 s 404910 171200 404966 172000 6 la_output[104]
port 419 nsew signal output
rlabel metal2 s 405554 171200 405610 172000 6 la_output[105]
port 420 nsew signal output
rlabel metal2 s 406198 171200 406254 172000 6 la_output[106]
port 421 nsew signal output
rlabel metal2 s 406842 171200 406898 172000 6 la_output[107]
port 422 nsew signal output
rlabel metal2 s 407486 171200 407542 172000 6 la_output[108]
port 423 nsew signal output
rlabel metal2 s 408130 171200 408186 172000 6 la_output[109]
port 424 nsew signal output
rlabel metal2 s 343822 171200 343878 172000 6 la_output[10]
port 425 nsew signal output
rlabel metal2 s 408866 171200 408922 172000 6 la_output[110]
port 426 nsew signal output
rlabel metal2 s 409510 171200 409566 172000 6 la_output[111]
port 427 nsew signal output
rlabel metal2 s 410154 171200 410210 172000 6 la_output[112]
port 428 nsew signal output
rlabel metal2 s 410798 171200 410854 172000 6 la_output[113]
port 429 nsew signal output
rlabel metal2 s 411442 171200 411498 172000 6 la_output[114]
port 430 nsew signal output
rlabel metal2 s 412086 171200 412142 172000 6 la_output[115]
port 431 nsew signal output
rlabel metal2 s 412730 171200 412786 172000 6 la_output[116]
port 432 nsew signal output
rlabel metal2 s 413374 171200 413430 172000 6 la_output[117]
port 433 nsew signal output
rlabel metal2 s 414018 171200 414074 172000 6 la_output[118]
port 434 nsew signal output
rlabel metal2 s 414662 171200 414718 172000 6 la_output[119]
port 435 nsew signal output
rlabel metal2 s 344558 171200 344614 172000 6 la_output[11]
port 436 nsew signal output
rlabel metal2 s 415306 171200 415362 172000 6 la_output[120]
port 437 nsew signal output
rlabel metal2 s 415950 171200 416006 172000 6 la_output[121]
port 438 nsew signal output
rlabel metal2 s 416594 171200 416650 172000 6 la_output[122]
port 439 nsew signal output
rlabel metal2 s 417238 171200 417294 172000 6 la_output[123]
port 440 nsew signal output
rlabel metal2 s 417882 171200 417938 172000 6 la_output[124]
port 441 nsew signal output
rlabel metal2 s 418526 171200 418582 172000 6 la_output[125]
port 442 nsew signal output
rlabel metal2 s 419170 171200 419226 172000 6 la_output[126]
port 443 nsew signal output
rlabel metal2 s 419906 171200 419962 172000 6 la_output[127]
port 444 nsew signal output
rlabel metal2 s 345202 171200 345258 172000 6 la_output[12]
port 445 nsew signal output
rlabel metal2 s 345846 171200 345902 172000 6 la_output[13]
port 446 nsew signal output
rlabel metal2 s 346490 171200 346546 172000 6 la_output[14]
port 447 nsew signal output
rlabel metal2 s 347134 171200 347190 172000 6 la_output[15]
port 448 nsew signal output
rlabel metal2 s 347778 171200 347834 172000 6 la_output[16]
port 449 nsew signal output
rlabel metal2 s 348422 171200 348478 172000 6 la_output[17]
port 450 nsew signal output
rlabel metal2 s 349066 171200 349122 172000 6 la_output[18]
port 451 nsew signal output
rlabel metal2 s 349710 171200 349766 172000 6 la_output[19]
port 452 nsew signal output
rlabel metal2 s 338026 171200 338082 172000 6 la_output[1]
port 453 nsew signal output
rlabel metal2 s 350354 171200 350410 172000 6 la_output[20]
port 454 nsew signal output
rlabel metal2 s 350998 171200 351054 172000 6 la_output[21]
port 455 nsew signal output
rlabel metal2 s 351642 171200 351698 172000 6 la_output[22]
port 456 nsew signal output
rlabel metal2 s 352286 171200 352342 172000 6 la_output[23]
port 457 nsew signal output
rlabel metal2 s 352930 171200 352986 172000 6 la_output[24]
port 458 nsew signal output
rlabel metal2 s 353574 171200 353630 172000 6 la_output[25]
port 459 nsew signal output
rlabel metal2 s 354218 171200 354274 172000 6 la_output[26]
port 460 nsew signal output
rlabel metal2 s 354862 171200 354918 172000 6 la_output[27]
port 461 nsew signal output
rlabel metal2 s 355598 171200 355654 172000 6 la_output[28]
port 462 nsew signal output
rlabel metal2 s 356242 171200 356298 172000 6 la_output[29]
port 463 nsew signal output
rlabel metal2 s 338670 171200 338726 172000 6 la_output[2]
port 464 nsew signal output
rlabel metal2 s 356886 171200 356942 172000 6 la_output[30]
port 465 nsew signal output
rlabel metal2 s 357530 171200 357586 172000 6 la_output[31]
port 466 nsew signal output
rlabel metal2 s 358174 171200 358230 172000 6 la_output[32]
port 467 nsew signal output
rlabel metal2 s 358818 171200 358874 172000 6 la_output[33]
port 468 nsew signal output
rlabel metal2 s 359462 171200 359518 172000 6 la_output[34]
port 469 nsew signal output
rlabel metal2 s 360106 171200 360162 172000 6 la_output[35]
port 470 nsew signal output
rlabel metal2 s 360750 171200 360806 172000 6 la_output[36]
port 471 nsew signal output
rlabel metal2 s 361394 171200 361450 172000 6 la_output[37]
port 472 nsew signal output
rlabel metal2 s 362038 171200 362094 172000 6 la_output[38]
port 473 nsew signal output
rlabel metal2 s 362682 171200 362738 172000 6 la_output[39]
port 474 nsew signal output
rlabel metal2 s 339314 171200 339370 172000 6 la_output[3]
port 475 nsew signal output
rlabel metal2 s 363326 171200 363382 172000 6 la_output[40]
port 476 nsew signal output
rlabel metal2 s 363970 171200 364026 172000 6 la_output[41]
port 477 nsew signal output
rlabel metal2 s 364614 171200 364670 172000 6 la_output[42]
port 478 nsew signal output
rlabel metal2 s 365258 171200 365314 172000 6 la_output[43]
port 479 nsew signal output
rlabel metal2 s 365994 171200 366050 172000 6 la_output[44]
port 480 nsew signal output
rlabel metal2 s 366638 171200 366694 172000 6 la_output[45]
port 481 nsew signal output
rlabel metal2 s 367282 171200 367338 172000 6 la_output[46]
port 482 nsew signal output
rlabel metal2 s 367926 171200 367982 172000 6 la_output[47]
port 483 nsew signal output
rlabel metal2 s 368570 171200 368626 172000 6 la_output[48]
port 484 nsew signal output
rlabel metal2 s 369214 171200 369270 172000 6 la_output[49]
port 485 nsew signal output
rlabel metal2 s 339958 171200 340014 172000 6 la_output[4]
port 486 nsew signal output
rlabel metal2 s 369858 171200 369914 172000 6 la_output[50]
port 487 nsew signal output
rlabel metal2 s 370502 171200 370558 172000 6 la_output[51]
port 488 nsew signal output
rlabel metal2 s 371146 171200 371202 172000 6 la_output[52]
port 489 nsew signal output
rlabel metal2 s 371790 171200 371846 172000 6 la_output[53]
port 490 nsew signal output
rlabel metal2 s 372434 171200 372490 172000 6 la_output[54]
port 491 nsew signal output
rlabel metal2 s 373078 171200 373134 172000 6 la_output[55]
port 492 nsew signal output
rlabel metal2 s 373722 171200 373778 172000 6 la_output[56]
port 493 nsew signal output
rlabel metal2 s 374366 171200 374422 172000 6 la_output[57]
port 494 nsew signal output
rlabel metal2 s 375010 171200 375066 172000 6 la_output[58]
port 495 nsew signal output
rlabel metal2 s 375654 171200 375710 172000 6 la_output[59]
port 496 nsew signal output
rlabel metal2 s 340602 171200 340658 172000 6 la_output[5]
port 497 nsew signal output
rlabel metal2 s 376298 171200 376354 172000 6 la_output[60]
port 498 nsew signal output
rlabel metal2 s 377034 171200 377090 172000 6 la_output[61]
port 499 nsew signal output
rlabel metal2 s 377678 171200 377734 172000 6 la_output[62]
port 500 nsew signal output
rlabel metal2 s 378322 171200 378378 172000 6 la_output[63]
port 501 nsew signal output
rlabel metal2 s 378966 171200 379022 172000 6 la_output[64]
port 502 nsew signal output
rlabel metal2 s 379610 171200 379666 172000 6 la_output[65]
port 503 nsew signal output
rlabel metal2 s 380254 171200 380310 172000 6 la_output[66]
port 504 nsew signal output
rlabel metal2 s 380898 171200 380954 172000 6 la_output[67]
port 505 nsew signal output
rlabel metal2 s 381542 171200 381598 172000 6 la_output[68]
port 506 nsew signal output
rlabel metal2 s 382186 171200 382242 172000 6 la_output[69]
port 507 nsew signal output
rlabel metal2 s 341246 171200 341302 172000 6 la_output[6]
port 508 nsew signal output
rlabel metal2 s 382830 171200 382886 172000 6 la_output[70]
port 509 nsew signal output
rlabel metal2 s 383474 171200 383530 172000 6 la_output[71]
port 510 nsew signal output
rlabel metal2 s 384118 171200 384174 172000 6 la_output[72]
port 511 nsew signal output
rlabel metal2 s 384762 171200 384818 172000 6 la_output[73]
port 512 nsew signal output
rlabel metal2 s 385406 171200 385462 172000 6 la_output[74]
port 513 nsew signal output
rlabel metal2 s 386050 171200 386106 172000 6 la_output[75]
port 514 nsew signal output
rlabel metal2 s 386694 171200 386750 172000 6 la_output[76]
port 515 nsew signal output
rlabel metal2 s 387430 171200 387486 172000 6 la_output[77]
port 516 nsew signal output
rlabel metal2 s 388074 171200 388130 172000 6 la_output[78]
port 517 nsew signal output
rlabel metal2 s 388718 171200 388774 172000 6 la_output[79]
port 518 nsew signal output
rlabel metal2 s 341890 171200 341946 172000 6 la_output[7]
port 519 nsew signal output
rlabel metal2 s 389362 171200 389418 172000 6 la_output[80]
port 520 nsew signal output
rlabel metal2 s 390006 171200 390062 172000 6 la_output[81]
port 521 nsew signal output
rlabel metal2 s 390650 171200 390706 172000 6 la_output[82]
port 522 nsew signal output
rlabel metal2 s 391294 171200 391350 172000 6 la_output[83]
port 523 nsew signal output
rlabel metal2 s 391938 171200 391994 172000 6 la_output[84]
port 524 nsew signal output
rlabel metal2 s 392582 171200 392638 172000 6 la_output[85]
port 525 nsew signal output
rlabel metal2 s 393226 171200 393282 172000 6 la_output[86]
port 526 nsew signal output
rlabel metal2 s 393870 171200 393926 172000 6 la_output[87]
port 527 nsew signal output
rlabel metal2 s 394514 171200 394570 172000 6 la_output[88]
port 528 nsew signal output
rlabel metal2 s 395158 171200 395214 172000 6 la_output[89]
port 529 nsew signal output
rlabel metal2 s 342534 171200 342590 172000 6 la_output[8]
port 530 nsew signal output
rlabel metal2 s 395802 171200 395858 172000 6 la_output[90]
port 531 nsew signal output
rlabel metal2 s 396446 171200 396502 172000 6 la_output[91]
port 532 nsew signal output
rlabel metal2 s 397090 171200 397146 172000 6 la_output[92]
port 533 nsew signal output
rlabel metal2 s 397734 171200 397790 172000 6 la_output[93]
port 534 nsew signal output
rlabel metal2 s 398470 171200 398526 172000 6 la_output[94]
port 535 nsew signal output
rlabel metal2 s 399114 171200 399170 172000 6 la_output[95]
port 536 nsew signal output
rlabel metal2 s 399758 171200 399814 172000 6 la_output[96]
port 537 nsew signal output
rlabel metal2 s 400402 171200 400458 172000 6 la_output[97]
port 538 nsew signal output
rlabel metal2 s 401046 171200 401102 172000 6 la_output[98]
port 539 nsew signal output
rlabel metal2 s 401690 171200 401746 172000 6 la_output[99]
port 540 nsew signal output
rlabel metal2 s 343178 171200 343234 172000 6 la_output[9]
port 541 nsew signal output
rlabel metal3 s 429200 960 430000 1080 6 mask_rev[0]
port 542 nsew signal input
rlabel metal3 s 429200 20272 430000 20392 6 mask_rev[10]
port 543 nsew signal input
rlabel metal3 s 429200 22176 430000 22296 6 mask_rev[11]
port 544 nsew signal input
rlabel metal3 s 429200 24080 430000 24200 6 mask_rev[12]
port 545 nsew signal input
rlabel metal3 s 429200 25984 430000 26104 6 mask_rev[13]
port 546 nsew signal input
rlabel metal3 s 429200 27888 430000 28008 6 mask_rev[14]
port 547 nsew signal input
rlabel metal3 s 429200 29928 430000 30048 6 mask_rev[15]
port 548 nsew signal input
rlabel metal3 s 429200 31832 430000 31952 6 mask_rev[16]
port 549 nsew signal input
rlabel metal3 s 429200 33736 430000 33856 6 mask_rev[17]
port 550 nsew signal input
rlabel metal3 s 429200 35640 430000 35760 6 mask_rev[18]
port 551 nsew signal input
rlabel metal3 s 429200 37680 430000 37800 6 mask_rev[19]
port 552 nsew signal input
rlabel metal3 s 429200 2864 430000 2984 6 mask_rev[1]
port 553 nsew signal input
rlabel metal3 s 429200 39584 430000 39704 6 mask_rev[20]
port 554 nsew signal input
rlabel metal3 s 429200 41488 430000 41608 6 mask_rev[21]
port 555 nsew signal input
rlabel metal3 s 429200 43392 430000 43512 6 mask_rev[22]
port 556 nsew signal input
rlabel metal3 s 429200 45296 430000 45416 6 mask_rev[23]
port 557 nsew signal input
rlabel metal3 s 429200 47336 430000 47456 6 mask_rev[24]
port 558 nsew signal input
rlabel metal3 s 429200 49240 430000 49360 6 mask_rev[25]
port 559 nsew signal input
rlabel metal3 s 429200 51144 430000 51264 6 mask_rev[26]
port 560 nsew signal input
rlabel metal3 s 429200 53048 430000 53168 6 mask_rev[27]
port 561 nsew signal input
rlabel metal3 s 429200 54952 430000 55072 6 mask_rev[28]
port 562 nsew signal input
rlabel metal3 s 429200 56992 430000 57112 6 mask_rev[29]
port 563 nsew signal input
rlabel metal3 s 429200 4768 430000 4888 6 mask_rev[2]
port 564 nsew signal input
rlabel metal3 s 429200 58896 430000 59016 6 mask_rev[30]
port 565 nsew signal input
rlabel metal3 s 429200 60800 430000 60920 6 mask_rev[31]
port 566 nsew signal input
rlabel metal3 s 429200 6672 430000 6792 6 mask_rev[3]
port 567 nsew signal input
rlabel metal3 s 429200 8576 430000 8696 6 mask_rev[4]
port 568 nsew signal input
rlabel metal3 s 429200 10616 430000 10736 6 mask_rev[5]
port 569 nsew signal input
rlabel metal3 s 429200 12520 430000 12640 6 mask_rev[6]
port 570 nsew signal input
rlabel metal3 s 429200 14424 430000 14544 6 mask_rev[7]
port 571 nsew signal input
rlabel metal3 s 429200 16328 430000 16448 6 mask_rev[8]
port 572 nsew signal input
rlabel metal3 s 429200 18232 430000 18352 6 mask_rev[9]
port 573 nsew signal input
rlabel metal3 s 0 416 800 536 6 mgmt_addr[0]
port 574 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 mgmt_addr[1]
port 575 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 mgmt_addr[2]
port 576 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 mgmt_addr[3]
port 577 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 mgmt_addr[4]
port 578 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 mgmt_addr[5]
port 579 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 mgmt_addr[6]
port 580 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 mgmt_addr[7]
port 581 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 mgmt_addr_ro[0]
port 582 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 mgmt_addr_ro[1]
port 583 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 mgmt_addr_ro[2]
port 584 nsew signal output
rlabel metal3 s 0 12112 800 12232 6 mgmt_addr_ro[3]
port 585 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 mgmt_addr_ro[4]
port 586 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 mgmt_addr_ro[5]
port 587 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 mgmt_addr_ro[6]
port 588 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 mgmt_addr_ro[7]
port 589 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 mgmt_ena[0]
port 590 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 mgmt_ena[1]
port 591 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 mgmt_ena_ro
port 592 nsew signal output
rlabel metal3 s 429200 76304 430000 76424 6 mgmt_in_data[0]
port 593 nsew signal input
rlabel metal3 s 429200 114928 430000 115048 6 mgmt_in_data[10]
port 594 nsew signal input
rlabel metal3 s 429200 118872 430000 118992 6 mgmt_in_data[11]
port 595 nsew signal input
rlabel metal3 s 429200 122680 430000 122800 6 mgmt_in_data[12]
port 596 nsew signal input
rlabel metal3 s 429200 126488 430000 126608 6 mgmt_in_data[13]
port 597 nsew signal input
rlabel metal3 s 429200 130432 430000 130552 6 mgmt_in_data[14]
port 598 nsew signal input
rlabel metal3 s 429200 134240 430000 134360 6 mgmt_in_data[15]
port 599 nsew signal input
rlabel metal3 s 429200 138184 430000 138304 6 mgmt_in_data[16]
port 600 nsew signal input
rlabel metal3 s 429200 141992 430000 142112 6 mgmt_in_data[17]
port 601 nsew signal input
rlabel metal3 s 429200 145936 430000 146056 6 mgmt_in_data[18]
port 602 nsew signal input
rlabel metal3 s 429200 149744 430000 149864 6 mgmt_in_data[19]
port 603 nsew signal input
rlabel metal3 s 429200 80112 430000 80232 6 mgmt_in_data[1]
port 604 nsew signal input
rlabel metal3 s 429200 153552 430000 153672 6 mgmt_in_data[20]
port 605 nsew signal input
rlabel metal3 s 429200 157496 430000 157616 6 mgmt_in_data[21]
port 606 nsew signal input
rlabel metal3 s 429200 161304 430000 161424 6 mgmt_in_data[22]
port 607 nsew signal input
rlabel metal3 s 429200 165248 430000 165368 6 mgmt_in_data[23]
port 608 nsew signal input
rlabel metal2 s 19062 171200 19118 172000 6 mgmt_in_data[24]
port 609 nsew signal input
rlabel metal2 s 17774 171200 17830 172000 6 mgmt_in_data[25]
port 610 nsew signal input
rlabel metal2 s 16486 171200 16542 172000 6 mgmt_in_data[26]
port 611 nsew signal input
rlabel metal2 s 15198 171200 15254 172000 6 mgmt_in_data[27]
port 612 nsew signal input
rlabel metal2 s 13910 171200 13966 172000 6 mgmt_in_data[28]
port 613 nsew signal input
rlabel metal2 s 12622 171200 12678 172000 6 mgmt_in_data[29]
port 614 nsew signal input
rlabel metal3 s 429200 84056 430000 84176 6 mgmt_in_data[2]
port 615 nsew signal input
rlabel metal2 s 11334 171200 11390 172000 6 mgmt_in_data[30]
port 616 nsew signal input
rlabel metal2 s 9954 171200 10010 172000 6 mgmt_in_data[31]
port 617 nsew signal input
rlabel metal2 s 8666 171200 8722 172000 6 mgmt_in_data[32]
port 618 nsew signal input
rlabel metal2 s 7378 171200 7434 172000 6 mgmt_in_data[33]
port 619 nsew signal input
rlabel metal2 s 6090 171200 6146 172000 6 mgmt_in_data[34]
port 620 nsew signal input
rlabel metal2 s 4802 171200 4858 172000 6 mgmt_in_data[35]
port 621 nsew signal input
rlabel metal2 s 3514 171200 3570 172000 6 mgmt_in_data[36]
port 622 nsew signal input
rlabel metal2 s 2226 171200 2282 172000 6 mgmt_in_data[37]
port 623 nsew signal input
rlabel metal3 s 429200 87864 430000 87984 6 mgmt_in_data[3]
port 624 nsew signal input
rlabel metal3 s 429200 91808 430000 91928 6 mgmt_in_data[4]
port 625 nsew signal input
rlabel metal3 s 429200 95616 430000 95736 6 mgmt_in_data[5]
port 626 nsew signal input
rlabel metal3 s 429200 99424 430000 99544 6 mgmt_in_data[6]
port 627 nsew signal input
rlabel metal3 s 429200 103368 430000 103488 6 mgmt_in_data[7]
port 628 nsew signal input
rlabel metal3 s 429200 107176 430000 107296 6 mgmt_in_data[8]
port 629 nsew signal input
rlabel metal3 s 429200 111120 430000 111240 6 mgmt_in_data[9]
port 630 nsew signal input
rlabel metal3 s 429200 78208 430000 78328 6 mgmt_out_data[0]
port 631 nsew signal output
rlabel metal3 s 429200 116832 430000 116952 6 mgmt_out_data[10]
port 632 nsew signal output
rlabel metal3 s 429200 120776 430000 120896 6 mgmt_out_data[11]
port 633 nsew signal output
rlabel metal3 s 429200 124584 430000 124704 6 mgmt_out_data[12]
port 634 nsew signal output
rlabel metal3 s 429200 128528 430000 128648 6 mgmt_out_data[13]
port 635 nsew signal output
rlabel metal3 s 429200 132336 430000 132456 6 mgmt_out_data[14]
port 636 nsew signal output
rlabel metal3 s 429200 136144 430000 136264 6 mgmt_out_data[15]
port 637 nsew signal output
rlabel metal3 s 429200 140088 430000 140208 6 mgmt_out_data[16]
port 638 nsew signal output
rlabel metal3 s 429200 143896 430000 144016 6 mgmt_out_data[17]
port 639 nsew signal output
rlabel metal3 s 429200 147840 430000 147960 6 mgmt_out_data[18]
port 640 nsew signal output
rlabel metal3 s 429200 151648 430000 151768 6 mgmt_out_data[19]
port 641 nsew signal output
rlabel metal3 s 429200 82016 430000 82136 6 mgmt_out_data[1]
port 642 nsew signal output
rlabel metal3 s 429200 155592 430000 155712 6 mgmt_out_data[20]
port 643 nsew signal output
rlabel metal3 s 429200 159400 430000 159520 6 mgmt_out_data[21]
port 644 nsew signal output
rlabel metal3 s 429200 163208 430000 163328 6 mgmt_out_data[22]
port 645 nsew signal output
rlabel metal3 s 429200 167152 430000 167272 6 mgmt_out_data[23]
port 646 nsew signal output
rlabel metal2 s 19706 171200 19762 172000 6 mgmt_out_data[24]
port 647 nsew signal output
rlabel metal2 s 18418 171200 18474 172000 6 mgmt_out_data[25]
port 648 nsew signal output
rlabel metal2 s 17130 171200 17186 172000 6 mgmt_out_data[26]
port 649 nsew signal output
rlabel metal2 s 15842 171200 15898 172000 6 mgmt_out_data[27]
port 650 nsew signal output
rlabel metal2 s 14554 171200 14610 172000 6 mgmt_out_data[28]
port 651 nsew signal output
rlabel metal2 s 13266 171200 13322 172000 6 mgmt_out_data[29]
port 652 nsew signal output
rlabel metal3 s 429200 85960 430000 86080 6 mgmt_out_data[2]
port 653 nsew signal output
rlabel metal2 s 11978 171200 12034 172000 6 mgmt_out_data[30]
port 654 nsew signal output
rlabel metal2 s 10598 171200 10654 172000 6 mgmt_out_data[31]
port 655 nsew signal output
rlabel metal2 s 9310 171200 9366 172000 6 mgmt_out_data[32]
port 656 nsew signal output
rlabel metal2 s 8022 171200 8078 172000 6 mgmt_out_data[33]
port 657 nsew signal output
rlabel metal2 s 6734 171200 6790 172000 6 mgmt_out_data[34]
port 658 nsew signal output
rlabel metal2 s 5446 171200 5502 172000 6 mgmt_out_data[35]
port 659 nsew signal output
rlabel metal2 s 4158 171200 4214 172000 6 mgmt_out_data[36]
port 660 nsew signal output
rlabel metal2 s 2870 171200 2926 172000 6 mgmt_out_data[37]
port 661 nsew signal output
rlabel metal3 s 429200 89768 430000 89888 6 mgmt_out_data[3]
port 662 nsew signal output
rlabel metal3 s 429200 93712 430000 93832 6 mgmt_out_data[4]
port 663 nsew signal output
rlabel metal3 s 429200 97520 430000 97640 6 mgmt_out_data[5]
port 664 nsew signal output
rlabel metal3 s 429200 101464 430000 101584 6 mgmt_out_data[6]
port 665 nsew signal output
rlabel metal3 s 429200 105272 430000 105392 6 mgmt_out_data[7]
port 666 nsew signal output
rlabel metal3 s 429200 109080 430000 109200 6 mgmt_out_data[8]
port 667 nsew signal output
rlabel metal3 s 429200 113024 430000 113144 6 mgmt_out_data[9]
port 668 nsew signal output
rlabel metal3 s 0 20816 800 20936 6 mgmt_rdata[0]
port 669 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 mgmt_rdata[10]
port 670 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 mgmt_rdata[11]
port 671 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 mgmt_rdata[12]
port 672 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 mgmt_rdata[13]
port 673 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 mgmt_rdata[14]
port 674 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 mgmt_rdata[15]
port 675 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 mgmt_rdata[16]
port 676 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 mgmt_rdata[17]
port 677 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 mgmt_rdata[18]
port 678 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 mgmt_rdata[19]
port 679 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 mgmt_rdata[1]
port 680 nsew signal input
rlabel metal3 s 0 42304 800 42424 6 mgmt_rdata[20]
port 681 nsew signal input
rlabel metal3 s 0 43392 800 43512 6 mgmt_rdata[21]
port 682 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 mgmt_rdata[22]
port 683 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 mgmt_rdata[23]
port 684 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 mgmt_rdata[24]
port 685 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 mgmt_rdata[25]
port 686 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 mgmt_rdata[26]
port 687 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 mgmt_rdata[27]
port 688 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 mgmt_rdata[28]
port 689 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 mgmt_rdata[29]
port 690 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 mgmt_rdata[2]
port 691 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 mgmt_rdata[30]
port 692 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 mgmt_rdata[31]
port 693 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 mgmt_rdata[32]
port 694 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 mgmt_rdata[33]
port 695 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 mgmt_rdata[34]
port 696 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 mgmt_rdata[35]
port 697 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 mgmt_rdata[36]
port 698 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 mgmt_rdata[37]
port 699 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 mgmt_rdata[38]
port 700 nsew signal input
rlabel metal3 s 0 62704 800 62824 6 mgmt_rdata[39]
port 701 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 mgmt_rdata[3]
port 702 nsew signal input
rlabel metal3 s 0 63792 800 63912 6 mgmt_rdata[40]
port 703 nsew signal input
rlabel metal3 s 0 64880 800 65000 6 mgmt_rdata[41]
port 704 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 mgmt_rdata[42]
port 705 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 mgmt_rdata[43]
port 706 nsew signal input
rlabel metal3 s 0 68144 800 68264 6 mgmt_rdata[44]
port 707 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 mgmt_rdata[45]
port 708 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 mgmt_rdata[46]
port 709 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 mgmt_rdata[47]
port 710 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 mgmt_rdata[48]
port 711 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 mgmt_rdata[49]
port 712 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 mgmt_rdata[4]
port 713 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 mgmt_rdata[50]
port 714 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 mgmt_rdata[51]
port 715 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 mgmt_rdata[52]
port 716 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 mgmt_rdata[53]
port 717 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 mgmt_rdata[54]
port 718 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 mgmt_rdata[55]
port 719 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 mgmt_rdata[56]
port 720 nsew signal input
rlabel metal3 s 0 82016 800 82136 6 mgmt_rdata[57]
port 721 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 mgmt_rdata[58]
port 722 nsew signal input
rlabel metal3 s 0 84192 800 84312 6 mgmt_rdata[59]
port 723 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 mgmt_rdata[5]
port 724 nsew signal input
rlabel metal3 s 0 85280 800 85400 6 mgmt_rdata[60]
port 725 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 mgmt_rdata[61]
port 726 nsew signal input
rlabel metal3 s 0 87456 800 87576 6 mgmt_rdata[62]
port 727 nsew signal input
rlabel metal3 s 0 88544 800 88664 6 mgmt_rdata[63]
port 728 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 mgmt_rdata[6]
port 729 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 mgmt_rdata[7]
port 730 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 mgmt_rdata[8]
port 731 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 mgmt_rdata[9]
port 732 nsew signal input
rlabel metal3 s 0 89632 800 89752 6 mgmt_rdata_ro[0]
port 733 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 mgmt_rdata_ro[10]
port 734 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 mgmt_rdata_ro[11]
port 735 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 mgmt_rdata_ro[12]
port 736 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 mgmt_rdata_ro[13]
port 737 nsew signal input
rlabel metal3 s 0 104592 800 104712 6 mgmt_rdata_ro[14]
port 738 nsew signal input
rlabel metal3 s 0 105680 800 105800 6 mgmt_rdata_ro[15]
port 739 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 mgmt_rdata_ro[16]
port 740 nsew signal input
rlabel metal3 s 0 107856 800 107976 6 mgmt_rdata_ro[17]
port 741 nsew signal input
rlabel metal3 s 0 108944 800 109064 6 mgmt_rdata_ro[18]
port 742 nsew signal input
rlabel metal3 s 0 110032 800 110152 6 mgmt_rdata_ro[19]
port 743 nsew signal input
rlabel metal3 s 0 90720 800 90840 6 mgmt_rdata_ro[1]
port 744 nsew signal input
rlabel metal3 s 0 111120 800 111240 6 mgmt_rdata_ro[20]
port 745 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 mgmt_rdata_ro[21]
port 746 nsew signal input
rlabel metal3 s 0 113296 800 113416 6 mgmt_rdata_ro[22]
port 747 nsew signal input
rlabel metal3 s 0 114384 800 114504 6 mgmt_rdata_ro[23]
port 748 nsew signal input
rlabel metal3 s 0 115336 800 115456 6 mgmt_rdata_ro[24]
port 749 nsew signal input
rlabel metal3 s 0 116424 800 116544 6 mgmt_rdata_ro[25]
port 750 nsew signal input
rlabel metal3 s 0 117512 800 117632 6 mgmt_rdata_ro[26]
port 751 nsew signal input
rlabel metal3 s 0 118600 800 118720 6 mgmt_rdata_ro[27]
port 752 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 mgmt_rdata_ro[28]
port 753 nsew signal input
rlabel metal3 s 0 120776 800 120896 6 mgmt_rdata_ro[29]
port 754 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 mgmt_rdata_ro[2]
port 755 nsew signal input
rlabel metal3 s 0 121864 800 121984 6 mgmt_rdata_ro[30]
port 756 nsew signal input
rlabel metal3 s 0 122952 800 123072 6 mgmt_rdata_ro[31]
port 757 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 mgmt_rdata_ro[3]
port 758 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 mgmt_rdata_ro[4]
port 759 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 mgmt_rdata_ro[5]
port 760 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 mgmt_rdata_ro[6]
port 761 nsew signal input
rlabel metal3 s 0 97112 800 97232 6 mgmt_rdata_ro[7]
port 762 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 mgmt_rdata_ro[8]
port 763 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 mgmt_rdata_ro[9]
port 764 nsew signal input
rlabel metal3 s 0 124040 800 124160 6 mgmt_wdata[0]
port 765 nsew signal output
rlabel metal3 s 0 134784 800 134904 6 mgmt_wdata[10]
port 766 nsew signal output
rlabel metal3 s 0 135872 800 135992 6 mgmt_wdata[11]
port 767 nsew signal output
rlabel metal3 s 0 136960 800 137080 6 mgmt_wdata[12]
port 768 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 mgmt_wdata[13]
port 769 nsew signal output
rlabel metal3 s 0 139000 800 139120 6 mgmt_wdata[14]
port 770 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 mgmt_wdata[15]
port 771 nsew signal output
rlabel metal3 s 0 141176 800 141296 6 mgmt_wdata[16]
port 772 nsew signal output
rlabel metal3 s 0 142264 800 142384 6 mgmt_wdata[17]
port 773 nsew signal output
rlabel metal3 s 0 143352 800 143472 6 mgmt_wdata[18]
port 774 nsew signal output
rlabel metal3 s 0 144440 800 144560 6 mgmt_wdata[19]
port 775 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 mgmt_wdata[1]
port 776 nsew signal output
rlabel metal3 s 0 145528 800 145648 6 mgmt_wdata[20]
port 777 nsew signal output
rlabel metal3 s 0 146616 800 146736 6 mgmt_wdata[21]
port 778 nsew signal output
rlabel metal3 s 0 147704 800 147824 6 mgmt_wdata[22]
port 779 nsew signal output
rlabel metal3 s 0 148792 800 148912 6 mgmt_wdata[23]
port 780 nsew signal output
rlabel metal3 s 0 149744 800 149864 6 mgmt_wdata[24]
port 781 nsew signal output
rlabel metal3 s 0 150832 800 150952 6 mgmt_wdata[25]
port 782 nsew signal output
rlabel metal3 s 0 151920 800 152040 6 mgmt_wdata[26]
port 783 nsew signal output
rlabel metal3 s 0 153008 800 153128 6 mgmt_wdata[27]
port 784 nsew signal output
rlabel metal3 s 0 154096 800 154216 6 mgmt_wdata[28]
port 785 nsew signal output
rlabel metal3 s 0 155184 800 155304 6 mgmt_wdata[29]
port 786 nsew signal output
rlabel metal3 s 0 126216 800 126336 6 mgmt_wdata[2]
port 787 nsew signal output
rlabel metal3 s 0 156272 800 156392 6 mgmt_wdata[30]
port 788 nsew signal output
rlabel metal3 s 0 157360 800 157480 6 mgmt_wdata[31]
port 789 nsew signal output
rlabel metal3 s 0 127168 800 127288 6 mgmt_wdata[3]
port 790 nsew signal output
rlabel metal3 s 0 128256 800 128376 6 mgmt_wdata[4]
port 791 nsew signal output
rlabel metal3 s 0 129344 800 129464 6 mgmt_wdata[5]
port 792 nsew signal output
rlabel metal3 s 0 130432 800 130552 6 mgmt_wdata[6]
port 793 nsew signal output
rlabel metal3 s 0 131520 800 131640 6 mgmt_wdata[7]
port 794 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 mgmt_wdata[8]
port 795 nsew signal output
rlabel metal3 s 0 133696 800 133816 6 mgmt_wdata[9]
port 796 nsew signal output
rlabel metal3 s 0 158448 800 158568 6 mgmt_wen[0]
port 797 nsew signal output
rlabel metal3 s 0 159536 800 159656 6 mgmt_wen[1]
port 798 nsew signal output
rlabel metal3 s 0 160624 800 160744 6 mgmt_wen_mask[0]
port 799 nsew signal output
rlabel metal3 s 0 161576 800 161696 6 mgmt_wen_mask[1]
port 800 nsew signal output
rlabel metal3 s 0 162664 800 162784 6 mgmt_wen_mask[2]
port 801 nsew signal output
rlabel metal3 s 0 163752 800 163872 6 mgmt_wen_mask[3]
port 802 nsew signal output
rlabel metal3 s 0 164840 800 164960 6 mgmt_wen_mask[4]
port 803 nsew signal output
rlabel metal3 s 0 165928 800 166048 6 mgmt_wen_mask[5]
port 804 nsew signal output
rlabel metal3 s 0 167016 800 167136 6 mgmt_wen_mask[6]
port 805 nsew signal output
rlabel metal3 s 0 168104 800 168224 6 mgmt_wen_mask[7]
port 806 nsew signal output
rlabel metal2 s 420550 171200 420606 172000 6 mprj2_vcc_pwrgood
port 807 nsew signal input
rlabel metal2 s 421194 171200 421250 172000 6 mprj2_vdd_pwrgood
port 808 nsew signal input
rlabel metal2 s 20350 171200 20406 172000 6 mprj_ack_i
port 809 nsew signal input
rlabel metal2 s 62578 171200 62634 172000 6 mprj_adr_o[0]
port 810 nsew signal output
rlabel metal2 s 69110 171200 69166 172000 6 mprj_adr_o[10]
port 811 nsew signal output
rlabel metal2 s 69754 171200 69810 172000 6 mprj_adr_o[11]
port 812 nsew signal output
rlabel metal2 s 70398 171200 70454 172000 6 mprj_adr_o[12]
port 813 nsew signal output
rlabel metal2 s 71042 171200 71098 172000 6 mprj_adr_o[13]
port 814 nsew signal output
rlabel metal2 s 71686 171200 71742 172000 6 mprj_adr_o[14]
port 815 nsew signal output
rlabel metal2 s 72330 171200 72386 172000 6 mprj_adr_o[15]
port 816 nsew signal output
rlabel metal2 s 72974 171200 73030 172000 6 mprj_adr_o[16]
port 817 nsew signal output
rlabel metal2 s 73618 171200 73674 172000 6 mprj_adr_o[17]
port 818 nsew signal output
rlabel metal2 s 74262 171200 74318 172000 6 mprj_adr_o[18]
port 819 nsew signal output
rlabel metal2 s 74906 171200 74962 172000 6 mprj_adr_o[19]
port 820 nsew signal output
rlabel metal2 s 63222 171200 63278 172000 6 mprj_adr_o[1]
port 821 nsew signal output
rlabel metal2 s 75642 171200 75698 172000 6 mprj_adr_o[20]
port 822 nsew signal output
rlabel metal2 s 76286 171200 76342 172000 6 mprj_adr_o[21]
port 823 nsew signal output
rlabel metal2 s 76930 171200 76986 172000 6 mprj_adr_o[22]
port 824 nsew signal output
rlabel metal2 s 77574 171200 77630 172000 6 mprj_adr_o[23]
port 825 nsew signal output
rlabel metal2 s 78218 171200 78274 172000 6 mprj_adr_o[24]
port 826 nsew signal output
rlabel metal2 s 78862 171200 78918 172000 6 mprj_adr_o[25]
port 827 nsew signal output
rlabel metal2 s 79506 171200 79562 172000 6 mprj_adr_o[26]
port 828 nsew signal output
rlabel metal2 s 80150 171200 80206 172000 6 mprj_adr_o[27]
port 829 nsew signal output
rlabel metal2 s 80794 171200 80850 172000 6 mprj_adr_o[28]
port 830 nsew signal output
rlabel metal2 s 81438 171200 81494 172000 6 mprj_adr_o[29]
port 831 nsew signal output
rlabel metal2 s 63866 171200 63922 172000 6 mprj_adr_o[2]
port 832 nsew signal output
rlabel metal2 s 82082 171200 82138 172000 6 mprj_adr_o[30]
port 833 nsew signal output
rlabel metal2 s 82726 171200 82782 172000 6 mprj_adr_o[31]
port 834 nsew signal output
rlabel metal2 s 64510 171200 64566 172000 6 mprj_adr_o[3]
port 835 nsew signal output
rlabel metal2 s 65246 171200 65302 172000 6 mprj_adr_o[4]
port 836 nsew signal output
rlabel metal2 s 65890 171200 65946 172000 6 mprj_adr_o[5]
port 837 nsew signal output
rlabel metal2 s 66534 171200 66590 172000 6 mprj_adr_o[6]
port 838 nsew signal output
rlabel metal2 s 67178 171200 67234 172000 6 mprj_adr_o[7]
port 839 nsew signal output
rlabel metal2 s 67822 171200 67878 172000 6 mprj_adr_o[8]
port 840 nsew signal output
rlabel metal2 s 68466 171200 68522 172000 6 mprj_adr_o[9]
port 841 nsew signal output
rlabel metal2 s 86682 171200 86738 172000 6 mprj_cyc_o
port 842 nsew signal output
rlabel metal2 s 20994 171200 21050 172000 6 mprj_dat_i[0]
port 843 nsew signal input
rlabel metal2 s 27526 171200 27582 172000 6 mprj_dat_i[10]
port 844 nsew signal input
rlabel metal2 s 28170 171200 28226 172000 6 mprj_dat_i[11]
port 845 nsew signal input
rlabel metal2 s 28814 171200 28870 172000 6 mprj_dat_i[12]
port 846 nsew signal input
rlabel metal2 s 29458 171200 29514 172000 6 mprj_dat_i[13]
port 847 nsew signal input
rlabel metal2 s 30102 171200 30158 172000 6 mprj_dat_i[14]
port 848 nsew signal input
rlabel metal2 s 30746 171200 30802 172000 6 mprj_dat_i[15]
port 849 nsew signal input
rlabel metal2 s 31390 171200 31446 172000 6 mprj_dat_i[16]
port 850 nsew signal input
rlabel metal2 s 32034 171200 32090 172000 6 mprj_dat_i[17]
port 851 nsew signal input
rlabel metal2 s 32770 171200 32826 172000 6 mprj_dat_i[18]
port 852 nsew signal input
rlabel metal2 s 33414 171200 33470 172000 6 mprj_dat_i[19]
port 853 nsew signal input
rlabel metal2 s 21638 171200 21694 172000 6 mprj_dat_i[1]
port 854 nsew signal input
rlabel metal2 s 34058 171200 34114 172000 6 mprj_dat_i[20]
port 855 nsew signal input
rlabel metal2 s 34702 171200 34758 172000 6 mprj_dat_i[21]
port 856 nsew signal input
rlabel metal2 s 35346 171200 35402 172000 6 mprj_dat_i[22]
port 857 nsew signal input
rlabel metal2 s 35990 171200 36046 172000 6 mprj_dat_i[23]
port 858 nsew signal input
rlabel metal2 s 36634 171200 36690 172000 6 mprj_dat_i[24]
port 859 nsew signal input
rlabel metal2 s 37278 171200 37334 172000 6 mprj_dat_i[25]
port 860 nsew signal input
rlabel metal2 s 37922 171200 37978 172000 6 mprj_dat_i[26]
port 861 nsew signal input
rlabel metal2 s 38566 171200 38622 172000 6 mprj_dat_i[27]
port 862 nsew signal input
rlabel metal2 s 39210 171200 39266 172000 6 mprj_dat_i[28]
port 863 nsew signal input
rlabel metal2 s 39854 171200 39910 172000 6 mprj_dat_i[29]
port 864 nsew signal input
rlabel metal2 s 22374 171200 22430 172000 6 mprj_dat_i[2]
port 865 nsew signal input
rlabel metal2 s 40498 171200 40554 172000 6 mprj_dat_i[30]
port 866 nsew signal input
rlabel metal2 s 41142 171200 41198 172000 6 mprj_dat_i[31]
port 867 nsew signal input
rlabel metal2 s 23018 171200 23074 172000 6 mprj_dat_i[3]
port 868 nsew signal input
rlabel metal2 s 23662 171200 23718 172000 6 mprj_dat_i[4]
port 869 nsew signal input
rlabel metal2 s 24306 171200 24362 172000 6 mprj_dat_i[5]
port 870 nsew signal input
rlabel metal2 s 24950 171200 25006 172000 6 mprj_dat_i[6]
port 871 nsew signal input
rlabel metal2 s 25594 171200 25650 172000 6 mprj_dat_i[7]
port 872 nsew signal input
rlabel metal2 s 26238 171200 26294 172000 6 mprj_dat_i[8]
port 873 nsew signal input
rlabel metal2 s 26882 171200 26938 172000 6 mprj_dat_i[9]
port 874 nsew signal input
rlabel metal2 s 41786 171200 41842 172000 6 mprj_dat_o[0]
port 875 nsew signal output
rlabel metal2 s 48318 171200 48374 172000 6 mprj_dat_o[10]
port 876 nsew signal output
rlabel metal2 s 48962 171200 49018 172000 6 mprj_dat_o[11]
port 877 nsew signal output
rlabel metal2 s 49606 171200 49662 172000 6 mprj_dat_o[12]
port 878 nsew signal output
rlabel metal2 s 50250 171200 50306 172000 6 mprj_dat_o[13]
port 879 nsew signal output
rlabel metal2 s 50894 171200 50950 172000 6 mprj_dat_o[14]
port 880 nsew signal output
rlabel metal2 s 51538 171200 51594 172000 6 mprj_dat_o[15]
port 881 nsew signal output
rlabel metal2 s 52182 171200 52238 172000 6 mprj_dat_o[16]
port 882 nsew signal output
rlabel metal2 s 52826 171200 52882 172000 6 mprj_dat_o[17]
port 883 nsew signal output
rlabel metal2 s 53470 171200 53526 172000 6 mprj_dat_o[18]
port 884 nsew signal output
rlabel metal2 s 54206 171200 54262 172000 6 mprj_dat_o[19]
port 885 nsew signal output
rlabel metal2 s 42430 171200 42486 172000 6 mprj_dat_o[1]
port 886 nsew signal output
rlabel metal2 s 54850 171200 54906 172000 6 mprj_dat_o[20]
port 887 nsew signal output
rlabel metal2 s 55494 171200 55550 172000 6 mprj_dat_o[21]
port 888 nsew signal output
rlabel metal2 s 56138 171200 56194 172000 6 mprj_dat_o[22]
port 889 nsew signal output
rlabel metal2 s 56782 171200 56838 172000 6 mprj_dat_o[23]
port 890 nsew signal output
rlabel metal2 s 57426 171200 57482 172000 6 mprj_dat_o[24]
port 891 nsew signal output
rlabel metal2 s 58070 171200 58126 172000 6 mprj_dat_o[25]
port 892 nsew signal output
rlabel metal2 s 58714 171200 58770 172000 6 mprj_dat_o[26]
port 893 nsew signal output
rlabel metal2 s 59358 171200 59414 172000 6 mprj_dat_o[27]
port 894 nsew signal output
rlabel metal2 s 60002 171200 60058 172000 6 mprj_dat_o[28]
port 895 nsew signal output
rlabel metal2 s 60646 171200 60702 172000 6 mprj_dat_o[29]
port 896 nsew signal output
rlabel metal2 s 43074 171200 43130 172000 6 mprj_dat_o[2]
port 897 nsew signal output
rlabel metal2 s 61290 171200 61346 172000 6 mprj_dat_o[30]
port 898 nsew signal output
rlabel metal2 s 61934 171200 61990 172000 6 mprj_dat_o[31]
port 899 nsew signal output
rlabel metal2 s 43810 171200 43866 172000 6 mprj_dat_o[3]
port 900 nsew signal output
rlabel metal2 s 44454 171200 44510 172000 6 mprj_dat_o[4]
port 901 nsew signal output
rlabel metal2 s 45098 171200 45154 172000 6 mprj_dat_o[5]
port 902 nsew signal output
rlabel metal2 s 45742 171200 45798 172000 6 mprj_dat_o[6]
port 903 nsew signal output
rlabel metal2 s 46386 171200 46442 172000 6 mprj_dat_o[7]
port 904 nsew signal output
rlabel metal2 s 47030 171200 47086 172000 6 mprj_dat_o[8]
port 905 nsew signal output
rlabel metal2 s 47674 171200 47730 172000 6 mprj_dat_o[9]
port 906 nsew signal output
rlabel metal3 s 429200 70456 430000 70576 6 mprj_io_loader_clock
port 907 nsew signal output
rlabel metal2 s 429566 171200 429622 172000 6 mprj_io_loader_data_1
port 908 nsew signal output
rlabel metal3 s 0 171368 800 171488 6 mprj_io_loader_data_2
port 909 nsew signal output
rlabel metal3 s 429200 68552 430000 68672 6 mprj_io_loader_resetn
port 910 nsew signal output
rlabel metal2 s 83370 171200 83426 172000 6 mprj_sel_o[0]
port 911 nsew signal output
rlabel metal2 s 84014 171200 84070 172000 6 mprj_sel_o[1]
port 912 nsew signal output
rlabel metal2 s 84658 171200 84714 172000 6 mprj_sel_o[2]
port 913 nsew signal output
rlabel metal2 s 85302 171200 85358 172000 6 mprj_sel_o[3]
port 914 nsew signal output
rlabel metal2 s 85946 171200 86002 172000 6 mprj_stb_o
port 915 nsew signal output
rlabel metal2 s 421838 171200 421894 172000 6 mprj_vcc_pwrgood
port 916 nsew signal input
rlabel metal2 s 422482 171200 422538 172000 6 mprj_vdd_pwrgood
port 917 nsew signal input
rlabel metal2 s 87326 171200 87382 172000 6 mprj_we_o
port 918 nsew signal output
rlabel metal3 s 429200 62704 430000 62824 6 porb
port 919 nsew signal input
rlabel metal2 s 423126 171200 423182 172000 6 pwr_ctrl_out[0]
port 920 nsew signal output
rlabel metal2 s 423770 171200 423826 172000 6 pwr_ctrl_out[1]
port 921 nsew signal output
rlabel metal2 s 424414 171200 424470 172000 6 pwr_ctrl_out[2]
port 922 nsew signal output
rlabel metal2 s 425058 171200 425114 172000 6 pwr_ctrl_out[3]
port 923 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 resetb
port 924 nsew signal input
rlabel metal3 s 429200 72360 430000 72480 6 sdo_out
port 925 nsew signal output
rlabel metal3 s 429200 74400 430000 74520 6 sdo_outenb
port 926 nsew signal output
rlabel metal2 s 1582 171200 1638 172000 6 user_clk
port 927 nsew signal output
rlabel metal2 s 425702 171200 425758 172000 6 user_irq[0]
port 928 nsew signal input
rlabel metal2 s 426346 171200 426402 172000 6 user_irq[1]
port 929 nsew signal input
rlabel metal2 s 426990 171200 427046 172000 6 user_irq[2]
port 930 nsew signal input
rlabel metal2 s 427634 171200 427690 172000 6 user_irq_ena[0]
port 931 nsew signal output
rlabel metal2 s 428278 171200 428334 172000 6 user_irq_ena[1]
port 932 nsew signal output
rlabel metal2 s 428922 171200 428978 172000 6 user_irq_ena[2]
port 933 nsew signal output
rlabel metal4 s 424208 2128 424528 169776 6 VPWR
port 934 nsew power bidirectional
rlabel metal4 s 414208 2128 414528 169776 6 VPWR
port 935 nsew power bidirectional
rlabel metal4 s 404208 2128 404528 169776 6 VPWR
port 936 nsew power bidirectional
rlabel metal4 s 394208 164296 394528 169776 6 VPWR
port 937 nsew power bidirectional
rlabel metal4 s 384208 2128 384528 169776 6 VPWR
port 938 nsew power bidirectional
rlabel metal4 s 374208 2128 374528 169776 6 VPWR
port 939 nsew power bidirectional
rlabel metal4 s 364208 2128 364528 169776 6 VPWR
port 940 nsew power bidirectional
rlabel metal4 s 354208 2128 354528 169776 6 VPWR
port 941 nsew power bidirectional
rlabel metal4 s 344208 2128 344528 169776 6 VPWR
port 942 nsew power bidirectional
rlabel metal4 s 334208 2128 334528 169776 6 VPWR
port 943 nsew power bidirectional
rlabel metal4 s 324208 2128 324528 169776 6 VPWR
port 944 nsew power bidirectional
rlabel metal4 s 314208 2128 314528 169776 6 VPWR
port 945 nsew power bidirectional
rlabel metal4 s 304208 2128 304528 169776 6 VPWR
port 946 nsew power bidirectional
rlabel metal4 s 294208 2128 294528 169776 6 VPWR
port 947 nsew power bidirectional
rlabel metal4 s 284208 2128 284528 169776 6 VPWR
port 948 nsew power bidirectional
rlabel metal4 s 274208 2128 274528 169776 6 VPWR
port 949 nsew power bidirectional
rlabel metal4 s 264208 2128 264528 169776 6 VPWR
port 950 nsew power bidirectional
rlabel metal4 s 254208 2128 254528 169776 6 VPWR
port 951 nsew power bidirectional
rlabel metal4 s 244208 2128 244528 169776 6 VPWR
port 952 nsew power bidirectional
rlabel metal4 s 234208 2128 234528 169776 6 VPWR
port 953 nsew power bidirectional
rlabel metal4 s 224208 2128 224528 169776 6 VPWR
port 954 nsew power bidirectional
rlabel metal4 s 214208 2128 214528 169776 6 VPWR
port 955 nsew power bidirectional
rlabel metal4 s 204208 2128 204528 169776 6 VPWR
port 956 nsew power bidirectional
rlabel metal4 s 194208 2128 194528 169776 6 VPWR
port 957 nsew power bidirectional
rlabel metal4 s 184208 2128 184528 169776 6 VPWR
port 958 nsew power bidirectional
rlabel metal4 s 174208 128152 174528 169776 6 VPWR
port 959 nsew power bidirectional
rlabel metal4 s 164208 128152 164528 169776 6 VPWR
port 960 nsew power bidirectional
rlabel metal4 s 154208 128152 154528 169776 6 VPWR
port 961 nsew power bidirectional
rlabel metal4 s 144208 128152 144528 169776 6 VPWR
port 962 nsew power bidirectional
rlabel metal4 s 134208 128152 134528 169776 6 VPWR
port 963 nsew power bidirectional
rlabel metal4 s 124208 128152 124528 169776 6 VPWR
port 964 nsew power bidirectional
rlabel metal4 s 114208 128152 114528 169776 6 VPWR
port 965 nsew power bidirectional
rlabel metal4 s 104208 128152 104528 169776 6 VPWR
port 966 nsew power bidirectional
rlabel metal4 s 94208 128152 94528 169776 6 VPWR
port 967 nsew power bidirectional
rlabel metal4 s 84208 128152 84528 169776 6 VPWR
port 968 nsew power bidirectional
rlabel metal4 s 74208 128152 74528 169776 6 VPWR
port 969 nsew power bidirectional
rlabel metal4 s 64208 128152 64528 169776 6 VPWR
port 970 nsew power bidirectional
rlabel metal4 s 54208 128152 54528 169776 6 VPWR
port 971 nsew power bidirectional
rlabel metal4 s 44208 128152 44528 169776 6 VPWR
port 972 nsew power bidirectional
rlabel metal4 s 34208 128152 34528 169776 6 VPWR
port 973 nsew power bidirectional
rlabel metal4 s 24208 128152 24528 169776 6 VPWR
port 974 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 169776 6 VPWR
port 975 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 169776 6 VPWR
port 976 nsew power bidirectional
rlabel metal4 s 394208 2128 394528 145392 6 VPWR
port 977 nsew power bidirectional
rlabel metal4 s 174208 2128 174528 21248 6 VPWR
port 978 nsew power bidirectional
rlabel metal4 s 164208 2128 164528 21248 6 VPWR
port 979 nsew power bidirectional
rlabel metal4 s 154208 2128 154528 21248 6 VPWR
port 980 nsew power bidirectional
rlabel metal4 s 144208 2128 144528 21248 6 VPWR
port 981 nsew power bidirectional
rlabel metal4 s 134208 2128 134528 21248 6 VPWR
port 982 nsew power bidirectional
rlabel metal4 s 124208 2128 124528 21248 6 VPWR
port 983 nsew power bidirectional
rlabel metal4 s 114208 2128 114528 21248 6 VPWR
port 984 nsew power bidirectional
rlabel metal4 s 104208 2128 104528 21248 6 VPWR
port 985 nsew power bidirectional
rlabel metal4 s 94208 2128 94528 21248 6 VPWR
port 986 nsew power bidirectional
rlabel metal4 s 84208 2128 84528 21248 6 VPWR
port 987 nsew power bidirectional
rlabel metal4 s 74208 2128 74528 21248 6 VPWR
port 988 nsew power bidirectional
rlabel metal4 s 64208 2128 64528 21248 6 VPWR
port 989 nsew power bidirectional
rlabel metal4 s 54208 2128 54528 21248 6 VPWR
port 990 nsew power bidirectional
rlabel metal4 s 44208 2128 44528 21248 6 VPWR
port 991 nsew power bidirectional
rlabel metal4 s 34208 2128 34528 21248 6 VPWR
port 992 nsew power bidirectional
rlabel metal4 s 24208 2128 24528 21248 6 VPWR
port 993 nsew power bidirectional
rlabel metal5 s 1104 161298 428812 161618 6 VPWR
port 994 nsew power bidirectional
rlabel metal5 s 1104 135298 428812 135618 6 VPWR
port 995 nsew power bidirectional
rlabel metal5 s 1104 109298 428812 109618 6 VPWR
port 996 nsew power bidirectional
rlabel metal5 s 1104 83298 428812 83618 6 VPWR
port 997 nsew power bidirectional
rlabel metal5 s 1104 57298 428812 57618 6 VPWR
port 998 nsew power bidirectional
rlabel metal5 s 1104 31298 428812 31618 6 VPWR
port 999 nsew power bidirectional
rlabel metal5 s 1104 5298 428812 5618 6 VPWR
port 1000 nsew power bidirectional
rlabel metal4 s 419208 2128 419528 169776 6 VGND
port 1001 nsew ground bidirectional
rlabel metal4 s 409208 2128 409528 169776 6 VGND
port 1002 nsew ground bidirectional
rlabel metal4 s 399208 164296 399528 169776 6 VGND
port 1003 nsew ground bidirectional
rlabel metal4 s 389208 164296 389528 169776 6 VGND
port 1004 nsew ground bidirectional
rlabel metal4 s 379208 2128 379528 169776 6 VGND
port 1005 nsew ground bidirectional
rlabel metal4 s 369208 2128 369528 169776 6 VGND
port 1006 nsew ground bidirectional
rlabel metal4 s 359208 2128 359528 169776 6 VGND
port 1007 nsew ground bidirectional
rlabel metal4 s 349208 2128 349528 169776 6 VGND
port 1008 nsew ground bidirectional
rlabel metal4 s 339208 2128 339528 169776 6 VGND
port 1009 nsew ground bidirectional
rlabel metal4 s 329208 2128 329528 169776 6 VGND
port 1010 nsew ground bidirectional
rlabel metal4 s 319208 2128 319528 169776 6 VGND
port 1011 nsew ground bidirectional
rlabel metal4 s 309208 2128 309528 169776 6 VGND
port 1012 nsew ground bidirectional
rlabel metal4 s 299208 2128 299528 169776 6 VGND
port 1013 nsew ground bidirectional
rlabel metal4 s 289208 2128 289528 169776 6 VGND
port 1014 nsew ground bidirectional
rlabel metal4 s 279208 2128 279528 169776 6 VGND
port 1015 nsew ground bidirectional
rlabel metal4 s 269208 2128 269528 169776 6 VGND
port 1016 nsew ground bidirectional
rlabel metal4 s 259208 2128 259528 169776 6 VGND
port 1017 nsew ground bidirectional
rlabel metal4 s 249208 2128 249528 169776 6 VGND
port 1018 nsew ground bidirectional
rlabel metal4 s 239208 2128 239528 169776 6 VGND
port 1019 nsew ground bidirectional
rlabel metal4 s 229208 2128 229528 169776 6 VGND
port 1020 nsew ground bidirectional
rlabel metal4 s 219208 2128 219528 169776 6 VGND
port 1021 nsew ground bidirectional
rlabel metal4 s 209208 2128 209528 169776 6 VGND
port 1022 nsew ground bidirectional
rlabel metal4 s 199208 2128 199528 169776 6 VGND
port 1023 nsew ground bidirectional
rlabel metal4 s 189208 2128 189528 169776 6 VGND
port 1024 nsew ground bidirectional
rlabel metal4 s 179208 2128 179528 169776 6 VGND
port 1025 nsew ground bidirectional
rlabel metal4 s 169208 128152 169528 169776 6 VGND
port 1026 nsew ground bidirectional
rlabel metal4 s 159208 128152 159528 169776 6 VGND
port 1027 nsew ground bidirectional
rlabel metal4 s 149208 128152 149528 169776 6 VGND
port 1028 nsew ground bidirectional
rlabel metal4 s 139208 128152 139528 169776 6 VGND
port 1029 nsew ground bidirectional
rlabel metal4 s 129208 128152 129528 169776 6 VGND
port 1030 nsew ground bidirectional
rlabel metal4 s 119208 128152 119528 169776 6 VGND
port 1031 nsew ground bidirectional
rlabel metal4 s 109208 128152 109528 169776 6 VGND
port 1032 nsew ground bidirectional
rlabel metal4 s 99208 128152 99528 169776 6 VGND
port 1033 nsew ground bidirectional
rlabel metal4 s 89208 128152 89528 169776 6 VGND
port 1034 nsew ground bidirectional
rlabel metal4 s 79208 128152 79528 169776 6 VGND
port 1035 nsew ground bidirectional
rlabel metal4 s 69208 128152 69528 169776 6 VGND
port 1036 nsew ground bidirectional
rlabel metal4 s 59208 128152 59528 169776 6 VGND
port 1037 nsew ground bidirectional
rlabel metal4 s 49208 128152 49528 169776 6 VGND
port 1038 nsew ground bidirectional
rlabel metal4 s 39208 128152 39528 169776 6 VGND
port 1039 nsew ground bidirectional
rlabel metal4 s 29208 128152 29528 169776 6 VGND
port 1040 nsew ground bidirectional
rlabel metal4 s 19208 2128 19528 169776 6 VGND
port 1041 nsew ground bidirectional
rlabel metal4 s 9208 2128 9528 169776 6 VGND
port 1042 nsew ground bidirectional
rlabel metal4 s 399208 2128 399528 145392 6 VGND
port 1043 nsew ground bidirectional
rlabel metal4 s 389208 2128 389528 145392 6 VGND
port 1044 nsew ground bidirectional
rlabel metal4 s 169208 2128 169528 21248 6 VGND
port 1045 nsew ground bidirectional
rlabel metal4 s 159208 2128 159528 21248 6 VGND
port 1046 nsew ground bidirectional
rlabel metal4 s 149208 2128 149528 21248 6 VGND
port 1047 nsew ground bidirectional
rlabel metal4 s 139208 2128 139528 21248 6 VGND
port 1048 nsew ground bidirectional
rlabel metal4 s 129208 2128 129528 21248 6 VGND
port 1049 nsew ground bidirectional
rlabel metal4 s 119208 2128 119528 21248 6 VGND
port 1050 nsew ground bidirectional
rlabel metal4 s 109208 2128 109528 21248 6 VGND
port 1051 nsew ground bidirectional
rlabel metal4 s 99208 2128 99528 21248 6 VGND
port 1052 nsew ground bidirectional
rlabel metal4 s 89208 2128 89528 21248 6 VGND
port 1053 nsew ground bidirectional
rlabel metal4 s 79208 2128 79528 21248 6 VGND
port 1054 nsew ground bidirectional
rlabel metal4 s 69208 2128 69528 21248 6 VGND
port 1055 nsew ground bidirectional
rlabel metal4 s 59208 2128 59528 21248 6 VGND
port 1056 nsew ground bidirectional
rlabel metal4 s 49208 2128 49528 21248 6 VGND
port 1057 nsew ground bidirectional
rlabel metal4 s 39208 2128 39528 21248 6 VGND
port 1058 nsew ground bidirectional
rlabel metal4 s 29208 2128 29528 21248 6 VGND
port 1059 nsew ground bidirectional
rlabel metal5 s 1104 148298 428812 148618 6 VGND
port 1060 nsew ground bidirectional
rlabel metal5 s 1104 122298 428812 122618 6 VGND
port 1061 nsew ground bidirectional
rlabel metal5 s 1104 96298 428812 96618 6 VGND
port 1062 nsew ground bidirectional
rlabel metal5 s 1104 70298 428812 70618 6 VGND
port 1063 nsew ground bidirectional
rlabel metal5 s 1104 44298 428812 44618 6 VGND
port 1064 nsew ground bidirectional
rlabel metal5 s 1104 18298 428812 18618 6 VGND
port 1065 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 430000 172000
string LEFview TRUE
string GDS_FILE /project/openlane/mgmt_core/runs/mgmt_core/results/magic/mgmt_core.gds
string GDS_END 182757822
string GDS_START 63832838
<< end >>

