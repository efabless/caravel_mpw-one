magic
tech sky130A
magscale 12 1
timestamp 1598785304
<< metal5 >>
rect 15 100 40 105
rect 5 95 45 100
rect 0 90 45 95
rect 60 90 75 95
rect 0 85 75 90
rect 0 80 15 85
rect 30 80 75 85
rect 30 75 70 80
rect 35 70 60 75
<< properties >>
string FIXED_BBOX 0 -30 90 105
<< end >>
