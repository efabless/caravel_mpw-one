* SPICE NETLIST
***************************************


***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808592 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.21 p=1.84
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808593 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.84 AS=0.84 PD=6.56 PS=6.56 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
.ENDS
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__res75only_small PAD ROUT
**
R0 PAD ROUT sky130_fd_pr__res_generic_po L=3.15 W=2 m=1
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808560 1 2 3 4 5
**
XM0 5 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=2.205 PD=7.28 PS=14.63 NRD=0 NRS=0.5586 m=1 sa=250000 sb=250005 a=3.5 p=15
XM1 3 2 5 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=1.225 AS=0.98 PD=7.35 PS=7.28 NRD=0.5586 NRS=0 m=1 sa=250001 sb=250004 a=3.5 p=15
XM2 5 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.225 PD=7.28 PS=7.35 NRD=0 NRS=0.5586 m=1 sa=250002 sb=250003 a=3.5 p=15
XM3 4 2 5 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=1.225 AS=0.98 PD=7.35 PS=7.28 NRD=0.5586 NRS=0 m=1 sa=250002 sb=250003 a=3.5 p=15
XM4 5 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.225 PD=7.28 PS=7.35 NRD=0 NRS=0.5586 m=1 sa=250003 sb=250002 a=3.5 p=15
XM5 4 2 5 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=1.225 AS=0.98 PD=7.35 PS=7.28 NRD=0.5586 NRS=0 m=1 sa=250004 sb=250001 a=3.5 p=15
XM6 5 2 4 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=1.96 AS=1.225 PD=14.56 PS=7.35 NRD=0 NRS=0.5586 m=1 sa=250005 sb=250000 a=3.5 p=15
.ENDS
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__amux_switch_1v2b VSSD 3 6 VDDIO VDDA PG_PAD_VDDIOQ_H_N PG_AMX_VDDA_H_N NG_AMX_VPMP_H NG_PAD_VPMP_H PAD_HV_P0 PAD_HV_P1 AMUXBUS_HV PAD_HV_N2 PAD_HV_N3 PAD_HV_N0 PAD_HV_N1
**
*.SEEDPROM
XM0 PAD_HV_N2 NG_PAD_VPMP_H 6 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=2.205 PD=7.28 PS=14.63 NRD=0 NRS=0.5586 m=1 sa=250000 sb=250006 a=3.5 p=15
XM1 6 NG_PAD_VPMP_H PAD_HV_N2 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=1.225 AS=0.98 PD=7.35 PS=7.28 NRD=0.5586 NRS=0 m=1 sa=250001 sb=250005 a=3.5 p=15
XM2 PAD_HV_N2 NG_PAD_VPMP_H 6 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.225 PD=7.28 PS=7.35 NRD=0 NRS=0.5586 m=1 sa=250002 sb=250004 a=3.5 p=15
XM3 6 NG_PAD_VPMP_H PAD_HV_N2 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=1.225 AS=0.98 PD=7.35 PS=7.28 NRD=0.5586 NRS=0 m=1 sa=250002 sb=250003 a=3.5 p=15
XM4 PAD_HV_N3 NG_PAD_VPMP_H 6 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.225 PD=7.28 PS=7.35 NRD=0 NRS=0.5586 m=1 sa=250003 sb=250002 a=3.5 p=15
XM5 6 NG_PAD_VPMP_H PAD_HV_N3 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=1.225 AS=0.98 PD=7.35 PS=7.28 NRD=0.5586 NRS=0 m=1 sa=250004 sb=250002 a=3.5 p=15
XM6 PAD_HV_N3 NG_PAD_VPMP_H 6 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.225 PD=7.28 PS=7.35 NRD=0 NRS=0.5586 m=1 sa=250005 sb=250001 a=3.5 p=15
XM7 6 NG_PAD_VPMP_H PAD_HV_N3 6 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=2.205 AS=0.98 PD=14.63 PS=7.28 NRD=0.5586 NRS=0 m=1 sa=250006 sb=250000 a=3.5 p=15
XM8 3 PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=2.205 PD=7.28 PS=14.63 NRD=0 NRS=0.9359 m=1 sa=250000 sb=250004 a=3.5 p=15
XM9 PAD_HV_P0 PG_PAD_VDDIOQ_H_N 3 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=1.225 AS=0.98 PD=7.35 PS=7.28 NRD=0.9359 NRS=0 m=1 sa=250001 sb=250003 a=3.5 p=15
XM10 3 PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.225 PD=7.28 PS=7.35 NRD=0 NRS=0.9359 m=1 sa=250002 sb=250002 a=3.5 p=15
XM11 PAD_HV_P1 PG_PAD_VDDIOQ_H_N 3 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=1.225 AS=0.98 PD=7.35 PS=7.28 NRD=0.9359 NRS=0 m=1 sa=250002 sb=250002 a=3.5 p=15
XM12 3 PG_PAD_VDDIOQ_H_N PAD_HV_P1 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.225 PD=7.28 PS=7.35 NRD=0 NRS=0.9359 m=1 sa=250003 sb=250001 a=3.5 p=15
XM13 PAD_HV_P1 PG_PAD_VDDIOQ_H_N 3 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=2.205 AS=0.98 PD=14.63 PS=7.28 NRD=0.9359 NRS=0 m=1 sa=250004 sb=250000 a=3.5 p=15
XM14 3 PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=1.225 AS=1.96 PD=7.35 PS=14.56 NRD=0.9359 NRS=0 m=1 sa=250000 sb=250003 a=3.5 p=15
XM15 AMUXBUS_HV PG_AMX_VDDA_H_N 3 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.225 PD=7.28 PS=7.35 NRD=0 NRS=0.9359 m=1 sa=250001 sb=250002 a=3.5 p=15
XM16 3 PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=1.225 AS=0.98 PD=7.35 PS=7.28 NRD=0.9359 NRS=0 m=1 sa=250002 sb=250002 a=3.5 p=15
XM17 AMUXBUS_HV PG_AMX_VDDA_H_N 3 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.225 PD=7.28 PS=7.35 NRD=0 NRS=0.9359 m=1 sa=250003 sb=250001 a=3.5 p=15
XM18 3 PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=2.205 AS=0.98 PD=14.63 PS=7.28 NRD=0.9359 NRS=0 m=1 sa=250003 sb=250000 a=3.5 p=15
X19 3 VDDA condiode a=1e-06 p=0.004 m=1
X20 6 VDDA condiode a=1e-06 p=0.004 m=1
X21 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw a=64.774 p=32.54 m=1
X22 VSSD VDDA sky130_fd_pr__model__parasitic__diode_ps2nw a=66.495 p=33.14 m=1
X23 3 VDDA sky130_fd_pr__model__parasitic__diode_pw2dn a=141.419 p=48.37 m=1
X24 6 VDDA sky130_fd_pr__model__parasitic__diode_pw2dn a=144.747 p=49.61 m=1
X30 3 NG_AMX_VPMP_H AMUXBUS_HV AMUXBUS_HV 3 sky130_fd_pr__nfet_01v8__example_55959141808560
X31 3 NG_PAD_VPMP_H PAD_HV_N0 PAD_HV_N1 3 sky130_fd_pr__nfet_01v8__example_55959141808560
X32 6 NG_AMX_VPMP_H 6 6 AMUXBUS_HV sky130_fd_pr__nfet_01v8__example_55959141808560
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls VGND VPWR_HV IN_B RST_H IN HLD_H_N OUT_H VPWR_LV OUT_H_N 10 11
**
XM0 10 IN_B VGND VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=75000.2 sb=75001.5 a=0.15 p=2.3
XM1 VGND IN_B 10 VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75000.6 sb=75001 a=0.15 p=2.3
XM2 11 IN VGND VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001 sb=75000.6 a=0.15 p=2.3
XM3 VGND IN 11 VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.5 sb=75000.2 a=0.15 p=2.3
XM4 VGND RST_H OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=0.75 p=4
XM5 OUT_H RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=0.75 p=4
XM6 19 HLD_H_N OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=0.75 p=4
XM7 OUT_H HLD_H_N 19 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=0.75 p=4
XM8 OUT_H_N HLD_H_N 18 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.75 p=4
XM9 18 HLD_H_N OUT_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.75 p=4
XM10 19 VPWR_LV 10 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=450000 sb=450001 a=0.9 p=3.8
XM11 10 VPWR_LV 19 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=450001 sb=450000 a=0.9 p=3.8
XM12 11 VPWR_LV 18 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=450000 sb=450001 a=0.9 p=3.8
XM13 18 VPWR_LV 11 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=450001 sb=450000 a=0.9 p=3.8
XM14 VPWR_HV OUT_H OUT_H_N VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM15 OUT_H OUT_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.42 p=2.6
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808568 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
.ENDS
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808567 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.5 p=3
XM1 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.5 p=3
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_drvr VSSD VSSA VDDA VSWITCH VCCD VDDIO_Q 9 10 11 12 13 14 AMUX_EN_VDDA_H_N 16 AMUX_EN_VDDA_H 18 AMUX_EN_VDDIO_H_N 20 21 PD_CSD_VSWITCH_H
+ PU_CSD_VDDIOQ_H_N PGA_AMX_VDDA_H_N PGB_AMX_VDDA_H_N PD_CSD_VSWITCH_H_N NGA_PAD_VSWITCH_H NGA_PAD_VSWITCH_H_N AMUX_EN_VSWITCH_H NGA_AMX_VSWITCH_H NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N D_B 35 36 NMIDA_ON_N NMIDA_VCCD NMIDA_VCCD_N AMUX_EN_VDDIO_H 41 42
+ 43 44 45 46 47 PGA_PAD_VDDIOQ_H_N PGB_PAD_VDDIOQ_H_N AMUXBUSA_ON_N AMUX_EN_VSWITCH_H_N AMUXBUSB_ON_N AMUXBUSA_ON AMUXBUSB_ON PU_ON_N PU_ON PD_ON_N PD_ON
**
*.SEEDPROM
XM0 VSSA PD_CSD_VSWITCH_H PD_CSD_VSWITCH_H_N VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.375 p=2.5
XM1 NGA_PAD_VSWITCH_H_N NGA_PAD_VSWITCH_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.375 p=2.5
XM2 PD_CSD_VSWITCH_H 13 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.75 p=4
XM3 VSSA VSSA PD_CSD_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.75 p=4
XM4 69 14 9 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250004 a=1.5 p=7
XM5 9 14 69 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250003 a=1.5 p=7
XM6 VSSA 9 PGA_AMX_VDDA_H_N VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.5 p=3
XM7 69 14 9 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=1.5 p=7
XM8 9 AMUX_EN_VDDA_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.5 p=3
XM9 11 16 69 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=1.5 p=7
XM10 NGA_AMX_VSWITCH_H 41 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 sa=300000 sb=300006 a=0.252 p=2.04
XM11 69 16 11 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250003 sb=250001 a=1.5 p=7
XM12 VSSA AMUX_EN_VDDA_H_N NGA_AMX_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.5 p=3
XM13 VSSA 41 NGA_AMX_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300001 sb=300005 a=0.252 p=2.04
XM14 11 16 69 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250004 sb=250000 a=1.5 p=7
XM15 NGB_AMX_VSWITCH_H AMUX_EN_VDDA_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.5 p=3
XM16 NGB_AMX_VSWITCH_H 43 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300002 sb=300004 a=0.252 p=2.04
XM17 VSSA 43 NGB_AMX_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300003 sb=300003 a=0.252 p=2.04
XM18 NGB_PAD_VSWITCH_H 43 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300003 sb=300003 a=0.252 p=2.04
XM19 VSSA AMUX_EN_VDDIO_H_N NGB_PAD_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.5 p=3
XM20 VSSA 43 NGB_PAD_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300004 sb=300002 a=0.252 p=2.04
XM21 NGA_PAD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.5 p=3
XM22 NGA_PAD_VSWITCH_H 41 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300005 sb=300001 a=0.252 p=2.04
XM23 70 18 12 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250004 a=1.5 p=7
XM24 VSSA 41 NGA_PAD_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 sa=300006 sb=300000 a=0.252 p=2.04
XM25 12 18 70 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250003 a=1.5 p=7
XM26 PD_CSD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.5 p=3
XM27 70 18 12 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=1.5 p=7
XM28 VSSA AMUX_EN_VDDA_H_N 10 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.5 p=3
XM29 10 20 70 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=1.5 p=7
XM30 PGB_AMX_VDDA_H_N 10 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.5 p=3
XM31 NGB_PAD_VSWITCH_H_N NGB_PAD_VSWITCH_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.375 p=2.5
XM32 70 20 10 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250003 sb=250001 a=1.5 p=7
XM33 10 20 70 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250004 sb=250000 a=1.5 p=7
XM34 VSSD 35 D_B VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300004 a=0.42 p=2.6
XM35 PGA_PAD_VDDIOQ_H_N 16 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 sa=300000 sb=300009 a=0.252 p=2.04
XM36 35 36 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.42 p=2.6
XM37 VSSD 16 PGA_PAD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300001 sb=300008 a=0.252 p=2.04
XM38 VSSD 36 35 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300003 a=0.42 p=2.6
XM39 PGB_PAD_VDDIOQ_H_N 18 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300002 sb=300007 a=0.252 p=2.04
XM40 NMIDA_VCCD NMIDA_ON_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300002 a=0.42 p=2.6
XM41 VSSD 18 PGB_PAD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300003 sb=300006 a=0.252 p=2.04
XM42 VSSD NMIDA_ON_N NMIDA_VCCD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.42 p=2.6
XM43 PU_CSD_VDDIOQ_H_N 21 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300003 sb=300005 a=0.252 p=2.04
XM44 NMIDA_VCCD_N NMIDA_VCCD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300004 sb=300000 a=0.42 p=2.6
XM45 VSSD 21 PU_CSD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300004 sb=300004 a=0.252 p=2.04
XM46 PU_CSD_VDDIOQ_H_N 21 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300005 sb=300003 a=0.252 p=2.04
XM47 VSSD 21 PU_CSD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300006 sb=300003 a=0.252 p=2.04
XM48 PU_CSD_VDDIOQ_H_N 21 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300007 sb=300002 a=0.252 p=2.04
XM49 VSSD 21 PU_CSD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=300008 sb=300001 a=0.252 p=2.04
XM50 PU_CSD_VDDIOQ_H_N 21 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 sa=300009 sb=300000 a=0.252 p=2.04
XM51 VSWITCH PD_CSD_VSWITCH_H PD_CSD_VSWITCH_H_N VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.75 p=4
XM52 NGA_PAD_VSWITCH_H_N NGA_PAD_VSWITCH_H VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.75 p=4
XM53 VDDA 11 9 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 sa=500000 sb=500001 a=0.42 p=2.84
XM54 VDDA 12 10 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 sa=500000 sb=500001 a=0.42 p=2.84
XM55 11 9 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 sa=500001 sb=500000 a=0.42 p=2.84
XM56 12 10 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 sa=500001 sb=500000 a=0.42 p=2.84
XM57 PD_CSD_VSWITCH_H 13 VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=2 W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 m=1 sa=999999 sb=1e+06 a=1.5 p=5.5
XM58 VSWITCH 13 PD_CSD_VSWITCH_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=2 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 m=1 sa=1e+06 sb=999999 a=1.5 p=5.5
XM59 NGA_AMX_VSWITCH_H 41 VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300006 a=0.6 p=3.2
XM60 VSWITCH 41 NGA_AMX_VSWITCH_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300005 a=0.6 p=3.2
XM61 NGB_AMX_VSWITCH_H 43 VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300004 a=0.6 p=3.2
XM62 VSWITCH 43 NGB_AMX_VSWITCH_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300003 a=0.6 p=3.2
XM63 NGB_PAD_VSWITCH_H 43 VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300003 a=0.6 p=3.2
XM64 VSWITCH 43 NGB_PAD_VSWITCH_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300002 a=0.6 p=3.2
XM65 NGA_PAD_VSWITCH_H 41 VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300005 sb=300001 a=0.6 p=3.2
XM66 VSWITCH 41 NGA_PAD_VSWITCH_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300006 sb=300000 a=0.6 p=3.2
XM67 NGB_PAD_VSWITCH_H_N NGB_PAD_VSWITCH_H VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.3975 PD=3.53 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.75 p=4
XM68 VCCD 35 D_B VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300004 a=0.6 p=3.2
XM69 VCCD 35 D_B VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300004 a=0.6 p=3.2
XM70 PGA_PAD_VDDIOQ_H_N 16 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300009 a=0.6 p=3.2
XM71 35 36 VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.6 p=3.2
XM72 35 36 VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.6 p=3.2
XM73 VDDIO_Q 16 PGA_PAD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300008 a=0.6 p=3.2
XM74 VCCD 36 35 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300003 a=0.6 p=3.2
XM75 VCCD 36 35 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300003 a=0.6 p=3.2
XM76 PGB_PAD_VDDIOQ_H_N 18 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300007 a=0.6 p=3.2
XM77 NMIDA_VCCD NMIDA_ON_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300002 a=0.6 p=3.2
XM78 NMIDA_VCCD NMIDA_ON_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300002 a=0.6 p=3.2
XM79 VDDIO_Q 18 PGB_PAD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300006 a=0.6 p=3.2
XM80 VCCD NMIDA_ON_N NMIDA_VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.6 p=3.2
XM81 VCCD NMIDA_ON_N NMIDA_VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.6 p=3.2
XM82 PU_CSD_VDDIOQ_H_N 21 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300005 a=0.6 p=3.2
XM83 NMIDA_VCCD_N NMIDA_VCCD VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300000 a=0.6 p=3.2
XM84 NMIDA_VCCD_N NMIDA_VCCD VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300000 a=0.6 p=3.2
XM85 VDDIO_Q 21 PU_CSD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300004 a=0.6 p=3.2
XM86 PU_CSD_VDDIOQ_H_N 21 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300005 sb=300003 a=0.6 p=3.2
XM87 VDDIO_Q 21 PU_CSD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300006 sb=300003 a=0.6 p=3.2
XM88 PU_CSD_VDDIOQ_H_N 21 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300007 sb=300002 a=0.6 p=3.2
XM89 VDDIO_Q 21 PU_CSD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300008 sb=300001 a=0.6 p=3.2
XM90 PU_CSD_VDDIOQ_H_N 21 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300009 sb=300000 a=0.6 p=3.2
X91 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=5.073 p=9.14 m=1
X92 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=23.245 p=25.57 m=1
X93 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=9.709 p=14.02 m=1
X94 VSSD VSWITCH sky130_fd_pr__model__parasitic__diode_ps2dn a=570.063 p=97.15 m=1
X95 VSSA VSWITCH sky130_fd_pr__model__parasitic__diode_pw2dn a=6.6852 p=10.51 m=1
X96 VSSA VSWITCH sky130_fd_pr__model__parasitic__diode_pw2dn a=51.6765 p=33.36 m=1
X97 VSSA VSWITCH sky130_fd_pr__model__parasitic__diode_pw2dn a=340.297 p=98.11 m=1
X98 VSSD VDDIO_Q AMUXBUSA_ON_N AMUX_EN_VDDIO_H_N AMUXBUSA_ON AMUX_EN_VDDIO_H 16 VCCD 14 71 72 sky130_fd_io__gpiov2_amux_drvr_ls
X99 VSSA VSWITCH AMUXBUSA_ON_N AMUX_EN_VSWITCH_H_N AMUXBUSA_ON AMUX_EN_VSWITCH_H 74 VCCD 41 42 73 sky130_fd_io__gpiov2_amux_drvr_ls
X100 VSSA VSWITCH AMUXBUSB_ON_N AMUX_EN_VSWITCH_H_N AMUXBUSB_ON AMUX_EN_VSWITCH_H 76 VCCD 43 44 75 sky130_fd_io__gpiov2_amux_drvr_ls
X101 VSSA VSWITCH PD_ON_N AMUX_EN_VSWITCH_H_N PD_ON AMUX_EN_VSWITCH_H 78 VCCD 13 45 77 sky130_fd_io__gpiov2_amux_drvr_ls
X102 VSSD VDDIO_Q AMUXBUSB_ON_N AMUX_EN_VDDIO_H_N AMUXBUSB_ON AMUX_EN_VDDIO_H 18 VCCD 20 46 79 sky130_fd_io__gpiov2_amux_drvr_ls
X103 VSSD VDDIO_Q PU_ON_N AMUX_EN_VDDIO_H_N PU_ON AMUX_EN_VDDIO_H 21 VCCD 80 47 81 sky130_fd_io__gpiov2_amux_drvr_ls
X129 VSSA AMUX_EN_VDDA_H 69 sky130_fd_pr__nfet_01v8__example_55959141808568
X130 VSSA AMUX_EN_VDDA_H 70 sky130_fd_pr__nfet_01v8__example_55959141808568
X139 VDDA 9 PGA_AMX_VDDA_H_N sky130_fd_pr__pfet_01v8__example_55959141808567
X140 VDDA 10 PGB_AMX_VDDA_H_N sky130_fd_pr__pfet_01v8__example_55959141808567
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808460 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.375 p=2.5
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_inv_1 VNB VPB IN VPWR OUT VGND
**
*.SEEDPROM
XM0 OUT IN VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 m=1 sa=75000.3 sb=75000.2 a=0.111 p=1.78
XM1 OUT IN VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=0.25 W=1 AD=0.295 AS=0.345 PD=2.59 PS=2.69 NRD=1.9503 NRS=11.8003 m=1 sa=125000 sb=125000 a=0.25 p=2.5
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808589 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
.ENDS
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_ls VSSA VSSD VSWITCH VDDA VDDIO_Q VCCD ENABLE_VDDA_H AMUX_EN_VDDIO_H 15 ENABLE_VSWITCH_H AMUX_EN_VDDIO_H_N 18 19 20 21 HLD_I_H_N HLD_I_H AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H AMUX_EN_VSWITCH_H_N
+ AMUX_EN_VSWITCH_H ANALOG_EN
**
*.SEEDPROM
XM0 35 32 34 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=75000.2 sb=75003.2 a=0.15 p=2.3
XM1 34 32 35 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75000.6 sb=75002.8 a=0.15 p=2.3
XM2 35 32 34 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001 sb=75002.3 a=0.15 p=2.3
XM3 34 32 35 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.5 sb=75001.9 a=0.15 p=2.3
XM4 36 33 34 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.9 sb=75001.5 a=0.15 p=2.3
XM5 34 33 36 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.3 sb=75001 a=0.15 p=2.3
XM6 36 33 34 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.8 sb=75000.6 a=0.15 p=2.3
XM7 34 33 36 VSSD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=75003.2 sb=75000.2 a=0.15 p=2.3
XM8 37 AMUX_EN_VDDIO_H 29 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250004 a=1.5 p=7
XM9 18 ENABLE_VDDA_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.5 p=3
XM10 VSSA ENABLE_VSWITCH_H 21 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.1855 PD=1.93 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.42 p=2.6
XM11 29 AMUX_EN_VDDIO_H 37 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250003 a=1.5 p=7
XM12 VSSA 15 AMUX_EN_VDDA_H_N VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.5 p=3
XM13 37 AMUX_EN_VDDIO_H 29 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=1.5 p=7
XM14 AMUX_EN_VDDA_H 29 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.5 p=3
XM15 15 AMUX_EN_VDDIO_H_N 37 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=1.5 p=7
XM16 37 AMUX_EN_VDDIO_H_N 15 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250003 sb=250001 a=1.5 p=7
XM17 15 18 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.5 p=3
XM18 15 AMUX_EN_VDDIO_H_N 37 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250004 sb=250000 a=1.5 p=7
XM19 VSSA 20 AMUX_EN_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.5 p=3
XM20 VSSA 19 AMUX_EN_VSWITCH_H_N VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.5 p=3
XM21 19 21 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.5 p=3
XM22 38 AMUX_EN_VDDIO_H 20 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250004 a=1.5 p=7
XM23 20 AMUX_EN_VDDIO_H 38 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250003 a=1.5 p=7
XM24 38 AMUX_EN_VDDIO_H 20 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=1.5 p=7
XM25 19 AMUX_EN_VDDIO_H_N 38 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=1.5 p=7
XM26 38 AMUX_EN_VDDIO_H_N 19 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250003 sb=250001 a=1.5 p=7
XM27 19 AMUX_EN_VDDIO_H_N 38 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250004 sb=250000 a=1.5 p=7
XM28 34 HLD_I_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=0.5 p=3
XM29 VSSD HLD_I_H_N 34 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=0.5 p=3
XM30 34 HLD_I_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=0.5 p=3
XM31 VSSD HLD_I_H_N 34 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=0.5 p=3
XM32 VSSD 31 AMUX_EN_VDDIO_H VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.5 p=3
XM33 30 HLD_I_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.5 p=3
XM34 AMUX_EN_VDDIO_H_N 30 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.5 p=3
XM35 30 VCCD 36 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=450000 sb=450003 a=0.9 p=3.8
XM36 31 VCCD 35 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=450000 sb=450003 a=0.9 p=3.8
XM37 36 VCCD 30 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=450001 sb=450002 a=0.9 p=3.8
XM38 35 VCCD 31 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=450001 sb=450002 a=0.9 p=3.8
XM39 30 VCCD 36 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=450002 sb=450001 a=0.9 p=3.8
XM40 31 VCCD 35 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=450002 sb=450001 a=0.9 p=3.8
XM41 36 VCCD 30 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=450003 sb=450000 a=0.9 p=3.8
XM42 35 VCCD 31 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=450003 sb=450000 a=0.9 p=3.8
XM43 18 ENABLE_VDDA_H VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.75 p=4
XM44 VDDA ENABLE_VDDA_H 18 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.75 p=4
XM45 21 ENABLE_VSWITCH_H VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM46 VDDA 15 AMUX_EN_VDDA_H_N VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.75 p=4
XM47 VSWITCH ENABLE_VSWITCH_H 21 VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM48 AMUX_EN_VDDA_H 29 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.75 p=4
XM49 VSWITCH 19 20 VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 sa=500000 sb=500001 a=0.42 p=2.84
XM50 VDDA 15 29 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 sa=500000 sb=500001 a=0.42 p=2.84
XM51 19 20 VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 sa=500001 sb=500000 a=0.42 p=2.84
XM52 15 29 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 sa=500001 sb=500000 a=0.42 p=2.84
XM53 VSWITCH 19 AMUX_EN_VSWITCH_H_N VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.75 p=4
XM54 AMUX_EN_VSWITCH_H 20 VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.75 p=4
XM55 VDDIO_Q 30 AMUX_EN_VDDIO_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.75 p=4
XM56 AMUX_EN_VDDIO_H 31 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.75 p=4
X57 VSSD VCCD sky130_fd_pr__model__parasitic__diode_ps2nw a=7.1653 p=11.43 m=1
X58 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=12.2407 p=15.81 m=1
X77 VDDIO_Q 31 30 sky130_fd_pr__pfet_01v8__example_55959141808460
X78 VDDIO_Q 30 31 sky130_fd_pr__pfet_01v8__example_55959141808460
X79 VSSD VCCD 33 VCCD 32 VSSD sky130_fd_io__gpiov2_amux_ctl_inv_1
X80 VSSD VCCD ANALOG_EN VCCD 33 VSSD sky130_fd_io__gpiov2_amux_ctl_inv_1
X84 VSSA ENABLE_VDDA_H 37 sky130_fd_pr__nfet_01v8__example_55959141808589
X85 VSSA ENABLE_VSWITCH_H 38 sky130_fd_pr__nfet_01v8__example_55959141808589
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_nand5 VGND VPWR OUT IN0 IN4 IN3 IN2 IN1
**
*.SEEDPROM
XM0 VGND 13 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 AD=0.101634 AS=0.1113 PD=0.7875 PS=1.37 NRD=24.4188 NRS=0 m=1 sa=250000 sb=250004 a=0.21 p=1.84
XM1 VGND OUT 13 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 AD=0.101634 AS=0.1113 PD=0.7875 PS=1.37 NRD=25.1028 NRS=0 m=1 sa=250000 sb=250004 a=0.21 p=1.84
XM2 14 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.20993 PD=5.28 PS=9.375 NRD=0 NRS=0 m=1 sa=250000 sb=250003 a=2.5 p=11
XM3 15 IN4 14 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=2.5 p=11
XM4 16 IN3 15 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=2.5 p=11
XM5 17 IN2 16 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250001 a=2.5 p=11
XM6 OUT IN1 17 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250000 a=2.5 p=11
XM7 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM8 VPWR IN0 OUT VPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM9 13 OUT VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM10 VPWR OUT 13 VPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.217676 AS=0.14 PD=1.92958 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM11 OUT 13 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 AD=0.1113 AS=0.0914239 PD=1.37 PS=0.810423 NRD=0 NRS=42.0582 m=1 sa=250004 sb=250000 a=0.21 p=1.84
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_nand4 VGND IN0 OUT IN3 IN2 IN1 15
**
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VPWR
XM0 VGND 15 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 AD=0.101634 AS=0.1113 PD=0.7875 PS=1.37 NRD=24.4188 NRS=0 m=1 sa=250000 sb=250003 a=0.21 p=1.84
XM1 VGND OUT 15 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 AD=0.101634 AS=0.1113 PD=0.7875 PS=1.37 NRD=25.1028 NRS=0 m=1 sa=250000 sb=250003 a=0.21 p=1.84
XM2 16 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.20993 PD=5.28 PS=9.375 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=2.5 p=11
XM3 17 IN3 16 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=2.5 p=11
XM4 18 IN2 17 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=2.5 p=11
XM5 OUT IN1 18 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250000 a=2.5 p=11
.ENDS
***************************************
.SUBCKT sky130_fd_io__inv_1 VNB VPB A VPWR Y VGND
**
*.SEEDPROM
XM0 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 m=1 sa=75000.3 sb=75000.2 a=0.111 p=1.78
XM1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.12 AD=0.3304 AS=0.3864 PD=2.83 PS=2.93 NRD=1.7533 NRS=10.5395 m=1 sa=75000.3 sb=75000.2 a=0.168 p=2.54
.ENDS
***************************************
.SUBCKT sky130_fd_io__nand2_1 VNB VPB B A VPWR Y VGND
**
*.SEEDPROM
XM0 8 B VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 m=1 sa=75000.2 sb=75000.6 a=0.111 p=1.78
XM1 Y A 8 VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 AD=0.2109 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 m=1 sa=75000.6 sb=75000.2 a=0.111 p=1.78
XM2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.12 AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 m=1 sa=75000.2 sb=75000.7 a=0.168 p=2.54
XM3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.12 AD=0.3192 AS=0.168 PD=2.81 PS=1.42 NRD=1.7533 NRS=1.7533 m=1 sa=75000.7 sb=75000.2 a=0.168 p=2.54
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__nor2_1 VNB VPB A B VPWR Y VGND
**
*.SEEDPROM
XM0 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 m=1 sa=75000.2 sb=75000.6 a=0.111 p=1.78
XM1 VGND B Y VNB sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 m=1 sa=75000.6 sb=75000.2 a=0.111 p=1.78
XM2 8 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.12 AD=0.1512 AS=0.3304 PD=1.39 PS=2.83 NRD=14.0658 NRS=1.7533 m=1 sa=75000.2 sb=75000.6 a=0.168 p=2.54
XM3 Y B 8 VPB sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.12 AD=0.3304 AS=0.1512 PD=2.83 PS=1.39 NRD=1.7533 NRS=14.0658 m=1 sa=75000.6 sb=75000.2 a=0.168 p=2.54
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_decoder VSSD VCCD 5 6 7 ANALOG_SEL 9 10 11 12 AMUXBUSA_ON_N AMUXBUSA_ON 15 PU_ON_N 17 NMIDA_ON_N PU_ON 20 ANALOG_EN D_B
+ 23 PD_ON AMUXBUSB_ON_N PGA_AMX_VDDA_H_N 27 AMUXBUSB_ON PD_ON_N PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N 32 33 PGB_PAD_VDDIOQ_H_N NGA_PAD_VSWITCH_H 36 OUT ANALOG_POL NGB_PAD_VSWITCH_H 40 41 NGB_PAD_VSWITCH_H_N
+ NGA_PAD_VSWITCH_H_N PU_VDDIOQ_H_N PD_VSWITCH_H_N 46 NMIDA_VCCD_N
**
*.SEEDPROM
XM0 48 5 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 m=1 sa=75000.2 sb=75002.5 a=0.126 p=1.98
XM1 VSSD 6 48 VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 m=1 sa=75000.6 sb=75002 a=0.126 p=1.98
XM2 51 6 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 AD=0.1008 AS=0.1176 PD=1.08 PS=1.12 NRD=9.276 NRS=0 m=1 sa=75001.1 sb=75001.6 a=0.126 p=1.98
XM3 7 5 51 VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 AD=0.2436 AS=0.1008 PD=1.42 PS=1.08 NRD=27.132 NRS=9.276 m=1 sa=75001.4 sb=75001.2 a=0.126 p=1.98
XM4 VSSD 48 7 VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 AD=0.4788 AS=0.2436 PD=2.82 PS=1.42 NRD=43.56 NRS=15.708 m=1 sa=75002.2 sb=75000.5 a=0.126 p=1.98
XM5 252 17 NMIDA_ON_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300003 a=0.42 p=2.6
XM6 VSSD 20 252 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300002 a=0.42 p=2.6
XM7 253 12 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=13.8396 NRS=0 m=1 sa=300002 sb=300001 a=0.42 p=2.6
XM8 D_B 23 253 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300003 sb=300000 a=0.42 p=2.6
XM9 254 PGA_AMX_VDDA_H_N 27 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM10 VSSD PGA_PAD_VDDIOQ_H_N 254 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM11 255 PGB_AMX_VDDA_H_N 32 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM12 VSSD PGB_PAD_VDDIOQ_H_N 255 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM13 17 NGA_PAD_VSWITCH_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM14 VSSD 27 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.196 AS=0.098 PD=1.96 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM15 23 32 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.196 PD=0.98 PS=1.96 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM16 VSSD NGB_PAD_VSWITCH_H 23 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM17 49 5 48 VCCD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.26 AD=0.1512 AS=0.3339 PD=1.5 PS=3.05 NRD=10.1455 NRS=0 m=1 sa=75000.2 sb=75001.6 a=0.189 p=2.82
XM18 VCCD 6 49 VCCD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.26 AD=0.189 AS=0.1512 PD=1.56 PS=1.5 NRD=0 NRS=10.1455 m=1 sa=75000.6 sb=75001.2 a=0.189 p=2.82
XM19 50 6 VCCD VCCD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.26 AD=0.1764 AS=0.189 PD=1.54 PS=1.56 NRD=0 NRS=3.1126 m=1 sa=75001 sb=75000.7 a=0.189 p=2.82
XM20 VCCD 5 50 VCCD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.26 AD=0.4786 AS=0.1764 PD=3.44 PS=1.54 NRD=15.6221 NRS=0 m=1 sa=75001.5 sb=75000.3 a=0.189 p=2.82
XM21 50 48 7 VCCD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.26 AD=0.3339 AS=0.3591 PD=3.05 PS=3.09 NRD=0 NRS=0 m=1 sa=75000.2 sb=75000.2 a=0.189 p=2.82
XM22 NMIDA_ON_N 17 VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM23 NMIDA_ON_N 17 VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM24 VCCD 20 NMIDA_ON_N VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM25 VCCD 20 NMIDA_ON_N VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM26 D_B 12 VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM27 D_B 12 VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM28 VCCD 23 D_B VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM29 VCCD 23 D_B VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM30 27 PGA_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM31 27 PGA_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM32 VCCD PGA_PAD_VDDIOQ_H_N 27 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM33 VCCD PGA_PAD_VDDIOQ_H_N 27 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM34 32 PGB_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM35 32 PGB_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM36 VCCD PGB_PAD_VDDIOQ_H_N 32 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM37 VCCD PGB_PAD_VDDIOQ_H_N 32 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM38 250 NGA_PAD_VSWITCH_H VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM39 250 NGA_PAD_VSWITCH_H VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM40 17 27 250 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM41 17 27 250 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM42 251 32 23 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM43 251 32 23 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM44 VCCD NGB_PAD_VSWITCH_H 251 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM45 VCCD NGB_PAD_VSWITCH_H 251 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM46 VCCD 248 AMUXBUSB_ON_N VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 AD=0.0914239 AS=0.1113 PD=0.810423 PS=1.37 NRD=42.0582 NRS=0 m=1 sa=250000 sb=250008 a=0.21 p=1.84
XM47 248 AMUXBUSB_ON_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.217676 PD=1.28 PS=1.92958 NRD=0 NRS=0 m=1 sa=300000 sb=300006 a=0.6 p=3.2
XM48 VCCD AMUXBUSB_ON_N 248 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300006 a=0.6 p=3.2
XM49 AMUXBUSB_ON_N 10 VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300005 a=0.6 p=3.2
XM50 VCCD 10 AMUXBUSB_ON_N VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300004 a=0.6 p=3.2
XM51 AMUXBUSA_ON_N 33 VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300003 a=0.6 p=3.2
XM52 VCCD 33 AMUXBUSA_ON_N VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300005 sb=300002 a=0.6 p=3.2
XM53 249 AMUXBUSA_ON_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300006 sb=300001 a=0.6 p=3.2
XM54 VCCD AMUXBUSA_ON_N 249 VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.217676 AS=0.14 PD=1.92958 PS=1.28 NRD=0 NRS=0 m=1 sa=300006 sb=300000 a=0.6 p=3.2
XM55 AMUXBUSA_ON_N 249 VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 AD=0.1113 AS=0.0914239 PD=1.37 PS=0.810423 NRD=0 NRS=42.0582 m=1 sa=250008 sb=250000 a=0.21 p=1.84
X56 VSSD VCCD sky130_fd_pr__model__parasitic__diode_ps2nw a=65.448 p=49.72 m=1
X57 VSSD VCCD sky130_fd_pr__model__parasitic__diode_ps2nw a=50.2164 p=38.54 m=1
X61 VSSD VCCD 40 41 NGB_PAD_VSWITCH_H_N NGA_PAD_VSWITCH_H_N PGB_PAD_VDDIOQ_H_N PGA_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_nand5
X62 VSSD VCCD 57 15 NGB_PAD_VSWITCH_H_N NGA_PAD_VSWITCH_H_N PGB_PAD_VDDIOQ_H_N PGA_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_nand5
X63 VSSD 10 AMUXBUSB_ON_N 46 PD_VSWITCH_H_N PU_VDDIOQ_H_N 248 sky130_fd_io__gpiov2_amux_nand4
X64 VSSD 33 AMUXBUSA_ON_N NMIDA_VCCD_N PD_VSWITCH_H_N PU_VDDIOQ_H_N 249 sky130_fd_io__gpiov2_amux_nand4
X65 VSSD VCCD ANALOG_SEL VCCD 52 VSSD sky130_fd_io__inv_1
X66 VSSD VCCD 52 VCCD 9 VSSD sky130_fd_io__inv_1
X67 VSSD VCCD 10 VCCD 12 VSSD sky130_fd_io__inv_1
X68 VSSD VCCD AMUXBUSA_ON_N VCCD AMUXBUSA_ON VSSD sky130_fd_io__inv_1
X69 VSSD VCCD PU_ON VCCD PU_ON_N VSSD sky130_fd_io__inv_1
X70 VSSD VCCD ANALOG_EN VCCD 53 VSSD sky130_fd_io__inv_1
X71 VSSD VCCD PD_ON VCCD PD_ON_N VSSD sky130_fd_io__inv_1
X72 VSSD VCCD AMUXBUSB_ON_N VCCD AMUXBUSB_ON VSSD sky130_fd_io__inv_1
X73 VSSD VCCD 57 VCCD PU_ON VSSD sky130_fd_io__inv_1
X74 VSSD VCCD 33 VCCD 20 VSSD sky130_fd_io__inv_1
X75 VSSD VCCD 36 VCCD 5 VSSD sky130_fd_io__inv_1
X76 VSSD VCCD 58 VCCD 6 VSSD sky130_fd_io__inv_1
X77 VSSD VCCD OUT VCCD 36 VSSD sky130_fd_io__inv_1
X78 VSSD VCCD ANALOG_POL VCCD 58 VSSD sky130_fd_io__inv_1
X79 VSSD VCCD 40 VCCD PD_ON VSSD sky130_fd_io__inv_1
X80 VSSD VCCD 7 52 VCCD 11 VSSD sky130_fd_io__nand2_1
X81 VSSD VCCD 9 7 VCCD 54 VSSD sky130_fd_io__nand2_1
X82 VSSD VCCD 5 6 VCCD 55 VSSD sky130_fd_io__nand2_1
X83 VSSD VCCD 36 58 VCCD 56 VSSD sky130_fd_io__nand2_1
X90 VSSD VCCD 53 54 VCCD 10 VSSD sky130_fd_io__nor2_1
X91 VSSD VCCD 53 55 VCCD 15 VSSD sky130_fd_io__nor2_1
X92 VSSD VCCD 53 56 VCCD 41 VSSD sky130_fd_io__nor2_1
X93 VSSD VCCD 53 11 VCCD 33 VSSD sky130_fd_io__nor2_1
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_logic VSSD VSSA VDDA VSWITCH VCCD 12 13 14 15 VDDIO_Q 17 PGA_AMX_VDDA_H_N NGB_PAD_VSWITCH_H NGA_PAD_VSWITCH_H AMUX_EN_VDDA_H_N PGB_AMX_VDDA_H_N 23 24 D_B 26
+ NMIDA_VCCD 28 ENABLE_VDDA_H ENABLE_VSWITCH_H 31 AMUX_EN_VDDIO_H_N 33 34 35 36 37 PGB_PAD_VDDIOQ_H_N 39 40 41 42 PGA_PAD_VDDIOQ_H_N 44 45 46
+ 47 48 49 50 51 52 PD_CSD_VSWITCH_H 54 55 56 NGA_AMX_VSWITCH_H NGB_AMX_VSWITCH_H 59 60 61 62 PU_CSD_VDDIOQ_H_N 64 65 66
+ ANALOG_EN HLD_I_H_N HLD_I_H ANALOG_SEL 71 72 73 74 75 76 77 78 79 OUT ANALOG_POL 82 83 84 85 86
**
X0 VSSD VSWITCH sky130_fd_pr__model__parasitic__diode_ps2nw a=2.8569 p=0 m=1
X1 VSSD VDDA sky130_fd_pr__model__parasitic__diode_ps2nw a=43.3597 p=31.46 m=1
X2 VSSD VCCD sky130_fd_pr__model__parasitic__diode_ps2nw a=70.2614 p=46.74 m=1
X3 VSSD VSSA VDDA VSWITCH VCCD VDDIO_Q 54 52 56 51 55 14 AMUX_EN_VDDA_H_N 17 89 61 AMUX_EN_VDDIO_H_N 62 65 PD_CSD_VSWITCH_H
+ PU_CSD_VDDIOQ_H_N PGA_AMX_VDDA_H_N PGB_AMX_VDDA_H_N 13 NGA_PAD_VSWITCH_H 39 34 NGA_AMX_VSWITCH_H NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H 23 24 D_B 12 26 NMIDA_VCCD 44 15 60 49
+ 84 50 59 64 66 PGA_PAD_VDDIOQ_H_N PGB_PAD_VDDIOQ_H_N 42 33 46 41 40 47 48 37 36
+ sky130_fd_io__gpiov2_amux_drvr
X4 VSSA VSSD VSWITCH VDDA VDDIO_Q VCCD ENABLE_VDDA_H 15 31 ENABLE_VSWITCH_H AMUX_EN_VDDIO_H_N 28 91 90 88 HLD_I_H_N HLD_I_H AMUX_EN_VDDA_H_N 89 33
+ 34 ANALOG_EN
+ sky130_fd_io__gpiov2_amux_ls
X5 VSSD VCCD 85 72 74 ANALOG_SEL 71 83 92 76 42 41 35 47 73 26 48 75 ANALOG_EN 12
+ 77 36 46 PGA_AMX_VDDA_H_N 78 40 37 PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N 79 45 PGB_PAD_VDDIOQ_H_N NGA_PAD_VSWITCH_H 86 OUT ANALOG_POL NGB_PAD_VSWITCH_H 82 87 23
+ 39 PU_CSD_VDDIOQ_H_N 13 24 44
+ sky130_fd_io__gpiov2_amux_decoder
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_amux VSSD VSSA VSSIO_Q 4 5 6 7 VSWITCH VDDIO_Q VDDA HLD_I_H PAD ENABLE_VDDA_H VCCD 16 ENABLE_VSWITCH_H AMUXBUS_B AMUXBUS_A ANALOG_SEL ANALOG_EN
+ OUT ANALOG_POL HLD_I_H_N
**
XM0 36 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 sa=250000 sb=250010 a=2.5 p=11
XM1 VSSIO_Q 27 36 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250009 a=2.5 p=11
XM2 36 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250009 a=2.5 p=11
XM3 VSSIO_Q 27 36 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250008 a=2.5 p=11
XM4 36 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250007 a=2.5 p=11
XM5 VSSIO_Q 27 36 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250004 sb=250006 a=2.5 p=11
XM6 37 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250005 a=2.5 p=11
XM7 VSSIO_Q 27 37 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250005 a=2.5 p=11
XM8 37 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250006 sb=250004 a=2.5 p=11
XM9 VSSIO_Q 27 37 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250007 sb=250003 a=2.5 p=11
XM10 37 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250008 sb=250002 a=2.5 p=11
XM11 VSSIO_Q 27 37 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250009 sb=250002 a=2.5 p=11
XM12 37 27 VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250009 sb=250001 a=2.5 p=11
XM13 VSSIO_Q 27 37 VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 sa=250010 sb=250000 a=2.5 p=11
XM14 37 25 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 AD=2.1 AS=4.2 PD=15.28 PS=30.56 NRD=0 NRS=0 m=1 sa=250000 sb=250005 a=7.5 p=31
XM15 VDDIO_Q 25 37 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 AD=2.1 AS=2.1 PD=15.28 PS=15.28 NRD=0 NRS=0 m=1 sa=250001 sb=250004 a=7.5 p=31
XM16 37 25 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 AD=2.1 AS=2.1 PD=15.28 PS=15.28 NRD=0 NRS=0 m=1 sa=250002 sb=250003 a=7.5 p=31
XM17 VDDIO_Q 25 37 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 AD=2.1 AS=2.1 PD=15.28 PS=15.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=7.5 p=31
XM18 36 25 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 AD=2.1 AS=2.1 PD=15.28 PS=15.28 NRD=0 NRS=0 m=1 sa=250003 sb=250002 a=7.5 p=31
XM19 VDDIO_Q 25 36 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 AD=2.1 AS=2.1 PD=15.28 PS=15.28 NRD=0 NRS=0 m=1 sa=250004 sb=250001 a=7.5 p=31
XM20 36 25 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 AD=4.2 AS=2.1 PD=30.56 PS=15.28 NRD=0 NRS=0 m=1 sa=250005 sb=250000 a=7.5 p=31
X21 VSSA VSWITCH condiode a=1e-06 p=0.004 m=1
X22 VSSA VSWITCH condiode a=1e-06 p=0.004 m=1
X23 VSSA VSWITCH condiode a=1e-06 p=0.004 m=1
X24 VSSIO_Q VDDA condiode a=1e-06 p=0.004 m=1
X25 VSSA VDDA condiode a=1e-06 p=0.004 m=1
X26 VSSIO_Q VDDA condiode a=1e-06 p=0.004 m=1
X27 VSSD VDDA sky130_fd_pr__model__parasitic__diode_ps2nw a=0.10455 p=0 m=1
X28 VSSD VDDA sky130_fd_pr__model__parasitic__diode_ps2nw a=0.10455 p=0 m=1
X29 VSSD VDDA sky130_fd_pr__model__parasitic__diode_ps2nw a=1.79917 p=0 m=1
X30 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=126.767 p=49.03 m=1
X31 VSSD VDDA sky130_fd_pr__model__parasitic__diode_ps2dn a=946.67 p=155.39 m=1
X32 VSSIO_Q VDDA sky130_fd_pr__model__parasitic__diode_pw2dn a=96.7472 p=41.01 m=1
X33 VSSA VDDA sky130_fd_pr__model__parasitic__diode_pw2dn a=48.208 p=27.82 m=1
X34 VSSA 28 7 VSSA sky130_fd_pr__nfet_01v8__example_55959141808592
X35 VSSA 28 5 VSSA sky130_fd_pr__nfet_01v8__example_55959141808592
X36 VSSA 28 VSSA 4 sky130_fd_pr__nfet_01v8__example_55959141808592
X37 VSSA 28 VSSA 6 sky130_fd_pr__nfet_01v8__example_55959141808592
X38 VSSA HLD_I_H 4 VSSA sky130_fd_pr__nfet_01v8__example_55959141808592
X39 VSSA HLD_I_H 6 VSSA sky130_fd_pr__nfet_01v8__example_55959141808592
X40 VSSA HLD_I_H VSSA 7 sky130_fd_pr__nfet_01v8__example_55959141808592
X41 VSSA HLD_I_H VSSA 5 sky130_fd_pr__nfet_01v8__example_55959141808592
X42 VSSA 26 41 5 sky130_fd_pr__nfet_01v8__example_55959141808593
X43 VSSA 26 39 6 sky130_fd_pr__nfet_01v8__example_55959141808593
X44 VSSA 29 4 40 sky130_fd_pr__nfet_01v8__example_55959141808593
X45 VSSA 29 38 7 sky130_fd_pr__nfet_01v8__example_55959141808593
X54 PAD 30 sky130_fd_io__res75only_small
X55 31 32 sky130_fd_io__res75only_small
X56 PAD PAD sky130_fd_io__res75only_small
X57 PAD 31 sky130_fd_io__res75only_small
X58 PAD 33 sky130_fd_io__res75only_small
X59 PAD PAD sky130_fd_io__res75only_small
X60 33 34 sky130_fd_io__res75only_small
X61 PAD 35 sky130_fd_io__res75only_small
X62 PAD 36 sky130_fd_io__res75only_small
X63 PAD 37 sky130_fd_io__res75only_small
X64 VSSA 38 sky130_fd_io__res75only_small
X65 VSSA 39 sky130_fd_io__res75only_small
X66 VSSA 40 sky130_fd_io__res75only_small
X67 VSSA 41 sky130_fd_io__res75only_small
X68 VSSD 5 6 VDDIO_Q VDDA 77 16 65 45 30 35 AMUXBUS_B 32 32 34 34 sky130_fd_io__amux_switch_1v2b
X69 VSSD 4 7 VDDIO_Q VDDA 73 57 64 46 30 35 AMUXBUS_A 32 32 34 34 sky130_fd_io__amux_switch_1v2b
X78 VSSD VSSA VDDA VSWITCH VCCD 75 72 42 43 VDDIO_Q 44 57 45 46 47 16 99 48 26 78
+ 29 28 ENABLE_VDDA_H ENABLE_VSWITCH_H 52 68 51 58 80 67 89 77 74 54 53 49 73 81 96 50
+ 79 97 55 56 59 60 27 61 62 63 64 65 66 69 70 71 25 90 92 95
+ ANALOG_EN HLD_I_H_N HLD_I_H ANALOG_SEL 76 82 83 84 85 86 87 88 91 OUT ANALOG_POL 93 94 98 100 101
+ sky130_fd_io__gpiov2_amux_ctl_logic
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em2s_cdns_55959141808438 2 3
**
R0 2 6 0.01 short m=1
R1 6 3 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1o_cdns_5595914180880 4
**
*.SEEDPROM
R0 7 4 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1s_cdns_5595914180882 1 2
**
R0 1 5 0.01 short m=1
R1 5 2 0.01 short m=1
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808430 2 3 4 5 6
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_01v8_hvt L=0.25 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=0.25 p=2.5
XM1 6 4 5 2 sky130_fd_pr__pfet_01v8_hvt L=0.25 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=0.25 p=2.5
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808623 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 m=1 sa=500000 sb=500000 a=0.75 p=3.5
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_5595914180822 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.375 p=2.5
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_ctl_lsv2 VGND VCC_IO VPWR HLD_H_N SET_H RST_H IN OUT_H OUT_H_N
**
*.SEEDPROM
XM0 VGND IN 12 VGND sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=0.25 p=2.5
XM1 13 12 VGND VGND sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=0.25 p=2.5
XM2 14 12 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=75000.2 sb=75003.2 a=0.15 p=2.3
XM3 VGND 12 14 VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75000.6 sb=75002.8 a=0.15 p=2.3
XM4 14 12 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001 sb=75002.3 a=0.15 p=2.3
XM5 VGND 12 14 VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.5 sb=75001.9 a=0.15 p=2.3
XM6 17 13 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.9 sb=75001.5 a=0.15 p=2.3
XM7 VGND 13 17 VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.3 sb=75001 a=0.15 p=2.3
XM8 17 13 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.8 sb=75000.6 a=0.15 p=2.3
XM9 VGND 13 17 VGND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=75003.2 sb=75000.2 a=0.15 p=2.3
XM10 VGND 10 OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM11 OUT_H_N 11 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM12 10 HLD_H_N 15 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=1.8 p=7.2
XM13 VGND SET_H 10 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=1.8 p=7.2
XM14 11 RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=1.8 p=7.2
XM15 16 HLD_H_N 11 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=1.8 p=7.2
XM16 16 VPWR 14 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=450000 sb=450002 a=0.9 p=3.8
XM17 17 VPWR 15 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=450000 sb=450003 a=0.9 p=3.8
XM18 14 VPWR 16 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=450001 sb=450001 a=0.9 p=3.8
XM19 15 VPWR 17 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=450001 sb=450002 a=0.9 p=3.8
XM20 16 VPWR 14 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=450002 sb=450000 a=0.9 p=3.8
XM21 17 VPWR 15 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=450002 sb=450001 a=0.9 p=3.8
XM22 16 VPWR 14 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=450000 sb=450000 a=0.9 p=3.8
XM23 15 VPWR 17 VGND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=450003 sb=450000 a=0.9 p=3.8
XM24 VCC_IO 11 OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM25 OUT_H 10 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
X28 VPWR IN 12 VPWR 13 sky130_fd_pr__pfet_01v8__example_55959141808430
X39 VGND 11 10 sky130_fd_pr__nfet_01v8__example_55959141808623
X40 VGND 10 11 sky130_fd_pr__nfet_01v8__example_55959141808623
X41 VCC_IO 11 10 sky130_fd_pr__pfet_01v8__example_5595914180822
X42 VCC_IO 10 11 sky130_fd_pr__pfet_01v8__example_5595914180822
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1o_cdns_5595914180879 1 2
**
R0 1 5 0.01 short m=1
R1 6 2 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1s_cdns_5595914180881 1 2
**
R0 1 5 0.01 short m=1
R1 5 2 0.01 short m=1
.ENDS
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808423 1 2 3 4
**
XM0 1 2 4 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=0.25 p=2.5
XM1 2 3 1 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=0.25 p=2.5
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808424 1 2 3
**
XM0 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 m=1 sa=500000 sb=500001 a=0.75 p=3.5
XM1 2 3 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 m=1 sa=500001 sb=500000 a=0.75 p=3.5
.ENDS
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808426 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=450000 sb=450001 a=0.9 p=3.8
XM1 3 2 4 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=450001 sb=450000 a=0.9 p=3.8
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808435 2 3 4
**
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.375 p=2.5
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808433 2 3 4
**
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.375 p=2.5
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_io__com_ctl_ls_1v2 1 VCC_IO VPB VPWR HLD_H_N IN RST_H SET_H OUT_H_N OUT_H
**
*.SEEDPROM
XM0 23 20 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=75000.2 sb=75003.2 a=0.15 p=2.3
XM1 1 20 23 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75000.6 sb=75002.8 a=0.15 p=2.3
XM2 23 20 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.1 sb=75002.3 a=0.15 p=2.3
XM3 1 20 23 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.5 sb=75001.9 a=0.15 p=2.3
XM4 25 21 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.9 sb=75001.5 a=0.15 p=2.3
XM5 1 21 25 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.4 sb=75001 a=0.15 p=2.3
XM6 25 21 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.8 sb=75000.6 a=0.15 p=2.3
XM7 1 21 25 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=75003.2 sb=75000.2 a=0.15 p=2.3
XM8 1 18 OUT_H_N 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM9 OUT_H 19 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM10 22 HLD_H_N 19 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=1.8 p=7.2
XM11 18 HLD_H_N 24 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=1.8 p=7.2
XM12 1 RST_H 18 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=1.8 p=7.2
XM13 19 SET_H 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=1.8 p=7.2
XM14 VCC_IO 19 OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM15 OUT_H_N 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
X16 VPB IN 21 VPWR 20 sky130_fd_pr__pfet_01v8__example_55959141808430
X19 1 21 IN 20 sky130_fd_pr__nfet_01v8__example_55959141808423
X21 1 19 18 sky130_fd_pr__nfet_01v8__example_55959141808424
X25 1 VPWR 23 22 sky130_fd_pr__nfet_01v8__example_55959141808426
X26 1 VPWR 23 22 sky130_fd_pr__nfet_01v8__example_55959141808426
X27 1 VPWR 25 24 sky130_fd_pr__nfet_01v8__example_55959141808426
X28 1 VPWR 25 24 sky130_fd_pr__nfet_01v8__example_55959141808426
X33 VCC_IO 18 19 sky130_fd_pr__pfet_01v8__example_55959141808435
X34 VCC_IO 19 18 sky130_fd_pr__pfet_01v8__example_55959141808433
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_ctl_ls_v2 1 VCC_IO VPB VPWR HLD_H_N IN RST_H SET_H OUT_H_N OUT_H
**
*.SEEDPROM
XM0 23 20 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=75000.2 sb=75003.2 a=0.15 p=2.3
XM1 1 20 23 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75000.6 sb=75002.8 a=0.15 p=2.3
XM2 23 20 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.1 sb=75002.3 a=0.15 p=2.3
XM3 1 20 23 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.5 sb=75001.9 a=0.15 p=2.3
XM4 25 21 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.9 sb=75001.5 a=0.15 p=2.3
XM5 1 21 25 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.4 sb=75001 a=0.15 p=2.3
XM6 25 21 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.8 sb=75000.6 a=0.15 p=2.3
XM7 1 21 25 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=75003.2 sb=75000.2 a=0.15 p=2.3
XM8 1 18 OUT_H_N 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM9 OUT_H 19 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM10 22 HLD_H_N 19 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=1.8 p=7.2
XM11 18 HLD_H_N 24 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=1.8 p=7.2
XM12 1 RST_H 18 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=1.8 p=7.2
XM13 19 SET_H 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=1.8 p=7.2
XM14 VCC_IO 19 OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM15 OUT_H_N 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
X16 1 VPB sky130_fd_pr__model__parasitic__diode_ps2nw a=3.1672 p=7.24 m=1
X17 VPB IN 21 VPWR 20 sky130_fd_pr__pfet_01v8__example_55959141808430
X20 1 21 IN 20 sky130_fd_pr__nfet_01v8__example_55959141808423
X22 1 19 18 sky130_fd_pr__nfet_01v8__example_55959141808424
X26 1 VPWR 23 22 sky130_fd_pr__nfet_01v8__example_55959141808426
X27 1 VPWR 23 22 sky130_fd_pr__nfet_01v8__example_55959141808426
X28 1 VPWR 25 24 sky130_fd_pr__nfet_01v8__example_55959141808426
X29 1 VPWR 25 24 sky130_fd_pr__nfet_01v8__example_55959141808426
X34 VCC_IO 18 19 sky130_fd_pr__pfet_01v8__example_55959141808435
X35 VCC_IO 19 18 sky130_fd_pr__pfet_01v8__example_55959141808433
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_io__com_ctl_ls_en_1_v2 1 VCC_IO 3 VPWR HLD_H_N DM[1] RST_H SET_H OUT_H_N OUT_H
**
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VPB
XM0 24 21 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=75000.2 sb=75003.2 a=0.15 p=2.3
XM1 1 21 24 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75000.6 sb=75002.8 a=0.15 p=2.3
XM2 24 21 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.1 sb=75002.3 a=0.15 p=2.3
XM3 1 21 24 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.5 sb=75001.9 a=0.15 p=2.3
XM4 26 22 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.9 sb=75001.5 a=0.15 p=2.3
XM5 1 22 26 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.4 sb=75001 a=0.15 p=2.3
XM6 26 22 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.8 sb=75000.6 a=0.15 p=2.3
XM7 1 22 26 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=75003.2 sb=75000.2 a=0.15 p=2.3
XM8 1 19 OUT_H_N 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM9 OUT_H 20 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM10 23 HLD_H_N 20 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=1.8 p=7.2
XM11 19 HLD_H_N 25 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=1.8 p=7.2
XM12 1 RST_H 19 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=1.8 p=7.2
XM13 20 SET_H 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=1.8 p=7.2
XM14 3 DM[1] 22 3 sky130_fd_pr__pfet_01v8_hvt L=0.25 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=0.25 p=2.5
XM15 21 22 3 3 sky130_fd_pr__pfet_01v8_hvt L=0.25 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=0.25 p=2.5
XM16 VCC_IO 20 OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM17 OUT_H_N 19 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
X18 1 3 sky130_fd_pr__model__parasitic__diode_ps2nw a=3.1008 p=7.28 m=1
X21 1 22 DM[1] 21 sky130_fd_pr__nfet_01v8__example_55959141808423
X23 1 20 19 sky130_fd_pr__nfet_01v8__example_55959141808424
X27 1 VPWR 24 23 sky130_fd_pr__nfet_01v8__example_55959141808426
X28 1 VPWR 24 23 sky130_fd_pr__nfet_01v8__example_55959141808426
X29 1 VPWR 26 25 sky130_fd_pr__nfet_01v8__example_55959141808426
X30 1 VPWR 26 25 sky130_fd_pr__nfet_01v8__example_55959141808426
X35 VCC_IO 19 20 sky130_fd_pr__pfet_01v8__example_55959141808435
X36 VCC_IO 20 19 sky130_fd_pr__pfet_01v8__example_55959141808433
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_ctl_lsbank VGND VCC_IO VPWR IB_MODE_SEL HLD_I_H_N OD_I_H DM_H[1] DM_H_N[1] DM_H_N[0] DM_H[0] STARTUP_RST_H DM[0] INP_DIS STARTUP_ST_H INP_DIS_H_N DM_H_N[2] DM_H[2] DM[2] VTRIP_SEL_H_N VTRIP_SEL_H
+ VTRIP_SEL IB_MODE_SEL_H IB_MODE_SEL_H_N DM[1]
**
*.SEEDPROM
X0 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw a=33.634 p=25.7 m=1
X1 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw a=33.634 p=25.7 m=1
X2 VGND VPWR sky130_fd_pr__model__parasitic__diode_ps2nw a=5.3636 p=10.47 m=1
R3 41 OD_I_H 0.01 short m=1
R4 43 STARTUP_RST_H 0.01 short m=1
R5 46 45 0.01 short m=1
R6 47 OD_I_H 0.01 short m=1
R7 49 OD_I_H 0.01 short m=1
R8 51 VGND 0.01 short m=1
R9 OD_I_H 52 0.01 short m=1
R10 53 40 0.01 short m=1
X11 39 OD_I_H sky130_fd_io__tk_em2s_cdns_55959141808438
X12 40 VGND sky130_fd_io__tk_em2s_cdns_55959141808438
X13 42 sky130_fd_io__tk_em1o_cdns_5595914180880
X14 44 sky130_fd_io__tk_em1o_cdns_5595914180880
X15 STARTUP_ST_H sky130_fd_io__tk_em1o_cdns_5595914180880
X16 48 sky130_fd_io__tk_em1o_cdns_5595914180880
X17 50 sky130_fd_io__tk_em1o_cdns_5595914180880
X18 39 sky130_fd_io__tk_em1o_cdns_5595914180880
X19 42 VGND sky130_fd_io__tk_em1s_cdns_5595914180882
X20 44 STARTUP_ST_H sky130_fd_io__tk_em1s_cdns_5595914180882
X21 STARTUP_RST_H 45 sky130_fd_io__tk_em1s_cdns_5595914180882
X22 48 VGND sky130_fd_io__tk_em1s_cdns_5595914180882
X23 VGND 50 sky130_fd_io__tk_em1s_cdns_5595914180882
X24 VGND VCC_IO VPWR HLD_I_H_N 40 39 IB_MODE_SEL IB_MODE_SEL_H IB_MODE_SEL_H_N sky130_fd_io__com_ctl_lsv2
X25 VGND 33 sky130_fd_io__tk_em1o_cdns_5595914180879
X26 STARTUP_ST_H 34 sky130_fd_io__tk_em1o_cdns_5595914180879
X27 35 STARTUP_RST_H sky130_fd_io__tk_em1o_cdns_5595914180879
X28 VGND 37 sky130_fd_io__tk_em1o_cdns_5595914180879
X29 VGND 38 sky130_fd_io__tk_em1o_cdns_5595914180879
X30 33 OD_I_H sky130_fd_io__tk_em1s_cdns_5595914180881
X31 34 STARTUP_RST_H sky130_fd_io__tk_em1s_cdns_5595914180881
X32 STARTUP_ST_H 35 sky130_fd_io__tk_em1s_cdns_5595914180881
X33 37 OD_I_H sky130_fd_io__tk_em1s_cdns_5595914180881
X34 OD_I_H 38 sky130_fd_io__tk_em1s_cdns_5595914180881
X35 VGND VCC_IO VPWR VPWR HLD_I_H_N VTRIP_SEL 38 50 VTRIP_SEL_H_N VTRIP_SEL_H sky130_fd_io__com_ctl_ls_1v2
X36 VGND VCC_IO VPWR VPWR HLD_I_H_N DM[0] 34 44 DM_H_N[0] DM_H[0] sky130_fd_io__com_ctl_ls_v2
X37 VGND VCC_IO VPWR VPWR HLD_I_H_N INP_DIS 35 45 INP_DIS_H_N INP_DIS_H sky130_fd_io__com_ctl_ls_v2
X38 VGND VCC_IO VPWR VPWR HLD_I_H_N DM[2] 37 48 DM_H_N[2] DM_H[2] sky130_fd_io__com_ctl_ls_v2
X39 VGND VCC_IO VPWR VPWR HLD_I_H_N DM[1] 33 42 DM_H_N[1] DM_H[1] sky130_fd_io__com_ctl_ls_en_1_v2
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_5595914180864 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po L=1.5 W=0.8 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1s_cdns_5595914180859 2 3
**
R0 2 6 0.01 short m=1
R1 6 3 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__res250only_small PAD ROUT
**
R0 PAD 6 sky130_fd_pr__res_generic_po L=0.17 W=2 m=1
R1 6 7 sky130_fd_pr__res_generic_po L=10.07 W=2 m=1
R2 7 ROUT sky130_fd_pr__res_generic_po L=0.17 W=2 m=1
R3 PAD 6 0.01 short m=1
R4 7 ROUT 0.01 short m=1
R5 PAD 6 0.01 short m=1
R6 7 ROUT 0.01 short m=1
.ENDS
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_5595914180862 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po L=6 W=0.8 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_5595914180850 1 2 3
**
XM0 1 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=3 p=11.2
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_pddrvr_weakv2 2 3 PD_H PAD
**
*.SEEDPROM
X0 2 3 sky130_fd_pr__model__parasitic__diode_pw2dn a=107.174 p=75.96 m=1
X1 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X2 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X3 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X4 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X5 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X6 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808654 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=3.5 p=15
XM1 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=3.5 p=15
XM2 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=3.5 p=15
XM3 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=3.5 p=15
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_pudrvr_strong_slowv2 2 PU_H_N PAD
**
*.SEEDPROM
X0 2 PU_H_N PAD sky130_fd_pr__pfet_01v8__example_55959141808654
X1 2 PU_H_N PAD sky130_fd_pr__pfet_01v8__example_55959141808654
.ENDS
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__gpio_pddrvr_strong_slowv2 2 3 PD_H PAD
**
*.SEEDPROM
X0 2 3 sky130_fd_pr__model__parasitic__diode_pw2dn a=72.759 p=53.54 m=1
X1 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X2 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X3 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
X4 2 PD_H PAD sky130_fd_pr__nfet_01v8__example_5595914180850
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em2o_cdns_55959141808653 2 3
**
R0 2 6 0.01 short m=1
R1 7 3 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em2s_cdns_55959141808652 2 3
**
R0 2 6 0.01 short m=1
R1 6 3 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_5595914180838 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po L=10.2 W=0.5 m=1
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__pfet_con_diff_wo_abt_270v2 1 2 3 4 5 6 7 8 9 10
**
XM0 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=4.325 PD=6.55 PS=11.73 NRD=17.381 NRS=17.381 m=1 sa=300002 sb=300020 a=3 p=11.2
XM1 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=4.325 PD=6.55 PS=11.73 NRD=17.381 NRS=17.381 m=1 sa=300002 sb=300020 a=3 p=11.2
XM2 2 3 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300004 sb=300020 a=3 p=11.2
XM3 2 3 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300004 sb=300020 a=3 p=11.2
XM4 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300007 sb=300020 a=3 p=11.2
XM5 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300007 sb=300020 a=3 p=11.2
XM6 2 3 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300009 sb=300020 a=3 p=11.2
XM7 2 3 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300009 sb=300020 a=3 p=11.2
XM8 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300012 sb=300020 a=3 p=11.2
XM9 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300012 sb=300020 a=3 p=11.2
XM10 2 3 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300014 sb=300020 a=3 p=11.2
XM11 2 3 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300014 sb=300020 a=3 p=11.2
XM12 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300017 sb=300020 a=3 p=11.2
XM13 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300017 sb=300020 a=3 p=11.2
XM14 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300019 sb=300020 a=3 p=11.2
XM15 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300019 sb=300020 a=3 p=11.2
XM16 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM17 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM18 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM19 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM20 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM21 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM22 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM23 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM24 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM25 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM26 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM27 2 4 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM28 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM29 10 4 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM30 2 5 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM31 2 5 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM32 10 5 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM33 10 5 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM34 2 5 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM35 2 5 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM36 10 6 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM37 10 6 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM38 2 6 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM39 2 6 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM40 10 6 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300018 a=3 p=11.2
XM41 10 6 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300018 a=3 p=11.2
XM42 2 7 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300016 a=3 p=11.2
XM43 2 7 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300016 a=3 p=11.2
XM44 10 7 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300013 a=3 p=11.2
XM45 10 7 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300013 a=3 p=11.2
XM46 2 7 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300011 a=3 p=11.2
XM47 2 7 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300011 a=3 p=11.2
XM48 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300008 a=3 p=11.2
XM49 10 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300008 a=3 p=11.2
XM50 2 8 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300006 a=3 p=11.2
XM51 2 8 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300006 a=3 p=11.2
XM52 10 9 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300003 a=3 p=11.2
XM53 10 9 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300003 a=3 p=11.2
XM54 2 9 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=4.3 AS=2.975 PD=11.72 PS=6.19 NRD=17.19 NRS=17.381 m=1 sa=300020 sb=300002 a=3 p=11.2
XM55 2 9 10 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=4.3 AS=2.975 PD=11.72 PS=6.19 NRD=17.19 NRS=17.381 m=1 sa=300020 sb=300002 a=3 p=11.2
X56 1 2 sky130_fd_pr__model__parasitic__diode_ps2nw a=1473.41 p=184.25 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_pudrvr_strongv2 VNB TIE_HI_ESD VCC_IO PAD PU_H_N[2] PU_H_N[3]
**
X0 TIE_HI_ESD 9 sky130_fd_io__tk_em2o_cdns_55959141808653
X1 PU_H_N[3] 9 sky130_fd_io__tk_em2o_cdns_55959141808653
X2 TIE_HI_ESD 10 sky130_fd_io__tk_em2o_cdns_55959141808653
X3 PU_H_N[2] 10 sky130_fd_io__tk_em2o_cdns_55959141808653
X4 PU_H_N[3] 11 sky130_fd_io__tk_em2o_cdns_55959141808653
X5 PU_H_N[2] 11 sky130_fd_io__tk_em2o_cdns_55959141808653
X6 TIE_HI_ESD 12 sky130_fd_io__tk_em2o_cdns_55959141808653
X7 PU_H_N[2] 12 sky130_fd_io__tk_em2o_cdns_55959141808653
X8 PU_H_N[3] 13 sky130_fd_io__tk_em2o_cdns_55959141808653
X9 PU_H_N[2] 13 sky130_fd_io__tk_em2o_cdns_55959141808653
X10 PU_H_N[2] 9 sky130_fd_io__tk_em2s_cdns_55959141808652
X11 PU_H_N[3] 10 sky130_fd_io__tk_em2s_cdns_55959141808652
X12 TIE_HI_ESD 11 sky130_fd_io__tk_em2s_cdns_55959141808652
X13 PU_H_N[3] 12 sky130_fd_io__tk_em2s_cdns_55959141808652
X14 TIE_HI_ESD 13 sky130_fd_io__tk_em2s_cdns_55959141808652
X15 TIE_HI_ESD VCC_IO sky130_fd_pr__res_generic_po__example_5595914180838
X16 VNB VCC_IO PU_H_N[2] PU_H_N[3] 9 10 11 12 13 PAD sky130_fd_io__pfet_con_diff_wo_abt_270v2
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__nfet_con_diff_wo_abt_270v2 VSSIO VCC_IO 4 5 6 7 8 9 10 11 12 13 PAD
**
*.SEEDPROM
XM0 PAD 4 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.425 PD=6.55 PS=11.37 NRD=10.374 NRS=8.7666 m=1 sa=300002 sb=300020 a=3 p=11.2
XM1 PAD 4 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.425 PD=6.55 PS=11.37 NRD=10.374 NRS=8.7666 m=1 sa=300002 sb=300020 a=3 p=11.2
XM2 VSSIO 4 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300004 sb=300020 a=3 p=11.2
XM3 VSSIO 4 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300004 sb=300020 a=3 p=11.2
XM4 PAD 4 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300007 sb=300020 a=3 p=11.2
XM5 PAD 4 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300007 sb=300020 a=3 p=11.2
XM6 VSSIO 4 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300009 sb=300020 a=3 p=11.2
XM7 VSSIO 4 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300009 sb=300020 a=3 p=11.2
XM8 PAD 5 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300011 sb=300020 a=3 p=11.2
XM9 PAD 5 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300011 sb=300020 a=3 p=11.2
XM10 VSSIO 5 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300014 sb=300020 a=3 p=11.2
XM11 VSSIO 5 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300014 sb=300020 a=3 p=11.2
XM12 PAD 5 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300016 sb=300020 a=3 p=11.2
XM13 PAD 5 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300016 sb=300020 a=3 p=11.2
XM14 VSSIO 6 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300019 sb=300020 a=3 p=11.2
XM15 VSSIO 6 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300019 sb=300020 a=3 p=11.2
XM16 PAD 6 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM17 PAD 6 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM18 VSSIO 6 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM19 VSSIO 6 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM20 PAD 7 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM21 PAD 7 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM22 VSSIO 7 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM23 VSSIO 7 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM24 PAD 7 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM25 PAD 7 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM26 VSSIO 8 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM27 VSSIO 8 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM28 PAD 9 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM29 PAD 9 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM30 VSSIO 9 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM31 VSSIO 9 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM32 PAD 9 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM33 PAD 9 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM34 VSSIO 10 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM35 VSSIO 10 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM36 PAD 10 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM37 PAD 10 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM38 VSSIO 10 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM39 VSSIO 10 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM40 PAD 10 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300018 a=3 p=11.2
XM41 PAD 10 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300018 a=3 p=11.2
XM42 VSSIO 10 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300016 a=3 p=11.2
XM43 VSSIO 10 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300016 a=3 p=11.2
XM44 PAD 10 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300013 a=3 p=11.2
XM45 PAD 10 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300013 a=3 p=11.2
XM46 VSSIO 11 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300011 a=3 p=11.2
XM47 VSSIO 11 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300011 a=3 p=11.2
XM48 PAD 12 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300008 a=3 p=11.2
XM49 PAD 12 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300008 a=3 p=11.2
XM50 VSSIO 13 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300006 a=3 p=11.2
XM51 VSSIO 13 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300006 a=3 p=11.2
XM52 PAD 13 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300003 a=3 p=11.2
XM53 PAD 13 VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300003 a=3 p=11.2
XM54 VSSIO 13 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.425 AS=2.975 PD=11.37 PS=6.19 NRD=8.7666 NRS=10.374 m=1 sa=300020 sb=300002 a=3 p=11.2
XM55 VSSIO 13 PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.425 AS=2.975 PD=11.37 PS=6.19 NRD=8.7666 NRS=10.374 m=1 sa=300020 sb=300002 a=3 p=11.2
X56 VSSIO VCC_IO sky130_fd_pr__model__parasitic__diode_pw2dn a=1576.75 p=188.14 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_pddrvr_strong VGND_IO VCC_IO TIE_LO_ESD PD_H[2] PD_H[3] PD_H_I2C PAD
**
*.SEEDPROM
*.CALIBRE ISOLATED NETS: FORCE_LO_H FORCE_LOVOL_H VSSIO_AMX
X0 VGND_IO VCC_IO condiode a=1e-06 p=0.004 m=1
X1 TIE_LO_ESD 26 sky130_fd_io__tk_em2o_cdns_55959141808653
X2 PD_H[2] 26 sky130_fd_io__tk_em2o_cdns_55959141808653
X3 PD_H[3] 25 sky130_fd_io__tk_em2o_cdns_55959141808653
X4 TIE_LO_ESD 25 sky130_fd_io__tk_em2o_cdns_55959141808653
X5 PD_H[2] 24 sky130_fd_io__tk_em2o_cdns_55959141808653
X6 TIE_LO_ESD 24 sky130_fd_io__tk_em2o_cdns_55959141808653
X7 PD_H[2] 23 sky130_fd_io__tk_em2o_cdns_55959141808653
X8 TIE_LO_ESD 23 sky130_fd_io__tk_em2o_cdns_55959141808653
X9 PD_H[2] 22 sky130_fd_io__tk_em2o_cdns_55959141808653
X10 TIE_LO_ESD 22 sky130_fd_io__tk_em2o_cdns_55959141808653
X11 PD_H[2] 21 sky130_fd_io__tk_em2o_cdns_55959141808653
X12 TIE_LO_ESD 21 sky130_fd_io__tk_em2o_cdns_55959141808653
X13 PD_H[2] 20 sky130_fd_io__tk_em2o_cdns_55959141808653
X14 PD_H[3] 20 sky130_fd_io__tk_em2o_cdns_55959141808653
X15 PD_H[3] 26 sky130_fd_io__tk_em2s_cdns_55959141808652
X16 PD_H[2] 25 sky130_fd_io__tk_em2s_cdns_55959141808652
X17 PD_H[3] 24 sky130_fd_io__tk_em2s_cdns_55959141808652
X18 PD_H[3] 23 sky130_fd_io__tk_em2s_cdns_55959141808652
X19 PD_H[3] 22 sky130_fd_io__tk_em2s_cdns_55959141808652
X20 PD_H[3] 21 sky130_fd_io__tk_em2s_cdns_55959141808652
X21 TIE_LO_ESD 20 sky130_fd_io__tk_em2s_cdns_55959141808652
X22 TIE_LO_ESD VGND_IO sky130_fd_pr__res_generic_po__example_5595914180838
X23 VGND_IO VCC_IO 20 21 22 23 24 PD_H[2] PD_H[3] PD_H_I2C 25 26 PAD sky130_fd_io__nfet_con_diff_wo_abt_270v2
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_odrvrv2 VGND VGND_IO VCC_IO PU_H_N[0] PD_H[1] PAD PD_H[0] PU_H_N[1] PU_H_N[3] TIE_HI_ESD PU_H_N[2] PD_H[2] PD_H[3] TIE_LO_ESD 25
**
*.SEEDPROM
*.CALIBRE ISOLATED NETS: FORCE_HI_H_N VSSIO_AMX FORCE_LOVOL_H FORCE_LO_H
XM0 26 PU_H_N[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=2.5 p=11
XM1 VCC_IO PU_H_N[0] 26 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=2.5 p=11
XM2 26 PU_H_N[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=2.5 p=11
XM3 VCC_IO PU_H_N[0] 26 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=2.5 p=11
X4 VGND_IO VCC_IO condiode a=1e-06 p=0.004 m=1
X5 VGND_IO VCC_IO condiode a=1e-06 p=0.004 m=1
X6 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw a=167.455 p=75.76 m=1
X7 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2dn a=2283.69 p=218.67 m=1
R8 26 27 sky130_fd_pr__res_generic_po L=50 W=0.8 m=1
R9 28 29 sky130_fd_pr__res_generic_po L=5 W=2 m=1
R10 29 31 sky130_fd_pr__res_generic_po L=3 W=2 m=1
R11 27 30 sky130_fd_pr__res_generic_po L=12 W=0.8 m=1
R12 31 32 sky130_fd_pr__res_generic_po L=2 W=2 m=1
R13 30 38 0.01 short m=1
R14 39 33 0.01 short m=1
R15 29 40 0.01 short m=1
R16 40 31 0.01 short m=1
X17 36 32 sky130_fd_pr__res_generic_po__example_5595914180864
X18 34 35 sky130_fd_pr__res_generic_po__example_5595914180864
X19 37 36 sky130_fd_pr__res_generic_po__example_5595914180864
X20 35 37 sky130_fd_pr__res_generic_po__example_5595914180864
X21 33 34 sky130_fd_io__tk_em1s_cdns_5595914180859
X22 36 32 sky130_fd_io__tk_em1s_cdns_5595914180859
X23 34 35 sky130_fd_io__tk_em1s_cdns_5595914180859
X24 35 37 sky130_fd_io__tk_em1s_cdns_5595914180859
X25 37 36 sky130_fd_io__tk_em1s_cdns_5595914180859
X26 PAD 32 sky130_fd_io__res250only_small
X35 33 30 sky130_fd_pr__res_bent_po__example_5595914180862
X36 34 33 sky130_fd_pr__res_bent_po__example_5595914180862
X37 VGND_IO VCC_IO PD_H[0] 26 sky130_fd_io__gpio_pddrvr_weakv2
X38 VCC_IO PU_H_N[0] 26 sky130_fd_pr__pfet_01v8__example_55959141808654
X39 VCC_IO PU_H_N[1] 28 sky130_fd_io__com_pudrvr_strong_slowv2
X45 VGND_IO VCC_IO PD_H[1] 28 sky130_fd_io__gpio_pddrvr_strong_slowv2
X46 VGND TIE_HI_ESD VCC_IO PAD PU_H_N[2] PU_H_N[3] sky130_fd_io__gpio_pudrvr_strongv2
X47 VGND_IO VCC_IO TIE_LO_ESD PD_H[2] PD_H[3] 25 PAD sky130_fd_io__gpiov2_pddrvr_strong
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__signal_5_sym_hv_local_5term NBODY NWELLRING GATE VGND IN 7
**
*.SEEDPROM
XM0 IN GATE VGND NBODY sky130_fd_pr__esd_nfet_g5v0d10v5 L=0.6 W=5.4 AD=3.65486 AS=3.65486 PD=11.6192 PS=11.6192 NRD=8.436 NRS=9.2796 m=1 sa=300000 sb=300000 a=3.24 p=12
R1 NWELLRING 7 0.01 short m=1
R2 NBODY 36 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_buf_localesd VSSD VDDIO_Q VTRIP_SEL_H OUT_VT OUT_H IN_H
**
*.SEEDPROM
XM0 OUT_H VTRIP_SEL_H OUT_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=500000 sb=500000 a=3 p=8
X1 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=5.32 p=17.88 m=1
X2 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=8.5092 p=29.27 m=1
X3 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=8.5092 p=29.27 m=1
X6 IN_H OUT_H sky130_fd_io__res250only_small
X7 VSSD VDDIO_Q VSSD VSSD OUT_H 10 sky130_fd_io__signal_5_sym_hv_local_5term
X8 VSSD VDDIO_Q VSSD OUT_H VDDIO_Q 9 sky130_fd_io__signal_5_sym_hv_local_5term
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__gpiov2_in_buf VSSD VDDIO_Q IN_H MODE_NORMAL_N IN_VT VTRIP_SEL_H_N OUT VTRIP_SEL_H
**
*.SEEDPROM
XM0 17 IN_H 11 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=400000 sb=400015 a=4 p=11.6
XM1 11 IN_H 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400001 sb=400014 a=4 p=11.6
XM2 17 IN_H 11 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400002 sb=400013 a=4 p=11.6
XM3 11 IN_H 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400003 sb=400012 a=4 p=11.6
XM4 17 IN_H 11 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400004 sb=400011 a=4 p=11.6
XM5 VSSD IN_VT 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400005 sb=400010 a=4 p=11.6
XM6 17 IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400006 sb=400009 a=4 p=11.6
XM7 VSSD IN_H 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400007 sb=400007 a=4 p=11.6
XM8 17 IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400009 sb=400006 a=4 p=11.6
XM9 VSSD IN_H 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400010 sb=400005 a=4 p=11.6
XM10 17 IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400011 sb=400004 a=4 p=11.6
XM11 19 11 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400012 sb=400003 a=4 p=11.6
XM12 17 11 19 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400013 sb=400002 a=4 p=11.6
XM13 19 11 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400014 sb=400001 a=4 p=11.6
XM14 17 11 19 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=400015 sb=400000 a=4 p=11.6
XM15 20 MODE_NORMAL_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.196 PD=0.98 PS=1.96 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.42 p=2.6
XM16 VSSD IN_H 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 sa=400000 sb=400000 a=4 p=11.6
XM17 VSSD VTRIP_SEL_H 20 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.42 p=2.6
XM18 10 20 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.42 p=2.6
XM19 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 sa=400000 sb=400000 a=4 p=11.6
XM20 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 sa=400000 sb=400000 a=4 p=11.6
XM21 18 11 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=400000 sb=400003 a=0.8 p=3.6
XM22 VSSD VTRIP_SEL_H_N IN_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=500000 sb=500003 a=3 p=8
XM23 12 MODE_NORMAL_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=1.5 p=7
XM24 17 11 18 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=400001 sb=400002 a=0.8 p=3.6
XM25 VSSD MODE_NORMAL_N 12 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=1.5 p=7
XM26 18 11 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=400002 sb=400001 a=0.8 p=3.6
XM27 12 11 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250003 sb=250001 a=1.5 p=7
XM28 17 11 18 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=400003 sb=400000 a=0.8 p=3.6
XM29 VSSD 11 12 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250004 sb=250000 a=1.5 p=7
XM30 VSSD 12 OUT_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=2.5 p=11
XM31 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=2.5 p=11
XM32 16 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=2.5 p=11
XM33 VDDIO_Q MODE_NORMAL_N 16 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=2.5 p=11
XM34 11 IN_H 16 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=400000 sb=400003 a=4 p=11.6
XM35 15 IN_H 11 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400001 sb=400001 a=4 p=11.6
XM36 VDDIO_Q 10 15 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=2.5 p=11
XM37 15 10 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250000 a=2.5 p=11
XM38 VDDIO_Q VDDIO_Q VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=400000 sb=400004 a=4 p=11.6
XM39 19 10 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250003 a=2.5 p=11
XM40 VDDIO_Q 10 19 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=2.5 p=11
XM41 18 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250002 a=2.5 p=11
XM42 VDDIO_Q MODE_NORMAL_N 18 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250001 a=2.5 p=11
XM43 14 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250004 sb=250000 a=2.5 p=11
XM44 12 11 14 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
XM45 VDDIO_Q 12 OUT_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=2.5 p=11
XM46 OUT OUT_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=2.5 p=11
XM47 858 MODE_NORMAL_N 20 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM48 858 MODE_NORMAL_N 20 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM49 VDDIO_Q VTRIP_SEL_H 858 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM50 VDDIO_Q VTRIP_SEL_H 858 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM51 10 20 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM52 10 20 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
.ENDS
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808600 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.3975 PD=3.53 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.75 p=4
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_io__gpiov2_ipath_hvls VSSD VDDIO_Q MODE_VCCHIB_N INB_VCCHIB MODE_VCCHIB MODE_NORMAL_N MODE_NORMAL IN_VDDIO IN_VCCHIB OUT
**
*.SEEDPROM
XM0 11 MODE_VCCHIB_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250005 a=2.5 p=11
XM1 18 INB_VCCHIB 11 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250005 a=2.5 p=11
XM2 11 INB_VCCHIB 18 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250004 a=2.5 p=11
XM3 18 INB_VCCHIB 11 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250003 a=2.5 p=11
XM4 VSSD MODE_VCCHIB 18 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250002 a=2.5 p=11
XM5 18 MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250004 sb=250002 a=2.5 p=11
XM6 VSSD MODE_VCCHIB 18 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250001 a=2.5 p=11
XM7 18 MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250000 a=2.5 p=11
XM8 VSSD MODE_VCCHIB 19 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250005 a=2.5 p=11
XM9 19 MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250004 a=2.5 p=11
XM10 20 13 OUT_B VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=1.5 p=7
XM11 VSSD MODE_VCCHIB 20 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=1.5 p=7
XM12 21 MODE_NORMAL VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=1.5 p=7
XM13 OUT_B IN_VDDIO 21 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=1.5 p=7
XM14 VSSD MODE_VCCHIB 19 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250003 a=2.5 p=11
XM15 19 MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=2.5 p=11
XM16 12 IN_VCCHIB 19 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250002 a=2.5 p=11
XM17 19 IN_VCCHIB 12 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250004 sb=250001 a=2.5 p=11
XM18 12 IN_VCCHIB 19 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250000 a=2.5 p=11
XM19 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=2.5 p=11
XM20 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250001 a=2.5 p=11
XM21 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=2.5 p=11
XM22 VDDIO_Q 11 12 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.75 p=4
XM23 11 12 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.75 p=4
XM24 13 12 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.3975 PD=3.53 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.75 p=4
XM25 OUT_B 13 16 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=2.5 p=11
XM26 16 13 OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=2.5 p=11
XM27 VDDIO_Q MODE_VCCHIB_N 16 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=2.5 p=11
XM28 16 MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=2.5 p=11
XM29 VDDIO_Q MODE_NORMAL_N 17 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=2.5 p=11
XM30 17 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=2.5 p=11
XM31 OUT_B IN_VDDIO 17 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=2.5 p=11
XM32 17 IN_VDDIO OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=2.5 p=11
XM33 15 MODE_VCCHIB OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=2.5 p=11
XM34 VDDIO_Q MODE_NORMAL 15 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=2.5 p=11
XM35 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250003 a=2.5 p=11
XM36 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=2.5 p=11
XM37 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250002 a=2.5 p=11
XM38 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=2.5 p=11
XM39 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250000 a=2.5 p=11
X62 VSSD 12 VSSD 13 sky130_fd_pr__nfet_01v8__example_55959141808600
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__gpiov2_vcchib_in_buf VSSD VCCHIB MODE_VCCHIB_LV_N OUT_N IN_H OUT
**
*.SEEDPROM
XM0 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=0.25 p=2.5
XM1 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.25 p=2.5
XM2 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=0.25 p=2.5
XM3 VSSD 7 OUT_N VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=125000 sb=125002 a=0.25 p=2.5
XM4 7 8 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=125001 sb=125002 a=0.25 p=2.5
XM5 VSSD 8 7 VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.25 p=2.5
XM6 7 MODE_VCCHIB_LV_N VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=125002 sb=125001 a=0.25 p=2.5
XM7 VSSD MODE_VCCHIB_LV_N 7 VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=125002 sb=125000 a=0.25 p=2.5
XM8 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=400000 sb=400000 a=0.8 p=3.6
XM9 12 8 11 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=400000 sb=400002 a=0.8 p=3.6
XM10 11 8 12 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=400001 sb=400001 a=0.8 p=3.6
XM11 12 8 11 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=400002 sb=400000 a=0.8 p=3.6
XM12 8 IN_H 12 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=400000 sb=400003 a=4 p=11.6
XM13 12 IN_H 8 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400001 sb=400002 a=4 p=11.6
XM14 VSSD IN_H 12 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400002 sb=400001 a=4 p=11.6
XM15 12 IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=400003 sb=400000 a=4 p=11.6
XM16 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 sa=400000 sb=400000 a=4 p=11.6
XM17 VCCHIB MODE_VCCHIB_LV_N 10 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=125000 sb=125000 a=0.75 p=6.5
XM18 VCCHIB MODE_VCCHIB_LV_N 9 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=125000 sb=125002 a=1.25 p=10.5
XM19 9 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=1.25 p=10.5
XM20 VCCHIB MODE_VCCHIB_LV_N 9 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=1.25 p=10.5
XM21 11 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=125002 sb=125000 a=1.25 p=10.5
XM22 VCCHIB 7 OUT_N VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=1.25 p=10.5
XM23 OUT OUT_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=1.25 p=10.5
XM24 7 8 10 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=0.25 p=2.5
XM25 10 8 7 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=0.25 p=2.5
XM26 8 IN_H 9 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=400000 sb=400001 a=4 p=11.6
XM27 9 IN_H 8 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=400001 sb=400000 a=4 p=11.6
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_inbuf_lvinv_x1 VGND VPWR IN OUT
**
*.SEEDPROM
XM0 VGND IN OUT VGND sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=125000 sb=125000 a=0.25 p=2.5
XM1 VPWR IN OUT VPWR sky130_fd_pr__pfet_01v8_hvt L=0.25 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=125000 sb=125000 a=0.75 p=6.5
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__gpiov2_ipath_lvls VSSD VCCHIB MODE_NORMAL_LV IN_VDDIO 5 MODE_NORMAL_LV_N OUT_B MODE_VCCHIB_LV_N IN_VCCHIB MODE_VCCHIB_LV OUT
**
*.SEEDPROM
XM0 VSSD MODE_NORMAL_LV 18 VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=0.75 p=6.5
XM1 5 12 VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=0.75 p=6.5
XM2 OUT_B 5 16 VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=125000 sb=125002 a=0.75 p=6.5
XM3 16 5 OUT_B VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.75 p=6.5
XM4 VSSD MODE_NORMAL_LV 16 VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.75 p=6.5
XM5 16 MODE_NORMAL_LV VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=125002 sb=125000 a=0.75 p=6.5
XM6 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=0.75 p=6.5
XM7 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=0.75 p=6.5
XM8 OUT_B IN_VCCHIB 17 VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=125000 sb=125002 a=0.75 p=6.5
XM9 17 IN_VCCHIB OUT_B VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.75 p=6.5
XM10 VSSD MODE_VCCHIB_LV 17 VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.75 p=6.5
XM11 17 MODE_VCCHIB_LV VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.25 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=125002 sb=125000 a=0.75 p=6.5
XM12 VCCHIB MODE_NORMAL_LV 12 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=1.25 p=10.5
XM13 5 12 VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=1.25 p=10.5
XM14 OUT_B 5 14 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=125000 sb=125002 a=0.75 p=6.5
XM15 14 5 OUT_B VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.75 p=6.5
XM16 VCCHIB MODE_NORMAL_LV_N 14 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.75 p=6.5
XM17 14 MODE_NORMAL_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=125002 sb=125000 a=0.75 p=6.5
XM18 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=125000 sb=125002 a=0.75 p=6.5
XM19 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.75 p=6.5
XM20 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.75 p=6.5
XM21 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=125002 sb=125000 a=0.75 p=6.5
XM22 VCCHIB MODE_VCCHIB_LV_N 15 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=125000 sb=125002 a=0.75 p=6.5
XM23 15 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.75 p=6.5
XM24 OUT_B IN_VCCHIB 15 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.75 p=6.5
XM25 15 IN_VCCHIB OUT_B VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=125002 sb=125000 a=0.75 p=6.5
XM26 13 MODE_NORMAL_LV OUT_B VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=0.75 p=6.5
XM27 VCCHIB MODE_VCCHIB_LV 13 VCCHIB sky130_fd_pr__pfet_01v8 L=0.25 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=0.75 p=6.5
XM28 12 IN_VDDIO VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=2.5 p=11
XM29 VCCHIB IN_VDDIO 12 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=2.5 p=11
X33 VSSD IN_VDDIO 12 18 sky130_fd_pr__nfet_01v8__example_55959141808600
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_ibuf_se VSSD VDDIO_Q VCCHIB MODE_NORMAL_N MODE_VCCHIB_N ENABLE_VDDIO_LV IN_H VTRIP_SEL_H VTRIP_SEL_H_N IN_VT IBUFMUX_OUT_H IBUFMUX_OUT 14
**
*.SEEDPROM
XM0 VSSD MODE_NORMAL_N 15 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM1 16 MODE_VCCHIB_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM2 127 16 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300003 a=0.42 p=2.6
XM3 VSSD ENABLE_VDDIO_LV 127 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300002 a=0.42 p=2.6
XM4 128 ENABLE_VDDIO_LV VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=13.8396 NRS=0 m=1 sa=300002 sb=300001 a=0.42 p=2.6
XM5 18 15 128 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300003 sb=300000 a=0.42 p=2.6
XM6 VDDIO_Q MODE_NORMAL_N 15 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM7 VDDIO_Q MODE_NORMAL_N 15 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM8 16 MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM9 16 MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM10 17 16 VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM11 17 16 VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM12 VCCHIB ENABLE_VDDIO_LV 17 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM13 VCCHIB ENABLE_VDDIO_LV 17 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM14 18 ENABLE_VDDIO_LV VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM15 18 ENABLE_VDDIO_LV VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM16 VCCHIB 15 18 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM17 VCCHIB 15 18 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
X18 VSSD VCCHIB sky130_fd_pr__model__parasitic__diode_ps2nw a=51.8546 p=44.62 m=1
X19 VSSD VCCHIB sky130_fd_pr__model__parasitic__diode_ps2nw a=98.14 p=57.76 m=1
X24 VSSD VDDIO_Q IN_H MODE_NORMAL_N IN_VT VTRIP_SEL_H_N 19 VTRIP_SEL_H sky130_fd_io__gpiov2_in_buf
X25 VSSD VDDIO_Q MODE_VCCHIB_N 21 16 MODE_NORMAL_N 15 19 20 IBUFMUX_OUT_H sky130_fd_io__gpiov2_ipath_hvls
X26 VSSD VCCHIB 17 21 IN_H 20 sky130_fd_io__gpiov2_vcchib_in_buf
X27 VSSD VCCHIB 17 22 sky130_fd_io__gpiov2_inbuf_lvinv_x1
X28 VSSD VCCHIB 18 23 sky130_fd_io__gpiov2_inbuf_lvinv_x1
X29 VSSD VCCHIB 23 19 14 18 24 17 20 22 IBUFMUX_OUT sky130_fd_io__gpiov2_ipath_lvls
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_ictl_logic VSSD VDDIO_Q DM_H_N[1] DM_H_N[0] DM_H_N[2] INP_DIS_H_N IB_MODE_SEL_H MODE_VCCHIB_N IB_MODE_SEL_H_N MODE_NORMAL_N TRIPSEL_I_H VTRIP_SEL_H_N TRIPSEL_I_H_N
**
*.SEEDPROM
XM0 16 DM_H_N[1] VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM1 15 DM_H_N[0] 16 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM2 VSSD 15 17 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.42 p=2.6
XM3 247 DM_H_N[2] VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=13.8396 NRS=0 m=1 sa=300001 sb=300001 a=0.42 p=2.6
XM4 18 17 247 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300002 sb=300000 a=0.42 p=2.6
XM5 248 INP_DIS_H_N INP_DIS_I_H VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300002 a=0.42 p=2.6
XM6 VSSD 18 248 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300001 a=0.42 p=2.6
XM7 INP_DIS_I_H_N INP_DIS_I_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.42 p=2.6
XM8 249 IB_MODE_SEL_H MODE_VCCHIB_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300003 a=0.42 p=2.6
XM9 VSSD INP_DIS_I_H_N 249 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300002 a=0.42 p=2.6
XM10 250 INP_DIS_I_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=13.8396 NRS=0 m=1 sa=300002 sb=300001 a=0.42 p=2.6
XM11 MODE_NORMAL_N IB_MODE_SEL_H_N 250 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300003 sb=300000 a=0.42 p=2.6
XM12 TRIPSEL_I_H MODE_NORMAL_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.196 PD=0.98 PS=1.96 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.42 p=2.6
XM13 VSSD VTRIP_SEL_H_N TRIPSEL_I_H VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.42 p=2.6
XM14 TRIPSEL_I_H_N TRIPSEL_I_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.42 p=2.6
XM15 15 DM_H_N[1] VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM16 15 DM_H_N[1] VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM17 VDDIO_Q DM_H_N[0] 15 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM18 VDDIO_Q DM_H_N[0] 15 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM19 VDDIO_Q 15 17 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM20 VDDIO_Q 15 17 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM21 18 DM_H_N[2] VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM22 18 DM_H_N[2] VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM23 VDDIO_Q 17 18 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM24 VDDIO_Q 17 18 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM25 INP_DIS_I_H INP_DIS_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM26 INP_DIS_I_H INP_DIS_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM27 VDDIO_Q 18 INP_DIS_I_H VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM28 VDDIO_Q 18 INP_DIS_I_H VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM29 INP_DIS_I_H_N INP_DIS_I_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM30 INP_DIS_I_H_N INP_DIS_I_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM31 MODE_VCCHIB_N IB_MODE_SEL_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM32 MODE_VCCHIB_N IB_MODE_SEL_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM33 VDDIO_Q INP_DIS_I_H_N MODE_VCCHIB_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM34 VDDIO_Q INP_DIS_I_H_N MODE_VCCHIB_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM35 MODE_NORMAL_N INP_DIS_I_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM36 MODE_NORMAL_N INP_DIS_I_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM37 VDDIO_Q IB_MODE_SEL_H_N MODE_NORMAL_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM38 VDDIO_Q IB_MODE_SEL_H_N MODE_NORMAL_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM39 246 MODE_NORMAL_N TRIPSEL_I_H VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM40 246 MODE_NORMAL_N TRIPSEL_I_H VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM41 VDDIO_Q VTRIP_SEL_H_N 246 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM42 VDDIO_Q VTRIP_SEL_H_N 246 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM43 TRIPSEL_I_H_N TRIPSEL_I_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM44 TRIPSEL_I_H_N TRIPSEL_I_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_ipath VSSD VDDIO_Q ENABLE_VDDIO_LV DM_H_N[0] 6 OUT_H 8 MODE_VCCHIB_N PAD 11 OUT VCCHIB DM_H_N[1] DM_H_N[2] INP_DIS_H_N IB_MODE_SEL_H IB_MODE_SEL_H_N VTRIP_SEL_H_N
**
*.SEEDPROM
X0 VSSD VDDIO_Q 8 22 21 PAD sky130_fd_io__gpiov2_buf_localesd
X1 VSSD VDDIO_Q VCCHIB 6 MODE_VCCHIB_N ENABLE_VDDIO_LV 21 8 11 22 OUT_H OUT 23 sky130_fd_io__gpiov2_ibuf_se
X2 VSSD VDDIO_Q DM_H_N[1] DM_H_N[0] DM_H_N[2] INP_DIS_H_N IB_MODE_SEL_H MODE_VCCHIB_N IB_MODE_SEL_H_N 6 8 VTRIP_SEL_H_N 11 sky130_fd_io__gpiov2_ictl_logic
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__tk_em1o_cdns_55959141808289 3 4
**
*.SEEDPROM
R0 3 8 0.01 short m=1
R1 9 4 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1s_cdns_55959141808288 2 3
**
*.SEEDPROM
R0 2 7 0.01 short m=1
R1 7 3 0.01 short m=1
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_55959141808285 2 3
**
*.SEEDPROM
R0 2 3 sky130_fd_pr__res_generic_po L=4 W=0.33 m=1
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808644 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 m=1 sa=2e+06 sb=2e+06 a=1.68 p=8.84
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_55959141808286 3 4
**
*.SEEDPROM
R0 3 4 sky130_fd_pr__res_generic_po L=11 W=0.33 m=1
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__feascom_pupredrvr_nbiasv2 VGND_IO VCC_IO EN_H NBIAS DRVHI_H PUEN_H 8 PU_H_N EN_H_N 11 12 13
**
*.SEEDPROM
XM0 VGND_IO DRVHI_H 33 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.259 AS=0.265 PD=1.612 PS=2.53 NRD=26.9724 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM1 NBIAS NBIAS 8 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=1.5 p=7
XM2 8 NBIAS NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=1.5 p=7
XM3 36 EN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.2025 AS=0.3885 PD=1.77 PS=2.418 NRD=6.0762 NRS=0 m=1 sa=250001 sb=250002 a=0.75 p=4
XM4 NBIAS NBIAS 8 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=1.5 p=7
XM5 37 31 36 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.2025 AS=0.2025 PD=1.77 PS=1.77 NRD=6.0762 NRS=6.0762 m=1 sa=250002 sb=250001 a=0.75 p=4
XM6 8 NBIAS NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=1.5 p=7
XM7 30 DRVHI_H 37 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.2025 PD=3.53 PS=1.77 NRD=0 NRS=6.0762 m=1 sa=250002 sb=250000 a=0.75 p=4
XM8 8 8 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250008 a=1.5 p=7
XM9 VGND_IO 8 8 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250007 a=1.5 p=7
XM10 8 8 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250006 a=1.5 p=7
XM11 VGND_IO 8 8 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250005 a=1.5 p=7
XM12 13 32 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250003 sb=250005 a=1.5 p=7
XM13 VGND_IO 30 38 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=4 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 sa=2e+06 sb=2.00001e+06 a=1.68 p=8.84
XM14 VGND_IO 32 13 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250004 sb=250004 a=1.5 p=7
XM15 13 32 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250005 sb=250003 a=1.5 p=7
XM16 VGND_IO 32 13 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250005 sb=250002 a=1.5 p=7
XM17 NBIAS EN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250006 sb=250002 a=1.5 p=7
XM18 VGND_IO 33 NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250007 sb=250001 a=1.5 p=7
XM19 32 33 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250008 sb=250000 a=1.5 p=7
XM20 11 11 12 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=1.5 p=7
XM21 12 11 11 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=1.5 p=7
XM22 32 12 12 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=1.5 p=7
XM23 12 12 32 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=1.5 p=7
XM24 32 VCC_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=8 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 sa=4e+06 sb=4e+06 a=3.36 p=16.84
XM25 33 DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250010 a=0.5 p=3
XM26 30 DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250006 a=0.5 p=3
XM27 VCC_IO DRVHI_H 33 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.1925 AS=0.14 PD=1.385 PS=1.28 NRD=20.055 NRS=0 m=1 sa=250001 sb=250009 a=0.5 p=3
XM28 VCC_IO EN_H 30 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250005 a=0.5 p=3
XM29 34 PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=250002 sb=250004 a=0.5 p=3
XM30 NBIAS 30 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.1925 PD=1.28 PS=1.385 NRD=0 NRS=0 m=1 sa=400002 sb=400007 a=0.8 p=3.6
XM31 VCC_IO DRVHI_H 34 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.260563 AS=0.14 PD=2.1338 PS=1.28 NRD=0 NRS=0 m=1 sa=250002 sb=250004 a=0.5 p=3
XM32 VCC_IO 30 NBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=400003 sb=400006 a=0.8 p=3.6
XM33 NBIAS 30 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=400004 sb=400005 a=0.8 p=3.6
XM34 VCC_IO 30 NBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=400005 sb=400004 a=0.8 p=3.6
XM35 39 30 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=400006 sb=400003 a=0.8 p=3.6
XM36 VCC_IO 30 39 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=400007 sb=400002 a=0.8 p=3.6
XM37 39 30 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=400008 sb=400001 a=0.8 p=3.6
XM38 VCC_IO 30 39 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=400009 sb=400000 a=0.8 p=3.6
XM39 34 31 31 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
XM40 35 PU_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=8 W=0.42 AD=0.1113 AS=0.109437 PD=1.37 PS=0.896197 NRD=0 NRS=106.864 m=1 sa=4e+06 sb=4e+06 a=3.36 p=16.84
XM41 30 34 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250004 a=1.5 p=7
XM42 VCC_IO 34 30 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250003 a=1.5 p=7
XM43 30 34 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250003 a=1.5 p=7
XM44 VCC_IO 34 30 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.778125 AS=0.42 PD=4.13625 PS=3.28 NRD=14.9553 NRS=0 m=1 sa=250002 sb=250002 a=1.5 p=7
XM45 11 30 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.29687 PD=5.28 PS=6.89375 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=2.5 p=11
XM46 VCC_IO 30 11 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250000 a=2.5 p=11
R47 EN_H 44 0.01 short m=1
R48 40 PU_H_N 0.01 short m=1
R49 40 31 0.01 short m=1
R50 41 8 0.01 short m=1
R51 42 31 0.01 short m=1
R52 43 34 0.01 short m=1
X60 31 sky130_fd_io__tk_em1o_cdns_5595914180880
X61 NBIAS sky130_fd_io__tk_em1o_cdns_5595914180880
X62 38 NBIAS sky130_fd_io__tk_em1s_cdns_5595914180882
X63 30 35 sky130_fd_io__tk_em1s_cdns_5595914180882
X64 NBIAS 39 sky130_fd_io__tk_em1s_cdns_5595914180881
X65 8 13 sky130_fd_io__tk_em1s_cdns_5595914180881
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_io__gpio_pupredrvr_strongv2 VGND_IO VCC_IO SLOW_H_N PUEN_H DRVHI_H PU_H_N[2] 8 PU_H_N[3] 10 11 12 13 14
**
*.SEEDPROM
XM0 57 SLOW_H_N 37 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=9.6786 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM1 VGND_IO PUEN_H 57 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=9.6786 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM2 46 37 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM3 51 DRVHI_H 40 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.1575 AS=0.3975 PD=1.71 PS=3.53 NRD=3.7962 NRS=0 m=1 sa=250000 sb=250003 a=0.75 p=4
XM4 52 DRVHI_H 40 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.1575 AS=0.3975 PD=1.71 PS=3.53 NRD=3.7962 NRS=0 m=1 sa=250000 sb=250003 a=0.75 p=4
XM5 VGND_IO 38 51 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.5 AD=0.21 AS=0.1575 PD=1.78 PS=1.71 NRD=0 NRS=3.7962 m=1 sa=500000 sb=500002 a=1.5 p=5
XM6 VGND_IO 38 52 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.5 AD=0.21 AS=0.1575 PD=1.78 PS=1.71 NRD=0 NRS=3.7962 m=1 sa=500000 sb=500002 a=1.5 p=5
XM7 47 38 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.5 AD=0.165 AS=0.21 PD=1.72 PS=1.78 NRD=4.1724 NRS=0 m=1 sa=500002 sb=500000 a=1.5 p=5
XM8 48 38 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.5 AD=0.165 AS=0.21 PD=1.72 PS=1.78 NRD=4.1724 NRS=0 m=1 sa=500002 sb=500000 a=1.5 p=5
XM9 40 DRVHI_H 47 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.165 PD=3.53 PS=1.72 NRD=0 NRS=4.1724 m=1 sa=250003 sb=250000 a=0.75 p=4
XM10 40 DRVHI_H 48 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.165 PD=3.53 PS=1.72 NRD=0 NRS=4.1724 m=1 sa=250003 sb=250000 a=0.75 p=4
XM11 PU_H_N[2] DRVHI_H 55 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=4 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 m=1 sa=2e+06 sb=2e+06 a=1.68 p=8.84
XM12 49 DRVHI_H 8 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.165 AS=0.3975 PD=1.72 PS=3.53 NRD=4.1724 NRS=0 m=1 sa=250000 sb=250003 a=0.75 p=4
XM13 50 DRVHI_H 8 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.165 AS=0.3975 PD=1.72 PS=3.53 NRD=4.1724 NRS=0 m=1 sa=250000 sb=250003 a=0.75 p=4
XM14 VGND_IO 42 49 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.5 AD=0.21 AS=0.165 PD=1.78 PS=1.72 NRD=0 NRS=4.1724 m=1 sa=500000 sb=500002 a=1.5 p=5
XM15 VGND_IO 43 50 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.5 AD=0.21 AS=0.165 PD=1.78 PS=1.72 NRD=0 NRS=4.1724 m=1 sa=500000 sb=500002 a=1.5 p=5
XM16 53 44 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.5 AD=0.1575 AS=0.21 PD=1.71 PS=1.78 NRD=3.7962 NRS=0 m=1 sa=500002 sb=500000 a=1.5 p=5
XM17 54 45 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.5 AD=0.1575 AS=0.21 PD=1.71 PS=1.78 NRD=3.7962 NRS=0 m=1 sa=500002 sb=500000 a=1.5 p=5
XM18 56 DRVHI_H PU_H_N[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=4 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 m=1 sa=2e+06 sb=2e+06 a=1.68 p=8.84
XM19 8 DRVHI_H 53 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.1575 PD=3.53 PS=1.71 NRD=0 NRS=3.7962 m=1 sa=250003 sb=250000 a=0.75 p=4
XM20 8 DRVHI_H 54 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.1575 PD=3.53 PS=1.71 NRD=0 NRS=3.7962 m=1 sa=250003 sb=250000 a=0.75 p=4
XM21 37 SLOW_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=1.8 p=7.2
XM22 VCC_IO PUEN_H 37 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=1.8 p=7.2
XM23 46 37 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=1.8 p=7.2
XM24 VCC_IO DRVHI_H PU_H_N[2] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=3 p=11.2
XM25 PU_H_N[2] DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=3 p=11.2
XM26 VCC_IO DRVHI_H PU_H_N[2] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=3 p=11.2
XM27 PU_H_N[2] PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=3 p=11.2
XM28 VCC_IO PUEN_H PU_H_N[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=3 p=11.2
XM29 PU_H_N[3] DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=3 p=11.2
XM30 VCC_IO DRVHI_H PU_H_N[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=3 p=11.2
XM31 PU_H_N[3] DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=3 p=11.2
R32 46 58 0.01 short m=1
R33 46 59 0.01 short m=1
X34 38 sky130_fd_io__tk_em1o_cdns_5595914180880
X35 44 sky130_fd_io__tk_em1o_cdns_5595914180880
X36 38 12 sky130_fd_io__tk_em1s_cdns_5595914180882
X37 40 PU_H_N[2] sky130_fd_io__tk_em1s_cdns_5595914180882
X38 44 12 sky130_fd_io__tk_em1s_cdns_5595914180882
X39 8 PU_H_N[3] sky130_fd_io__tk_em1s_cdns_5595914180882
X55 42 VGND_IO sky130_fd_io__tk_em1o_cdns_55959141808289
X56 43 44 sky130_fd_io__tk_em1o_cdns_55959141808289
X57 45 44 sky130_fd_io__tk_em1o_cdns_55959141808289
X58 42 44 sky130_fd_io__tk_em1s_cdns_55959141808288
X59 VGND_IO 43 sky130_fd_io__tk_em1s_cdns_55959141808288
X60 VGND_IO 45 sky130_fd_io__tk_em1s_cdns_55959141808288
X74 39 PU_H_N[2] sky130_fd_pr__res_generic_po__example_55959141808285
X75 41 PU_H_N[3] sky130_fd_pr__res_generic_po__example_55959141808285
X78 VGND_IO PUEN_H 55 sky130_fd_pr__nfet_01v8__example_55959141808644
X79 VGND_IO PUEN_H 56 sky130_fd_pr__nfet_01v8__example_55959141808644
X80 39 40 sky130_fd_pr__res_generic_po__example_55959141808286
X81 41 8 sky130_fd_pr__res_generic_po__example_55959141808286
X82 VGND_IO VCC_IO 46 12 DRVHI_H PUEN_H 10 PU_H_N[2] 37 14 13 11 sky130_fd_io__feascom_pupredrvr_nbiasv2
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808630 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=4 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 m=1 sa=2e+06 sb=2e+06 a=1.68 p=8.84
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808354 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__pfet_g5v0d10v5 L=4 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 m=1 sa=2e+06 sb=2e+06 a=1.68 p=8.84
.ENDS
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr2 VGND_IO VCC_IO I2C_MODE_H DRVLO_H_N EN_FAST_N[0] EN_FAST_N[1] PDEN_H_N PD_H PD_I2C_H
**
*.SEEDPROM
XM0 PD_H I2C_MODE_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300005 a=1.8 p=7.2
XM1 VGND_IO DRVLO_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300004 a=1.8 p=7.2
XM2 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300003 a=1.8 p=7.2
XM3 VGND_IO PDEN_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300003 sb=300003 a=1.8 p=7.2
XM4 PD_I2C_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300003 sb=300002 a=1.8 p=7.2
XM5 VGND_IO DRVLO_H_N PD_I2C_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300004 sb=300001 a=1.8 p=7.2
XM6 PD_I2C_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300005 sb=300000 a=1.8 p=7.2
XM7 12 I2C_MODE_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=1.5 p=7
XM8 VCC_IO I2C_MODE_H 12 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250001 a=1.5 p=7
XM9 12 I2C_MODE_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=1.5 p=7
XM10 14 DRVLO_H_N PD_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=1.5 p=7
XM11 PD_H DRVLO_H_N 14 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=1.5 p=7
XM12 15 DRVLO_H_N PD_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=1.5 p=7
XM13 PD_H DRVLO_H_N 15 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=1.5 p=7
XM14 12 EN_FAST_N[0] 14 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=1.5 p=7
XM15 15 EN_FAST_N[1] 12 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=1.5 p=7
XM16 VCC_IO EN_FAST_N[1] 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 m=1 sa=500000 sb=500000 a=0.42 p=2.84
XM17 13 DRVLO_H_N PD_I2C_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 sa=500000 sb=500001 a=0.42 p=2.84
XM18 PD_I2C_H DRVLO_H_N 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 sa=500001 sb=500000 a=0.42 p=2.84
X26 VCC_IO PDEN_H_N VCC_IO 17 sky130_fd_pr__pfet_01v8__example_55959141808630
X27 VCC_IO DRVLO_H_N 17 PD_I2C_H sky130_fd_pr__pfet_01v8__example_55959141808630
X33 VCC_IO PDEN_H_N 16 18 sky130_fd_pr__pfet_01v8__example_55959141808354
X34 VCC_IO PDEN_H_N 12 18 sky130_fd_pr__pfet_01v8__example_55959141808354
X35 VCC_IO DRVLO_H_N 16 PD_H sky130_fd_pr__pfet_01v8__example_55959141808354
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808330 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=3 p=11.2
.ENDS
***************************************
***************************************
.SUBCKT sky130_fd_io__com_pdpredrvr_pbiasv2 VGND_IO VCC_IO PD_H DRVLO_H_N PDEN_H_N EN_H_N EN_H 9 PBIAS 11 12 13 14 15
**
*.SEEDPROM
XM0 59 53 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=500000 sb=500008 a=1 p=4
XM1 VGND_IO 53 59 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=500001 sb=500007 a=1 p=4
XM2 54 52 52 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
XM3 PBIAS 53 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=500002 sb=500005 a=1 p=4
XM4 VGND_IO PD_H 14 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=4 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 m=1 sa=2e+06 sb=2e+06 a=1.68 p=8.84
XM5 VGND_IO 53 PBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=500004 sb=500004 a=1 p=4
XM6 60 PD_H 14 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=4 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 m=1 sa=2e+06 sb=2e+06 a=1.68 p=8.84
XM7 54 DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300005 sb=300003 a=0.6 p=3.2
XM8 VGND_IO PDEN_H_N 54 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300006 sb=300003 a=0.6 p=3.2
XM9 53 DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300007 sb=300002 a=0.6 p=3.2
XM10 VGND_IO EN_H_N 53 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300008 sb=300001 a=0.6 p=3.2
XM11 55 DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300009 sb=300000 a=0.6 p=3.2
XM12 56 53 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 m=1 sa=2e+06 sb=2e+06 a=1.68 p=8.84
XM13 57 DRVLO_H_N 53 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.315 AS=0.795 PD=3.21 PS=6.53 NRD=3.1706 NRS=0 m=1 sa=250000 sb=250001 a=1.5 p=7
XM14 55 DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.5 p=3
XM15 58 52 57 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.315 AS=0.315 PD=3.21 PS=3.21 NRD=3.1706 NRS=3.1706 m=1 sa=250001 sb=250001 a=1.5 p=7
XM16 VCC_IO EN_H_N 58 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.315 PD=6.53 PS=3.21 NRD=0 NRS=3.1706 m=1 sa=250001 sb=250000 a=1.5 p=7
XM17 VCC_IO DRVLO_H_N 55 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.5 p=3
XM18 VCC_IO EN_H PBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250006 a=2.5 p=11
XM19 9 9 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250005 a=2.5 p=11
XM20 VCC_IO 9 9 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250005 a=2.5 p=11
XM21 9 9 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250004 a=2.5 p=11
XM22 VCC_IO 9 9 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250003 a=2.5 p=11
XM23 9 9 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250004 sb=250002 a=2.5 p=11
XM24 VCC_IO 9 9 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250002 a=2.5 p=11
XM25 9 9 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250001 a=2.5 p=11
XM26 VCC_IO 9 9 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250006 sb=250000 a=2.5 p=11
XM27 PBIAS PBIAS 9 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250005 a=2.5 p=11
XM28 9 PBIAS PBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250005 a=2.5 p=11
XM29 PBIAS PBIAS 9 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250004 a=2.5 p=11
XM30 9 PBIAS PBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250003 a=2.5 p=11
XM31 PBIAS PBIAS 9 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250002 a=2.5 p=11
XM32 9 PBIAS PBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250004 sb=250002 a=2.5 p=11
XM33 PBIAS PBIAS 9 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250001 a=2.5 p=11
XM34 9 PBIAS PBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250000 a=2.5 p=11
XM35 15 11 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250005 a=2.5 p=11
XM36 VCC_IO 11 15 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250005 a=2.5 p=11
XM37 15 11 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250004 a=2.5 p=11
XM38 VCC_IO 11 15 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250003 a=2.5 p=11
XM39 15 11 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250002 a=2.5 p=11
XM40 VCC_IO 11 15 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250004 sb=250002 a=2.5 p=11
XM41 15 11 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250001 a=2.5 p=11
XM42 VCC_IO 11 15 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250000 a=2.5 p=11
XM43 12 12 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250005 a=2.5 p=11
XM44 13 12 12 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250005 a=2.5 p=11
XM45 12 12 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250004 a=2.5 p=11
XM46 13 12 12 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250003 a=2.5 p=11
XM47 11 13 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250002 a=2.5 p=11
XM48 13 13 11 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250004 sb=250002 a=2.5 p=11
XM49 11 13 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250001 a=2.5 p=11
XM50 11 VGND_IO VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=8 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 m=1 sa=4e+06 sb=4e+06 a=3.36 p=16.84
XM51 13 13 11 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250000 a=2.5 p=11
XM52 VCC_IO 55 11 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=2.5 p=11
XM53 PBIAS 55 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=2.5 p=11
R54 61 52 0.01 short m=1
R55 62 54 0.01 short m=1
R56 52 63 0.01 short m=1
R57 64 EN_H_N 0.01 short m=1
X58 52 PD_H sky130_fd_io__tk_em1s_cdns_5595914180882
X59 59 PBIAS sky130_fd_io__tk_em1s_cdns_5595914180882
X60 PBIAS 9 sky130_fd_io__tk_em1o_cdns_5595914180879
X61 9 15 sky130_fd_io__tk_em1s_cdns_5595914180881
X64 60 53 sky130_fd_io__tk_em1s_cdns_55959141808288
X65 PBIAS 56 sky130_fd_io__tk_em1s_cdns_55959141808288
X85 VGND_IO 53 12 sky130_fd_pr__nfet_01v8__example_55959141808330
X86 VGND_IO 54 53 sky130_fd_pr__nfet_01v8__example_55959141808330
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong VGND VGND_IO VCC_IO PD_H[4] I2C_MODE_H_N PDEN_H_N 7 PD_H[3] DRVLO_H_N SLOW_H 11 12 13 14 15 16 17 PD_H[2]
**
*.SEEDPROM
XM0 VGND PD_H[4] 65 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.21 p=1.84
XM1 VGND 74 60 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.42 p=2.6
XM2 VGND 75 62 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.42 p=2.6
XM3 567 I2C_MODE_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=13.8396 NRS=0 m=1 sa=300001 sb=300001 a=0.42 p=2.6
XM4 568 59 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=13.8396 NRS=0 m=1 sa=300001 sb=300001 a=0.42 p=2.6
XM5 59 I2C_MODE_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.1855 PD=1.93 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.42 p=2.6
XM6 74 SLOW_H 567 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300002 sb=300000 a=0.42 p=2.6
XM7 75 SLOW_H 568 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300002 sb=300000 a=0.42 p=2.6
XM8 7 59 65 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=1.5 p=7
XM9 DRVLO_H_N I2C_MODE_H_N 7 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=1.5 p=7
XM10 61 PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.335 PD=1.28 PS=2.67 NRD=0 NRS=7.9686 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM11 VGND_IO 60 61 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.21 AS=0.14 PD=1.42 PS=1.28 NRD=7.9686 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM12 66 61 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.21 PD=2.53 PS=1.42 NRD=0 NRS=7.9686 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM13 VGND_IO 7 PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300005 a=1.8 p=7.2
XM14 PD_H[3] 7 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300004 a=1.8 p=7.2
XM15 VGND_IO 7 PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300003 a=1.8 p=7.2
XM16 PD_H[3] 7 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300003 sb=300003 a=1.8 p=7.2
XM17 VGND_IO 7 PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300003 sb=300002 a=1.8 p=7.2
XM18 PD_H[3] PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300004 sb=300001 a=1.8 p=7.2
XM19 VGND_IO PDEN_H_N PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300005 sb=300000 a=1.8 p=7.2
XM20 VCC_IO PD_H[4] 65 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
XM21 VCC_IO 74 60 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM22 VCC_IO 74 60 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM23 VCC_IO 75 62 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM24 VCC_IO 75 62 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM25 74 I2C_MODE_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM26 74 I2C_MODE_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM27 75 59 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM28 75 59 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM29 59 I2C_MODE_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.6 p=3.2
XM30 59 I2C_MODE_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.6 p=3.2
XM31 VCC_IO SLOW_H 74 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM32 VCC_IO SLOW_H 74 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM33 VCC_IO SLOW_H 75 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM34 VCC_IO SLOW_H 75 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM35 7 59 DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=1.5 p=7
XM36 65 I2C_MODE_H_N 7 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=1.5 p=7
XM37 73 PDEN_H_N 61 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=1.005 PD=3.28 PS=6.67 NRD=5.4053 NRS=4.4503 m=1 sa=300000 sb=300002 a=1.8 p=7.2
XM38 VCC_IO 60 73 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.63 AS=0.42 PD=3.42 PS=3.28 NRD=4.4503 NRS=5.4053 m=1 sa=300001 sb=300001 a=1.8 p=7.2
XM39 66 61 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.63 PD=6.53 PS=3.42 NRD=0 NRS=4.4503 m=1 sa=300002 sb=300000 a=1.8 p=7.2
XM40 VCC_IO 62 67 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.5 p=3
XM41 67 62 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.5 p=3
XM42 PD_H[3] 7 69 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=0.75 p=4
XM43 70 7 PD_H[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=0.75 p=4
XM44 VCC_IO 63 70 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=0.75 p=4
XM45 68 63 67 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.21 p=1.84
XM46 69 64 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=0.75 p=4
XM47 67 64 68 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.21 p=1.84
XM48 PD_H[3] 7 71 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=2 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 sa=999999 sb=1e+06 a=0.84 p=4.84
XM49 PD_H[3] 7 68 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.21 p=1.84
XM50 68 7 PD_H[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.21 p=1.84
XM51 72 7 PD_H[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=2 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 sa=1e+06 sb=1e+06 a=0.84 p=4.84
XM52 67 PDEN_H_N 72 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=2 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 sa=1e+06 sb=999999 a=0.84 p=4.84
R53 77 66 0.01 short m=1
R54 66 78 0.01 short m=1
R55 79 64 0.01 short m=1
X72 76 sky130_fd_io__tk_em1o_cdns_5595914180880
X73 63 sky130_fd_io__tk_em1o_cdns_5595914180880
X74 63 sky130_fd_io__tk_em1o_cdns_5595914180880
X75 76 11 sky130_fd_io__tk_em1s_cdns_5595914180882
X76 63 11 sky130_fd_io__tk_em1s_cdns_5595914180882
X77 64 VCC_IO sky130_fd_io__tk_em1s_cdns_5595914180882
X89 VCC_IO PDEN_H_N VCC_IO 71 sky130_fd_pr__pfet_01v8__example_55959141808630
X96 VGND_IO VCC_IO 62 DRVLO_H_N 11 11 PDEN_H_N PD_H[2] PD_H[4] sky130_fd_io__gpiov2_pdpredrvr_strong_nr2
X99 VGND_IO VCC_IO PD_H[4] DRVLO_H_N PDEN_H_N 66 61 13 11 17 16 15 12 14 sky130_fd_io__com_pdpredrvr_pbiasv2
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_obpredrvr VGND VGND_IO VCC_IO DRVHI_H PUEN_H[0] DRVLO_H_N PDEN_H_N[0] PDEN_H_N[1] PUEN_H[1] PD_H[0] PU_H_N[1] PU_H_N[0] 13 PD_H[1] PD_H[3] 16 17 18 19 20
+ PU_H_N[2] 22 23 24 25 26 27 28 29 SLOW_H_N PU_H_N[3] I2C_MODE_H_N SLOW_H PD_H[2] PD_H[4] 36
**
*.SEEDPROM
XM0 104 DRVHI_H PU_H_N[0] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM1 VGND_IO PUEN_H[0] 104 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
XM2 PD_H[0] DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM3 VGND_IO PDEN_H_N[0] PD_H[0] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
XM4 PD_H[1] PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM5 VGND_IO DRVLO_H_N PD_H[1] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
XM6 PU_H_N[1] DRVHI_H 13 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=1.8 p=7.2
XM7 13 DRVHI_H PU_H_N[1] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=1.8 p=7.2
XM8 VGND_IO PUEN_H[1] 13 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=1.8 p=7.2
XM9 13 PUEN_H[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=1.8 p=7.2
XM10 PU_H_N[0] DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=3 p=11.2
XM11 VCC_IO DRVHI_H PU_H_N[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=3 p=11.2
XM12 PU_H_N[0] PUEN_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=3 p=11.2
XM13 102 DRVLO_H_N PD_H[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=1.8 p=7.2
XM14 VCC_IO PDEN_H_N[0] 102 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=1.8 p=7.2
XM15 102 PDEN_H_N[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=1.8 p=7.2
XM16 VCC_IO PDEN_H_N[1] 103 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=1.5 p=7
XM17 103 PDEN_H_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=1.5 p=7
XM18 PD_H[1] DRVLO_H_N 103 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=1.5 p=7
XM19 103 DRVLO_H_N PD_H[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=1.5 p=7
XM20 VCC_IO DRVHI_H PU_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=1.5 p=7
XM21 PU_H_N[1] DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=1.5 p=7
XM22 VCC_IO DRVHI_H PU_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=1.5 p=7
XM23 PU_H_N[1] PUEN_H[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=1.5 p=7
X24 VGND_IO VCC_IO condiode a=1e-06 p=0.004 m=1
X25 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2dn a=1211.58 p=164.72 m=1
X26 VGND_IO VCC_IO sky130_fd_pr__model__parasitic__diode_pw2dn a=453.842 p=155.65 m=1
X52 VGND_IO VCC_IO SLOW_H_N PUEN_H[1] DRVHI_H PU_H_N[2] 22 PU_H_N[3] 16 17 18 19 20 sky130_fd_io__gpio_pupredrvr_strongv2
X53 VGND VGND_IO VCC_IO PD_H[4] I2C_MODE_H_N PDEN_H_N[1] 36 PD_H[3] DRVLO_H_N SLOW_H 23 29 28 27 25 26 24 PD_H[2] sky130_fd_io__gpiov2_pdpredrvr_strong
.ENDS
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__com_ctl_ls_octl SET_H VCC_IO VPB 4 HLD_H_N IN RST_H OUT_H_N OUT_H
**
*.SEEDPROM
XM0 14 12 SET_H SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=75000.2 sb=75003.2 a=0.15 p=2.3
XM1 SET_H 12 14 SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75000.6 sb=75002.8 a=0.15 p=2.3
XM2 14 12 SET_H SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.1 sb=75002.3 a=0.15 p=2.3
XM3 SET_H 12 14 SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.5 sb=75001.9 a=0.15 p=2.3
XM4 16 4 SET_H SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.9 sb=75001.5 a=0.15 p=2.3
XM5 SET_H 4 16 SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.4 sb=75001 a=0.15 p=2.3
XM6 16 4 SET_H SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.8 sb=75000.6 a=0.15 p=2.3
XM7 SET_H 4 16 SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=75003.2 sb=75000.2 a=0.15 p=2.3
XM8 SET_H 10 OUT_H_N SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM9 OUT_H 11 SET_H SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM10 13 HLD_H_N 11 SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=1.8 p=7.2
XM11 10 HLD_H_N 15 SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=1.8 p=7.2
XM12 SET_H RST_H 10 SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=1.8 p=7.2
XM13 11 SET_H SET_H SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=1.8 p=7.2
XM14 VCC_IO 11 OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM15 OUT_H_N 10 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
X16 SET_H VPB sky130_fd_pr__model__parasitic__diode_ps2nw a=3.1672 p=7.24 m=1
X17 VPB IN 4 VPB 12 sky130_fd_pr__pfet_01v8__example_55959141808430
X20 SET_H 4 IN 12 sky130_fd_pr__nfet_01v8__example_55959141808423
X22 SET_H 11 10 sky130_fd_pr__nfet_01v8__example_55959141808424
X26 SET_H VPB 14 13 sky130_fd_pr__nfet_01v8__example_55959141808426
X27 SET_H VPB 14 13 sky130_fd_pr__nfet_01v8__example_55959141808426
X28 SET_H VPB 16 15 sky130_fd_pr__nfet_01v8__example_55959141808426
X29 SET_H VPB 16 15 sky130_fd_pr__nfet_01v8__example_55959141808426
X34 VCC_IO 10 11 sky130_fd_pr__pfet_01v8__example_55959141808435
X35 VCC_IO 11 10 sky130_fd_pr__pfet_01v8__example_55959141808433
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_octl VGND VCC_IO DM_H[2] DM_H[0] 6 DM_H[1] 8 DM_H_N[1] DM_H_N[2] DM_H_N[0] 12 13 PDEN_H_N[0] PDEN_H_N[1] VPWR SLOW_H SLOW_H_N HLD_I_H_N SLOW OD_H
**
*.SEEDPROM
XM0 35 DM_H[0] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.196 PD=0.98 PS=1.96 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.42 p=2.6
XM1 VGND DM_H[1] 35 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.42 p=2.6
XM2 718 DM_H[2] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=13.8396 NRS=0 m=1 sa=300002 sb=300001 a=0.42 p=2.6
XM3 8 35 718 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300003 sb=300000 a=0.42 p=2.6
XM4 36 DM_H_N[1] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.196 PD=0.98 PS=1.96 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM5 719 VCC_IO 37 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM6 VGND DM_H[2] 23 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300004 a=0.42 p=2.6
XM7 VGND DM_H[2] 24 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300004 a=0.42 p=2.6
XM8 VGND DM_H_N[2] 36 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM9 VGND PUEN_2OR1_H 719 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM10 31 DM_H[2] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.42 p=2.6
XM11 32 DM_H[2] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.42 p=2.6
XM12 26 DM_H[0] 31 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300003 a=0.42 p=2.6
XM13 28 DM_H[1] 32 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300003 a=0.42 p=2.6
XM14 720 36 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM15 721 DM_H[0] 39 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300003 a=0.42 p=2.6
XM16 33 6 26 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300002 a=0.42 p=2.6
XM17 34 22 28 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300002 a=0.42 p=2.6
XM18 40 DM_H_N[0] 720 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM19 VGND DM_H[1] 721 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300002 a=0.42 p=2.6
XM20 VGND 23 33 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.42 p=2.6
XM21 VGND 24 34 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.42 p=2.6
XM22 722 DM_H_N[2] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=13.8396 NRS=0 m=1 sa=300002 sb=300001 a=0.42 p=2.6
XM23 6 DM_H[0] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300004 sb=300000 a=0.42 p=2.6
XM24 723 40 PUEN_2OR1_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300003 a=0.42 p=2.6
XM25 22 DM_H[1] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300004 sb=300000 a=0.42 p=2.6
XM26 41 DM_H_N[1] 722 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300003 sb=300000 a=0.42 p=2.6
XM27 VGND 42 723 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300002 a=0.42 p=2.6
XM28 724 28 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=13.8396 NRS=0 m=1 sa=300002 sb=300001 a=0.42 p=2.6
XM29 725 41 44 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM30 43 DM_H_N[1] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.196 PD=0.98 PS=1.96 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.42 p=2.6
XM31 45 37 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.1855 PD=1.93 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.42 p=2.6
XM32 42 DM_H[0] 724 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300003 sb=300000 a=0.42 p=2.6
XM33 VGND DM_H_N[0] 725 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM34 VGND 26 43 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.42 p=2.6
XM35 12 48 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.42 p=2.6
XM36 VGND 39 46 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.42 p=2.6
XM37 VGND 44 47 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.42 p=2.6
XM38 13 49 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300002 a=0.42 p=2.6
XM39 VGND 48 12 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.42 p=2.6
XM40 PDEN_H_N[0] 46 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.42 p=2.6
XM41 PDEN_H_N[1] 47 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.42 p=2.6
XM42 VGND 49 13 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.42 p=2.6
XM43 48 45 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.42 p=2.6
XM44 VGND 46 PDEN_H_N[0] VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.42 p=2.6
XM45 VGND 47 PDEN_H_N[1] VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.42 p=2.6
XM46 49 43 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300004 sb=300000 a=0.42 p=2.6
XM47 715 DM_H[0] 35 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM48 715 DM_H[0] 35 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM49 VCC_IO DM_H[1] 715 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM50 VCC_IO DM_H[1] 715 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM51 8 DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM52 8 DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM53 VCC_IO 35 8 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM54 VCC_IO 35 8 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM55 716 DM_H_N[1] 36 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM56 716 DM_H_N[1] 36 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM57 37 VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM58 37 VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM59 VCC_IO DM_H[2] 23 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300004 a=0.6 p=3.2
XM60 VCC_IO DM_H[2] 23 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300004 a=0.6 p=3.2
XM61 VCC_IO DM_H[2] 24 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300004 a=0.6 p=3.2
XM62 VCC_IO DM_H[2] 24 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300004 a=0.6 p=3.2
XM63 VCC_IO DM_H_N[2] 716 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM64 VCC_IO DM_H_N[2] 716 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM65 VCC_IO PUEN_2OR1_H 37 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM66 VCC_IO PUEN_2OR1_H 37 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM67 25 DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.6 p=3.2
XM68 25 DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.6 p=3.2
XM69 27 DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.6 p=3.2
XM70 27 DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.6 p=3.2
XM71 26 6 25 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300003 a=0.6 p=3.2
XM72 26 6 25 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300003 a=0.6 p=3.2
XM73 28 22 27 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300003 a=0.6 p=3.2
XM74 28 22 27 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300003 a=0.6 p=3.2
XM75 40 36 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM76 40 36 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM77 39 DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM78 39 DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM79 29 23 26 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300002 a=0.6 p=3.2
XM80 29 23 26 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300002 a=0.6 p=3.2
XM81 30 24 28 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300002 a=0.6 p=3.2
XM82 30 24 28 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300002 a=0.6 p=3.2
XM83 VCC_IO DM_H_N[0] 40 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM84 VCC_IO DM_H_N[0] 40 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM85 VCC_IO DM_H[1] 39 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM86 VCC_IO DM_H[1] 39 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM87 VCC_IO DM_H[0] 29 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.6 p=3.2
XM88 VCC_IO DM_H[0] 29 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.6 p=3.2
XM89 VCC_IO DM_H[1] 30 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.6 p=3.2
XM90 VCC_IO DM_H[1] 30 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.6 p=3.2
XM91 41 DM_H_N[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM92 41 DM_H_N[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM93 6 DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300000 a=0.6 p=3.2
XM94 6 DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300000 a=0.6 p=3.2
XM95 PUEN_2OR1_H 40 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM96 PUEN_2OR1_H 40 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM97 22 DM_H[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300000 a=0.6 p=3.2
XM98 22 DM_H[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300000 a=0.6 p=3.2
XM99 VCC_IO DM_H_N[1] 41 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM100 VCC_IO DM_H_N[1] 41 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM101 VCC_IO 42 PUEN_2OR1_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM102 VCC_IO 42 PUEN_2OR1_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM103 42 28 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM104 42 28 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM105 44 41 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM106 44 41 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM107 717 DM_H_N[1] 43 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM108 717 DM_H_N[1] 43 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM109 45 37 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.6 p=3.2
XM110 45 37 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.6 p=3.2
XM111 VCC_IO DM_H[0] 42 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM112 VCC_IO DM_H[0] 42 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM113 VCC_IO DM_H_N[0] 44 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM114 VCC_IO DM_H_N[0] 44 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM115 VCC_IO 26 717 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.6 p=3.2
XM116 VCC_IO 26 717 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.6 p=3.2
XM117 12 48 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM118 12 48 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM119 VCC_IO 39 46 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM120 VCC_IO 39 46 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM121 VCC_IO 44 47 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM122 VCC_IO 44 47 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM123 13 49 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300002 a=0.6 p=3.2
XM124 13 49 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300002 a=0.6 p=3.2
XM125 VCC_IO 48 12 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM126 VCC_IO 48 12 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM127 PDEN_H_N[0] 46 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM128 PDEN_H_N[0] 46 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM129 PDEN_H_N[1] 47 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM130 PDEN_H_N[1] 47 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM131 VCC_IO 49 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.6 p=3.2
XM132 VCC_IO 49 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.6 p=3.2
XM133 48 45 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM134 48 45 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM135 VCC_IO 46 PDEN_H_N[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM136 VCC_IO 46 PDEN_H_N[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM137 VCC_IO 47 PDEN_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM138 VCC_IO 47 PDEN_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM139 49 43 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM140 49 43 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
X189 VGND VCC_IO VPWR 50 HLD_I_H_N SLOW OD_H SLOW_H_N SLOW_H sky130_fd_io__com_ctl_ls_octl
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808389 2 3 4 5
**
*.SEEDPROM
XM0 2 3 5 2 sky130_fd_pr__pfet_01v8_hvt L=0.25 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=125000 sb=125001 a=0.75 p=6.5
XM1 3 4 2 2 sky130_fd_pr__pfet_01v8_hvt L=0.25 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=125001 sb=125000 a=0.75 p=6.5
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808375 1 2 3 4
**
XM0 4 2 1 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=125000 sb=125002 a=0.25 p=2.5
XM1 1 2 4 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.25 p=2.5
XM2 2 3 1 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=125001 sb=125001 a=0.25 p=2.5
XM3 1 3 2 1 sky130_fd_pr__nfet_01v8 L=0.25 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=125002 sb=125000 a=0.25 p=2.5
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808387 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=450000 sb=450000 a=0.9 p=3.8
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808388 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=75000.2 sb=75000.6 a=0.15 p=2.3
XM1 1 2 3 1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=75000.6 sb=75000.2 a=0.15 p=2.3
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6
**
X0 1 2 4 5 sky130_fd_pr__nfet_01v8__example_55959141808387
X1 1 3 6 sky130_fd_pr__nfet_01v8__example_55959141808388
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808376 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=2.5 p=11
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808377 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=1.4 PD=10.53 PS=10.56 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=2.5 p=11
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808386 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=450000 sb=450001 a=0.9 p=3.8
XM1 3 2 4 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=450001 sb=450000 a=0.9 p=3.8
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808391 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.5 p=3
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808390 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.5 p=3
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_dat_lsv2 VGND VCC_IO VPWR_KA 4 RST_H SET_H HLD_H_N IN OUT_H OUT_H_N
**
*.SEEDPROM
XM0 VGND 22 OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM1 OUT_H_N 4 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM2 VGND 22 4 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM3 VGND RST_H 4 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM4 22 4 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM5 22 SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
XM6 VCC_IO 4 OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=1.5 p=7
XM7 OUT_H 22 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=1.5 p=7
X14 VPWR_KA 24 IN 23 sky130_fd_pr__pfet_01v8__example_55959141808389
X15 VGND 24 IN 23 sky130_fd_pr__nfet_01v8__example_55959141808375
X16 VGND VPWR_KA 23 27 28 26 ICV_8
X17 VGND VPWR_KA 23 27 28 26 ICV_8
X18 VGND VPWR_KA 23 27 28 26 ICV_8
X19 VGND VPWR_KA 23 27 28 26 ICV_8
X20 VGND VPWR_KA 24 27 28 28 ICV_8
X21 VGND VPWR_KA 24 27 28 28 ICV_8
X22 VGND VPWR_KA 24 27 28 28 ICV_8
X23 VGND VPWR_KA 24 27 28 28 ICV_8
X24 VGND HLD_H_N 4 27 sky130_fd_pr__nfet_01v8__example_55959141808376
X25 VGND HLD_H_N 25 22 sky130_fd_pr__nfet_01v8__example_55959141808377
X26 VGND VPWR_KA 25 26 sky130_fd_pr__nfet_01v8__example_55959141808386
X27 VGND VPWR_KA 25 26 sky130_fd_pr__nfet_01v8__example_55959141808386
X28 VGND VPWR_KA 25 26 sky130_fd_pr__nfet_01v8__example_55959141808386
X29 VGND VPWR_KA 25 26 sky130_fd_pr__nfet_01v8__example_55959141808386
X35 VCC_IO 22 4 sky130_fd_pr__pfet_01v8__example_55959141808391
X36 VCC_IO 4 22 sky130_fd_pr__pfet_01v8__example_55959141808390
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_dat_ls_1v2 VGND VCC_IO VPWR_KA RST_H SET_H HLD_H_N IN OUT_H OUT_H_N
**
*.SEEDPROM
XM0 VGND 20 OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM1 OUT_H_N 21 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM2 VGND 20 21 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM3 VGND RST_H 21 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM4 20 21 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM5 20 SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
XM6 VCC_IO 21 OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=1.5 p=7
XM7 OUT_H 20 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=1.5 p=7
X14 VPWR_KA 23 IN 22 sky130_fd_pr__pfet_01v8__example_55959141808389
X15 VGND 23 IN 22 sky130_fd_pr__nfet_01v8__example_55959141808375
X16 VGND VPWR_KA 22 26 27 25 ICV_8
X17 VGND VPWR_KA 22 26 27 25 ICV_8
X18 VGND VPWR_KA 22 26 27 25 ICV_8
X19 VGND VPWR_KA 22 26 27 25 ICV_8
X20 VGND VPWR_KA 23 26 27 27 ICV_8
X21 VGND VPWR_KA 23 26 27 27 ICV_8
X22 VGND VPWR_KA 23 26 27 27 ICV_8
X23 VGND VPWR_KA 23 26 27 27 ICV_8
X24 VGND HLD_H_N 21 26 sky130_fd_pr__nfet_01v8__example_55959141808376
X25 VGND HLD_H_N 24 20 sky130_fd_pr__nfet_01v8__example_55959141808377
X26 VGND VPWR_KA 24 25 sky130_fd_pr__nfet_01v8__example_55959141808386
X27 VGND VPWR_KA 24 25 sky130_fd_pr__nfet_01v8__example_55959141808386
X28 VGND VPWR_KA 24 25 sky130_fd_pr__nfet_01v8__example_55959141808386
X29 VGND VPWR_KA 24 25 sky130_fd_pr__nfet_01v8__example_55959141808386
X35 VCC_IO 20 21 sky130_fd_pr__pfet_01v8__example_55959141808391
X36 VCC_IO 21 20 sky130_fd_pr__pfet_01v8__example_55959141808390
.ENDS
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__com_cclat VGND VCC_IO OE_H_N PU_DIS_H DRVLO_H_N DRVHI_H PD_DIS_H
**
*.SEEDPROM
XM0 VGND OE_H_N 12 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM1 16 12 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
XM2 VGND PU_DIS_H 13 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=1.8 p=7.2
XM3 19 12 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=1.8 p=7.2
XM4 VGND 12 19 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300002 a=1.8 p=7.2
XM5 19 12 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=1.8 p=7.2
XM6 VGND 12 19 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=1.8 p=7.2
XM7 19 DRVLO_H_N 20 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=1.8 p=7.2
XM8 20 DRVLO_H_N 19 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=1.8 p=7.2
XM9 14 13 20 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=1.8 p=7.2
XM10 20 13 14 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=1.8 p=7.2
XM11 DRVLO_H_N 15 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300015 a=1.8 p=7.2
XM12 VGND 15 DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300014 a=1.8 p=7.2
XM13 DRVLO_H_N 15 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300013 a=1.8 p=7.2
XM14 VGND 15 DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300003 sb=300012 a=1.8 p=7.2
XM15 DRVLO_H_N 15 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300003 sb=300011 a=1.8 p=7.2
XM16 VGND 15 DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300004 sb=300011 a=1.8 p=7.2
XM17 DRVHI_H 14 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300005 sb=300010 a=1.8 p=7.2
XM18 VGND 14 DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300006 sb=300009 a=1.8 p=7.2
XM19 DRVHI_H 14 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300007 sb=300008 a=1.8 p=7.2
XM20 VGND 14 DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300008 sb=300007 a=1.8 p=7.2
XM21 DRVHI_H 14 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300009 sb=300006 a=1.8 p=7.2
XM22 VGND 14 DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300010 sb=300005 a=1.8 p=7.2
XM23 15 16 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300011 sb=300004 a=1.8 p=7.2
XM24 VGND 16 15 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300011 sb=300003 a=1.8 p=7.2
XM25 15 DRVHI_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300012 sb=300003 a=1.8 p=7.2
XM26 VGND DRVHI_H 15 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300013 sb=300002 a=1.8 p=7.2
XM27 15 PD_DIS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300014 sb=300001 a=1.8 p=7.2
XM28 VGND PD_DIS_H 15 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300015 sb=300000 a=1.8 p=7.2
XM29 VCC_IO OE_H_N 12 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=2.5 p=11
XM30 16 12 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=2.5 p=11
XM31 VCC_IO PU_DIS_H 13 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=2.5 p=11
XM32 14 12 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=2.5 p=11
XM33 VCC_IO 13 14 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=2.5 p=11
XM34 14 DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=2.5 p=11
XM35 DRVHI_H 14 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250016 a=2.5 p=11
XM36 VCC_IO 14 DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250015 a=2.5 p=11
XM37 DRVHI_H 14 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250014 a=2.5 p=11
XM38 VCC_IO 14 DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250013 a=2.5 p=11
XM39 DRVHI_H 14 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250013 a=2.5 p=11
XM40 VCC_IO 14 DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250004 sb=250012 a=2.5 p=11
XM41 DRVLO_H_N 15 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250011 a=2.5 p=11
XM42 VCC_IO 15 DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250010 a=2.5 p=11
XM43 DRVLO_H_N 15 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250006 sb=250009 a=2.5 p=11
XM44 VCC_IO 15 DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250007 sb=250009 a=2.5 p=11
XM45 DRVLO_H_N 15 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250008 sb=250008 a=2.5 p=11
XM46 VCC_IO 15 DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250009 sb=250007 a=2.5 p=11
XM47 17 16 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300009 sb=300006 a=3 p=11.2
XM48 VCC_IO 16 17 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300010 sb=300005 a=3 p=11.2
XM49 17 16 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300011 sb=300004 a=3 p=11.2
XM50 VCC_IO 16 17 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300012 sb=300003 a=3 p=11.2
XM51 17 16 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300013 sb=300003 a=3 p=11.2
XM52 VCC_IO 16 17 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300014 sb=300002 a=3 p=11.2
XM53 17 16 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=300015 sb=300001 a=3 p=11.2
XM54 VCC_IO 16 17 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=300015 sb=300000 a=3 p=11.2
XM55 17 DRVHI_H 18 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250005 a=2.5 p=11
XM56 18 DRVHI_H 17 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250005 a=2.5 p=11
XM57 17 DRVHI_H 18 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250004 a=2.5 p=11
XM58 18 DRVHI_H 17 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250003 a=2.5 p=11
XM59 15 PD_DIS_H 18 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250003 sb=250002 a=2.5 p=11
XM60 18 PD_DIS_H 15 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250004 sb=250002 a=2.5 p=11
XM61 15 PD_DIS_H 18 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250001 a=2.5 p=11
XM62 18 PD_DIS_H 15 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250005 sb=250000 a=2.5 p=11
.ENDS
***************************************
.SUBCKT sky130_fd_io__com_opath_datoev2 VGND VCC_IO VPWR_KA HLD_I_OVR_H OD_H 6 OE_N DRVHI_H DRVLO_H_N OUT
**
*.SEEDPROM
X0 VGND VPWR_KA sky130_fd_pr__model__parasitic__diode_ps2nw a=13.8768 p=14.98 m=1
X1 VGND VCC_IO VPWR_KA 11 VGND OD_H HLD_I_OVR_H OE_N 12 OE_H sky130_fd_io__gpio_dat_lsv2
X2 VGND VCC_IO VPWR_KA VGND OD_H HLD_I_OVR_H OUT 6 13 sky130_fd_io__gpio_dat_ls_1v2
X5 VGND VCC_IO 12 13 DRVLO_H_N DRVHI_H 6 sky130_fd_io__com_cclat
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpiov2_octl_dat VGND VGND_IO VCC_IO 5 PD_H[3] OD_H 8 9 10 11 12 13 14 15 16 17 18 PU_H_N[2] 20 PU_H_N[0]
+ PD_H[0] 23 PD_H[1] PU_H_N[1] DM_H[0] DM_H[1] DM_H[2] PU_H_N[3] PD_H[2] PD_H[4] DM_H_N[1] VPWR HLD_I_H_N SLOW VPWR_KA OE_N HLD_I_OVR_H DM_H_N[0] DM_H_N[2] OUT
+ 42
**
*.SEEDPROM
X0 VGND VGND_IO VCC_IO DRVHI_H 109 DRVLO_H_N 110 111 116 PD_H[0] PU_H_N[1] PU_H_N[0] 5 PD_H[1] PD_H[3] 12 13 15 16 18
+ PU_H_N[2] 20 8 9 10 11 14 17 23 SLOW_H_N PU_H_N[3] 117 113 PD_H[2] PD_H[4] 42
+ sky130_fd_io__gpiov2_obpredrvr
X1 VGND VCC_IO DM_H[2] DM_H[0] 108 DM_H[1] 117 DM_H_N[1] DM_H_N[2] DM_H_N[0] 116 109 110 111 VPWR 113 SLOW_H_N HLD_I_H_N SLOW OD_H sky130_fd_io__gpiov2_octl
X2 VGND VCC_IO VPWR_KA HLD_I_OVR_H OD_H 114 OE_N DRVHI_H DRVLO_H_N OUT sky130_fd_io__com_opath_datoev2
.ENDS
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__com_ctl_ls SET_H VCC_IO VPB VPWR HLD_H_N IN RST_H OUT_H
**
*.SEEDPROM
XM0 22 18 SET_H SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=75000.2 sb=75003.2 a=0.15 p=2.3
XM1 SET_H 18 22 SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75000.6 sb=75002.8 a=0.15 p=2.3
XM2 22 18 SET_H SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.1 sb=75002.3 a=0.15 p=2.3
XM3 SET_H 18 22 SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.5 sb=75001.9 a=0.15 p=2.3
XM4 24 19 SET_H SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75001.9 sb=75001.5 a=0.15 p=2.3
XM5 SET_H 19 24 SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.4 sb=75001 a=0.15 p=2.3
XM6 24 19 SET_H SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=75002.8 sb=75000.6 a=0.15 p=2.3
XM7 SET_H 19 24 SET_H sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=75003.2 sb=75000.2 a=0.15 p=2.3
XM8 SET_H 16 OUT_H_N SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM9 OUT_H 17 SET_H SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM10 20 HLD_H_N 17 SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=1.8 p=7.2
XM11 16 HLD_H_N 23 SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=1.8 p=7.2
XM12 SET_H RST_H 16 SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=1.8 p=7.2
XM13 17 SET_H SET_H SET_H sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=1.8 p=7.2
XM14 VCC_IO 17 OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=1.8 p=7.2
XM15 OUT_H_N 16 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=1.8 p=7.2
X16 SET_H VPB sky130_fd_pr__model__parasitic__diode_ps2nw a=3.1672 p=7.24 m=1
X17 VPB IN 19 VPWR 18 sky130_fd_pr__pfet_01v8__example_55959141808430
X20 SET_H 19 IN 18 sky130_fd_pr__nfet_01v8__example_55959141808423
X22 SET_H 17 16 sky130_fd_pr__nfet_01v8__example_55959141808424
X26 SET_H VPWR 22 20 sky130_fd_pr__nfet_01v8__example_55959141808426
X27 SET_H VPWR 22 20 sky130_fd_pr__nfet_01v8__example_55959141808426
X28 SET_H VPWR 24 23 sky130_fd_pr__nfet_01v8__example_55959141808426
X29 SET_H VPWR 24 23 sky130_fd_pr__nfet_01v8__example_55959141808426
X34 VCC_IO 16 17 sky130_fd_pr__pfet_01v8__example_55959141808435
X35 VCC_IO 17 16 sky130_fd_pr__pfet_01v8__example_55959141808433
.ENDS
***************************************
***************************************
***************************************
.SUBCKT sky130_fd_io__com_ctl_hldv2 VGND VCC_IO 3 4 5 OD_I_H HLD_I_H HLD_OVR HLD_I_H_N VPWR
**
*.SEEDPROM
XM0 VGND 3 19 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.42 p=2.6
XM1 508 3 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=13.8396 NRS=0 m=1 sa=300001 sb=300001 a=0.42 p=2.6
XM2 20 4 508 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300002 sb=300000 a=0.42 p=2.6
XM3 21 20 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.1855 PD=1.93 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.42 p=2.6
XM4 18 21 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300017 a=0.42 p=2.6
XM5 VGND 21 18 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300016 a=0.42 p=2.6
XM6 18 21 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300015 a=0.42 p=2.6
XM7 VGND 21 18 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300014 a=0.42 p=2.6
XM8 22 18 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300013 a=0.42 p=2.6
XM9 VGND 18 22 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300004 sb=300012 a=0.42 p=2.6
XM10 22 18 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300005 sb=300011 a=0.42 p=2.6
XM11 VGND 18 22 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300006 sb=300011 a=0.42 p=2.6
XM12 22 18 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300007 sb=300010 a=0.42 p=2.6
XM13 VGND 18 22 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300008 sb=300009 a=0.42 p=2.6
XM14 22 18 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300009 sb=300008 a=0.42 p=2.6
XM15 VGND 18 22 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300010 sb=300007 a=0.42 p=2.6
XM16 23 18 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300011 sb=300006 a=0.42 p=2.6
XM17 VGND 18 23 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300011 sb=300005 a=0.42 p=2.6
XM18 23 18 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300012 sb=300004 a=0.42 p=2.6
XM19 VGND 18 23 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300013 sb=300003 a=0.42 p=2.6
XM20 23 18 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300014 sb=300003 a=0.42 p=2.6
XM21 VGND 18 23 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300015 sb=300002 a=0.42 p=2.6
XM22 23 18 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300016 sb=300001 a=0.42 p=2.6
XM23 VGND 18 23 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300017 sb=300000 a=0.42 p=2.6
XM24 VGND 19 24 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.42 p=2.6
XM25 OD_I_H 24 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.42 p=2.6
XM26 VGND 24 OD_I_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300002 a=0.42 p=2.6
XM27 OD_I_H 24 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.42 p=2.6
XM28 VGND 24 OD_I_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.42 p=2.6
XM29 5 25 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.196 PD=0.98 PS=1.96 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.42 p=2.6
XM30 VGND OD_I_H 5 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.42 p=2.6
XM31 25 21 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.42 p=2.6
XM32 VGND 26 25 VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.196 AS=0.098 PD=1.96 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.42 p=2.6
XM33 VCC_IO 3 19 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM34 VCC_IO 3 19 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM35 20 3 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM36 20 3 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM37 VCC_IO 4 20 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM38 VCC_IO 4 20 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM39 21 20 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.6 p=3.2
XM40 21 20 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.6 p=3.2
XM41 18 21 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300017 a=0.6 p=3.2
XM42 18 21 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300017 a=0.6 p=3.2
XM43 VCC_IO 21 18 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300016 a=0.6 p=3.2
XM44 VCC_IO 21 18 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300016 a=0.6 p=3.2
XM45 18 21 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300015 a=0.6 p=3.2
XM46 18 21 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300015 a=0.6 p=3.2
XM47 VCC_IO 21 18 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300014 a=0.6 p=3.2
XM48 VCC_IO 21 18 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300014 a=0.6 p=3.2
XM49 22 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300013 a=0.6 p=3.2
XM50 22 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300013 a=0.6 p=3.2
XM51 VCC_IO 18 22 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300012 a=0.6 p=3.2
XM52 VCC_IO 18 22 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300012 a=0.6 p=3.2
XM53 22 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300005 sb=300011 a=0.6 p=3.2
XM54 22 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300005 sb=300011 a=0.6 p=3.2
XM55 VCC_IO 18 22 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300006 sb=300011 a=0.6 p=3.2
XM56 VCC_IO 18 22 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300006 sb=300011 a=0.6 p=3.2
XM57 22 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300007 sb=300010 a=0.6 p=3.2
XM58 22 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300007 sb=300010 a=0.6 p=3.2
XM59 VCC_IO 18 22 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300008 sb=300009 a=0.6 p=3.2
XM60 VCC_IO 18 22 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300008 sb=300009 a=0.6 p=3.2
XM61 22 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300009 sb=300008 a=0.6 p=3.2
XM62 22 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300009 sb=300008 a=0.6 p=3.2
XM63 VCC_IO 18 22 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300010 sb=300007 a=0.6 p=3.2
XM64 VCC_IO 18 22 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300010 sb=300007 a=0.6 p=3.2
XM65 23 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300011 sb=300006 a=0.6 p=3.2
XM66 23 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300011 sb=300006 a=0.6 p=3.2
XM67 VCC_IO 18 23 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300011 sb=300005 a=0.6 p=3.2
XM68 VCC_IO 18 23 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300011 sb=300005 a=0.6 p=3.2
XM69 23 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300012 sb=300004 a=0.6 p=3.2
XM70 23 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300012 sb=300004 a=0.6 p=3.2
XM71 VCC_IO 18 23 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300013 sb=300003 a=0.6 p=3.2
XM72 VCC_IO 18 23 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300013 sb=300003 a=0.6 p=3.2
XM73 23 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300014 sb=300003 a=0.6 p=3.2
XM74 23 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300014 sb=300003 a=0.6 p=3.2
XM75 VCC_IO 18 23 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300015 sb=300002 a=0.6 p=3.2
XM76 VCC_IO 18 23 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300015 sb=300002 a=0.6 p=3.2
XM77 23 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300016 sb=300001 a=0.6 p=3.2
XM78 23 18 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300016 sb=300001 a=0.6 p=3.2
XM79 VCC_IO 18 23 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300017 sb=300000 a=0.6 p=3.2
XM80 VCC_IO 18 23 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300017 sb=300000 a=0.6 p=3.2
XM81 VCC_IO 19 24 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM82 VCC_IO 19 24 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM83 OD_I_H 24 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.6 p=3.2
XM84 OD_I_H 24 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300003 a=0.6 p=3.2
XM85 VCC_IO 24 OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300002 a=0.6 p=3.2
XM86 VCC_IO 24 OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300002 a=0.6 p=3.2
XM87 OD_I_H 24 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.6 p=3.2
XM88 OD_I_H 24 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300001 a=0.6 p=3.2
XM89 VCC_IO 24 OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM90 VCC_IO 24 OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM91 506 25 5 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM92 506 25 5 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM93 VCC_IO OD_I_H 506 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM94 VCC_IO OD_I_H 506 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM95 507 21 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM96 507 21 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM97 25 26 507 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM98 25 26 507 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
R99 HLD_I_H 18 0.01 short m=1
R100 22 HLD_I_H_N 0.01 short m=1
R101 HLD_I_H_N 23 0.01 short m=1
X110 VGND VCC_IO VPWR VPWR 21 HLD_OVR 19 26 sky130_fd_io__com_ctl_ls
.ENDS
***************************************
.SUBCKT sky130_ef_io__gpiov2_pad_wrapped  VSSD VSSIO VSSA VSSIO_Q VDDIO VDDIO_Q PAD_A_ESD_1_H PAD PAD_A_ESD_0_H IB_MODE_SEL ENABLE_INP_H ENABLE_H VDDA ENABLE_VDDA_H VCCD OE_N VTRIP_SEL VCCHIB ENABLE_VSWITCH_H OUT
+ HLD_OVR DM[2] ANALOG_SEL HLD_H_N ANALOG_EN INP_DIS ANALOG_POL DM[0] PAD_A_NOESD_H DM[1] SLOW TIE_HI_ESD IN IN_H ENABLE_VDDIO TIE_LO_ESD VSWITCH AMUXBUS_A AMUXBUS_B
**
XM0 4111 ENABLE_INP_H 33 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300002 a=0.42 p=2.6
XM1 VSSD 34 4111 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300001 a=0.42 p=2.6
XM2 35 33 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.42 p=2.6
XM3 37 ENABLE_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.196 PD=0.98 PS=1.96 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM4 VSSD ENABLE_INP_H 37 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM5 33 ENABLE_INP_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM6 33 ENABLE_INP_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300002 a=0.6 p=3.2
XM7 VDDIO_Q 34 33 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM8 VDDIO_Q 34 33 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300001 a=0.6 p=3.2
XM9 35 33 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM10 35 33 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300000 a=0.6 p=3.2
XM11 4110 ENABLE_H 37 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM12 4110 ENABLE_H 37 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM13 VDDIO_Q ENABLE_INP_H 4110 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM14 VDDIO_Q ENABLE_INP_H 4110 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
X15 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw a=384.91 p=0 m=1
X16 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw a=560.026 p=0 m=1
X17 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=12.9015 p=14.37 m=1
X18 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=67.5428 p=62.24 m=1
X19 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=33.634 p=25.7 m=1
X20 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=237.836 p=101.02 m=1
X21 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=215.42 p=130.01 m=1
X22 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw a=785.678 p=181.15 m=1
R23 PAD_A_NOESD_H PAD 0.01 short m=1
R24 PAD_A_NOESD_H PAD 0.01 short m=1
R25 PAD_A_NOESD_H PAD 0.01 short m=1
X26 PAD_A_ESD_1_H 12 sky130_fd_io__res75only_small
X27 12 PAD sky130_fd_io__res75only_small
X28 14 PAD sky130_fd_io__res75only_small
X29 PAD_A_ESD_0_H 14 sky130_fd_io__res75only_small
X33 VSSD VSSA VSSIO_Q 3 2 6 8 VSWITCH VDDIO_Q VDDA 60 PAD ENABLE_VDDA_H VCCD 85 ENABLE_VSWITCH_H AMUXBUS_B AMUXBUS_A ANALOG_SEL ANALOG_EN
+ OUT ANALOG_POL 56
+ sky130_fd_io__gpiov2_amux
X34 VSSD VDDIO_Q VCCD IB_MODE_SEL 56 34 75 73 39 71 37 DM[0] INP_DIS 35 70 63 65 DM[2] 55 90
+ VTRIP_SEL 47 48 DM[1]
+ sky130_fd_io__gpiov2_ctl_lsbank
X35 VSSD VSSIO VDDIO 43 45 PAD 44 46 76 TIE_HI_ESD 30 69 17 TIE_LO_ESD 81 sky130_fd_io__gpio_odrvrv2
X36 VSSD VDDIO_Q ENABLE_VDDIO 39 83 IN_H 82 49 PAD 84 IN VCCHIB 73 63 70 47 48 55 sky130_fd_io__gpiov2_ipath
X37 VSSD VSSIO VDDIO 16 17 34 19 20 21 22 23 24 25 26 27 29 28 30 31 43
+ 44 38 45 46 71 75 65 76 69 81 73 VCCD 56 SLOW VCCHIB OE_N 50 39 63 OUT
+ 91
+ sky130_fd_io__gpiov2_octl_dat
X38 VSSD VDDIO_Q ENABLE_H HLD_H_N 50 34 60 HLD_OVR 56 VCCD sky130_fd_io__com_ctl_hldv2
.ENDS
***************************************
