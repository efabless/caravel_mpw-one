VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3481.340 2.400 3482.540 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3182.140 2.400 3183.340 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2882.260 2.400 2883.460 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2583.060 2.400 2584.260 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2283.180 2.400 2284.380 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2433.460 2924.800 2434.660 ;
    END
  END io_in[10]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2903.340 2924.800 2904.540 ;
    END
  END io_in[12]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3406.540 2.400 3407.740 ;
    END
  END io_in[24]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3331.740 2.400 3332.940 ;
    END
  END io_out[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3107.340 2.400 3108.540 ;
    END
  END io_in[25]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3032.540 2.400 3033.740 ;
    END
  END io_out[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2807.460 2.400 2808.660 ;
    END
  END io_in[26]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2732.660 2.400 2733.860 ;
    END
  END io_out[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_in[27]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2433.460 2.400 2434.660 ;
    END
  END io_out[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2208.380 2.400 2209.580 ;
    END
  END io_in[28]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2133.580 2.400 2134.780 ;
    END
  END io_out[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1983.980 2.400 1985.180 ;
    END
  END io_in[29]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1909.180 2.400 1910.380 ;
    END
  END io_out[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END io_in[30]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1684.100 2.400 1685.300 ;
    END
  END io_out[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1534.500 2.400 1535.700 ;
    END
  END io_in[31]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1459.700 2.400 1460.900 ;
    END
  END io_out[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1310.100 2.400 1311.300 ;
    END
  END io_in[32]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1235.300 2.400 1236.500 ;
    END
  END io_out[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1085.020 2.400 1086.220 ;
    END
  END io_in[33]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1010.220 2.400 1011.420 ;
    END
  END io_out[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 860.620 2.400 861.820 ;
    END
  END io_in[34]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 785.820 2.400 787.020 ;
    END
  END io_out[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 636.220 2.400 637.420 ;
    END
  END io_in[35]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 560.740 2.400 561.940 ;
    END
  END io_out[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 411.140 2.400 412.340 ;
    END
  END io_in[36]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 336.340 2.400 337.540 ;
    END
  END io_out[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 186.740 2.400 187.940 ;
    END
  END io_in[37]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 111.940 2.400 113.140 ;
    END
  END io_out[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1964.260 2924.800 1965.460 ;
    END
  END io_in[8]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2198.860 2924.800 2200.060 ;
    END
  END io_in[9]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3256.940 2.400 3258.140 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2957.060 2.400 2958.260 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2657.860 2.400 2659.060 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2357.980 2.400 2359.180 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2058.780 2.400 2059.980 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1834.380 2.400 1835.580 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1609.300 2.400 1610.500 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1384.900 2.400 1386.100 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1159.820 2.400 1161.020 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 935.420 2.400 936.620 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 711.020 2.400 712.220 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 485.940 2.400 487.140 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 261.540 2.400 262.740 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 37.140 2.400 38.340 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 9.020 -9.320 12.020 3529.000 ;
        RECT 189.020 -9.320 192.020 3529.000 ;
        RECT 369.020 -9.320 372.020 3529.000 ;
        RECT 549.020 -9.320 552.020 3529.000 ;
        RECT 729.020 -9.320 732.020 3529.000 ;
        RECT 909.020 -9.320 912.020 3529.000 ;
        RECT 1089.020 -9.320 1092.020 3529.000 ;
        RECT 1269.020 -9.320 1272.020 3529.000 ;
        RECT 1449.020 -9.320 1452.020 3529.000 ;
        RECT 1629.020 -9.320 1632.020 3529.000 ;
        RECT 1809.020 -9.320 1812.020 3529.000 ;
        RECT 1989.020 -9.320 1992.020 3529.000 ;
        RECT 2169.020 -9.320 2172.020 3529.000 ;
        RECT 2349.020 -9.320 2352.020 3529.000 ;
        RECT 2529.020 -9.320 2532.020 3529.000 ;
        RECT 2709.020 -9.320 2712.020 3529.000 ;
        RECT 2889.020 -9.320 2892.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3436.090 -7.890 3437.270 ;
        RECT -9.070 3434.490 -7.890 3435.670 ;
        RECT -9.070 3256.090 -7.890 3257.270 ;
        RECT -9.070 3254.490 -7.890 3255.670 ;
        RECT -9.070 3076.090 -7.890 3077.270 ;
        RECT -9.070 3074.490 -7.890 3075.670 ;
        RECT -9.070 2896.090 -7.890 2897.270 ;
        RECT -9.070 2894.490 -7.890 2895.670 ;
        RECT -9.070 2716.090 -7.890 2717.270 ;
        RECT -9.070 2714.490 -7.890 2715.670 ;
        RECT -9.070 2536.090 -7.890 2537.270 ;
        RECT -9.070 2534.490 -7.890 2535.670 ;
        RECT -9.070 2356.090 -7.890 2357.270 ;
        RECT -9.070 2354.490 -7.890 2355.670 ;
        RECT -9.070 2176.090 -7.890 2177.270 ;
        RECT -9.070 2174.490 -7.890 2175.670 ;
        RECT -9.070 1996.090 -7.890 1997.270 ;
        RECT -9.070 1994.490 -7.890 1995.670 ;
        RECT -9.070 1816.090 -7.890 1817.270 ;
        RECT -9.070 1814.490 -7.890 1815.670 ;
        RECT -9.070 1636.090 -7.890 1637.270 ;
        RECT -9.070 1634.490 -7.890 1635.670 ;
        RECT -9.070 1456.090 -7.890 1457.270 ;
        RECT -9.070 1454.490 -7.890 1455.670 ;
        RECT -9.070 1276.090 -7.890 1277.270 ;
        RECT -9.070 1274.490 -7.890 1275.670 ;
        RECT -9.070 1096.090 -7.890 1097.270 ;
        RECT -9.070 1094.490 -7.890 1095.670 ;
        RECT -9.070 916.090 -7.890 917.270 ;
        RECT -9.070 914.490 -7.890 915.670 ;
        RECT -9.070 736.090 -7.890 737.270 ;
        RECT -9.070 734.490 -7.890 735.670 ;
        RECT -9.070 556.090 -7.890 557.270 ;
        RECT -9.070 554.490 -7.890 555.670 ;
        RECT -9.070 376.090 -7.890 377.270 ;
        RECT -9.070 374.490 -7.890 375.670 ;
        RECT -9.070 196.090 -7.890 197.270 ;
        RECT -9.070 194.490 -7.890 195.670 ;
        RECT -9.070 16.090 -7.890 17.270 ;
        RECT -9.070 14.490 -7.890 15.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 9.930 3523.010 11.110 3524.190 ;
        RECT 9.930 3521.410 11.110 3522.590 ;
        RECT 9.930 3436.090 11.110 3437.270 ;
        RECT 9.930 3434.490 11.110 3435.670 ;
        RECT 9.930 3256.090 11.110 3257.270 ;
        RECT 9.930 3254.490 11.110 3255.670 ;
        RECT 9.930 3076.090 11.110 3077.270 ;
        RECT 9.930 3074.490 11.110 3075.670 ;
        RECT 9.930 2896.090 11.110 2897.270 ;
        RECT 9.930 2894.490 11.110 2895.670 ;
        RECT 9.930 2716.090 11.110 2717.270 ;
        RECT 9.930 2714.490 11.110 2715.670 ;
        RECT 9.930 2536.090 11.110 2537.270 ;
        RECT 9.930 2534.490 11.110 2535.670 ;
        RECT 9.930 2356.090 11.110 2357.270 ;
        RECT 9.930 2354.490 11.110 2355.670 ;
        RECT 9.930 2176.090 11.110 2177.270 ;
        RECT 9.930 2174.490 11.110 2175.670 ;
        RECT 9.930 1996.090 11.110 1997.270 ;
        RECT 9.930 1994.490 11.110 1995.670 ;
        RECT 9.930 1816.090 11.110 1817.270 ;
        RECT 9.930 1814.490 11.110 1815.670 ;
        RECT 9.930 1636.090 11.110 1637.270 ;
        RECT 9.930 1634.490 11.110 1635.670 ;
        RECT 9.930 1456.090 11.110 1457.270 ;
        RECT 9.930 1454.490 11.110 1455.670 ;
        RECT 9.930 1276.090 11.110 1277.270 ;
        RECT 9.930 1274.490 11.110 1275.670 ;
        RECT 9.930 1096.090 11.110 1097.270 ;
        RECT 9.930 1094.490 11.110 1095.670 ;
        RECT 9.930 916.090 11.110 917.270 ;
        RECT 9.930 914.490 11.110 915.670 ;
        RECT 9.930 736.090 11.110 737.270 ;
        RECT 9.930 734.490 11.110 735.670 ;
        RECT 9.930 556.090 11.110 557.270 ;
        RECT 9.930 554.490 11.110 555.670 ;
        RECT 9.930 376.090 11.110 377.270 ;
        RECT 9.930 374.490 11.110 375.670 ;
        RECT 9.930 196.090 11.110 197.270 ;
        RECT 9.930 194.490 11.110 195.670 ;
        RECT 9.930 16.090 11.110 17.270 ;
        RECT 9.930 14.490 11.110 15.670 ;
        RECT 9.930 -2.910 11.110 -1.730 ;
        RECT 9.930 -4.510 11.110 -3.330 ;
        RECT 189.930 3523.010 191.110 3524.190 ;
        RECT 189.930 3521.410 191.110 3522.590 ;
        RECT 189.930 3436.090 191.110 3437.270 ;
        RECT 189.930 3434.490 191.110 3435.670 ;
        RECT 189.930 3256.090 191.110 3257.270 ;
        RECT 189.930 3254.490 191.110 3255.670 ;
        RECT 189.930 3076.090 191.110 3077.270 ;
        RECT 189.930 3074.490 191.110 3075.670 ;
        RECT 189.930 2896.090 191.110 2897.270 ;
        RECT 189.930 2894.490 191.110 2895.670 ;
        RECT 189.930 2716.090 191.110 2717.270 ;
        RECT 189.930 2714.490 191.110 2715.670 ;
        RECT 189.930 2536.090 191.110 2537.270 ;
        RECT 189.930 2534.490 191.110 2535.670 ;
        RECT 189.930 2356.090 191.110 2357.270 ;
        RECT 189.930 2354.490 191.110 2355.670 ;
        RECT 189.930 2176.090 191.110 2177.270 ;
        RECT 189.930 2174.490 191.110 2175.670 ;
        RECT 189.930 1996.090 191.110 1997.270 ;
        RECT 189.930 1994.490 191.110 1995.670 ;
        RECT 189.930 1816.090 191.110 1817.270 ;
        RECT 189.930 1814.490 191.110 1815.670 ;
        RECT 189.930 1636.090 191.110 1637.270 ;
        RECT 189.930 1634.490 191.110 1635.670 ;
        RECT 189.930 1456.090 191.110 1457.270 ;
        RECT 189.930 1454.490 191.110 1455.670 ;
        RECT 189.930 1276.090 191.110 1277.270 ;
        RECT 189.930 1274.490 191.110 1275.670 ;
        RECT 189.930 1096.090 191.110 1097.270 ;
        RECT 189.930 1094.490 191.110 1095.670 ;
        RECT 189.930 916.090 191.110 917.270 ;
        RECT 189.930 914.490 191.110 915.670 ;
        RECT 189.930 736.090 191.110 737.270 ;
        RECT 189.930 734.490 191.110 735.670 ;
        RECT 189.930 556.090 191.110 557.270 ;
        RECT 189.930 554.490 191.110 555.670 ;
        RECT 189.930 376.090 191.110 377.270 ;
        RECT 189.930 374.490 191.110 375.670 ;
        RECT 189.930 196.090 191.110 197.270 ;
        RECT 189.930 194.490 191.110 195.670 ;
        RECT 189.930 16.090 191.110 17.270 ;
        RECT 189.930 14.490 191.110 15.670 ;
        RECT 189.930 -2.910 191.110 -1.730 ;
        RECT 189.930 -4.510 191.110 -3.330 ;
        RECT 369.930 3523.010 371.110 3524.190 ;
        RECT 369.930 3521.410 371.110 3522.590 ;
        RECT 369.930 3436.090 371.110 3437.270 ;
        RECT 369.930 3434.490 371.110 3435.670 ;
        RECT 369.930 3256.090 371.110 3257.270 ;
        RECT 369.930 3254.490 371.110 3255.670 ;
        RECT 369.930 3076.090 371.110 3077.270 ;
        RECT 369.930 3074.490 371.110 3075.670 ;
        RECT 369.930 2896.090 371.110 2897.270 ;
        RECT 369.930 2894.490 371.110 2895.670 ;
        RECT 369.930 2716.090 371.110 2717.270 ;
        RECT 369.930 2714.490 371.110 2715.670 ;
        RECT 369.930 2536.090 371.110 2537.270 ;
        RECT 369.930 2534.490 371.110 2535.670 ;
        RECT 369.930 2356.090 371.110 2357.270 ;
        RECT 369.930 2354.490 371.110 2355.670 ;
        RECT 369.930 2176.090 371.110 2177.270 ;
        RECT 369.930 2174.490 371.110 2175.670 ;
        RECT 369.930 1996.090 371.110 1997.270 ;
        RECT 369.930 1994.490 371.110 1995.670 ;
        RECT 369.930 1816.090 371.110 1817.270 ;
        RECT 369.930 1814.490 371.110 1815.670 ;
        RECT 369.930 1636.090 371.110 1637.270 ;
        RECT 369.930 1634.490 371.110 1635.670 ;
        RECT 369.930 1456.090 371.110 1457.270 ;
        RECT 369.930 1454.490 371.110 1455.670 ;
        RECT 369.930 1276.090 371.110 1277.270 ;
        RECT 369.930 1274.490 371.110 1275.670 ;
        RECT 369.930 1096.090 371.110 1097.270 ;
        RECT 369.930 1094.490 371.110 1095.670 ;
        RECT 369.930 916.090 371.110 917.270 ;
        RECT 369.930 914.490 371.110 915.670 ;
        RECT 369.930 736.090 371.110 737.270 ;
        RECT 369.930 734.490 371.110 735.670 ;
        RECT 369.930 556.090 371.110 557.270 ;
        RECT 369.930 554.490 371.110 555.670 ;
        RECT 369.930 376.090 371.110 377.270 ;
        RECT 369.930 374.490 371.110 375.670 ;
        RECT 369.930 196.090 371.110 197.270 ;
        RECT 369.930 194.490 371.110 195.670 ;
        RECT 369.930 16.090 371.110 17.270 ;
        RECT 369.930 14.490 371.110 15.670 ;
        RECT 369.930 -2.910 371.110 -1.730 ;
        RECT 369.930 -4.510 371.110 -3.330 ;
        RECT 549.930 3523.010 551.110 3524.190 ;
        RECT 549.930 3521.410 551.110 3522.590 ;
        RECT 549.930 3436.090 551.110 3437.270 ;
        RECT 549.930 3434.490 551.110 3435.670 ;
        RECT 549.930 3256.090 551.110 3257.270 ;
        RECT 549.930 3254.490 551.110 3255.670 ;
        RECT 549.930 3076.090 551.110 3077.270 ;
        RECT 549.930 3074.490 551.110 3075.670 ;
        RECT 549.930 2896.090 551.110 2897.270 ;
        RECT 549.930 2894.490 551.110 2895.670 ;
        RECT 549.930 2716.090 551.110 2717.270 ;
        RECT 549.930 2714.490 551.110 2715.670 ;
        RECT 549.930 2536.090 551.110 2537.270 ;
        RECT 549.930 2534.490 551.110 2535.670 ;
        RECT 549.930 2356.090 551.110 2357.270 ;
        RECT 549.930 2354.490 551.110 2355.670 ;
        RECT 549.930 2176.090 551.110 2177.270 ;
        RECT 549.930 2174.490 551.110 2175.670 ;
        RECT 549.930 1996.090 551.110 1997.270 ;
        RECT 549.930 1994.490 551.110 1995.670 ;
        RECT 549.930 1816.090 551.110 1817.270 ;
        RECT 549.930 1814.490 551.110 1815.670 ;
        RECT 549.930 1636.090 551.110 1637.270 ;
        RECT 549.930 1634.490 551.110 1635.670 ;
        RECT 549.930 1456.090 551.110 1457.270 ;
        RECT 549.930 1454.490 551.110 1455.670 ;
        RECT 549.930 1276.090 551.110 1277.270 ;
        RECT 549.930 1274.490 551.110 1275.670 ;
        RECT 549.930 1096.090 551.110 1097.270 ;
        RECT 549.930 1094.490 551.110 1095.670 ;
        RECT 549.930 916.090 551.110 917.270 ;
        RECT 549.930 914.490 551.110 915.670 ;
        RECT 549.930 736.090 551.110 737.270 ;
        RECT 549.930 734.490 551.110 735.670 ;
        RECT 549.930 556.090 551.110 557.270 ;
        RECT 549.930 554.490 551.110 555.670 ;
        RECT 549.930 376.090 551.110 377.270 ;
        RECT 549.930 374.490 551.110 375.670 ;
        RECT 549.930 196.090 551.110 197.270 ;
        RECT 549.930 194.490 551.110 195.670 ;
        RECT 549.930 16.090 551.110 17.270 ;
        RECT 549.930 14.490 551.110 15.670 ;
        RECT 549.930 -2.910 551.110 -1.730 ;
        RECT 549.930 -4.510 551.110 -3.330 ;
        RECT 729.930 3523.010 731.110 3524.190 ;
        RECT 729.930 3521.410 731.110 3522.590 ;
        RECT 729.930 3436.090 731.110 3437.270 ;
        RECT 729.930 3434.490 731.110 3435.670 ;
        RECT 729.930 3256.090 731.110 3257.270 ;
        RECT 729.930 3254.490 731.110 3255.670 ;
        RECT 729.930 3076.090 731.110 3077.270 ;
        RECT 729.930 3074.490 731.110 3075.670 ;
        RECT 729.930 2896.090 731.110 2897.270 ;
        RECT 729.930 2894.490 731.110 2895.670 ;
        RECT 729.930 2716.090 731.110 2717.270 ;
        RECT 729.930 2714.490 731.110 2715.670 ;
        RECT 729.930 2536.090 731.110 2537.270 ;
        RECT 729.930 2534.490 731.110 2535.670 ;
        RECT 729.930 2356.090 731.110 2357.270 ;
        RECT 729.930 2354.490 731.110 2355.670 ;
        RECT 729.930 2176.090 731.110 2177.270 ;
        RECT 729.930 2174.490 731.110 2175.670 ;
        RECT 729.930 1996.090 731.110 1997.270 ;
        RECT 729.930 1994.490 731.110 1995.670 ;
        RECT 729.930 1816.090 731.110 1817.270 ;
        RECT 729.930 1814.490 731.110 1815.670 ;
        RECT 729.930 1636.090 731.110 1637.270 ;
        RECT 729.930 1634.490 731.110 1635.670 ;
        RECT 729.930 1456.090 731.110 1457.270 ;
        RECT 729.930 1454.490 731.110 1455.670 ;
        RECT 729.930 1276.090 731.110 1277.270 ;
        RECT 729.930 1274.490 731.110 1275.670 ;
        RECT 729.930 1096.090 731.110 1097.270 ;
        RECT 729.930 1094.490 731.110 1095.670 ;
        RECT 729.930 916.090 731.110 917.270 ;
        RECT 729.930 914.490 731.110 915.670 ;
        RECT 729.930 736.090 731.110 737.270 ;
        RECT 729.930 734.490 731.110 735.670 ;
        RECT 729.930 556.090 731.110 557.270 ;
        RECT 729.930 554.490 731.110 555.670 ;
        RECT 729.930 376.090 731.110 377.270 ;
        RECT 729.930 374.490 731.110 375.670 ;
        RECT 729.930 196.090 731.110 197.270 ;
        RECT 729.930 194.490 731.110 195.670 ;
        RECT 729.930 16.090 731.110 17.270 ;
        RECT 729.930 14.490 731.110 15.670 ;
        RECT 729.930 -2.910 731.110 -1.730 ;
        RECT 729.930 -4.510 731.110 -3.330 ;
        RECT 909.930 3523.010 911.110 3524.190 ;
        RECT 909.930 3521.410 911.110 3522.590 ;
        RECT 909.930 3436.090 911.110 3437.270 ;
        RECT 909.930 3434.490 911.110 3435.670 ;
        RECT 909.930 3256.090 911.110 3257.270 ;
        RECT 909.930 3254.490 911.110 3255.670 ;
        RECT 909.930 3076.090 911.110 3077.270 ;
        RECT 909.930 3074.490 911.110 3075.670 ;
        RECT 909.930 2896.090 911.110 2897.270 ;
        RECT 909.930 2894.490 911.110 2895.670 ;
        RECT 909.930 2716.090 911.110 2717.270 ;
        RECT 909.930 2714.490 911.110 2715.670 ;
        RECT 909.930 2536.090 911.110 2537.270 ;
        RECT 909.930 2534.490 911.110 2535.670 ;
        RECT 909.930 2356.090 911.110 2357.270 ;
        RECT 909.930 2354.490 911.110 2355.670 ;
        RECT 909.930 2176.090 911.110 2177.270 ;
        RECT 909.930 2174.490 911.110 2175.670 ;
        RECT 909.930 1996.090 911.110 1997.270 ;
        RECT 909.930 1994.490 911.110 1995.670 ;
        RECT 909.930 1816.090 911.110 1817.270 ;
        RECT 909.930 1814.490 911.110 1815.670 ;
        RECT 909.930 1636.090 911.110 1637.270 ;
        RECT 909.930 1634.490 911.110 1635.670 ;
        RECT 909.930 1456.090 911.110 1457.270 ;
        RECT 909.930 1454.490 911.110 1455.670 ;
        RECT 909.930 1276.090 911.110 1277.270 ;
        RECT 909.930 1274.490 911.110 1275.670 ;
        RECT 909.930 1096.090 911.110 1097.270 ;
        RECT 909.930 1094.490 911.110 1095.670 ;
        RECT 909.930 916.090 911.110 917.270 ;
        RECT 909.930 914.490 911.110 915.670 ;
        RECT 909.930 736.090 911.110 737.270 ;
        RECT 909.930 734.490 911.110 735.670 ;
        RECT 909.930 556.090 911.110 557.270 ;
        RECT 909.930 554.490 911.110 555.670 ;
        RECT 909.930 376.090 911.110 377.270 ;
        RECT 909.930 374.490 911.110 375.670 ;
        RECT 909.930 196.090 911.110 197.270 ;
        RECT 909.930 194.490 911.110 195.670 ;
        RECT 909.930 16.090 911.110 17.270 ;
        RECT 909.930 14.490 911.110 15.670 ;
        RECT 909.930 -2.910 911.110 -1.730 ;
        RECT 909.930 -4.510 911.110 -3.330 ;
        RECT 1089.930 3523.010 1091.110 3524.190 ;
        RECT 1089.930 3521.410 1091.110 3522.590 ;
        RECT 1089.930 3436.090 1091.110 3437.270 ;
        RECT 1089.930 3434.490 1091.110 3435.670 ;
        RECT 1089.930 3256.090 1091.110 3257.270 ;
        RECT 1089.930 3254.490 1091.110 3255.670 ;
        RECT 1089.930 3076.090 1091.110 3077.270 ;
        RECT 1089.930 3074.490 1091.110 3075.670 ;
        RECT 1089.930 2896.090 1091.110 2897.270 ;
        RECT 1089.930 2894.490 1091.110 2895.670 ;
        RECT 1089.930 2716.090 1091.110 2717.270 ;
        RECT 1089.930 2714.490 1091.110 2715.670 ;
        RECT 1089.930 2536.090 1091.110 2537.270 ;
        RECT 1089.930 2534.490 1091.110 2535.670 ;
        RECT 1089.930 2356.090 1091.110 2357.270 ;
        RECT 1089.930 2354.490 1091.110 2355.670 ;
        RECT 1089.930 2176.090 1091.110 2177.270 ;
        RECT 1089.930 2174.490 1091.110 2175.670 ;
        RECT 1089.930 1996.090 1091.110 1997.270 ;
        RECT 1089.930 1994.490 1091.110 1995.670 ;
        RECT 1089.930 1816.090 1091.110 1817.270 ;
        RECT 1089.930 1814.490 1091.110 1815.670 ;
        RECT 1089.930 1636.090 1091.110 1637.270 ;
        RECT 1089.930 1634.490 1091.110 1635.670 ;
        RECT 1089.930 1456.090 1091.110 1457.270 ;
        RECT 1089.930 1454.490 1091.110 1455.670 ;
        RECT 1089.930 1276.090 1091.110 1277.270 ;
        RECT 1089.930 1274.490 1091.110 1275.670 ;
        RECT 1089.930 1096.090 1091.110 1097.270 ;
        RECT 1089.930 1094.490 1091.110 1095.670 ;
        RECT 1089.930 916.090 1091.110 917.270 ;
        RECT 1089.930 914.490 1091.110 915.670 ;
        RECT 1089.930 736.090 1091.110 737.270 ;
        RECT 1089.930 734.490 1091.110 735.670 ;
        RECT 1089.930 556.090 1091.110 557.270 ;
        RECT 1089.930 554.490 1091.110 555.670 ;
        RECT 1089.930 376.090 1091.110 377.270 ;
        RECT 1089.930 374.490 1091.110 375.670 ;
        RECT 1089.930 196.090 1091.110 197.270 ;
        RECT 1089.930 194.490 1091.110 195.670 ;
        RECT 1089.930 16.090 1091.110 17.270 ;
        RECT 1089.930 14.490 1091.110 15.670 ;
        RECT 1089.930 -2.910 1091.110 -1.730 ;
        RECT 1089.930 -4.510 1091.110 -3.330 ;
        RECT 1269.930 3523.010 1271.110 3524.190 ;
        RECT 1269.930 3521.410 1271.110 3522.590 ;
        RECT 1269.930 3436.090 1271.110 3437.270 ;
        RECT 1269.930 3434.490 1271.110 3435.670 ;
        RECT 1269.930 3256.090 1271.110 3257.270 ;
        RECT 1269.930 3254.490 1271.110 3255.670 ;
        RECT 1269.930 3076.090 1271.110 3077.270 ;
        RECT 1269.930 3074.490 1271.110 3075.670 ;
        RECT 1269.930 2896.090 1271.110 2897.270 ;
        RECT 1269.930 2894.490 1271.110 2895.670 ;
        RECT 1269.930 2716.090 1271.110 2717.270 ;
        RECT 1269.930 2714.490 1271.110 2715.670 ;
        RECT 1269.930 2536.090 1271.110 2537.270 ;
        RECT 1269.930 2534.490 1271.110 2535.670 ;
        RECT 1269.930 2356.090 1271.110 2357.270 ;
        RECT 1269.930 2354.490 1271.110 2355.670 ;
        RECT 1269.930 2176.090 1271.110 2177.270 ;
        RECT 1269.930 2174.490 1271.110 2175.670 ;
        RECT 1269.930 1996.090 1271.110 1997.270 ;
        RECT 1269.930 1994.490 1271.110 1995.670 ;
        RECT 1269.930 1816.090 1271.110 1817.270 ;
        RECT 1269.930 1814.490 1271.110 1815.670 ;
        RECT 1269.930 1636.090 1271.110 1637.270 ;
        RECT 1269.930 1634.490 1271.110 1635.670 ;
        RECT 1269.930 1456.090 1271.110 1457.270 ;
        RECT 1269.930 1454.490 1271.110 1455.670 ;
        RECT 1269.930 1276.090 1271.110 1277.270 ;
        RECT 1269.930 1274.490 1271.110 1275.670 ;
        RECT 1269.930 1096.090 1271.110 1097.270 ;
        RECT 1269.930 1094.490 1271.110 1095.670 ;
        RECT 1269.930 916.090 1271.110 917.270 ;
        RECT 1269.930 914.490 1271.110 915.670 ;
        RECT 1269.930 736.090 1271.110 737.270 ;
        RECT 1269.930 734.490 1271.110 735.670 ;
        RECT 1269.930 556.090 1271.110 557.270 ;
        RECT 1269.930 554.490 1271.110 555.670 ;
        RECT 1269.930 376.090 1271.110 377.270 ;
        RECT 1269.930 374.490 1271.110 375.670 ;
        RECT 1269.930 196.090 1271.110 197.270 ;
        RECT 1269.930 194.490 1271.110 195.670 ;
        RECT 1269.930 16.090 1271.110 17.270 ;
        RECT 1269.930 14.490 1271.110 15.670 ;
        RECT 1269.930 -2.910 1271.110 -1.730 ;
        RECT 1269.930 -4.510 1271.110 -3.330 ;
        RECT 1449.930 3523.010 1451.110 3524.190 ;
        RECT 1449.930 3521.410 1451.110 3522.590 ;
        RECT 1449.930 3436.090 1451.110 3437.270 ;
        RECT 1449.930 3434.490 1451.110 3435.670 ;
        RECT 1449.930 3256.090 1451.110 3257.270 ;
        RECT 1449.930 3254.490 1451.110 3255.670 ;
        RECT 1449.930 3076.090 1451.110 3077.270 ;
        RECT 1449.930 3074.490 1451.110 3075.670 ;
        RECT 1449.930 2896.090 1451.110 2897.270 ;
        RECT 1449.930 2894.490 1451.110 2895.670 ;
        RECT 1449.930 2716.090 1451.110 2717.270 ;
        RECT 1449.930 2714.490 1451.110 2715.670 ;
        RECT 1449.930 2536.090 1451.110 2537.270 ;
        RECT 1449.930 2534.490 1451.110 2535.670 ;
        RECT 1449.930 2356.090 1451.110 2357.270 ;
        RECT 1449.930 2354.490 1451.110 2355.670 ;
        RECT 1449.930 2176.090 1451.110 2177.270 ;
        RECT 1449.930 2174.490 1451.110 2175.670 ;
        RECT 1449.930 1996.090 1451.110 1997.270 ;
        RECT 1449.930 1994.490 1451.110 1995.670 ;
        RECT 1449.930 1816.090 1451.110 1817.270 ;
        RECT 1449.930 1814.490 1451.110 1815.670 ;
        RECT 1449.930 1636.090 1451.110 1637.270 ;
        RECT 1449.930 1634.490 1451.110 1635.670 ;
        RECT 1449.930 1456.090 1451.110 1457.270 ;
        RECT 1449.930 1454.490 1451.110 1455.670 ;
        RECT 1449.930 1276.090 1451.110 1277.270 ;
        RECT 1449.930 1274.490 1451.110 1275.670 ;
        RECT 1449.930 1096.090 1451.110 1097.270 ;
        RECT 1449.930 1094.490 1451.110 1095.670 ;
        RECT 1449.930 916.090 1451.110 917.270 ;
        RECT 1449.930 914.490 1451.110 915.670 ;
        RECT 1449.930 736.090 1451.110 737.270 ;
        RECT 1449.930 734.490 1451.110 735.670 ;
        RECT 1449.930 556.090 1451.110 557.270 ;
        RECT 1449.930 554.490 1451.110 555.670 ;
        RECT 1449.930 376.090 1451.110 377.270 ;
        RECT 1449.930 374.490 1451.110 375.670 ;
        RECT 1449.930 196.090 1451.110 197.270 ;
        RECT 1449.930 194.490 1451.110 195.670 ;
        RECT 1449.930 16.090 1451.110 17.270 ;
        RECT 1449.930 14.490 1451.110 15.670 ;
        RECT 1449.930 -2.910 1451.110 -1.730 ;
        RECT 1449.930 -4.510 1451.110 -3.330 ;
        RECT 1629.930 3523.010 1631.110 3524.190 ;
        RECT 1629.930 3521.410 1631.110 3522.590 ;
        RECT 1629.930 3436.090 1631.110 3437.270 ;
        RECT 1629.930 3434.490 1631.110 3435.670 ;
        RECT 1629.930 3256.090 1631.110 3257.270 ;
        RECT 1629.930 3254.490 1631.110 3255.670 ;
        RECT 1629.930 3076.090 1631.110 3077.270 ;
        RECT 1629.930 3074.490 1631.110 3075.670 ;
        RECT 1629.930 2896.090 1631.110 2897.270 ;
        RECT 1629.930 2894.490 1631.110 2895.670 ;
        RECT 1629.930 2716.090 1631.110 2717.270 ;
        RECT 1629.930 2714.490 1631.110 2715.670 ;
        RECT 1629.930 2536.090 1631.110 2537.270 ;
        RECT 1629.930 2534.490 1631.110 2535.670 ;
        RECT 1629.930 2356.090 1631.110 2357.270 ;
        RECT 1629.930 2354.490 1631.110 2355.670 ;
        RECT 1629.930 2176.090 1631.110 2177.270 ;
        RECT 1629.930 2174.490 1631.110 2175.670 ;
        RECT 1629.930 1996.090 1631.110 1997.270 ;
        RECT 1629.930 1994.490 1631.110 1995.670 ;
        RECT 1629.930 1816.090 1631.110 1817.270 ;
        RECT 1629.930 1814.490 1631.110 1815.670 ;
        RECT 1629.930 1636.090 1631.110 1637.270 ;
        RECT 1629.930 1634.490 1631.110 1635.670 ;
        RECT 1629.930 1456.090 1631.110 1457.270 ;
        RECT 1629.930 1454.490 1631.110 1455.670 ;
        RECT 1629.930 1276.090 1631.110 1277.270 ;
        RECT 1629.930 1274.490 1631.110 1275.670 ;
        RECT 1629.930 1096.090 1631.110 1097.270 ;
        RECT 1629.930 1094.490 1631.110 1095.670 ;
        RECT 1629.930 916.090 1631.110 917.270 ;
        RECT 1629.930 914.490 1631.110 915.670 ;
        RECT 1629.930 736.090 1631.110 737.270 ;
        RECT 1629.930 734.490 1631.110 735.670 ;
        RECT 1629.930 556.090 1631.110 557.270 ;
        RECT 1629.930 554.490 1631.110 555.670 ;
        RECT 1629.930 376.090 1631.110 377.270 ;
        RECT 1629.930 374.490 1631.110 375.670 ;
        RECT 1629.930 196.090 1631.110 197.270 ;
        RECT 1629.930 194.490 1631.110 195.670 ;
        RECT 1629.930 16.090 1631.110 17.270 ;
        RECT 1629.930 14.490 1631.110 15.670 ;
        RECT 1629.930 -2.910 1631.110 -1.730 ;
        RECT 1629.930 -4.510 1631.110 -3.330 ;
        RECT 1809.930 3523.010 1811.110 3524.190 ;
        RECT 1809.930 3521.410 1811.110 3522.590 ;
        RECT 1809.930 3436.090 1811.110 3437.270 ;
        RECT 1809.930 3434.490 1811.110 3435.670 ;
        RECT 1809.930 3256.090 1811.110 3257.270 ;
        RECT 1809.930 3254.490 1811.110 3255.670 ;
        RECT 1809.930 3076.090 1811.110 3077.270 ;
        RECT 1809.930 3074.490 1811.110 3075.670 ;
        RECT 1809.930 2896.090 1811.110 2897.270 ;
        RECT 1809.930 2894.490 1811.110 2895.670 ;
        RECT 1809.930 2716.090 1811.110 2717.270 ;
        RECT 1809.930 2714.490 1811.110 2715.670 ;
        RECT 1809.930 2536.090 1811.110 2537.270 ;
        RECT 1809.930 2534.490 1811.110 2535.670 ;
        RECT 1809.930 2356.090 1811.110 2357.270 ;
        RECT 1809.930 2354.490 1811.110 2355.670 ;
        RECT 1809.930 2176.090 1811.110 2177.270 ;
        RECT 1809.930 2174.490 1811.110 2175.670 ;
        RECT 1809.930 1996.090 1811.110 1997.270 ;
        RECT 1809.930 1994.490 1811.110 1995.670 ;
        RECT 1809.930 1816.090 1811.110 1817.270 ;
        RECT 1809.930 1814.490 1811.110 1815.670 ;
        RECT 1809.930 1636.090 1811.110 1637.270 ;
        RECT 1809.930 1634.490 1811.110 1635.670 ;
        RECT 1809.930 1456.090 1811.110 1457.270 ;
        RECT 1809.930 1454.490 1811.110 1455.670 ;
        RECT 1809.930 1276.090 1811.110 1277.270 ;
        RECT 1809.930 1274.490 1811.110 1275.670 ;
        RECT 1809.930 1096.090 1811.110 1097.270 ;
        RECT 1809.930 1094.490 1811.110 1095.670 ;
        RECT 1809.930 916.090 1811.110 917.270 ;
        RECT 1809.930 914.490 1811.110 915.670 ;
        RECT 1809.930 736.090 1811.110 737.270 ;
        RECT 1809.930 734.490 1811.110 735.670 ;
        RECT 1809.930 556.090 1811.110 557.270 ;
        RECT 1809.930 554.490 1811.110 555.670 ;
        RECT 1809.930 376.090 1811.110 377.270 ;
        RECT 1809.930 374.490 1811.110 375.670 ;
        RECT 1809.930 196.090 1811.110 197.270 ;
        RECT 1809.930 194.490 1811.110 195.670 ;
        RECT 1809.930 16.090 1811.110 17.270 ;
        RECT 1809.930 14.490 1811.110 15.670 ;
        RECT 1809.930 -2.910 1811.110 -1.730 ;
        RECT 1809.930 -4.510 1811.110 -3.330 ;
        RECT 1989.930 3523.010 1991.110 3524.190 ;
        RECT 1989.930 3521.410 1991.110 3522.590 ;
        RECT 1989.930 3436.090 1991.110 3437.270 ;
        RECT 1989.930 3434.490 1991.110 3435.670 ;
        RECT 1989.930 3256.090 1991.110 3257.270 ;
        RECT 1989.930 3254.490 1991.110 3255.670 ;
        RECT 1989.930 3076.090 1991.110 3077.270 ;
        RECT 1989.930 3074.490 1991.110 3075.670 ;
        RECT 1989.930 2896.090 1991.110 2897.270 ;
        RECT 1989.930 2894.490 1991.110 2895.670 ;
        RECT 1989.930 2716.090 1991.110 2717.270 ;
        RECT 1989.930 2714.490 1991.110 2715.670 ;
        RECT 1989.930 2536.090 1991.110 2537.270 ;
        RECT 1989.930 2534.490 1991.110 2535.670 ;
        RECT 1989.930 2356.090 1991.110 2357.270 ;
        RECT 1989.930 2354.490 1991.110 2355.670 ;
        RECT 1989.930 2176.090 1991.110 2177.270 ;
        RECT 1989.930 2174.490 1991.110 2175.670 ;
        RECT 1989.930 1996.090 1991.110 1997.270 ;
        RECT 1989.930 1994.490 1991.110 1995.670 ;
        RECT 1989.930 1816.090 1991.110 1817.270 ;
        RECT 1989.930 1814.490 1991.110 1815.670 ;
        RECT 1989.930 1636.090 1991.110 1637.270 ;
        RECT 1989.930 1634.490 1991.110 1635.670 ;
        RECT 1989.930 1456.090 1991.110 1457.270 ;
        RECT 1989.930 1454.490 1991.110 1455.670 ;
        RECT 1989.930 1276.090 1991.110 1277.270 ;
        RECT 1989.930 1274.490 1991.110 1275.670 ;
        RECT 1989.930 1096.090 1991.110 1097.270 ;
        RECT 1989.930 1094.490 1991.110 1095.670 ;
        RECT 1989.930 916.090 1991.110 917.270 ;
        RECT 1989.930 914.490 1991.110 915.670 ;
        RECT 1989.930 736.090 1991.110 737.270 ;
        RECT 1989.930 734.490 1991.110 735.670 ;
        RECT 1989.930 556.090 1991.110 557.270 ;
        RECT 1989.930 554.490 1991.110 555.670 ;
        RECT 1989.930 376.090 1991.110 377.270 ;
        RECT 1989.930 374.490 1991.110 375.670 ;
        RECT 1989.930 196.090 1991.110 197.270 ;
        RECT 1989.930 194.490 1991.110 195.670 ;
        RECT 1989.930 16.090 1991.110 17.270 ;
        RECT 1989.930 14.490 1991.110 15.670 ;
        RECT 1989.930 -2.910 1991.110 -1.730 ;
        RECT 1989.930 -4.510 1991.110 -3.330 ;
        RECT 2169.930 3523.010 2171.110 3524.190 ;
        RECT 2169.930 3521.410 2171.110 3522.590 ;
        RECT 2169.930 3436.090 2171.110 3437.270 ;
        RECT 2169.930 3434.490 2171.110 3435.670 ;
        RECT 2169.930 3256.090 2171.110 3257.270 ;
        RECT 2169.930 3254.490 2171.110 3255.670 ;
        RECT 2169.930 3076.090 2171.110 3077.270 ;
        RECT 2169.930 3074.490 2171.110 3075.670 ;
        RECT 2169.930 2896.090 2171.110 2897.270 ;
        RECT 2169.930 2894.490 2171.110 2895.670 ;
        RECT 2169.930 2716.090 2171.110 2717.270 ;
        RECT 2169.930 2714.490 2171.110 2715.670 ;
        RECT 2169.930 2536.090 2171.110 2537.270 ;
        RECT 2169.930 2534.490 2171.110 2535.670 ;
        RECT 2169.930 2356.090 2171.110 2357.270 ;
        RECT 2169.930 2354.490 2171.110 2355.670 ;
        RECT 2169.930 2176.090 2171.110 2177.270 ;
        RECT 2169.930 2174.490 2171.110 2175.670 ;
        RECT 2169.930 1996.090 2171.110 1997.270 ;
        RECT 2169.930 1994.490 2171.110 1995.670 ;
        RECT 2169.930 1816.090 2171.110 1817.270 ;
        RECT 2169.930 1814.490 2171.110 1815.670 ;
        RECT 2169.930 1636.090 2171.110 1637.270 ;
        RECT 2169.930 1634.490 2171.110 1635.670 ;
        RECT 2169.930 1456.090 2171.110 1457.270 ;
        RECT 2169.930 1454.490 2171.110 1455.670 ;
        RECT 2169.930 1276.090 2171.110 1277.270 ;
        RECT 2169.930 1274.490 2171.110 1275.670 ;
        RECT 2169.930 1096.090 2171.110 1097.270 ;
        RECT 2169.930 1094.490 2171.110 1095.670 ;
        RECT 2169.930 916.090 2171.110 917.270 ;
        RECT 2169.930 914.490 2171.110 915.670 ;
        RECT 2169.930 736.090 2171.110 737.270 ;
        RECT 2169.930 734.490 2171.110 735.670 ;
        RECT 2169.930 556.090 2171.110 557.270 ;
        RECT 2169.930 554.490 2171.110 555.670 ;
        RECT 2169.930 376.090 2171.110 377.270 ;
        RECT 2169.930 374.490 2171.110 375.670 ;
        RECT 2169.930 196.090 2171.110 197.270 ;
        RECT 2169.930 194.490 2171.110 195.670 ;
        RECT 2169.930 16.090 2171.110 17.270 ;
        RECT 2169.930 14.490 2171.110 15.670 ;
        RECT 2169.930 -2.910 2171.110 -1.730 ;
        RECT 2169.930 -4.510 2171.110 -3.330 ;
        RECT 2349.930 3523.010 2351.110 3524.190 ;
        RECT 2349.930 3521.410 2351.110 3522.590 ;
        RECT 2349.930 3436.090 2351.110 3437.270 ;
        RECT 2349.930 3434.490 2351.110 3435.670 ;
        RECT 2349.930 3256.090 2351.110 3257.270 ;
        RECT 2349.930 3254.490 2351.110 3255.670 ;
        RECT 2349.930 3076.090 2351.110 3077.270 ;
        RECT 2349.930 3074.490 2351.110 3075.670 ;
        RECT 2349.930 2896.090 2351.110 2897.270 ;
        RECT 2349.930 2894.490 2351.110 2895.670 ;
        RECT 2349.930 2716.090 2351.110 2717.270 ;
        RECT 2349.930 2714.490 2351.110 2715.670 ;
        RECT 2349.930 2536.090 2351.110 2537.270 ;
        RECT 2349.930 2534.490 2351.110 2535.670 ;
        RECT 2349.930 2356.090 2351.110 2357.270 ;
        RECT 2349.930 2354.490 2351.110 2355.670 ;
        RECT 2349.930 2176.090 2351.110 2177.270 ;
        RECT 2349.930 2174.490 2351.110 2175.670 ;
        RECT 2349.930 1996.090 2351.110 1997.270 ;
        RECT 2349.930 1994.490 2351.110 1995.670 ;
        RECT 2349.930 1816.090 2351.110 1817.270 ;
        RECT 2349.930 1814.490 2351.110 1815.670 ;
        RECT 2349.930 1636.090 2351.110 1637.270 ;
        RECT 2349.930 1634.490 2351.110 1635.670 ;
        RECT 2349.930 1456.090 2351.110 1457.270 ;
        RECT 2349.930 1454.490 2351.110 1455.670 ;
        RECT 2349.930 1276.090 2351.110 1277.270 ;
        RECT 2349.930 1274.490 2351.110 1275.670 ;
        RECT 2349.930 1096.090 2351.110 1097.270 ;
        RECT 2349.930 1094.490 2351.110 1095.670 ;
        RECT 2349.930 916.090 2351.110 917.270 ;
        RECT 2349.930 914.490 2351.110 915.670 ;
        RECT 2349.930 736.090 2351.110 737.270 ;
        RECT 2349.930 734.490 2351.110 735.670 ;
        RECT 2349.930 556.090 2351.110 557.270 ;
        RECT 2349.930 554.490 2351.110 555.670 ;
        RECT 2349.930 376.090 2351.110 377.270 ;
        RECT 2349.930 374.490 2351.110 375.670 ;
        RECT 2349.930 196.090 2351.110 197.270 ;
        RECT 2349.930 194.490 2351.110 195.670 ;
        RECT 2349.930 16.090 2351.110 17.270 ;
        RECT 2349.930 14.490 2351.110 15.670 ;
        RECT 2349.930 -2.910 2351.110 -1.730 ;
        RECT 2349.930 -4.510 2351.110 -3.330 ;
        RECT 2529.930 3523.010 2531.110 3524.190 ;
        RECT 2529.930 3521.410 2531.110 3522.590 ;
        RECT 2529.930 3436.090 2531.110 3437.270 ;
        RECT 2529.930 3434.490 2531.110 3435.670 ;
        RECT 2529.930 3256.090 2531.110 3257.270 ;
        RECT 2529.930 3254.490 2531.110 3255.670 ;
        RECT 2529.930 3076.090 2531.110 3077.270 ;
        RECT 2529.930 3074.490 2531.110 3075.670 ;
        RECT 2529.930 2896.090 2531.110 2897.270 ;
        RECT 2529.930 2894.490 2531.110 2895.670 ;
        RECT 2529.930 2716.090 2531.110 2717.270 ;
        RECT 2529.930 2714.490 2531.110 2715.670 ;
        RECT 2529.930 2536.090 2531.110 2537.270 ;
        RECT 2529.930 2534.490 2531.110 2535.670 ;
        RECT 2529.930 2356.090 2531.110 2357.270 ;
        RECT 2529.930 2354.490 2531.110 2355.670 ;
        RECT 2529.930 2176.090 2531.110 2177.270 ;
        RECT 2529.930 2174.490 2531.110 2175.670 ;
        RECT 2529.930 1996.090 2531.110 1997.270 ;
        RECT 2529.930 1994.490 2531.110 1995.670 ;
        RECT 2529.930 1816.090 2531.110 1817.270 ;
        RECT 2529.930 1814.490 2531.110 1815.670 ;
        RECT 2529.930 1636.090 2531.110 1637.270 ;
        RECT 2529.930 1634.490 2531.110 1635.670 ;
        RECT 2529.930 1456.090 2531.110 1457.270 ;
        RECT 2529.930 1454.490 2531.110 1455.670 ;
        RECT 2529.930 1276.090 2531.110 1277.270 ;
        RECT 2529.930 1274.490 2531.110 1275.670 ;
        RECT 2529.930 1096.090 2531.110 1097.270 ;
        RECT 2529.930 1094.490 2531.110 1095.670 ;
        RECT 2529.930 916.090 2531.110 917.270 ;
        RECT 2529.930 914.490 2531.110 915.670 ;
        RECT 2529.930 736.090 2531.110 737.270 ;
        RECT 2529.930 734.490 2531.110 735.670 ;
        RECT 2529.930 556.090 2531.110 557.270 ;
        RECT 2529.930 554.490 2531.110 555.670 ;
        RECT 2529.930 376.090 2531.110 377.270 ;
        RECT 2529.930 374.490 2531.110 375.670 ;
        RECT 2529.930 196.090 2531.110 197.270 ;
        RECT 2529.930 194.490 2531.110 195.670 ;
        RECT 2529.930 16.090 2531.110 17.270 ;
        RECT 2529.930 14.490 2531.110 15.670 ;
        RECT 2529.930 -2.910 2531.110 -1.730 ;
        RECT 2529.930 -4.510 2531.110 -3.330 ;
        RECT 2709.930 3523.010 2711.110 3524.190 ;
        RECT 2709.930 3521.410 2711.110 3522.590 ;
        RECT 2709.930 3436.090 2711.110 3437.270 ;
        RECT 2709.930 3434.490 2711.110 3435.670 ;
        RECT 2709.930 3256.090 2711.110 3257.270 ;
        RECT 2709.930 3254.490 2711.110 3255.670 ;
        RECT 2709.930 3076.090 2711.110 3077.270 ;
        RECT 2709.930 3074.490 2711.110 3075.670 ;
        RECT 2709.930 2896.090 2711.110 2897.270 ;
        RECT 2709.930 2894.490 2711.110 2895.670 ;
        RECT 2709.930 2716.090 2711.110 2717.270 ;
        RECT 2709.930 2714.490 2711.110 2715.670 ;
        RECT 2709.930 2536.090 2711.110 2537.270 ;
        RECT 2709.930 2534.490 2711.110 2535.670 ;
        RECT 2709.930 2356.090 2711.110 2357.270 ;
        RECT 2709.930 2354.490 2711.110 2355.670 ;
        RECT 2709.930 2176.090 2711.110 2177.270 ;
        RECT 2709.930 2174.490 2711.110 2175.670 ;
        RECT 2709.930 1996.090 2711.110 1997.270 ;
        RECT 2709.930 1994.490 2711.110 1995.670 ;
        RECT 2709.930 1816.090 2711.110 1817.270 ;
        RECT 2709.930 1814.490 2711.110 1815.670 ;
        RECT 2709.930 1636.090 2711.110 1637.270 ;
        RECT 2709.930 1634.490 2711.110 1635.670 ;
        RECT 2709.930 1456.090 2711.110 1457.270 ;
        RECT 2709.930 1454.490 2711.110 1455.670 ;
        RECT 2709.930 1276.090 2711.110 1277.270 ;
        RECT 2709.930 1274.490 2711.110 1275.670 ;
        RECT 2709.930 1096.090 2711.110 1097.270 ;
        RECT 2709.930 1094.490 2711.110 1095.670 ;
        RECT 2709.930 916.090 2711.110 917.270 ;
        RECT 2709.930 914.490 2711.110 915.670 ;
        RECT 2709.930 736.090 2711.110 737.270 ;
        RECT 2709.930 734.490 2711.110 735.670 ;
        RECT 2709.930 556.090 2711.110 557.270 ;
        RECT 2709.930 554.490 2711.110 555.670 ;
        RECT 2709.930 376.090 2711.110 377.270 ;
        RECT 2709.930 374.490 2711.110 375.670 ;
        RECT 2709.930 196.090 2711.110 197.270 ;
        RECT 2709.930 194.490 2711.110 195.670 ;
        RECT 2709.930 16.090 2711.110 17.270 ;
        RECT 2709.930 14.490 2711.110 15.670 ;
        RECT 2709.930 -2.910 2711.110 -1.730 ;
        RECT 2709.930 -4.510 2711.110 -3.330 ;
        RECT 2889.930 3523.010 2891.110 3524.190 ;
        RECT 2889.930 3521.410 2891.110 3522.590 ;
        RECT 2889.930 3436.090 2891.110 3437.270 ;
        RECT 2889.930 3434.490 2891.110 3435.670 ;
        RECT 2889.930 3256.090 2891.110 3257.270 ;
        RECT 2889.930 3254.490 2891.110 3255.670 ;
        RECT 2889.930 3076.090 2891.110 3077.270 ;
        RECT 2889.930 3074.490 2891.110 3075.670 ;
        RECT 2889.930 2896.090 2891.110 2897.270 ;
        RECT 2889.930 2894.490 2891.110 2895.670 ;
        RECT 2889.930 2716.090 2891.110 2717.270 ;
        RECT 2889.930 2714.490 2891.110 2715.670 ;
        RECT 2889.930 2536.090 2891.110 2537.270 ;
        RECT 2889.930 2534.490 2891.110 2535.670 ;
        RECT 2889.930 2356.090 2891.110 2357.270 ;
        RECT 2889.930 2354.490 2891.110 2355.670 ;
        RECT 2889.930 2176.090 2891.110 2177.270 ;
        RECT 2889.930 2174.490 2891.110 2175.670 ;
        RECT 2889.930 1996.090 2891.110 1997.270 ;
        RECT 2889.930 1994.490 2891.110 1995.670 ;
        RECT 2889.930 1816.090 2891.110 1817.270 ;
        RECT 2889.930 1814.490 2891.110 1815.670 ;
        RECT 2889.930 1636.090 2891.110 1637.270 ;
        RECT 2889.930 1634.490 2891.110 1635.670 ;
        RECT 2889.930 1456.090 2891.110 1457.270 ;
        RECT 2889.930 1454.490 2891.110 1455.670 ;
        RECT 2889.930 1276.090 2891.110 1277.270 ;
        RECT 2889.930 1274.490 2891.110 1275.670 ;
        RECT 2889.930 1096.090 2891.110 1097.270 ;
        RECT 2889.930 1094.490 2891.110 1095.670 ;
        RECT 2889.930 916.090 2891.110 917.270 ;
        RECT 2889.930 914.490 2891.110 915.670 ;
        RECT 2889.930 736.090 2891.110 737.270 ;
        RECT 2889.930 734.490 2891.110 735.670 ;
        RECT 2889.930 556.090 2891.110 557.270 ;
        RECT 2889.930 554.490 2891.110 555.670 ;
        RECT 2889.930 376.090 2891.110 377.270 ;
        RECT 2889.930 374.490 2891.110 375.670 ;
        RECT 2889.930 196.090 2891.110 197.270 ;
        RECT 2889.930 194.490 2891.110 195.670 ;
        RECT 2889.930 16.090 2891.110 17.270 ;
        RECT 2889.930 14.490 2891.110 15.670 ;
        RECT 2889.930 -2.910 2891.110 -1.730 ;
        RECT 2889.930 -4.510 2891.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3436.090 2928.690 3437.270 ;
        RECT 2927.510 3434.490 2928.690 3435.670 ;
        RECT 2927.510 3256.090 2928.690 3257.270 ;
        RECT 2927.510 3254.490 2928.690 3255.670 ;
        RECT 2927.510 3076.090 2928.690 3077.270 ;
        RECT 2927.510 3074.490 2928.690 3075.670 ;
        RECT 2927.510 2896.090 2928.690 2897.270 ;
        RECT 2927.510 2894.490 2928.690 2895.670 ;
        RECT 2927.510 2716.090 2928.690 2717.270 ;
        RECT 2927.510 2714.490 2928.690 2715.670 ;
        RECT 2927.510 2536.090 2928.690 2537.270 ;
        RECT 2927.510 2534.490 2928.690 2535.670 ;
        RECT 2927.510 2356.090 2928.690 2357.270 ;
        RECT 2927.510 2354.490 2928.690 2355.670 ;
        RECT 2927.510 2176.090 2928.690 2177.270 ;
        RECT 2927.510 2174.490 2928.690 2175.670 ;
        RECT 2927.510 1996.090 2928.690 1997.270 ;
        RECT 2927.510 1994.490 2928.690 1995.670 ;
        RECT 2927.510 1816.090 2928.690 1817.270 ;
        RECT 2927.510 1814.490 2928.690 1815.670 ;
        RECT 2927.510 1636.090 2928.690 1637.270 ;
        RECT 2927.510 1634.490 2928.690 1635.670 ;
        RECT 2927.510 1456.090 2928.690 1457.270 ;
        RECT 2927.510 1454.490 2928.690 1455.670 ;
        RECT 2927.510 1276.090 2928.690 1277.270 ;
        RECT 2927.510 1274.490 2928.690 1275.670 ;
        RECT 2927.510 1096.090 2928.690 1097.270 ;
        RECT 2927.510 1094.490 2928.690 1095.670 ;
        RECT 2927.510 916.090 2928.690 917.270 ;
        RECT 2927.510 914.490 2928.690 915.670 ;
        RECT 2927.510 736.090 2928.690 737.270 ;
        RECT 2927.510 734.490 2928.690 735.670 ;
        RECT 2927.510 556.090 2928.690 557.270 ;
        RECT 2927.510 554.490 2928.690 555.670 ;
        RECT 2927.510 376.090 2928.690 377.270 ;
        RECT 2927.510 374.490 2928.690 375.670 ;
        RECT 2927.510 196.090 2928.690 197.270 ;
        RECT 2927.510 194.490 2928.690 195.670 ;
        RECT 2927.510 16.090 2928.690 17.270 ;
        RECT 2927.510 14.490 2928.690 15.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 9.020 3524.300 12.020 3524.310 ;
        RECT 189.020 3524.300 192.020 3524.310 ;
        RECT 369.020 3524.300 372.020 3524.310 ;
        RECT 549.020 3524.300 552.020 3524.310 ;
        RECT 729.020 3524.300 732.020 3524.310 ;
        RECT 909.020 3524.300 912.020 3524.310 ;
        RECT 1089.020 3524.300 1092.020 3524.310 ;
        RECT 1269.020 3524.300 1272.020 3524.310 ;
        RECT 1449.020 3524.300 1452.020 3524.310 ;
        RECT 1629.020 3524.300 1632.020 3524.310 ;
        RECT 1809.020 3524.300 1812.020 3524.310 ;
        RECT 1989.020 3524.300 1992.020 3524.310 ;
        RECT 2169.020 3524.300 2172.020 3524.310 ;
        RECT 2349.020 3524.300 2352.020 3524.310 ;
        RECT 2529.020 3524.300 2532.020 3524.310 ;
        RECT 2709.020 3524.300 2712.020 3524.310 ;
        RECT 2889.020 3524.300 2892.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 9.020 3521.290 12.020 3521.300 ;
        RECT 189.020 3521.290 192.020 3521.300 ;
        RECT 369.020 3521.290 372.020 3521.300 ;
        RECT 549.020 3521.290 552.020 3521.300 ;
        RECT 729.020 3521.290 732.020 3521.300 ;
        RECT 909.020 3521.290 912.020 3521.300 ;
        RECT 1089.020 3521.290 1092.020 3521.300 ;
        RECT 1269.020 3521.290 1272.020 3521.300 ;
        RECT 1449.020 3521.290 1452.020 3521.300 ;
        RECT 1629.020 3521.290 1632.020 3521.300 ;
        RECT 1809.020 3521.290 1812.020 3521.300 ;
        RECT 1989.020 3521.290 1992.020 3521.300 ;
        RECT 2169.020 3521.290 2172.020 3521.300 ;
        RECT 2349.020 3521.290 2352.020 3521.300 ;
        RECT 2529.020 3521.290 2532.020 3521.300 ;
        RECT 2709.020 3521.290 2712.020 3521.300 ;
        RECT 2889.020 3521.290 2892.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3437.380 -6.980 3437.390 ;
        RECT 9.020 3437.380 12.020 3437.390 ;
        RECT 189.020 3437.380 192.020 3437.390 ;
        RECT 369.020 3437.380 372.020 3437.390 ;
        RECT 549.020 3437.380 552.020 3437.390 ;
        RECT 729.020 3437.380 732.020 3437.390 ;
        RECT 909.020 3437.380 912.020 3437.390 ;
        RECT 1089.020 3437.380 1092.020 3437.390 ;
        RECT 1269.020 3437.380 1272.020 3437.390 ;
        RECT 1449.020 3437.380 1452.020 3437.390 ;
        RECT 1629.020 3437.380 1632.020 3437.390 ;
        RECT 1809.020 3437.380 1812.020 3437.390 ;
        RECT 1989.020 3437.380 1992.020 3437.390 ;
        RECT 2169.020 3437.380 2172.020 3437.390 ;
        RECT 2349.020 3437.380 2352.020 3437.390 ;
        RECT 2529.020 3437.380 2532.020 3437.390 ;
        RECT 2709.020 3437.380 2712.020 3437.390 ;
        RECT 2889.020 3437.380 2892.020 3437.390 ;
        RECT 2926.600 3437.380 2929.600 3437.390 ;
        RECT -14.680 3434.380 2934.300 3437.380 ;
        RECT -9.980 3434.370 -6.980 3434.380 ;
        RECT 9.020 3434.370 12.020 3434.380 ;
        RECT 189.020 3434.370 192.020 3434.380 ;
        RECT 369.020 3434.370 372.020 3434.380 ;
        RECT 549.020 3434.370 552.020 3434.380 ;
        RECT 729.020 3434.370 732.020 3434.380 ;
        RECT 909.020 3434.370 912.020 3434.380 ;
        RECT 1089.020 3434.370 1092.020 3434.380 ;
        RECT 1269.020 3434.370 1272.020 3434.380 ;
        RECT 1449.020 3434.370 1452.020 3434.380 ;
        RECT 1629.020 3434.370 1632.020 3434.380 ;
        RECT 1809.020 3434.370 1812.020 3434.380 ;
        RECT 1989.020 3434.370 1992.020 3434.380 ;
        RECT 2169.020 3434.370 2172.020 3434.380 ;
        RECT 2349.020 3434.370 2352.020 3434.380 ;
        RECT 2529.020 3434.370 2532.020 3434.380 ;
        RECT 2709.020 3434.370 2712.020 3434.380 ;
        RECT 2889.020 3434.370 2892.020 3434.380 ;
        RECT 2926.600 3434.370 2929.600 3434.380 ;
        RECT -9.980 3257.380 -6.980 3257.390 ;
        RECT 9.020 3257.380 12.020 3257.390 ;
        RECT 189.020 3257.380 192.020 3257.390 ;
        RECT 369.020 3257.380 372.020 3257.390 ;
        RECT 549.020 3257.380 552.020 3257.390 ;
        RECT 729.020 3257.380 732.020 3257.390 ;
        RECT 909.020 3257.380 912.020 3257.390 ;
        RECT 1089.020 3257.380 1092.020 3257.390 ;
        RECT 1269.020 3257.380 1272.020 3257.390 ;
        RECT 1449.020 3257.380 1452.020 3257.390 ;
        RECT 1629.020 3257.380 1632.020 3257.390 ;
        RECT 1809.020 3257.380 1812.020 3257.390 ;
        RECT 1989.020 3257.380 1992.020 3257.390 ;
        RECT 2169.020 3257.380 2172.020 3257.390 ;
        RECT 2349.020 3257.380 2352.020 3257.390 ;
        RECT 2529.020 3257.380 2532.020 3257.390 ;
        RECT 2709.020 3257.380 2712.020 3257.390 ;
        RECT 2889.020 3257.380 2892.020 3257.390 ;
        RECT 2926.600 3257.380 2929.600 3257.390 ;
        RECT -14.680 3254.380 2934.300 3257.380 ;
        RECT -9.980 3254.370 -6.980 3254.380 ;
        RECT 9.020 3254.370 12.020 3254.380 ;
        RECT 189.020 3254.370 192.020 3254.380 ;
        RECT 369.020 3254.370 372.020 3254.380 ;
        RECT 549.020 3254.370 552.020 3254.380 ;
        RECT 729.020 3254.370 732.020 3254.380 ;
        RECT 909.020 3254.370 912.020 3254.380 ;
        RECT 1089.020 3254.370 1092.020 3254.380 ;
        RECT 1269.020 3254.370 1272.020 3254.380 ;
        RECT 1449.020 3254.370 1452.020 3254.380 ;
        RECT 1629.020 3254.370 1632.020 3254.380 ;
        RECT 1809.020 3254.370 1812.020 3254.380 ;
        RECT 1989.020 3254.370 1992.020 3254.380 ;
        RECT 2169.020 3254.370 2172.020 3254.380 ;
        RECT 2349.020 3254.370 2352.020 3254.380 ;
        RECT 2529.020 3254.370 2532.020 3254.380 ;
        RECT 2709.020 3254.370 2712.020 3254.380 ;
        RECT 2889.020 3254.370 2892.020 3254.380 ;
        RECT 2926.600 3254.370 2929.600 3254.380 ;
        RECT -9.980 3077.380 -6.980 3077.390 ;
        RECT 9.020 3077.380 12.020 3077.390 ;
        RECT 189.020 3077.380 192.020 3077.390 ;
        RECT 369.020 3077.380 372.020 3077.390 ;
        RECT 549.020 3077.380 552.020 3077.390 ;
        RECT 729.020 3077.380 732.020 3077.390 ;
        RECT 909.020 3077.380 912.020 3077.390 ;
        RECT 1089.020 3077.380 1092.020 3077.390 ;
        RECT 1269.020 3077.380 1272.020 3077.390 ;
        RECT 1449.020 3077.380 1452.020 3077.390 ;
        RECT 1629.020 3077.380 1632.020 3077.390 ;
        RECT 1809.020 3077.380 1812.020 3077.390 ;
        RECT 1989.020 3077.380 1992.020 3077.390 ;
        RECT 2169.020 3077.380 2172.020 3077.390 ;
        RECT 2349.020 3077.380 2352.020 3077.390 ;
        RECT 2529.020 3077.380 2532.020 3077.390 ;
        RECT 2709.020 3077.380 2712.020 3077.390 ;
        RECT 2889.020 3077.380 2892.020 3077.390 ;
        RECT 2926.600 3077.380 2929.600 3077.390 ;
        RECT -14.680 3074.380 2934.300 3077.380 ;
        RECT -9.980 3074.370 -6.980 3074.380 ;
        RECT 9.020 3074.370 12.020 3074.380 ;
        RECT 189.020 3074.370 192.020 3074.380 ;
        RECT 369.020 3074.370 372.020 3074.380 ;
        RECT 549.020 3074.370 552.020 3074.380 ;
        RECT 729.020 3074.370 732.020 3074.380 ;
        RECT 909.020 3074.370 912.020 3074.380 ;
        RECT 1089.020 3074.370 1092.020 3074.380 ;
        RECT 1269.020 3074.370 1272.020 3074.380 ;
        RECT 1449.020 3074.370 1452.020 3074.380 ;
        RECT 1629.020 3074.370 1632.020 3074.380 ;
        RECT 1809.020 3074.370 1812.020 3074.380 ;
        RECT 1989.020 3074.370 1992.020 3074.380 ;
        RECT 2169.020 3074.370 2172.020 3074.380 ;
        RECT 2349.020 3074.370 2352.020 3074.380 ;
        RECT 2529.020 3074.370 2532.020 3074.380 ;
        RECT 2709.020 3074.370 2712.020 3074.380 ;
        RECT 2889.020 3074.370 2892.020 3074.380 ;
        RECT 2926.600 3074.370 2929.600 3074.380 ;
        RECT -9.980 2897.380 -6.980 2897.390 ;
        RECT 9.020 2897.380 12.020 2897.390 ;
        RECT 189.020 2897.380 192.020 2897.390 ;
        RECT 369.020 2897.380 372.020 2897.390 ;
        RECT 549.020 2897.380 552.020 2897.390 ;
        RECT 729.020 2897.380 732.020 2897.390 ;
        RECT 909.020 2897.380 912.020 2897.390 ;
        RECT 1089.020 2897.380 1092.020 2897.390 ;
        RECT 1269.020 2897.380 1272.020 2897.390 ;
        RECT 1449.020 2897.380 1452.020 2897.390 ;
        RECT 1629.020 2897.380 1632.020 2897.390 ;
        RECT 1809.020 2897.380 1812.020 2897.390 ;
        RECT 1989.020 2897.380 1992.020 2897.390 ;
        RECT 2169.020 2897.380 2172.020 2897.390 ;
        RECT 2349.020 2897.380 2352.020 2897.390 ;
        RECT 2529.020 2897.380 2532.020 2897.390 ;
        RECT 2709.020 2897.380 2712.020 2897.390 ;
        RECT 2889.020 2897.380 2892.020 2897.390 ;
        RECT 2926.600 2897.380 2929.600 2897.390 ;
        RECT -14.680 2894.380 2934.300 2897.380 ;
        RECT -9.980 2894.370 -6.980 2894.380 ;
        RECT 9.020 2894.370 12.020 2894.380 ;
        RECT 189.020 2894.370 192.020 2894.380 ;
        RECT 369.020 2894.370 372.020 2894.380 ;
        RECT 549.020 2894.370 552.020 2894.380 ;
        RECT 729.020 2894.370 732.020 2894.380 ;
        RECT 909.020 2894.370 912.020 2894.380 ;
        RECT 1089.020 2894.370 1092.020 2894.380 ;
        RECT 1269.020 2894.370 1272.020 2894.380 ;
        RECT 1449.020 2894.370 1452.020 2894.380 ;
        RECT 1629.020 2894.370 1632.020 2894.380 ;
        RECT 1809.020 2894.370 1812.020 2894.380 ;
        RECT 1989.020 2894.370 1992.020 2894.380 ;
        RECT 2169.020 2894.370 2172.020 2894.380 ;
        RECT 2349.020 2894.370 2352.020 2894.380 ;
        RECT 2529.020 2894.370 2532.020 2894.380 ;
        RECT 2709.020 2894.370 2712.020 2894.380 ;
        RECT 2889.020 2894.370 2892.020 2894.380 ;
        RECT 2926.600 2894.370 2929.600 2894.380 ;
        RECT -9.980 2717.380 -6.980 2717.390 ;
        RECT 9.020 2717.380 12.020 2717.390 ;
        RECT 189.020 2717.380 192.020 2717.390 ;
        RECT 369.020 2717.380 372.020 2717.390 ;
        RECT 549.020 2717.380 552.020 2717.390 ;
        RECT 729.020 2717.380 732.020 2717.390 ;
        RECT 909.020 2717.380 912.020 2717.390 ;
        RECT 1089.020 2717.380 1092.020 2717.390 ;
        RECT 1269.020 2717.380 1272.020 2717.390 ;
        RECT 1449.020 2717.380 1452.020 2717.390 ;
        RECT 1629.020 2717.380 1632.020 2717.390 ;
        RECT 1809.020 2717.380 1812.020 2717.390 ;
        RECT 1989.020 2717.380 1992.020 2717.390 ;
        RECT 2169.020 2717.380 2172.020 2717.390 ;
        RECT 2349.020 2717.380 2352.020 2717.390 ;
        RECT 2529.020 2717.380 2532.020 2717.390 ;
        RECT 2709.020 2717.380 2712.020 2717.390 ;
        RECT 2889.020 2717.380 2892.020 2717.390 ;
        RECT 2926.600 2717.380 2929.600 2717.390 ;
        RECT -14.680 2714.380 2934.300 2717.380 ;
        RECT -9.980 2714.370 -6.980 2714.380 ;
        RECT 9.020 2714.370 12.020 2714.380 ;
        RECT 189.020 2714.370 192.020 2714.380 ;
        RECT 369.020 2714.370 372.020 2714.380 ;
        RECT 549.020 2714.370 552.020 2714.380 ;
        RECT 729.020 2714.370 732.020 2714.380 ;
        RECT 909.020 2714.370 912.020 2714.380 ;
        RECT 1089.020 2714.370 1092.020 2714.380 ;
        RECT 1269.020 2714.370 1272.020 2714.380 ;
        RECT 1449.020 2714.370 1452.020 2714.380 ;
        RECT 1629.020 2714.370 1632.020 2714.380 ;
        RECT 1809.020 2714.370 1812.020 2714.380 ;
        RECT 1989.020 2714.370 1992.020 2714.380 ;
        RECT 2169.020 2714.370 2172.020 2714.380 ;
        RECT 2349.020 2714.370 2352.020 2714.380 ;
        RECT 2529.020 2714.370 2532.020 2714.380 ;
        RECT 2709.020 2714.370 2712.020 2714.380 ;
        RECT 2889.020 2714.370 2892.020 2714.380 ;
        RECT 2926.600 2714.370 2929.600 2714.380 ;
        RECT -9.980 2537.380 -6.980 2537.390 ;
        RECT 9.020 2537.380 12.020 2537.390 ;
        RECT 189.020 2537.380 192.020 2537.390 ;
        RECT 369.020 2537.380 372.020 2537.390 ;
        RECT 549.020 2537.380 552.020 2537.390 ;
        RECT 729.020 2537.380 732.020 2537.390 ;
        RECT 909.020 2537.380 912.020 2537.390 ;
        RECT 1089.020 2537.380 1092.020 2537.390 ;
        RECT 1269.020 2537.380 1272.020 2537.390 ;
        RECT 1449.020 2537.380 1452.020 2537.390 ;
        RECT 1629.020 2537.380 1632.020 2537.390 ;
        RECT 1809.020 2537.380 1812.020 2537.390 ;
        RECT 1989.020 2537.380 1992.020 2537.390 ;
        RECT 2169.020 2537.380 2172.020 2537.390 ;
        RECT 2349.020 2537.380 2352.020 2537.390 ;
        RECT 2529.020 2537.380 2532.020 2537.390 ;
        RECT 2709.020 2537.380 2712.020 2537.390 ;
        RECT 2889.020 2537.380 2892.020 2537.390 ;
        RECT 2926.600 2537.380 2929.600 2537.390 ;
        RECT -14.680 2534.380 2934.300 2537.380 ;
        RECT -9.980 2534.370 -6.980 2534.380 ;
        RECT 9.020 2534.370 12.020 2534.380 ;
        RECT 189.020 2534.370 192.020 2534.380 ;
        RECT 369.020 2534.370 372.020 2534.380 ;
        RECT 549.020 2534.370 552.020 2534.380 ;
        RECT 729.020 2534.370 732.020 2534.380 ;
        RECT 909.020 2534.370 912.020 2534.380 ;
        RECT 1089.020 2534.370 1092.020 2534.380 ;
        RECT 1269.020 2534.370 1272.020 2534.380 ;
        RECT 1449.020 2534.370 1452.020 2534.380 ;
        RECT 1629.020 2534.370 1632.020 2534.380 ;
        RECT 1809.020 2534.370 1812.020 2534.380 ;
        RECT 1989.020 2534.370 1992.020 2534.380 ;
        RECT 2169.020 2534.370 2172.020 2534.380 ;
        RECT 2349.020 2534.370 2352.020 2534.380 ;
        RECT 2529.020 2534.370 2532.020 2534.380 ;
        RECT 2709.020 2534.370 2712.020 2534.380 ;
        RECT 2889.020 2534.370 2892.020 2534.380 ;
        RECT 2926.600 2534.370 2929.600 2534.380 ;
        RECT -9.980 2357.380 -6.980 2357.390 ;
        RECT 9.020 2357.380 12.020 2357.390 ;
        RECT 189.020 2357.380 192.020 2357.390 ;
        RECT 369.020 2357.380 372.020 2357.390 ;
        RECT 549.020 2357.380 552.020 2357.390 ;
        RECT 729.020 2357.380 732.020 2357.390 ;
        RECT 909.020 2357.380 912.020 2357.390 ;
        RECT 1089.020 2357.380 1092.020 2357.390 ;
        RECT 1269.020 2357.380 1272.020 2357.390 ;
        RECT 1449.020 2357.380 1452.020 2357.390 ;
        RECT 1629.020 2357.380 1632.020 2357.390 ;
        RECT 1809.020 2357.380 1812.020 2357.390 ;
        RECT 1989.020 2357.380 1992.020 2357.390 ;
        RECT 2169.020 2357.380 2172.020 2357.390 ;
        RECT 2349.020 2357.380 2352.020 2357.390 ;
        RECT 2529.020 2357.380 2532.020 2357.390 ;
        RECT 2709.020 2357.380 2712.020 2357.390 ;
        RECT 2889.020 2357.380 2892.020 2357.390 ;
        RECT 2926.600 2357.380 2929.600 2357.390 ;
        RECT -14.680 2354.380 2934.300 2357.380 ;
        RECT -9.980 2354.370 -6.980 2354.380 ;
        RECT 9.020 2354.370 12.020 2354.380 ;
        RECT 189.020 2354.370 192.020 2354.380 ;
        RECT 369.020 2354.370 372.020 2354.380 ;
        RECT 549.020 2354.370 552.020 2354.380 ;
        RECT 729.020 2354.370 732.020 2354.380 ;
        RECT 909.020 2354.370 912.020 2354.380 ;
        RECT 1089.020 2354.370 1092.020 2354.380 ;
        RECT 1269.020 2354.370 1272.020 2354.380 ;
        RECT 1449.020 2354.370 1452.020 2354.380 ;
        RECT 1629.020 2354.370 1632.020 2354.380 ;
        RECT 1809.020 2354.370 1812.020 2354.380 ;
        RECT 1989.020 2354.370 1992.020 2354.380 ;
        RECT 2169.020 2354.370 2172.020 2354.380 ;
        RECT 2349.020 2354.370 2352.020 2354.380 ;
        RECT 2529.020 2354.370 2532.020 2354.380 ;
        RECT 2709.020 2354.370 2712.020 2354.380 ;
        RECT 2889.020 2354.370 2892.020 2354.380 ;
        RECT 2926.600 2354.370 2929.600 2354.380 ;
        RECT -9.980 2177.380 -6.980 2177.390 ;
        RECT 9.020 2177.380 12.020 2177.390 ;
        RECT 189.020 2177.380 192.020 2177.390 ;
        RECT 369.020 2177.380 372.020 2177.390 ;
        RECT 549.020 2177.380 552.020 2177.390 ;
        RECT 729.020 2177.380 732.020 2177.390 ;
        RECT 909.020 2177.380 912.020 2177.390 ;
        RECT 1089.020 2177.380 1092.020 2177.390 ;
        RECT 1269.020 2177.380 1272.020 2177.390 ;
        RECT 1449.020 2177.380 1452.020 2177.390 ;
        RECT 1629.020 2177.380 1632.020 2177.390 ;
        RECT 1809.020 2177.380 1812.020 2177.390 ;
        RECT 1989.020 2177.380 1992.020 2177.390 ;
        RECT 2169.020 2177.380 2172.020 2177.390 ;
        RECT 2349.020 2177.380 2352.020 2177.390 ;
        RECT 2529.020 2177.380 2532.020 2177.390 ;
        RECT 2709.020 2177.380 2712.020 2177.390 ;
        RECT 2889.020 2177.380 2892.020 2177.390 ;
        RECT 2926.600 2177.380 2929.600 2177.390 ;
        RECT -14.680 2174.380 2934.300 2177.380 ;
        RECT -9.980 2174.370 -6.980 2174.380 ;
        RECT 9.020 2174.370 12.020 2174.380 ;
        RECT 189.020 2174.370 192.020 2174.380 ;
        RECT 369.020 2174.370 372.020 2174.380 ;
        RECT 549.020 2174.370 552.020 2174.380 ;
        RECT 729.020 2174.370 732.020 2174.380 ;
        RECT 909.020 2174.370 912.020 2174.380 ;
        RECT 1089.020 2174.370 1092.020 2174.380 ;
        RECT 1269.020 2174.370 1272.020 2174.380 ;
        RECT 1449.020 2174.370 1452.020 2174.380 ;
        RECT 1629.020 2174.370 1632.020 2174.380 ;
        RECT 1809.020 2174.370 1812.020 2174.380 ;
        RECT 1989.020 2174.370 1992.020 2174.380 ;
        RECT 2169.020 2174.370 2172.020 2174.380 ;
        RECT 2349.020 2174.370 2352.020 2174.380 ;
        RECT 2529.020 2174.370 2532.020 2174.380 ;
        RECT 2709.020 2174.370 2712.020 2174.380 ;
        RECT 2889.020 2174.370 2892.020 2174.380 ;
        RECT 2926.600 2174.370 2929.600 2174.380 ;
        RECT -9.980 1997.380 -6.980 1997.390 ;
        RECT 9.020 1997.380 12.020 1997.390 ;
        RECT 189.020 1997.380 192.020 1997.390 ;
        RECT 369.020 1997.380 372.020 1997.390 ;
        RECT 549.020 1997.380 552.020 1997.390 ;
        RECT 729.020 1997.380 732.020 1997.390 ;
        RECT 909.020 1997.380 912.020 1997.390 ;
        RECT 1089.020 1997.380 1092.020 1997.390 ;
        RECT 1269.020 1997.380 1272.020 1997.390 ;
        RECT 1449.020 1997.380 1452.020 1997.390 ;
        RECT 1629.020 1997.380 1632.020 1997.390 ;
        RECT 1809.020 1997.380 1812.020 1997.390 ;
        RECT 1989.020 1997.380 1992.020 1997.390 ;
        RECT 2169.020 1997.380 2172.020 1997.390 ;
        RECT 2349.020 1997.380 2352.020 1997.390 ;
        RECT 2529.020 1997.380 2532.020 1997.390 ;
        RECT 2709.020 1997.380 2712.020 1997.390 ;
        RECT 2889.020 1997.380 2892.020 1997.390 ;
        RECT 2926.600 1997.380 2929.600 1997.390 ;
        RECT -14.680 1994.380 2934.300 1997.380 ;
        RECT -9.980 1994.370 -6.980 1994.380 ;
        RECT 9.020 1994.370 12.020 1994.380 ;
        RECT 189.020 1994.370 192.020 1994.380 ;
        RECT 369.020 1994.370 372.020 1994.380 ;
        RECT 549.020 1994.370 552.020 1994.380 ;
        RECT 729.020 1994.370 732.020 1994.380 ;
        RECT 909.020 1994.370 912.020 1994.380 ;
        RECT 1089.020 1994.370 1092.020 1994.380 ;
        RECT 1269.020 1994.370 1272.020 1994.380 ;
        RECT 1449.020 1994.370 1452.020 1994.380 ;
        RECT 1629.020 1994.370 1632.020 1994.380 ;
        RECT 1809.020 1994.370 1812.020 1994.380 ;
        RECT 1989.020 1994.370 1992.020 1994.380 ;
        RECT 2169.020 1994.370 2172.020 1994.380 ;
        RECT 2349.020 1994.370 2352.020 1994.380 ;
        RECT 2529.020 1994.370 2532.020 1994.380 ;
        RECT 2709.020 1994.370 2712.020 1994.380 ;
        RECT 2889.020 1994.370 2892.020 1994.380 ;
        RECT 2926.600 1994.370 2929.600 1994.380 ;
        RECT -9.980 1817.380 -6.980 1817.390 ;
        RECT 9.020 1817.380 12.020 1817.390 ;
        RECT 189.020 1817.380 192.020 1817.390 ;
        RECT 369.020 1817.380 372.020 1817.390 ;
        RECT 549.020 1817.380 552.020 1817.390 ;
        RECT 729.020 1817.380 732.020 1817.390 ;
        RECT 909.020 1817.380 912.020 1817.390 ;
        RECT 1089.020 1817.380 1092.020 1817.390 ;
        RECT 1269.020 1817.380 1272.020 1817.390 ;
        RECT 1449.020 1817.380 1452.020 1817.390 ;
        RECT 1629.020 1817.380 1632.020 1817.390 ;
        RECT 1809.020 1817.380 1812.020 1817.390 ;
        RECT 1989.020 1817.380 1992.020 1817.390 ;
        RECT 2169.020 1817.380 2172.020 1817.390 ;
        RECT 2349.020 1817.380 2352.020 1817.390 ;
        RECT 2529.020 1817.380 2532.020 1817.390 ;
        RECT 2709.020 1817.380 2712.020 1817.390 ;
        RECT 2889.020 1817.380 2892.020 1817.390 ;
        RECT 2926.600 1817.380 2929.600 1817.390 ;
        RECT -14.680 1814.380 2934.300 1817.380 ;
        RECT -9.980 1814.370 -6.980 1814.380 ;
        RECT 9.020 1814.370 12.020 1814.380 ;
        RECT 189.020 1814.370 192.020 1814.380 ;
        RECT 369.020 1814.370 372.020 1814.380 ;
        RECT 549.020 1814.370 552.020 1814.380 ;
        RECT 729.020 1814.370 732.020 1814.380 ;
        RECT 909.020 1814.370 912.020 1814.380 ;
        RECT 1089.020 1814.370 1092.020 1814.380 ;
        RECT 1269.020 1814.370 1272.020 1814.380 ;
        RECT 1449.020 1814.370 1452.020 1814.380 ;
        RECT 1629.020 1814.370 1632.020 1814.380 ;
        RECT 1809.020 1814.370 1812.020 1814.380 ;
        RECT 1989.020 1814.370 1992.020 1814.380 ;
        RECT 2169.020 1814.370 2172.020 1814.380 ;
        RECT 2349.020 1814.370 2352.020 1814.380 ;
        RECT 2529.020 1814.370 2532.020 1814.380 ;
        RECT 2709.020 1814.370 2712.020 1814.380 ;
        RECT 2889.020 1814.370 2892.020 1814.380 ;
        RECT 2926.600 1814.370 2929.600 1814.380 ;
        RECT -9.980 1637.380 -6.980 1637.390 ;
        RECT 9.020 1637.380 12.020 1637.390 ;
        RECT 189.020 1637.380 192.020 1637.390 ;
        RECT 369.020 1637.380 372.020 1637.390 ;
        RECT 549.020 1637.380 552.020 1637.390 ;
        RECT 729.020 1637.380 732.020 1637.390 ;
        RECT 909.020 1637.380 912.020 1637.390 ;
        RECT 1089.020 1637.380 1092.020 1637.390 ;
        RECT 1269.020 1637.380 1272.020 1637.390 ;
        RECT 1449.020 1637.380 1452.020 1637.390 ;
        RECT 1629.020 1637.380 1632.020 1637.390 ;
        RECT 1809.020 1637.380 1812.020 1637.390 ;
        RECT 1989.020 1637.380 1992.020 1637.390 ;
        RECT 2169.020 1637.380 2172.020 1637.390 ;
        RECT 2349.020 1637.380 2352.020 1637.390 ;
        RECT 2529.020 1637.380 2532.020 1637.390 ;
        RECT 2709.020 1637.380 2712.020 1637.390 ;
        RECT 2889.020 1637.380 2892.020 1637.390 ;
        RECT 2926.600 1637.380 2929.600 1637.390 ;
        RECT -14.680 1634.380 2934.300 1637.380 ;
        RECT -9.980 1634.370 -6.980 1634.380 ;
        RECT 9.020 1634.370 12.020 1634.380 ;
        RECT 189.020 1634.370 192.020 1634.380 ;
        RECT 369.020 1634.370 372.020 1634.380 ;
        RECT 549.020 1634.370 552.020 1634.380 ;
        RECT 729.020 1634.370 732.020 1634.380 ;
        RECT 909.020 1634.370 912.020 1634.380 ;
        RECT 1089.020 1634.370 1092.020 1634.380 ;
        RECT 1269.020 1634.370 1272.020 1634.380 ;
        RECT 1449.020 1634.370 1452.020 1634.380 ;
        RECT 1629.020 1634.370 1632.020 1634.380 ;
        RECT 1809.020 1634.370 1812.020 1634.380 ;
        RECT 1989.020 1634.370 1992.020 1634.380 ;
        RECT 2169.020 1634.370 2172.020 1634.380 ;
        RECT 2349.020 1634.370 2352.020 1634.380 ;
        RECT 2529.020 1634.370 2532.020 1634.380 ;
        RECT 2709.020 1634.370 2712.020 1634.380 ;
        RECT 2889.020 1634.370 2892.020 1634.380 ;
        RECT 2926.600 1634.370 2929.600 1634.380 ;
        RECT -9.980 1457.380 -6.980 1457.390 ;
        RECT 9.020 1457.380 12.020 1457.390 ;
        RECT 189.020 1457.380 192.020 1457.390 ;
        RECT 369.020 1457.380 372.020 1457.390 ;
        RECT 549.020 1457.380 552.020 1457.390 ;
        RECT 729.020 1457.380 732.020 1457.390 ;
        RECT 909.020 1457.380 912.020 1457.390 ;
        RECT 1089.020 1457.380 1092.020 1457.390 ;
        RECT 1269.020 1457.380 1272.020 1457.390 ;
        RECT 1449.020 1457.380 1452.020 1457.390 ;
        RECT 1629.020 1457.380 1632.020 1457.390 ;
        RECT 1809.020 1457.380 1812.020 1457.390 ;
        RECT 1989.020 1457.380 1992.020 1457.390 ;
        RECT 2169.020 1457.380 2172.020 1457.390 ;
        RECT 2349.020 1457.380 2352.020 1457.390 ;
        RECT 2529.020 1457.380 2532.020 1457.390 ;
        RECT 2709.020 1457.380 2712.020 1457.390 ;
        RECT 2889.020 1457.380 2892.020 1457.390 ;
        RECT 2926.600 1457.380 2929.600 1457.390 ;
        RECT -14.680 1454.380 2934.300 1457.380 ;
        RECT -9.980 1454.370 -6.980 1454.380 ;
        RECT 9.020 1454.370 12.020 1454.380 ;
        RECT 189.020 1454.370 192.020 1454.380 ;
        RECT 369.020 1454.370 372.020 1454.380 ;
        RECT 549.020 1454.370 552.020 1454.380 ;
        RECT 729.020 1454.370 732.020 1454.380 ;
        RECT 909.020 1454.370 912.020 1454.380 ;
        RECT 1089.020 1454.370 1092.020 1454.380 ;
        RECT 1269.020 1454.370 1272.020 1454.380 ;
        RECT 1449.020 1454.370 1452.020 1454.380 ;
        RECT 1629.020 1454.370 1632.020 1454.380 ;
        RECT 1809.020 1454.370 1812.020 1454.380 ;
        RECT 1989.020 1454.370 1992.020 1454.380 ;
        RECT 2169.020 1454.370 2172.020 1454.380 ;
        RECT 2349.020 1454.370 2352.020 1454.380 ;
        RECT 2529.020 1454.370 2532.020 1454.380 ;
        RECT 2709.020 1454.370 2712.020 1454.380 ;
        RECT 2889.020 1454.370 2892.020 1454.380 ;
        RECT 2926.600 1454.370 2929.600 1454.380 ;
        RECT -9.980 1277.380 -6.980 1277.390 ;
        RECT 9.020 1277.380 12.020 1277.390 ;
        RECT 189.020 1277.380 192.020 1277.390 ;
        RECT 369.020 1277.380 372.020 1277.390 ;
        RECT 549.020 1277.380 552.020 1277.390 ;
        RECT 729.020 1277.380 732.020 1277.390 ;
        RECT 909.020 1277.380 912.020 1277.390 ;
        RECT 1089.020 1277.380 1092.020 1277.390 ;
        RECT 1269.020 1277.380 1272.020 1277.390 ;
        RECT 1449.020 1277.380 1452.020 1277.390 ;
        RECT 1629.020 1277.380 1632.020 1277.390 ;
        RECT 1809.020 1277.380 1812.020 1277.390 ;
        RECT 1989.020 1277.380 1992.020 1277.390 ;
        RECT 2169.020 1277.380 2172.020 1277.390 ;
        RECT 2349.020 1277.380 2352.020 1277.390 ;
        RECT 2529.020 1277.380 2532.020 1277.390 ;
        RECT 2709.020 1277.380 2712.020 1277.390 ;
        RECT 2889.020 1277.380 2892.020 1277.390 ;
        RECT 2926.600 1277.380 2929.600 1277.390 ;
        RECT -14.680 1274.380 2934.300 1277.380 ;
        RECT -9.980 1274.370 -6.980 1274.380 ;
        RECT 9.020 1274.370 12.020 1274.380 ;
        RECT 189.020 1274.370 192.020 1274.380 ;
        RECT 369.020 1274.370 372.020 1274.380 ;
        RECT 549.020 1274.370 552.020 1274.380 ;
        RECT 729.020 1274.370 732.020 1274.380 ;
        RECT 909.020 1274.370 912.020 1274.380 ;
        RECT 1089.020 1274.370 1092.020 1274.380 ;
        RECT 1269.020 1274.370 1272.020 1274.380 ;
        RECT 1449.020 1274.370 1452.020 1274.380 ;
        RECT 1629.020 1274.370 1632.020 1274.380 ;
        RECT 1809.020 1274.370 1812.020 1274.380 ;
        RECT 1989.020 1274.370 1992.020 1274.380 ;
        RECT 2169.020 1274.370 2172.020 1274.380 ;
        RECT 2349.020 1274.370 2352.020 1274.380 ;
        RECT 2529.020 1274.370 2532.020 1274.380 ;
        RECT 2709.020 1274.370 2712.020 1274.380 ;
        RECT 2889.020 1274.370 2892.020 1274.380 ;
        RECT 2926.600 1274.370 2929.600 1274.380 ;
        RECT -9.980 1097.380 -6.980 1097.390 ;
        RECT 9.020 1097.380 12.020 1097.390 ;
        RECT 189.020 1097.380 192.020 1097.390 ;
        RECT 369.020 1097.380 372.020 1097.390 ;
        RECT 549.020 1097.380 552.020 1097.390 ;
        RECT 729.020 1097.380 732.020 1097.390 ;
        RECT 909.020 1097.380 912.020 1097.390 ;
        RECT 1089.020 1097.380 1092.020 1097.390 ;
        RECT 1269.020 1097.380 1272.020 1097.390 ;
        RECT 1449.020 1097.380 1452.020 1097.390 ;
        RECT 1629.020 1097.380 1632.020 1097.390 ;
        RECT 1809.020 1097.380 1812.020 1097.390 ;
        RECT 1989.020 1097.380 1992.020 1097.390 ;
        RECT 2169.020 1097.380 2172.020 1097.390 ;
        RECT 2349.020 1097.380 2352.020 1097.390 ;
        RECT 2529.020 1097.380 2532.020 1097.390 ;
        RECT 2709.020 1097.380 2712.020 1097.390 ;
        RECT 2889.020 1097.380 2892.020 1097.390 ;
        RECT 2926.600 1097.380 2929.600 1097.390 ;
        RECT -14.680 1094.380 2934.300 1097.380 ;
        RECT -9.980 1094.370 -6.980 1094.380 ;
        RECT 9.020 1094.370 12.020 1094.380 ;
        RECT 189.020 1094.370 192.020 1094.380 ;
        RECT 369.020 1094.370 372.020 1094.380 ;
        RECT 549.020 1094.370 552.020 1094.380 ;
        RECT 729.020 1094.370 732.020 1094.380 ;
        RECT 909.020 1094.370 912.020 1094.380 ;
        RECT 1089.020 1094.370 1092.020 1094.380 ;
        RECT 1269.020 1094.370 1272.020 1094.380 ;
        RECT 1449.020 1094.370 1452.020 1094.380 ;
        RECT 1629.020 1094.370 1632.020 1094.380 ;
        RECT 1809.020 1094.370 1812.020 1094.380 ;
        RECT 1989.020 1094.370 1992.020 1094.380 ;
        RECT 2169.020 1094.370 2172.020 1094.380 ;
        RECT 2349.020 1094.370 2352.020 1094.380 ;
        RECT 2529.020 1094.370 2532.020 1094.380 ;
        RECT 2709.020 1094.370 2712.020 1094.380 ;
        RECT 2889.020 1094.370 2892.020 1094.380 ;
        RECT 2926.600 1094.370 2929.600 1094.380 ;
        RECT -9.980 917.380 -6.980 917.390 ;
        RECT 9.020 917.380 12.020 917.390 ;
        RECT 189.020 917.380 192.020 917.390 ;
        RECT 369.020 917.380 372.020 917.390 ;
        RECT 549.020 917.380 552.020 917.390 ;
        RECT 729.020 917.380 732.020 917.390 ;
        RECT 909.020 917.380 912.020 917.390 ;
        RECT 1089.020 917.380 1092.020 917.390 ;
        RECT 1269.020 917.380 1272.020 917.390 ;
        RECT 1449.020 917.380 1452.020 917.390 ;
        RECT 1629.020 917.380 1632.020 917.390 ;
        RECT 1809.020 917.380 1812.020 917.390 ;
        RECT 1989.020 917.380 1992.020 917.390 ;
        RECT 2169.020 917.380 2172.020 917.390 ;
        RECT 2349.020 917.380 2352.020 917.390 ;
        RECT 2529.020 917.380 2532.020 917.390 ;
        RECT 2709.020 917.380 2712.020 917.390 ;
        RECT 2889.020 917.380 2892.020 917.390 ;
        RECT 2926.600 917.380 2929.600 917.390 ;
        RECT -14.680 914.380 2934.300 917.380 ;
        RECT -9.980 914.370 -6.980 914.380 ;
        RECT 9.020 914.370 12.020 914.380 ;
        RECT 189.020 914.370 192.020 914.380 ;
        RECT 369.020 914.370 372.020 914.380 ;
        RECT 549.020 914.370 552.020 914.380 ;
        RECT 729.020 914.370 732.020 914.380 ;
        RECT 909.020 914.370 912.020 914.380 ;
        RECT 1089.020 914.370 1092.020 914.380 ;
        RECT 1269.020 914.370 1272.020 914.380 ;
        RECT 1449.020 914.370 1452.020 914.380 ;
        RECT 1629.020 914.370 1632.020 914.380 ;
        RECT 1809.020 914.370 1812.020 914.380 ;
        RECT 1989.020 914.370 1992.020 914.380 ;
        RECT 2169.020 914.370 2172.020 914.380 ;
        RECT 2349.020 914.370 2352.020 914.380 ;
        RECT 2529.020 914.370 2532.020 914.380 ;
        RECT 2709.020 914.370 2712.020 914.380 ;
        RECT 2889.020 914.370 2892.020 914.380 ;
        RECT 2926.600 914.370 2929.600 914.380 ;
        RECT -9.980 737.380 -6.980 737.390 ;
        RECT 9.020 737.380 12.020 737.390 ;
        RECT 189.020 737.380 192.020 737.390 ;
        RECT 369.020 737.380 372.020 737.390 ;
        RECT 549.020 737.380 552.020 737.390 ;
        RECT 729.020 737.380 732.020 737.390 ;
        RECT 909.020 737.380 912.020 737.390 ;
        RECT 1089.020 737.380 1092.020 737.390 ;
        RECT 1269.020 737.380 1272.020 737.390 ;
        RECT 1449.020 737.380 1452.020 737.390 ;
        RECT 1629.020 737.380 1632.020 737.390 ;
        RECT 1809.020 737.380 1812.020 737.390 ;
        RECT 1989.020 737.380 1992.020 737.390 ;
        RECT 2169.020 737.380 2172.020 737.390 ;
        RECT 2349.020 737.380 2352.020 737.390 ;
        RECT 2529.020 737.380 2532.020 737.390 ;
        RECT 2709.020 737.380 2712.020 737.390 ;
        RECT 2889.020 737.380 2892.020 737.390 ;
        RECT 2926.600 737.380 2929.600 737.390 ;
        RECT -14.680 734.380 2934.300 737.380 ;
        RECT -9.980 734.370 -6.980 734.380 ;
        RECT 9.020 734.370 12.020 734.380 ;
        RECT 189.020 734.370 192.020 734.380 ;
        RECT 369.020 734.370 372.020 734.380 ;
        RECT 549.020 734.370 552.020 734.380 ;
        RECT 729.020 734.370 732.020 734.380 ;
        RECT 909.020 734.370 912.020 734.380 ;
        RECT 1089.020 734.370 1092.020 734.380 ;
        RECT 1269.020 734.370 1272.020 734.380 ;
        RECT 1449.020 734.370 1452.020 734.380 ;
        RECT 1629.020 734.370 1632.020 734.380 ;
        RECT 1809.020 734.370 1812.020 734.380 ;
        RECT 1989.020 734.370 1992.020 734.380 ;
        RECT 2169.020 734.370 2172.020 734.380 ;
        RECT 2349.020 734.370 2352.020 734.380 ;
        RECT 2529.020 734.370 2532.020 734.380 ;
        RECT 2709.020 734.370 2712.020 734.380 ;
        RECT 2889.020 734.370 2892.020 734.380 ;
        RECT 2926.600 734.370 2929.600 734.380 ;
        RECT -9.980 557.380 -6.980 557.390 ;
        RECT 9.020 557.380 12.020 557.390 ;
        RECT 189.020 557.380 192.020 557.390 ;
        RECT 369.020 557.380 372.020 557.390 ;
        RECT 549.020 557.380 552.020 557.390 ;
        RECT 729.020 557.380 732.020 557.390 ;
        RECT 909.020 557.380 912.020 557.390 ;
        RECT 1089.020 557.380 1092.020 557.390 ;
        RECT 1269.020 557.380 1272.020 557.390 ;
        RECT 1449.020 557.380 1452.020 557.390 ;
        RECT 1629.020 557.380 1632.020 557.390 ;
        RECT 1809.020 557.380 1812.020 557.390 ;
        RECT 1989.020 557.380 1992.020 557.390 ;
        RECT 2169.020 557.380 2172.020 557.390 ;
        RECT 2349.020 557.380 2352.020 557.390 ;
        RECT 2529.020 557.380 2532.020 557.390 ;
        RECT 2709.020 557.380 2712.020 557.390 ;
        RECT 2889.020 557.380 2892.020 557.390 ;
        RECT 2926.600 557.380 2929.600 557.390 ;
        RECT -14.680 554.380 2934.300 557.380 ;
        RECT -9.980 554.370 -6.980 554.380 ;
        RECT 9.020 554.370 12.020 554.380 ;
        RECT 189.020 554.370 192.020 554.380 ;
        RECT 369.020 554.370 372.020 554.380 ;
        RECT 549.020 554.370 552.020 554.380 ;
        RECT 729.020 554.370 732.020 554.380 ;
        RECT 909.020 554.370 912.020 554.380 ;
        RECT 1089.020 554.370 1092.020 554.380 ;
        RECT 1269.020 554.370 1272.020 554.380 ;
        RECT 1449.020 554.370 1452.020 554.380 ;
        RECT 1629.020 554.370 1632.020 554.380 ;
        RECT 1809.020 554.370 1812.020 554.380 ;
        RECT 1989.020 554.370 1992.020 554.380 ;
        RECT 2169.020 554.370 2172.020 554.380 ;
        RECT 2349.020 554.370 2352.020 554.380 ;
        RECT 2529.020 554.370 2532.020 554.380 ;
        RECT 2709.020 554.370 2712.020 554.380 ;
        RECT 2889.020 554.370 2892.020 554.380 ;
        RECT 2926.600 554.370 2929.600 554.380 ;
        RECT -9.980 377.380 -6.980 377.390 ;
        RECT 9.020 377.380 12.020 377.390 ;
        RECT 189.020 377.380 192.020 377.390 ;
        RECT 369.020 377.380 372.020 377.390 ;
        RECT 549.020 377.380 552.020 377.390 ;
        RECT 729.020 377.380 732.020 377.390 ;
        RECT 909.020 377.380 912.020 377.390 ;
        RECT 1089.020 377.380 1092.020 377.390 ;
        RECT 1269.020 377.380 1272.020 377.390 ;
        RECT 1449.020 377.380 1452.020 377.390 ;
        RECT 1629.020 377.380 1632.020 377.390 ;
        RECT 1809.020 377.380 1812.020 377.390 ;
        RECT 1989.020 377.380 1992.020 377.390 ;
        RECT 2169.020 377.380 2172.020 377.390 ;
        RECT 2349.020 377.380 2352.020 377.390 ;
        RECT 2529.020 377.380 2532.020 377.390 ;
        RECT 2709.020 377.380 2712.020 377.390 ;
        RECT 2889.020 377.380 2892.020 377.390 ;
        RECT 2926.600 377.380 2929.600 377.390 ;
        RECT -14.680 374.380 2934.300 377.380 ;
        RECT -9.980 374.370 -6.980 374.380 ;
        RECT 9.020 374.370 12.020 374.380 ;
        RECT 189.020 374.370 192.020 374.380 ;
        RECT 369.020 374.370 372.020 374.380 ;
        RECT 549.020 374.370 552.020 374.380 ;
        RECT 729.020 374.370 732.020 374.380 ;
        RECT 909.020 374.370 912.020 374.380 ;
        RECT 1089.020 374.370 1092.020 374.380 ;
        RECT 1269.020 374.370 1272.020 374.380 ;
        RECT 1449.020 374.370 1452.020 374.380 ;
        RECT 1629.020 374.370 1632.020 374.380 ;
        RECT 1809.020 374.370 1812.020 374.380 ;
        RECT 1989.020 374.370 1992.020 374.380 ;
        RECT 2169.020 374.370 2172.020 374.380 ;
        RECT 2349.020 374.370 2352.020 374.380 ;
        RECT 2529.020 374.370 2532.020 374.380 ;
        RECT 2709.020 374.370 2712.020 374.380 ;
        RECT 2889.020 374.370 2892.020 374.380 ;
        RECT 2926.600 374.370 2929.600 374.380 ;
        RECT -9.980 197.380 -6.980 197.390 ;
        RECT 9.020 197.380 12.020 197.390 ;
        RECT 189.020 197.380 192.020 197.390 ;
        RECT 369.020 197.380 372.020 197.390 ;
        RECT 549.020 197.380 552.020 197.390 ;
        RECT 729.020 197.380 732.020 197.390 ;
        RECT 909.020 197.380 912.020 197.390 ;
        RECT 1089.020 197.380 1092.020 197.390 ;
        RECT 1269.020 197.380 1272.020 197.390 ;
        RECT 1449.020 197.380 1452.020 197.390 ;
        RECT 1629.020 197.380 1632.020 197.390 ;
        RECT 1809.020 197.380 1812.020 197.390 ;
        RECT 1989.020 197.380 1992.020 197.390 ;
        RECT 2169.020 197.380 2172.020 197.390 ;
        RECT 2349.020 197.380 2352.020 197.390 ;
        RECT 2529.020 197.380 2532.020 197.390 ;
        RECT 2709.020 197.380 2712.020 197.390 ;
        RECT 2889.020 197.380 2892.020 197.390 ;
        RECT 2926.600 197.380 2929.600 197.390 ;
        RECT -14.680 194.380 2934.300 197.380 ;
        RECT -9.980 194.370 -6.980 194.380 ;
        RECT 9.020 194.370 12.020 194.380 ;
        RECT 189.020 194.370 192.020 194.380 ;
        RECT 369.020 194.370 372.020 194.380 ;
        RECT 549.020 194.370 552.020 194.380 ;
        RECT 729.020 194.370 732.020 194.380 ;
        RECT 909.020 194.370 912.020 194.380 ;
        RECT 1089.020 194.370 1092.020 194.380 ;
        RECT 1269.020 194.370 1272.020 194.380 ;
        RECT 1449.020 194.370 1452.020 194.380 ;
        RECT 1629.020 194.370 1632.020 194.380 ;
        RECT 1809.020 194.370 1812.020 194.380 ;
        RECT 1989.020 194.370 1992.020 194.380 ;
        RECT 2169.020 194.370 2172.020 194.380 ;
        RECT 2349.020 194.370 2352.020 194.380 ;
        RECT 2529.020 194.370 2532.020 194.380 ;
        RECT 2709.020 194.370 2712.020 194.380 ;
        RECT 2889.020 194.370 2892.020 194.380 ;
        RECT 2926.600 194.370 2929.600 194.380 ;
        RECT -9.980 17.380 -6.980 17.390 ;
        RECT 9.020 17.380 12.020 17.390 ;
        RECT 189.020 17.380 192.020 17.390 ;
        RECT 369.020 17.380 372.020 17.390 ;
        RECT 549.020 17.380 552.020 17.390 ;
        RECT 729.020 17.380 732.020 17.390 ;
        RECT 909.020 17.380 912.020 17.390 ;
        RECT 1089.020 17.380 1092.020 17.390 ;
        RECT 1269.020 17.380 1272.020 17.390 ;
        RECT 1449.020 17.380 1452.020 17.390 ;
        RECT 1629.020 17.380 1632.020 17.390 ;
        RECT 1809.020 17.380 1812.020 17.390 ;
        RECT 1989.020 17.380 1992.020 17.390 ;
        RECT 2169.020 17.380 2172.020 17.390 ;
        RECT 2349.020 17.380 2352.020 17.390 ;
        RECT 2529.020 17.380 2532.020 17.390 ;
        RECT 2709.020 17.380 2712.020 17.390 ;
        RECT 2889.020 17.380 2892.020 17.390 ;
        RECT 2926.600 17.380 2929.600 17.390 ;
        RECT -14.680 14.380 2934.300 17.380 ;
        RECT -9.980 14.370 -6.980 14.380 ;
        RECT 9.020 14.370 12.020 14.380 ;
        RECT 189.020 14.370 192.020 14.380 ;
        RECT 369.020 14.370 372.020 14.380 ;
        RECT 549.020 14.370 552.020 14.380 ;
        RECT 729.020 14.370 732.020 14.380 ;
        RECT 909.020 14.370 912.020 14.380 ;
        RECT 1089.020 14.370 1092.020 14.380 ;
        RECT 1269.020 14.370 1272.020 14.380 ;
        RECT 1449.020 14.370 1452.020 14.380 ;
        RECT 1629.020 14.370 1632.020 14.380 ;
        RECT 1809.020 14.370 1812.020 14.380 ;
        RECT 1989.020 14.370 1992.020 14.380 ;
        RECT 2169.020 14.370 2172.020 14.380 ;
        RECT 2349.020 14.370 2352.020 14.380 ;
        RECT 2529.020 14.370 2532.020 14.380 ;
        RECT 2709.020 14.370 2712.020 14.380 ;
        RECT 2889.020 14.370 2892.020 14.380 ;
        RECT 2926.600 14.370 2929.600 14.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 9.020 -1.620 12.020 -1.610 ;
        RECT 189.020 -1.620 192.020 -1.610 ;
        RECT 369.020 -1.620 372.020 -1.610 ;
        RECT 549.020 -1.620 552.020 -1.610 ;
        RECT 729.020 -1.620 732.020 -1.610 ;
        RECT 909.020 -1.620 912.020 -1.610 ;
        RECT 1089.020 -1.620 1092.020 -1.610 ;
        RECT 1269.020 -1.620 1272.020 -1.610 ;
        RECT 1449.020 -1.620 1452.020 -1.610 ;
        RECT 1629.020 -1.620 1632.020 -1.610 ;
        RECT 1809.020 -1.620 1812.020 -1.610 ;
        RECT 1989.020 -1.620 1992.020 -1.610 ;
        RECT 2169.020 -1.620 2172.020 -1.610 ;
        RECT 2349.020 -1.620 2352.020 -1.610 ;
        RECT 2529.020 -1.620 2532.020 -1.610 ;
        RECT 2709.020 -1.620 2712.020 -1.610 ;
        RECT 2889.020 -1.620 2892.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 9.020 -4.630 12.020 -4.620 ;
        RECT 189.020 -4.630 192.020 -4.620 ;
        RECT 369.020 -4.630 372.020 -4.620 ;
        RECT 549.020 -4.630 552.020 -4.620 ;
        RECT 729.020 -4.630 732.020 -4.620 ;
        RECT 909.020 -4.630 912.020 -4.620 ;
        RECT 1089.020 -4.630 1092.020 -4.620 ;
        RECT 1269.020 -4.630 1272.020 -4.620 ;
        RECT 1449.020 -4.630 1452.020 -4.620 ;
        RECT 1629.020 -4.630 1632.020 -4.620 ;
        RECT 1809.020 -4.630 1812.020 -4.620 ;
        RECT 1989.020 -4.630 1992.020 -4.620 ;
        RECT 2169.020 -4.630 2172.020 -4.620 ;
        RECT 2349.020 -4.630 2352.020 -4.620 ;
        RECT 2529.020 -4.630 2532.020 -4.620 ;
        RECT 2709.020 -4.630 2712.020 -4.620 ;
        RECT 2889.020 -4.630 2892.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 99.020 -9.320 102.020 3529.000 ;
        RECT 279.020 -9.320 282.020 3529.000 ;
        RECT 459.020 -9.320 462.020 3529.000 ;
        RECT 639.020 -9.320 642.020 3529.000 ;
        RECT 819.020 -9.320 822.020 3529.000 ;
        RECT 999.020 -9.320 1002.020 3529.000 ;
        RECT 1179.020 -9.320 1182.020 3529.000 ;
        RECT 1359.020 -9.320 1362.020 3529.000 ;
        RECT 1539.020 -9.320 1542.020 3529.000 ;
        RECT 1719.020 -9.320 1722.020 3529.000 ;
        RECT 1899.020 -9.320 1902.020 3529.000 ;
        RECT 2079.020 -9.320 2082.020 3529.000 ;
        RECT 2259.020 -9.320 2262.020 3529.000 ;
        RECT 2439.020 -9.320 2442.020 3529.000 ;
        RECT 2619.020 -9.320 2622.020 3529.000 ;
        RECT 2799.020 -9.320 2802.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3346.090 -12.590 3347.270 ;
        RECT -13.770 3344.490 -12.590 3345.670 ;
        RECT -13.770 3166.090 -12.590 3167.270 ;
        RECT -13.770 3164.490 -12.590 3165.670 ;
        RECT -13.770 2986.090 -12.590 2987.270 ;
        RECT -13.770 2984.490 -12.590 2985.670 ;
        RECT -13.770 2806.090 -12.590 2807.270 ;
        RECT -13.770 2804.490 -12.590 2805.670 ;
        RECT -13.770 2626.090 -12.590 2627.270 ;
        RECT -13.770 2624.490 -12.590 2625.670 ;
        RECT -13.770 2446.090 -12.590 2447.270 ;
        RECT -13.770 2444.490 -12.590 2445.670 ;
        RECT -13.770 2266.090 -12.590 2267.270 ;
        RECT -13.770 2264.490 -12.590 2265.670 ;
        RECT -13.770 2086.090 -12.590 2087.270 ;
        RECT -13.770 2084.490 -12.590 2085.670 ;
        RECT -13.770 1906.090 -12.590 1907.270 ;
        RECT -13.770 1904.490 -12.590 1905.670 ;
        RECT -13.770 1726.090 -12.590 1727.270 ;
        RECT -13.770 1724.490 -12.590 1725.670 ;
        RECT -13.770 1546.090 -12.590 1547.270 ;
        RECT -13.770 1544.490 -12.590 1545.670 ;
        RECT -13.770 1366.090 -12.590 1367.270 ;
        RECT -13.770 1364.490 -12.590 1365.670 ;
        RECT -13.770 1186.090 -12.590 1187.270 ;
        RECT -13.770 1184.490 -12.590 1185.670 ;
        RECT -13.770 1006.090 -12.590 1007.270 ;
        RECT -13.770 1004.490 -12.590 1005.670 ;
        RECT -13.770 826.090 -12.590 827.270 ;
        RECT -13.770 824.490 -12.590 825.670 ;
        RECT -13.770 646.090 -12.590 647.270 ;
        RECT -13.770 644.490 -12.590 645.670 ;
        RECT -13.770 466.090 -12.590 467.270 ;
        RECT -13.770 464.490 -12.590 465.670 ;
        RECT -13.770 286.090 -12.590 287.270 ;
        RECT -13.770 284.490 -12.590 285.670 ;
        RECT -13.770 106.090 -12.590 107.270 ;
        RECT -13.770 104.490 -12.590 105.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 99.930 3527.710 101.110 3528.890 ;
        RECT 99.930 3526.110 101.110 3527.290 ;
        RECT 99.930 3346.090 101.110 3347.270 ;
        RECT 99.930 3344.490 101.110 3345.670 ;
        RECT 99.930 3166.090 101.110 3167.270 ;
        RECT 99.930 3164.490 101.110 3165.670 ;
        RECT 99.930 2986.090 101.110 2987.270 ;
        RECT 99.930 2984.490 101.110 2985.670 ;
        RECT 99.930 2806.090 101.110 2807.270 ;
        RECT 99.930 2804.490 101.110 2805.670 ;
        RECT 99.930 2626.090 101.110 2627.270 ;
        RECT 99.930 2624.490 101.110 2625.670 ;
        RECT 99.930 2446.090 101.110 2447.270 ;
        RECT 99.930 2444.490 101.110 2445.670 ;
        RECT 99.930 2266.090 101.110 2267.270 ;
        RECT 99.930 2264.490 101.110 2265.670 ;
        RECT 99.930 2086.090 101.110 2087.270 ;
        RECT 99.930 2084.490 101.110 2085.670 ;
        RECT 99.930 1906.090 101.110 1907.270 ;
        RECT 99.930 1904.490 101.110 1905.670 ;
        RECT 99.930 1726.090 101.110 1727.270 ;
        RECT 99.930 1724.490 101.110 1725.670 ;
        RECT 99.930 1546.090 101.110 1547.270 ;
        RECT 99.930 1544.490 101.110 1545.670 ;
        RECT 99.930 1366.090 101.110 1367.270 ;
        RECT 99.930 1364.490 101.110 1365.670 ;
        RECT 99.930 1186.090 101.110 1187.270 ;
        RECT 99.930 1184.490 101.110 1185.670 ;
        RECT 99.930 1006.090 101.110 1007.270 ;
        RECT 99.930 1004.490 101.110 1005.670 ;
        RECT 99.930 826.090 101.110 827.270 ;
        RECT 99.930 824.490 101.110 825.670 ;
        RECT 99.930 646.090 101.110 647.270 ;
        RECT 99.930 644.490 101.110 645.670 ;
        RECT 99.930 466.090 101.110 467.270 ;
        RECT 99.930 464.490 101.110 465.670 ;
        RECT 99.930 286.090 101.110 287.270 ;
        RECT 99.930 284.490 101.110 285.670 ;
        RECT 99.930 106.090 101.110 107.270 ;
        RECT 99.930 104.490 101.110 105.670 ;
        RECT 99.930 -7.610 101.110 -6.430 ;
        RECT 99.930 -9.210 101.110 -8.030 ;
        RECT 279.930 3527.710 281.110 3528.890 ;
        RECT 279.930 3526.110 281.110 3527.290 ;
        RECT 279.930 3346.090 281.110 3347.270 ;
        RECT 279.930 3344.490 281.110 3345.670 ;
        RECT 279.930 3166.090 281.110 3167.270 ;
        RECT 279.930 3164.490 281.110 3165.670 ;
        RECT 279.930 2986.090 281.110 2987.270 ;
        RECT 279.930 2984.490 281.110 2985.670 ;
        RECT 279.930 2806.090 281.110 2807.270 ;
        RECT 279.930 2804.490 281.110 2805.670 ;
        RECT 279.930 2626.090 281.110 2627.270 ;
        RECT 279.930 2624.490 281.110 2625.670 ;
        RECT 279.930 2446.090 281.110 2447.270 ;
        RECT 279.930 2444.490 281.110 2445.670 ;
        RECT 279.930 2266.090 281.110 2267.270 ;
        RECT 279.930 2264.490 281.110 2265.670 ;
        RECT 279.930 2086.090 281.110 2087.270 ;
        RECT 279.930 2084.490 281.110 2085.670 ;
        RECT 279.930 1906.090 281.110 1907.270 ;
        RECT 279.930 1904.490 281.110 1905.670 ;
        RECT 279.930 1726.090 281.110 1727.270 ;
        RECT 279.930 1724.490 281.110 1725.670 ;
        RECT 279.930 1546.090 281.110 1547.270 ;
        RECT 279.930 1544.490 281.110 1545.670 ;
        RECT 279.930 1366.090 281.110 1367.270 ;
        RECT 279.930 1364.490 281.110 1365.670 ;
        RECT 279.930 1186.090 281.110 1187.270 ;
        RECT 279.930 1184.490 281.110 1185.670 ;
        RECT 279.930 1006.090 281.110 1007.270 ;
        RECT 279.930 1004.490 281.110 1005.670 ;
        RECT 279.930 826.090 281.110 827.270 ;
        RECT 279.930 824.490 281.110 825.670 ;
        RECT 279.930 646.090 281.110 647.270 ;
        RECT 279.930 644.490 281.110 645.670 ;
        RECT 279.930 466.090 281.110 467.270 ;
        RECT 279.930 464.490 281.110 465.670 ;
        RECT 279.930 286.090 281.110 287.270 ;
        RECT 279.930 284.490 281.110 285.670 ;
        RECT 279.930 106.090 281.110 107.270 ;
        RECT 279.930 104.490 281.110 105.670 ;
        RECT 279.930 -7.610 281.110 -6.430 ;
        RECT 279.930 -9.210 281.110 -8.030 ;
        RECT 459.930 3527.710 461.110 3528.890 ;
        RECT 459.930 3526.110 461.110 3527.290 ;
        RECT 459.930 3346.090 461.110 3347.270 ;
        RECT 459.930 3344.490 461.110 3345.670 ;
        RECT 459.930 3166.090 461.110 3167.270 ;
        RECT 459.930 3164.490 461.110 3165.670 ;
        RECT 459.930 2986.090 461.110 2987.270 ;
        RECT 459.930 2984.490 461.110 2985.670 ;
        RECT 459.930 2806.090 461.110 2807.270 ;
        RECT 459.930 2804.490 461.110 2805.670 ;
        RECT 459.930 2626.090 461.110 2627.270 ;
        RECT 459.930 2624.490 461.110 2625.670 ;
        RECT 459.930 2446.090 461.110 2447.270 ;
        RECT 459.930 2444.490 461.110 2445.670 ;
        RECT 459.930 2266.090 461.110 2267.270 ;
        RECT 459.930 2264.490 461.110 2265.670 ;
        RECT 459.930 2086.090 461.110 2087.270 ;
        RECT 459.930 2084.490 461.110 2085.670 ;
        RECT 459.930 1906.090 461.110 1907.270 ;
        RECT 459.930 1904.490 461.110 1905.670 ;
        RECT 459.930 1726.090 461.110 1727.270 ;
        RECT 459.930 1724.490 461.110 1725.670 ;
        RECT 459.930 1546.090 461.110 1547.270 ;
        RECT 459.930 1544.490 461.110 1545.670 ;
        RECT 459.930 1366.090 461.110 1367.270 ;
        RECT 459.930 1364.490 461.110 1365.670 ;
        RECT 459.930 1186.090 461.110 1187.270 ;
        RECT 459.930 1184.490 461.110 1185.670 ;
        RECT 459.930 1006.090 461.110 1007.270 ;
        RECT 459.930 1004.490 461.110 1005.670 ;
        RECT 459.930 826.090 461.110 827.270 ;
        RECT 459.930 824.490 461.110 825.670 ;
        RECT 459.930 646.090 461.110 647.270 ;
        RECT 459.930 644.490 461.110 645.670 ;
        RECT 459.930 466.090 461.110 467.270 ;
        RECT 459.930 464.490 461.110 465.670 ;
        RECT 459.930 286.090 461.110 287.270 ;
        RECT 459.930 284.490 461.110 285.670 ;
        RECT 459.930 106.090 461.110 107.270 ;
        RECT 459.930 104.490 461.110 105.670 ;
        RECT 459.930 -7.610 461.110 -6.430 ;
        RECT 459.930 -9.210 461.110 -8.030 ;
        RECT 639.930 3527.710 641.110 3528.890 ;
        RECT 639.930 3526.110 641.110 3527.290 ;
        RECT 639.930 3346.090 641.110 3347.270 ;
        RECT 639.930 3344.490 641.110 3345.670 ;
        RECT 639.930 3166.090 641.110 3167.270 ;
        RECT 639.930 3164.490 641.110 3165.670 ;
        RECT 639.930 2986.090 641.110 2987.270 ;
        RECT 639.930 2984.490 641.110 2985.670 ;
        RECT 639.930 2806.090 641.110 2807.270 ;
        RECT 639.930 2804.490 641.110 2805.670 ;
        RECT 639.930 2626.090 641.110 2627.270 ;
        RECT 639.930 2624.490 641.110 2625.670 ;
        RECT 639.930 2446.090 641.110 2447.270 ;
        RECT 639.930 2444.490 641.110 2445.670 ;
        RECT 639.930 2266.090 641.110 2267.270 ;
        RECT 639.930 2264.490 641.110 2265.670 ;
        RECT 639.930 2086.090 641.110 2087.270 ;
        RECT 639.930 2084.490 641.110 2085.670 ;
        RECT 639.930 1906.090 641.110 1907.270 ;
        RECT 639.930 1904.490 641.110 1905.670 ;
        RECT 639.930 1726.090 641.110 1727.270 ;
        RECT 639.930 1724.490 641.110 1725.670 ;
        RECT 639.930 1546.090 641.110 1547.270 ;
        RECT 639.930 1544.490 641.110 1545.670 ;
        RECT 639.930 1366.090 641.110 1367.270 ;
        RECT 639.930 1364.490 641.110 1365.670 ;
        RECT 639.930 1186.090 641.110 1187.270 ;
        RECT 639.930 1184.490 641.110 1185.670 ;
        RECT 639.930 1006.090 641.110 1007.270 ;
        RECT 639.930 1004.490 641.110 1005.670 ;
        RECT 639.930 826.090 641.110 827.270 ;
        RECT 639.930 824.490 641.110 825.670 ;
        RECT 639.930 646.090 641.110 647.270 ;
        RECT 639.930 644.490 641.110 645.670 ;
        RECT 639.930 466.090 641.110 467.270 ;
        RECT 639.930 464.490 641.110 465.670 ;
        RECT 639.930 286.090 641.110 287.270 ;
        RECT 639.930 284.490 641.110 285.670 ;
        RECT 639.930 106.090 641.110 107.270 ;
        RECT 639.930 104.490 641.110 105.670 ;
        RECT 639.930 -7.610 641.110 -6.430 ;
        RECT 639.930 -9.210 641.110 -8.030 ;
        RECT 819.930 3527.710 821.110 3528.890 ;
        RECT 819.930 3526.110 821.110 3527.290 ;
        RECT 819.930 3346.090 821.110 3347.270 ;
        RECT 819.930 3344.490 821.110 3345.670 ;
        RECT 819.930 3166.090 821.110 3167.270 ;
        RECT 819.930 3164.490 821.110 3165.670 ;
        RECT 819.930 2986.090 821.110 2987.270 ;
        RECT 819.930 2984.490 821.110 2985.670 ;
        RECT 819.930 2806.090 821.110 2807.270 ;
        RECT 819.930 2804.490 821.110 2805.670 ;
        RECT 819.930 2626.090 821.110 2627.270 ;
        RECT 819.930 2624.490 821.110 2625.670 ;
        RECT 819.930 2446.090 821.110 2447.270 ;
        RECT 819.930 2444.490 821.110 2445.670 ;
        RECT 819.930 2266.090 821.110 2267.270 ;
        RECT 819.930 2264.490 821.110 2265.670 ;
        RECT 819.930 2086.090 821.110 2087.270 ;
        RECT 819.930 2084.490 821.110 2085.670 ;
        RECT 819.930 1906.090 821.110 1907.270 ;
        RECT 819.930 1904.490 821.110 1905.670 ;
        RECT 819.930 1726.090 821.110 1727.270 ;
        RECT 819.930 1724.490 821.110 1725.670 ;
        RECT 819.930 1546.090 821.110 1547.270 ;
        RECT 819.930 1544.490 821.110 1545.670 ;
        RECT 819.930 1366.090 821.110 1367.270 ;
        RECT 819.930 1364.490 821.110 1365.670 ;
        RECT 819.930 1186.090 821.110 1187.270 ;
        RECT 819.930 1184.490 821.110 1185.670 ;
        RECT 819.930 1006.090 821.110 1007.270 ;
        RECT 819.930 1004.490 821.110 1005.670 ;
        RECT 819.930 826.090 821.110 827.270 ;
        RECT 819.930 824.490 821.110 825.670 ;
        RECT 819.930 646.090 821.110 647.270 ;
        RECT 819.930 644.490 821.110 645.670 ;
        RECT 819.930 466.090 821.110 467.270 ;
        RECT 819.930 464.490 821.110 465.670 ;
        RECT 819.930 286.090 821.110 287.270 ;
        RECT 819.930 284.490 821.110 285.670 ;
        RECT 819.930 106.090 821.110 107.270 ;
        RECT 819.930 104.490 821.110 105.670 ;
        RECT 819.930 -7.610 821.110 -6.430 ;
        RECT 819.930 -9.210 821.110 -8.030 ;
        RECT 999.930 3527.710 1001.110 3528.890 ;
        RECT 999.930 3526.110 1001.110 3527.290 ;
        RECT 999.930 3346.090 1001.110 3347.270 ;
        RECT 999.930 3344.490 1001.110 3345.670 ;
        RECT 999.930 3166.090 1001.110 3167.270 ;
        RECT 999.930 3164.490 1001.110 3165.670 ;
        RECT 999.930 2986.090 1001.110 2987.270 ;
        RECT 999.930 2984.490 1001.110 2985.670 ;
        RECT 999.930 2806.090 1001.110 2807.270 ;
        RECT 999.930 2804.490 1001.110 2805.670 ;
        RECT 999.930 2626.090 1001.110 2627.270 ;
        RECT 999.930 2624.490 1001.110 2625.670 ;
        RECT 999.930 2446.090 1001.110 2447.270 ;
        RECT 999.930 2444.490 1001.110 2445.670 ;
        RECT 999.930 2266.090 1001.110 2267.270 ;
        RECT 999.930 2264.490 1001.110 2265.670 ;
        RECT 999.930 2086.090 1001.110 2087.270 ;
        RECT 999.930 2084.490 1001.110 2085.670 ;
        RECT 999.930 1906.090 1001.110 1907.270 ;
        RECT 999.930 1904.490 1001.110 1905.670 ;
        RECT 999.930 1726.090 1001.110 1727.270 ;
        RECT 999.930 1724.490 1001.110 1725.670 ;
        RECT 999.930 1546.090 1001.110 1547.270 ;
        RECT 999.930 1544.490 1001.110 1545.670 ;
        RECT 999.930 1366.090 1001.110 1367.270 ;
        RECT 999.930 1364.490 1001.110 1365.670 ;
        RECT 999.930 1186.090 1001.110 1187.270 ;
        RECT 999.930 1184.490 1001.110 1185.670 ;
        RECT 999.930 1006.090 1001.110 1007.270 ;
        RECT 999.930 1004.490 1001.110 1005.670 ;
        RECT 999.930 826.090 1001.110 827.270 ;
        RECT 999.930 824.490 1001.110 825.670 ;
        RECT 999.930 646.090 1001.110 647.270 ;
        RECT 999.930 644.490 1001.110 645.670 ;
        RECT 999.930 466.090 1001.110 467.270 ;
        RECT 999.930 464.490 1001.110 465.670 ;
        RECT 999.930 286.090 1001.110 287.270 ;
        RECT 999.930 284.490 1001.110 285.670 ;
        RECT 999.930 106.090 1001.110 107.270 ;
        RECT 999.930 104.490 1001.110 105.670 ;
        RECT 999.930 -7.610 1001.110 -6.430 ;
        RECT 999.930 -9.210 1001.110 -8.030 ;
        RECT 1179.930 3527.710 1181.110 3528.890 ;
        RECT 1179.930 3526.110 1181.110 3527.290 ;
        RECT 1179.930 3346.090 1181.110 3347.270 ;
        RECT 1179.930 3344.490 1181.110 3345.670 ;
        RECT 1179.930 3166.090 1181.110 3167.270 ;
        RECT 1179.930 3164.490 1181.110 3165.670 ;
        RECT 1179.930 2986.090 1181.110 2987.270 ;
        RECT 1179.930 2984.490 1181.110 2985.670 ;
        RECT 1179.930 2806.090 1181.110 2807.270 ;
        RECT 1179.930 2804.490 1181.110 2805.670 ;
        RECT 1179.930 2626.090 1181.110 2627.270 ;
        RECT 1179.930 2624.490 1181.110 2625.670 ;
        RECT 1179.930 2446.090 1181.110 2447.270 ;
        RECT 1179.930 2444.490 1181.110 2445.670 ;
        RECT 1179.930 2266.090 1181.110 2267.270 ;
        RECT 1179.930 2264.490 1181.110 2265.670 ;
        RECT 1179.930 2086.090 1181.110 2087.270 ;
        RECT 1179.930 2084.490 1181.110 2085.670 ;
        RECT 1179.930 1906.090 1181.110 1907.270 ;
        RECT 1179.930 1904.490 1181.110 1905.670 ;
        RECT 1179.930 1726.090 1181.110 1727.270 ;
        RECT 1179.930 1724.490 1181.110 1725.670 ;
        RECT 1179.930 1546.090 1181.110 1547.270 ;
        RECT 1179.930 1544.490 1181.110 1545.670 ;
        RECT 1179.930 1366.090 1181.110 1367.270 ;
        RECT 1179.930 1364.490 1181.110 1365.670 ;
        RECT 1179.930 1186.090 1181.110 1187.270 ;
        RECT 1179.930 1184.490 1181.110 1185.670 ;
        RECT 1179.930 1006.090 1181.110 1007.270 ;
        RECT 1179.930 1004.490 1181.110 1005.670 ;
        RECT 1179.930 826.090 1181.110 827.270 ;
        RECT 1179.930 824.490 1181.110 825.670 ;
        RECT 1179.930 646.090 1181.110 647.270 ;
        RECT 1179.930 644.490 1181.110 645.670 ;
        RECT 1179.930 466.090 1181.110 467.270 ;
        RECT 1179.930 464.490 1181.110 465.670 ;
        RECT 1179.930 286.090 1181.110 287.270 ;
        RECT 1179.930 284.490 1181.110 285.670 ;
        RECT 1179.930 106.090 1181.110 107.270 ;
        RECT 1179.930 104.490 1181.110 105.670 ;
        RECT 1179.930 -7.610 1181.110 -6.430 ;
        RECT 1179.930 -9.210 1181.110 -8.030 ;
        RECT 1359.930 3527.710 1361.110 3528.890 ;
        RECT 1359.930 3526.110 1361.110 3527.290 ;
        RECT 1359.930 3346.090 1361.110 3347.270 ;
        RECT 1359.930 3344.490 1361.110 3345.670 ;
        RECT 1359.930 3166.090 1361.110 3167.270 ;
        RECT 1359.930 3164.490 1361.110 3165.670 ;
        RECT 1359.930 2986.090 1361.110 2987.270 ;
        RECT 1359.930 2984.490 1361.110 2985.670 ;
        RECT 1359.930 2806.090 1361.110 2807.270 ;
        RECT 1359.930 2804.490 1361.110 2805.670 ;
        RECT 1359.930 2626.090 1361.110 2627.270 ;
        RECT 1359.930 2624.490 1361.110 2625.670 ;
        RECT 1359.930 2446.090 1361.110 2447.270 ;
        RECT 1359.930 2444.490 1361.110 2445.670 ;
        RECT 1359.930 2266.090 1361.110 2267.270 ;
        RECT 1359.930 2264.490 1361.110 2265.670 ;
        RECT 1359.930 2086.090 1361.110 2087.270 ;
        RECT 1359.930 2084.490 1361.110 2085.670 ;
        RECT 1359.930 1906.090 1361.110 1907.270 ;
        RECT 1359.930 1904.490 1361.110 1905.670 ;
        RECT 1359.930 1726.090 1361.110 1727.270 ;
        RECT 1359.930 1724.490 1361.110 1725.670 ;
        RECT 1359.930 1546.090 1361.110 1547.270 ;
        RECT 1359.930 1544.490 1361.110 1545.670 ;
        RECT 1359.930 1366.090 1361.110 1367.270 ;
        RECT 1359.930 1364.490 1361.110 1365.670 ;
        RECT 1359.930 1186.090 1361.110 1187.270 ;
        RECT 1359.930 1184.490 1361.110 1185.670 ;
        RECT 1359.930 1006.090 1361.110 1007.270 ;
        RECT 1359.930 1004.490 1361.110 1005.670 ;
        RECT 1359.930 826.090 1361.110 827.270 ;
        RECT 1359.930 824.490 1361.110 825.670 ;
        RECT 1359.930 646.090 1361.110 647.270 ;
        RECT 1359.930 644.490 1361.110 645.670 ;
        RECT 1359.930 466.090 1361.110 467.270 ;
        RECT 1359.930 464.490 1361.110 465.670 ;
        RECT 1359.930 286.090 1361.110 287.270 ;
        RECT 1359.930 284.490 1361.110 285.670 ;
        RECT 1359.930 106.090 1361.110 107.270 ;
        RECT 1359.930 104.490 1361.110 105.670 ;
        RECT 1359.930 -7.610 1361.110 -6.430 ;
        RECT 1359.930 -9.210 1361.110 -8.030 ;
        RECT 1539.930 3527.710 1541.110 3528.890 ;
        RECT 1539.930 3526.110 1541.110 3527.290 ;
        RECT 1539.930 3346.090 1541.110 3347.270 ;
        RECT 1539.930 3344.490 1541.110 3345.670 ;
        RECT 1539.930 3166.090 1541.110 3167.270 ;
        RECT 1539.930 3164.490 1541.110 3165.670 ;
        RECT 1539.930 2986.090 1541.110 2987.270 ;
        RECT 1539.930 2984.490 1541.110 2985.670 ;
        RECT 1539.930 2806.090 1541.110 2807.270 ;
        RECT 1539.930 2804.490 1541.110 2805.670 ;
        RECT 1539.930 2626.090 1541.110 2627.270 ;
        RECT 1539.930 2624.490 1541.110 2625.670 ;
        RECT 1539.930 2446.090 1541.110 2447.270 ;
        RECT 1539.930 2444.490 1541.110 2445.670 ;
        RECT 1539.930 2266.090 1541.110 2267.270 ;
        RECT 1539.930 2264.490 1541.110 2265.670 ;
        RECT 1539.930 2086.090 1541.110 2087.270 ;
        RECT 1539.930 2084.490 1541.110 2085.670 ;
        RECT 1539.930 1906.090 1541.110 1907.270 ;
        RECT 1539.930 1904.490 1541.110 1905.670 ;
        RECT 1539.930 1726.090 1541.110 1727.270 ;
        RECT 1539.930 1724.490 1541.110 1725.670 ;
        RECT 1539.930 1546.090 1541.110 1547.270 ;
        RECT 1539.930 1544.490 1541.110 1545.670 ;
        RECT 1539.930 1366.090 1541.110 1367.270 ;
        RECT 1539.930 1364.490 1541.110 1365.670 ;
        RECT 1539.930 1186.090 1541.110 1187.270 ;
        RECT 1539.930 1184.490 1541.110 1185.670 ;
        RECT 1539.930 1006.090 1541.110 1007.270 ;
        RECT 1539.930 1004.490 1541.110 1005.670 ;
        RECT 1539.930 826.090 1541.110 827.270 ;
        RECT 1539.930 824.490 1541.110 825.670 ;
        RECT 1539.930 646.090 1541.110 647.270 ;
        RECT 1539.930 644.490 1541.110 645.670 ;
        RECT 1539.930 466.090 1541.110 467.270 ;
        RECT 1539.930 464.490 1541.110 465.670 ;
        RECT 1539.930 286.090 1541.110 287.270 ;
        RECT 1539.930 284.490 1541.110 285.670 ;
        RECT 1539.930 106.090 1541.110 107.270 ;
        RECT 1539.930 104.490 1541.110 105.670 ;
        RECT 1539.930 -7.610 1541.110 -6.430 ;
        RECT 1539.930 -9.210 1541.110 -8.030 ;
        RECT 1719.930 3527.710 1721.110 3528.890 ;
        RECT 1719.930 3526.110 1721.110 3527.290 ;
        RECT 1719.930 3346.090 1721.110 3347.270 ;
        RECT 1719.930 3344.490 1721.110 3345.670 ;
        RECT 1719.930 3166.090 1721.110 3167.270 ;
        RECT 1719.930 3164.490 1721.110 3165.670 ;
        RECT 1719.930 2986.090 1721.110 2987.270 ;
        RECT 1719.930 2984.490 1721.110 2985.670 ;
        RECT 1719.930 2806.090 1721.110 2807.270 ;
        RECT 1719.930 2804.490 1721.110 2805.670 ;
        RECT 1719.930 2626.090 1721.110 2627.270 ;
        RECT 1719.930 2624.490 1721.110 2625.670 ;
        RECT 1719.930 2446.090 1721.110 2447.270 ;
        RECT 1719.930 2444.490 1721.110 2445.670 ;
        RECT 1719.930 2266.090 1721.110 2267.270 ;
        RECT 1719.930 2264.490 1721.110 2265.670 ;
        RECT 1719.930 2086.090 1721.110 2087.270 ;
        RECT 1719.930 2084.490 1721.110 2085.670 ;
        RECT 1719.930 1906.090 1721.110 1907.270 ;
        RECT 1719.930 1904.490 1721.110 1905.670 ;
        RECT 1719.930 1726.090 1721.110 1727.270 ;
        RECT 1719.930 1724.490 1721.110 1725.670 ;
        RECT 1719.930 1546.090 1721.110 1547.270 ;
        RECT 1719.930 1544.490 1721.110 1545.670 ;
        RECT 1719.930 1366.090 1721.110 1367.270 ;
        RECT 1719.930 1364.490 1721.110 1365.670 ;
        RECT 1719.930 1186.090 1721.110 1187.270 ;
        RECT 1719.930 1184.490 1721.110 1185.670 ;
        RECT 1719.930 1006.090 1721.110 1007.270 ;
        RECT 1719.930 1004.490 1721.110 1005.670 ;
        RECT 1719.930 826.090 1721.110 827.270 ;
        RECT 1719.930 824.490 1721.110 825.670 ;
        RECT 1719.930 646.090 1721.110 647.270 ;
        RECT 1719.930 644.490 1721.110 645.670 ;
        RECT 1719.930 466.090 1721.110 467.270 ;
        RECT 1719.930 464.490 1721.110 465.670 ;
        RECT 1719.930 286.090 1721.110 287.270 ;
        RECT 1719.930 284.490 1721.110 285.670 ;
        RECT 1719.930 106.090 1721.110 107.270 ;
        RECT 1719.930 104.490 1721.110 105.670 ;
        RECT 1719.930 -7.610 1721.110 -6.430 ;
        RECT 1719.930 -9.210 1721.110 -8.030 ;
        RECT 1899.930 3527.710 1901.110 3528.890 ;
        RECT 1899.930 3526.110 1901.110 3527.290 ;
        RECT 1899.930 3346.090 1901.110 3347.270 ;
        RECT 1899.930 3344.490 1901.110 3345.670 ;
        RECT 1899.930 3166.090 1901.110 3167.270 ;
        RECT 1899.930 3164.490 1901.110 3165.670 ;
        RECT 1899.930 2986.090 1901.110 2987.270 ;
        RECT 1899.930 2984.490 1901.110 2985.670 ;
        RECT 1899.930 2806.090 1901.110 2807.270 ;
        RECT 1899.930 2804.490 1901.110 2805.670 ;
        RECT 1899.930 2626.090 1901.110 2627.270 ;
        RECT 1899.930 2624.490 1901.110 2625.670 ;
        RECT 1899.930 2446.090 1901.110 2447.270 ;
        RECT 1899.930 2444.490 1901.110 2445.670 ;
        RECT 1899.930 2266.090 1901.110 2267.270 ;
        RECT 1899.930 2264.490 1901.110 2265.670 ;
        RECT 1899.930 2086.090 1901.110 2087.270 ;
        RECT 1899.930 2084.490 1901.110 2085.670 ;
        RECT 1899.930 1906.090 1901.110 1907.270 ;
        RECT 1899.930 1904.490 1901.110 1905.670 ;
        RECT 1899.930 1726.090 1901.110 1727.270 ;
        RECT 1899.930 1724.490 1901.110 1725.670 ;
        RECT 1899.930 1546.090 1901.110 1547.270 ;
        RECT 1899.930 1544.490 1901.110 1545.670 ;
        RECT 1899.930 1366.090 1901.110 1367.270 ;
        RECT 1899.930 1364.490 1901.110 1365.670 ;
        RECT 1899.930 1186.090 1901.110 1187.270 ;
        RECT 1899.930 1184.490 1901.110 1185.670 ;
        RECT 1899.930 1006.090 1901.110 1007.270 ;
        RECT 1899.930 1004.490 1901.110 1005.670 ;
        RECT 1899.930 826.090 1901.110 827.270 ;
        RECT 1899.930 824.490 1901.110 825.670 ;
        RECT 1899.930 646.090 1901.110 647.270 ;
        RECT 1899.930 644.490 1901.110 645.670 ;
        RECT 1899.930 466.090 1901.110 467.270 ;
        RECT 1899.930 464.490 1901.110 465.670 ;
        RECT 1899.930 286.090 1901.110 287.270 ;
        RECT 1899.930 284.490 1901.110 285.670 ;
        RECT 1899.930 106.090 1901.110 107.270 ;
        RECT 1899.930 104.490 1901.110 105.670 ;
        RECT 1899.930 -7.610 1901.110 -6.430 ;
        RECT 1899.930 -9.210 1901.110 -8.030 ;
        RECT 2079.930 3527.710 2081.110 3528.890 ;
        RECT 2079.930 3526.110 2081.110 3527.290 ;
        RECT 2079.930 3346.090 2081.110 3347.270 ;
        RECT 2079.930 3344.490 2081.110 3345.670 ;
        RECT 2079.930 3166.090 2081.110 3167.270 ;
        RECT 2079.930 3164.490 2081.110 3165.670 ;
        RECT 2079.930 2986.090 2081.110 2987.270 ;
        RECT 2079.930 2984.490 2081.110 2985.670 ;
        RECT 2079.930 2806.090 2081.110 2807.270 ;
        RECT 2079.930 2804.490 2081.110 2805.670 ;
        RECT 2079.930 2626.090 2081.110 2627.270 ;
        RECT 2079.930 2624.490 2081.110 2625.670 ;
        RECT 2079.930 2446.090 2081.110 2447.270 ;
        RECT 2079.930 2444.490 2081.110 2445.670 ;
        RECT 2079.930 2266.090 2081.110 2267.270 ;
        RECT 2079.930 2264.490 2081.110 2265.670 ;
        RECT 2079.930 2086.090 2081.110 2087.270 ;
        RECT 2079.930 2084.490 2081.110 2085.670 ;
        RECT 2079.930 1906.090 2081.110 1907.270 ;
        RECT 2079.930 1904.490 2081.110 1905.670 ;
        RECT 2079.930 1726.090 2081.110 1727.270 ;
        RECT 2079.930 1724.490 2081.110 1725.670 ;
        RECT 2079.930 1546.090 2081.110 1547.270 ;
        RECT 2079.930 1544.490 2081.110 1545.670 ;
        RECT 2079.930 1366.090 2081.110 1367.270 ;
        RECT 2079.930 1364.490 2081.110 1365.670 ;
        RECT 2079.930 1186.090 2081.110 1187.270 ;
        RECT 2079.930 1184.490 2081.110 1185.670 ;
        RECT 2079.930 1006.090 2081.110 1007.270 ;
        RECT 2079.930 1004.490 2081.110 1005.670 ;
        RECT 2079.930 826.090 2081.110 827.270 ;
        RECT 2079.930 824.490 2081.110 825.670 ;
        RECT 2079.930 646.090 2081.110 647.270 ;
        RECT 2079.930 644.490 2081.110 645.670 ;
        RECT 2079.930 466.090 2081.110 467.270 ;
        RECT 2079.930 464.490 2081.110 465.670 ;
        RECT 2079.930 286.090 2081.110 287.270 ;
        RECT 2079.930 284.490 2081.110 285.670 ;
        RECT 2079.930 106.090 2081.110 107.270 ;
        RECT 2079.930 104.490 2081.110 105.670 ;
        RECT 2079.930 -7.610 2081.110 -6.430 ;
        RECT 2079.930 -9.210 2081.110 -8.030 ;
        RECT 2259.930 3527.710 2261.110 3528.890 ;
        RECT 2259.930 3526.110 2261.110 3527.290 ;
        RECT 2259.930 3346.090 2261.110 3347.270 ;
        RECT 2259.930 3344.490 2261.110 3345.670 ;
        RECT 2259.930 3166.090 2261.110 3167.270 ;
        RECT 2259.930 3164.490 2261.110 3165.670 ;
        RECT 2259.930 2986.090 2261.110 2987.270 ;
        RECT 2259.930 2984.490 2261.110 2985.670 ;
        RECT 2259.930 2806.090 2261.110 2807.270 ;
        RECT 2259.930 2804.490 2261.110 2805.670 ;
        RECT 2259.930 2626.090 2261.110 2627.270 ;
        RECT 2259.930 2624.490 2261.110 2625.670 ;
        RECT 2259.930 2446.090 2261.110 2447.270 ;
        RECT 2259.930 2444.490 2261.110 2445.670 ;
        RECT 2259.930 2266.090 2261.110 2267.270 ;
        RECT 2259.930 2264.490 2261.110 2265.670 ;
        RECT 2259.930 2086.090 2261.110 2087.270 ;
        RECT 2259.930 2084.490 2261.110 2085.670 ;
        RECT 2259.930 1906.090 2261.110 1907.270 ;
        RECT 2259.930 1904.490 2261.110 1905.670 ;
        RECT 2259.930 1726.090 2261.110 1727.270 ;
        RECT 2259.930 1724.490 2261.110 1725.670 ;
        RECT 2259.930 1546.090 2261.110 1547.270 ;
        RECT 2259.930 1544.490 2261.110 1545.670 ;
        RECT 2259.930 1366.090 2261.110 1367.270 ;
        RECT 2259.930 1364.490 2261.110 1365.670 ;
        RECT 2259.930 1186.090 2261.110 1187.270 ;
        RECT 2259.930 1184.490 2261.110 1185.670 ;
        RECT 2259.930 1006.090 2261.110 1007.270 ;
        RECT 2259.930 1004.490 2261.110 1005.670 ;
        RECT 2259.930 826.090 2261.110 827.270 ;
        RECT 2259.930 824.490 2261.110 825.670 ;
        RECT 2259.930 646.090 2261.110 647.270 ;
        RECT 2259.930 644.490 2261.110 645.670 ;
        RECT 2259.930 466.090 2261.110 467.270 ;
        RECT 2259.930 464.490 2261.110 465.670 ;
        RECT 2259.930 286.090 2261.110 287.270 ;
        RECT 2259.930 284.490 2261.110 285.670 ;
        RECT 2259.930 106.090 2261.110 107.270 ;
        RECT 2259.930 104.490 2261.110 105.670 ;
        RECT 2259.930 -7.610 2261.110 -6.430 ;
        RECT 2259.930 -9.210 2261.110 -8.030 ;
        RECT 2439.930 3527.710 2441.110 3528.890 ;
        RECT 2439.930 3526.110 2441.110 3527.290 ;
        RECT 2439.930 3346.090 2441.110 3347.270 ;
        RECT 2439.930 3344.490 2441.110 3345.670 ;
        RECT 2439.930 3166.090 2441.110 3167.270 ;
        RECT 2439.930 3164.490 2441.110 3165.670 ;
        RECT 2439.930 2986.090 2441.110 2987.270 ;
        RECT 2439.930 2984.490 2441.110 2985.670 ;
        RECT 2439.930 2806.090 2441.110 2807.270 ;
        RECT 2439.930 2804.490 2441.110 2805.670 ;
        RECT 2439.930 2626.090 2441.110 2627.270 ;
        RECT 2439.930 2624.490 2441.110 2625.670 ;
        RECT 2439.930 2446.090 2441.110 2447.270 ;
        RECT 2439.930 2444.490 2441.110 2445.670 ;
        RECT 2439.930 2266.090 2441.110 2267.270 ;
        RECT 2439.930 2264.490 2441.110 2265.670 ;
        RECT 2439.930 2086.090 2441.110 2087.270 ;
        RECT 2439.930 2084.490 2441.110 2085.670 ;
        RECT 2439.930 1906.090 2441.110 1907.270 ;
        RECT 2439.930 1904.490 2441.110 1905.670 ;
        RECT 2439.930 1726.090 2441.110 1727.270 ;
        RECT 2439.930 1724.490 2441.110 1725.670 ;
        RECT 2439.930 1546.090 2441.110 1547.270 ;
        RECT 2439.930 1544.490 2441.110 1545.670 ;
        RECT 2439.930 1366.090 2441.110 1367.270 ;
        RECT 2439.930 1364.490 2441.110 1365.670 ;
        RECT 2439.930 1186.090 2441.110 1187.270 ;
        RECT 2439.930 1184.490 2441.110 1185.670 ;
        RECT 2439.930 1006.090 2441.110 1007.270 ;
        RECT 2439.930 1004.490 2441.110 1005.670 ;
        RECT 2439.930 826.090 2441.110 827.270 ;
        RECT 2439.930 824.490 2441.110 825.670 ;
        RECT 2439.930 646.090 2441.110 647.270 ;
        RECT 2439.930 644.490 2441.110 645.670 ;
        RECT 2439.930 466.090 2441.110 467.270 ;
        RECT 2439.930 464.490 2441.110 465.670 ;
        RECT 2439.930 286.090 2441.110 287.270 ;
        RECT 2439.930 284.490 2441.110 285.670 ;
        RECT 2439.930 106.090 2441.110 107.270 ;
        RECT 2439.930 104.490 2441.110 105.670 ;
        RECT 2439.930 -7.610 2441.110 -6.430 ;
        RECT 2439.930 -9.210 2441.110 -8.030 ;
        RECT 2619.930 3527.710 2621.110 3528.890 ;
        RECT 2619.930 3526.110 2621.110 3527.290 ;
        RECT 2619.930 3346.090 2621.110 3347.270 ;
        RECT 2619.930 3344.490 2621.110 3345.670 ;
        RECT 2619.930 3166.090 2621.110 3167.270 ;
        RECT 2619.930 3164.490 2621.110 3165.670 ;
        RECT 2619.930 2986.090 2621.110 2987.270 ;
        RECT 2619.930 2984.490 2621.110 2985.670 ;
        RECT 2619.930 2806.090 2621.110 2807.270 ;
        RECT 2619.930 2804.490 2621.110 2805.670 ;
        RECT 2619.930 2626.090 2621.110 2627.270 ;
        RECT 2619.930 2624.490 2621.110 2625.670 ;
        RECT 2619.930 2446.090 2621.110 2447.270 ;
        RECT 2619.930 2444.490 2621.110 2445.670 ;
        RECT 2619.930 2266.090 2621.110 2267.270 ;
        RECT 2619.930 2264.490 2621.110 2265.670 ;
        RECT 2619.930 2086.090 2621.110 2087.270 ;
        RECT 2619.930 2084.490 2621.110 2085.670 ;
        RECT 2619.930 1906.090 2621.110 1907.270 ;
        RECT 2619.930 1904.490 2621.110 1905.670 ;
        RECT 2619.930 1726.090 2621.110 1727.270 ;
        RECT 2619.930 1724.490 2621.110 1725.670 ;
        RECT 2619.930 1546.090 2621.110 1547.270 ;
        RECT 2619.930 1544.490 2621.110 1545.670 ;
        RECT 2619.930 1366.090 2621.110 1367.270 ;
        RECT 2619.930 1364.490 2621.110 1365.670 ;
        RECT 2619.930 1186.090 2621.110 1187.270 ;
        RECT 2619.930 1184.490 2621.110 1185.670 ;
        RECT 2619.930 1006.090 2621.110 1007.270 ;
        RECT 2619.930 1004.490 2621.110 1005.670 ;
        RECT 2619.930 826.090 2621.110 827.270 ;
        RECT 2619.930 824.490 2621.110 825.670 ;
        RECT 2619.930 646.090 2621.110 647.270 ;
        RECT 2619.930 644.490 2621.110 645.670 ;
        RECT 2619.930 466.090 2621.110 467.270 ;
        RECT 2619.930 464.490 2621.110 465.670 ;
        RECT 2619.930 286.090 2621.110 287.270 ;
        RECT 2619.930 284.490 2621.110 285.670 ;
        RECT 2619.930 106.090 2621.110 107.270 ;
        RECT 2619.930 104.490 2621.110 105.670 ;
        RECT 2619.930 -7.610 2621.110 -6.430 ;
        RECT 2619.930 -9.210 2621.110 -8.030 ;
        RECT 2799.930 3527.710 2801.110 3528.890 ;
        RECT 2799.930 3526.110 2801.110 3527.290 ;
        RECT 2799.930 3346.090 2801.110 3347.270 ;
        RECT 2799.930 3344.490 2801.110 3345.670 ;
        RECT 2799.930 3166.090 2801.110 3167.270 ;
        RECT 2799.930 3164.490 2801.110 3165.670 ;
        RECT 2799.930 2986.090 2801.110 2987.270 ;
        RECT 2799.930 2984.490 2801.110 2985.670 ;
        RECT 2799.930 2806.090 2801.110 2807.270 ;
        RECT 2799.930 2804.490 2801.110 2805.670 ;
        RECT 2799.930 2626.090 2801.110 2627.270 ;
        RECT 2799.930 2624.490 2801.110 2625.670 ;
        RECT 2799.930 2446.090 2801.110 2447.270 ;
        RECT 2799.930 2444.490 2801.110 2445.670 ;
        RECT 2799.930 2266.090 2801.110 2267.270 ;
        RECT 2799.930 2264.490 2801.110 2265.670 ;
        RECT 2799.930 2086.090 2801.110 2087.270 ;
        RECT 2799.930 2084.490 2801.110 2085.670 ;
        RECT 2799.930 1906.090 2801.110 1907.270 ;
        RECT 2799.930 1904.490 2801.110 1905.670 ;
        RECT 2799.930 1726.090 2801.110 1727.270 ;
        RECT 2799.930 1724.490 2801.110 1725.670 ;
        RECT 2799.930 1546.090 2801.110 1547.270 ;
        RECT 2799.930 1544.490 2801.110 1545.670 ;
        RECT 2799.930 1366.090 2801.110 1367.270 ;
        RECT 2799.930 1364.490 2801.110 1365.670 ;
        RECT 2799.930 1186.090 2801.110 1187.270 ;
        RECT 2799.930 1184.490 2801.110 1185.670 ;
        RECT 2799.930 1006.090 2801.110 1007.270 ;
        RECT 2799.930 1004.490 2801.110 1005.670 ;
        RECT 2799.930 826.090 2801.110 827.270 ;
        RECT 2799.930 824.490 2801.110 825.670 ;
        RECT 2799.930 646.090 2801.110 647.270 ;
        RECT 2799.930 644.490 2801.110 645.670 ;
        RECT 2799.930 466.090 2801.110 467.270 ;
        RECT 2799.930 464.490 2801.110 465.670 ;
        RECT 2799.930 286.090 2801.110 287.270 ;
        RECT 2799.930 284.490 2801.110 285.670 ;
        RECT 2799.930 106.090 2801.110 107.270 ;
        RECT 2799.930 104.490 2801.110 105.670 ;
        RECT 2799.930 -7.610 2801.110 -6.430 ;
        RECT 2799.930 -9.210 2801.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3346.090 2933.390 3347.270 ;
        RECT 2932.210 3344.490 2933.390 3345.670 ;
        RECT 2932.210 3166.090 2933.390 3167.270 ;
        RECT 2932.210 3164.490 2933.390 3165.670 ;
        RECT 2932.210 2986.090 2933.390 2987.270 ;
        RECT 2932.210 2984.490 2933.390 2985.670 ;
        RECT 2932.210 2806.090 2933.390 2807.270 ;
        RECT 2932.210 2804.490 2933.390 2805.670 ;
        RECT 2932.210 2626.090 2933.390 2627.270 ;
        RECT 2932.210 2624.490 2933.390 2625.670 ;
        RECT 2932.210 2446.090 2933.390 2447.270 ;
        RECT 2932.210 2444.490 2933.390 2445.670 ;
        RECT 2932.210 2266.090 2933.390 2267.270 ;
        RECT 2932.210 2264.490 2933.390 2265.670 ;
        RECT 2932.210 2086.090 2933.390 2087.270 ;
        RECT 2932.210 2084.490 2933.390 2085.670 ;
        RECT 2932.210 1906.090 2933.390 1907.270 ;
        RECT 2932.210 1904.490 2933.390 1905.670 ;
        RECT 2932.210 1726.090 2933.390 1727.270 ;
        RECT 2932.210 1724.490 2933.390 1725.670 ;
        RECT 2932.210 1546.090 2933.390 1547.270 ;
        RECT 2932.210 1544.490 2933.390 1545.670 ;
        RECT 2932.210 1366.090 2933.390 1367.270 ;
        RECT 2932.210 1364.490 2933.390 1365.670 ;
        RECT 2932.210 1186.090 2933.390 1187.270 ;
        RECT 2932.210 1184.490 2933.390 1185.670 ;
        RECT 2932.210 1006.090 2933.390 1007.270 ;
        RECT 2932.210 1004.490 2933.390 1005.670 ;
        RECT 2932.210 826.090 2933.390 827.270 ;
        RECT 2932.210 824.490 2933.390 825.670 ;
        RECT 2932.210 646.090 2933.390 647.270 ;
        RECT 2932.210 644.490 2933.390 645.670 ;
        RECT 2932.210 466.090 2933.390 467.270 ;
        RECT 2932.210 464.490 2933.390 465.670 ;
        RECT 2932.210 286.090 2933.390 287.270 ;
        RECT 2932.210 284.490 2933.390 285.670 ;
        RECT 2932.210 106.090 2933.390 107.270 ;
        RECT 2932.210 104.490 2933.390 105.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 99.020 3529.000 102.020 3529.010 ;
        RECT 279.020 3529.000 282.020 3529.010 ;
        RECT 459.020 3529.000 462.020 3529.010 ;
        RECT 639.020 3529.000 642.020 3529.010 ;
        RECT 819.020 3529.000 822.020 3529.010 ;
        RECT 999.020 3529.000 1002.020 3529.010 ;
        RECT 1179.020 3529.000 1182.020 3529.010 ;
        RECT 1359.020 3529.000 1362.020 3529.010 ;
        RECT 1539.020 3529.000 1542.020 3529.010 ;
        RECT 1719.020 3529.000 1722.020 3529.010 ;
        RECT 1899.020 3529.000 1902.020 3529.010 ;
        RECT 2079.020 3529.000 2082.020 3529.010 ;
        RECT 2259.020 3529.000 2262.020 3529.010 ;
        RECT 2439.020 3529.000 2442.020 3529.010 ;
        RECT 2619.020 3529.000 2622.020 3529.010 ;
        RECT 2799.020 3529.000 2802.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 99.020 3525.990 102.020 3526.000 ;
        RECT 279.020 3525.990 282.020 3526.000 ;
        RECT 459.020 3525.990 462.020 3526.000 ;
        RECT 639.020 3525.990 642.020 3526.000 ;
        RECT 819.020 3525.990 822.020 3526.000 ;
        RECT 999.020 3525.990 1002.020 3526.000 ;
        RECT 1179.020 3525.990 1182.020 3526.000 ;
        RECT 1359.020 3525.990 1362.020 3526.000 ;
        RECT 1539.020 3525.990 1542.020 3526.000 ;
        RECT 1719.020 3525.990 1722.020 3526.000 ;
        RECT 1899.020 3525.990 1902.020 3526.000 ;
        RECT 2079.020 3525.990 2082.020 3526.000 ;
        RECT 2259.020 3525.990 2262.020 3526.000 ;
        RECT 2439.020 3525.990 2442.020 3526.000 ;
        RECT 2619.020 3525.990 2622.020 3526.000 ;
        RECT 2799.020 3525.990 2802.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3347.380 -11.680 3347.390 ;
        RECT 99.020 3347.380 102.020 3347.390 ;
        RECT 279.020 3347.380 282.020 3347.390 ;
        RECT 459.020 3347.380 462.020 3347.390 ;
        RECT 639.020 3347.380 642.020 3347.390 ;
        RECT 819.020 3347.380 822.020 3347.390 ;
        RECT 999.020 3347.380 1002.020 3347.390 ;
        RECT 1179.020 3347.380 1182.020 3347.390 ;
        RECT 1359.020 3347.380 1362.020 3347.390 ;
        RECT 1539.020 3347.380 1542.020 3347.390 ;
        RECT 1719.020 3347.380 1722.020 3347.390 ;
        RECT 1899.020 3347.380 1902.020 3347.390 ;
        RECT 2079.020 3347.380 2082.020 3347.390 ;
        RECT 2259.020 3347.380 2262.020 3347.390 ;
        RECT 2439.020 3347.380 2442.020 3347.390 ;
        RECT 2619.020 3347.380 2622.020 3347.390 ;
        RECT 2799.020 3347.380 2802.020 3347.390 ;
        RECT 2931.300 3347.380 2934.300 3347.390 ;
        RECT -14.680 3344.380 2934.300 3347.380 ;
        RECT -14.680 3344.370 -11.680 3344.380 ;
        RECT 99.020 3344.370 102.020 3344.380 ;
        RECT 279.020 3344.370 282.020 3344.380 ;
        RECT 459.020 3344.370 462.020 3344.380 ;
        RECT 639.020 3344.370 642.020 3344.380 ;
        RECT 819.020 3344.370 822.020 3344.380 ;
        RECT 999.020 3344.370 1002.020 3344.380 ;
        RECT 1179.020 3344.370 1182.020 3344.380 ;
        RECT 1359.020 3344.370 1362.020 3344.380 ;
        RECT 1539.020 3344.370 1542.020 3344.380 ;
        RECT 1719.020 3344.370 1722.020 3344.380 ;
        RECT 1899.020 3344.370 1902.020 3344.380 ;
        RECT 2079.020 3344.370 2082.020 3344.380 ;
        RECT 2259.020 3344.370 2262.020 3344.380 ;
        RECT 2439.020 3344.370 2442.020 3344.380 ;
        RECT 2619.020 3344.370 2622.020 3344.380 ;
        RECT 2799.020 3344.370 2802.020 3344.380 ;
        RECT 2931.300 3344.370 2934.300 3344.380 ;
        RECT -14.680 3167.380 -11.680 3167.390 ;
        RECT 99.020 3167.380 102.020 3167.390 ;
        RECT 279.020 3167.380 282.020 3167.390 ;
        RECT 459.020 3167.380 462.020 3167.390 ;
        RECT 639.020 3167.380 642.020 3167.390 ;
        RECT 819.020 3167.380 822.020 3167.390 ;
        RECT 999.020 3167.380 1002.020 3167.390 ;
        RECT 1179.020 3167.380 1182.020 3167.390 ;
        RECT 1359.020 3167.380 1362.020 3167.390 ;
        RECT 1539.020 3167.380 1542.020 3167.390 ;
        RECT 1719.020 3167.380 1722.020 3167.390 ;
        RECT 1899.020 3167.380 1902.020 3167.390 ;
        RECT 2079.020 3167.380 2082.020 3167.390 ;
        RECT 2259.020 3167.380 2262.020 3167.390 ;
        RECT 2439.020 3167.380 2442.020 3167.390 ;
        RECT 2619.020 3167.380 2622.020 3167.390 ;
        RECT 2799.020 3167.380 2802.020 3167.390 ;
        RECT 2931.300 3167.380 2934.300 3167.390 ;
        RECT -14.680 3164.380 2934.300 3167.380 ;
        RECT -14.680 3164.370 -11.680 3164.380 ;
        RECT 99.020 3164.370 102.020 3164.380 ;
        RECT 279.020 3164.370 282.020 3164.380 ;
        RECT 459.020 3164.370 462.020 3164.380 ;
        RECT 639.020 3164.370 642.020 3164.380 ;
        RECT 819.020 3164.370 822.020 3164.380 ;
        RECT 999.020 3164.370 1002.020 3164.380 ;
        RECT 1179.020 3164.370 1182.020 3164.380 ;
        RECT 1359.020 3164.370 1362.020 3164.380 ;
        RECT 1539.020 3164.370 1542.020 3164.380 ;
        RECT 1719.020 3164.370 1722.020 3164.380 ;
        RECT 1899.020 3164.370 1902.020 3164.380 ;
        RECT 2079.020 3164.370 2082.020 3164.380 ;
        RECT 2259.020 3164.370 2262.020 3164.380 ;
        RECT 2439.020 3164.370 2442.020 3164.380 ;
        RECT 2619.020 3164.370 2622.020 3164.380 ;
        RECT 2799.020 3164.370 2802.020 3164.380 ;
        RECT 2931.300 3164.370 2934.300 3164.380 ;
        RECT -14.680 2987.380 -11.680 2987.390 ;
        RECT 99.020 2987.380 102.020 2987.390 ;
        RECT 279.020 2987.380 282.020 2987.390 ;
        RECT 459.020 2987.380 462.020 2987.390 ;
        RECT 639.020 2987.380 642.020 2987.390 ;
        RECT 819.020 2987.380 822.020 2987.390 ;
        RECT 999.020 2987.380 1002.020 2987.390 ;
        RECT 1179.020 2987.380 1182.020 2987.390 ;
        RECT 1359.020 2987.380 1362.020 2987.390 ;
        RECT 1539.020 2987.380 1542.020 2987.390 ;
        RECT 1719.020 2987.380 1722.020 2987.390 ;
        RECT 1899.020 2987.380 1902.020 2987.390 ;
        RECT 2079.020 2987.380 2082.020 2987.390 ;
        RECT 2259.020 2987.380 2262.020 2987.390 ;
        RECT 2439.020 2987.380 2442.020 2987.390 ;
        RECT 2619.020 2987.380 2622.020 2987.390 ;
        RECT 2799.020 2987.380 2802.020 2987.390 ;
        RECT 2931.300 2987.380 2934.300 2987.390 ;
        RECT -14.680 2984.380 2934.300 2987.380 ;
        RECT -14.680 2984.370 -11.680 2984.380 ;
        RECT 99.020 2984.370 102.020 2984.380 ;
        RECT 279.020 2984.370 282.020 2984.380 ;
        RECT 459.020 2984.370 462.020 2984.380 ;
        RECT 639.020 2984.370 642.020 2984.380 ;
        RECT 819.020 2984.370 822.020 2984.380 ;
        RECT 999.020 2984.370 1002.020 2984.380 ;
        RECT 1179.020 2984.370 1182.020 2984.380 ;
        RECT 1359.020 2984.370 1362.020 2984.380 ;
        RECT 1539.020 2984.370 1542.020 2984.380 ;
        RECT 1719.020 2984.370 1722.020 2984.380 ;
        RECT 1899.020 2984.370 1902.020 2984.380 ;
        RECT 2079.020 2984.370 2082.020 2984.380 ;
        RECT 2259.020 2984.370 2262.020 2984.380 ;
        RECT 2439.020 2984.370 2442.020 2984.380 ;
        RECT 2619.020 2984.370 2622.020 2984.380 ;
        RECT 2799.020 2984.370 2802.020 2984.380 ;
        RECT 2931.300 2984.370 2934.300 2984.380 ;
        RECT -14.680 2807.380 -11.680 2807.390 ;
        RECT 99.020 2807.380 102.020 2807.390 ;
        RECT 279.020 2807.380 282.020 2807.390 ;
        RECT 459.020 2807.380 462.020 2807.390 ;
        RECT 639.020 2807.380 642.020 2807.390 ;
        RECT 819.020 2807.380 822.020 2807.390 ;
        RECT 999.020 2807.380 1002.020 2807.390 ;
        RECT 1179.020 2807.380 1182.020 2807.390 ;
        RECT 1359.020 2807.380 1362.020 2807.390 ;
        RECT 1539.020 2807.380 1542.020 2807.390 ;
        RECT 1719.020 2807.380 1722.020 2807.390 ;
        RECT 1899.020 2807.380 1902.020 2807.390 ;
        RECT 2079.020 2807.380 2082.020 2807.390 ;
        RECT 2259.020 2807.380 2262.020 2807.390 ;
        RECT 2439.020 2807.380 2442.020 2807.390 ;
        RECT 2619.020 2807.380 2622.020 2807.390 ;
        RECT 2799.020 2807.380 2802.020 2807.390 ;
        RECT 2931.300 2807.380 2934.300 2807.390 ;
        RECT -14.680 2804.380 2934.300 2807.380 ;
        RECT -14.680 2804.370 -11.680 2804.380 ;
        RECT 99.020 2804.370 102.020 2804.380 ;
        RECT 279.020 2804.370 282.020 2804.380 ;
        RECT 459.020 2804.370 462.020 2804.380 ;
        RECT 639.020 2804.370 642.020 2804.380 ;
        RECT 819.020 2804.370 822.020 2804.380 ;
        RECT 999.020 2804.370 1002.020 2804.380 ;
        RECT 1179.020 2804.370 1182.020 2804.380 ;
        RECT 1359.020 2804.370 1362.020 2804.380 ;
        RECT 1539.020 2804.370 1542.020 2804.380 ;
        RECT 1719.020 2804.370 1722.020 2804.380 ;
        RECT 1899.020 2804.370 1902.020 2804.380 ;
        RECT 2079.020 2804.370 2082.020 2804.380 ;
        RECT 2259.020 2804.370 2262.020 2804.380 ;
        RECT 2439.020 2804.370 2442.020 2804.380 ;
        RECT 2619.020 2804.370 2622.020 2804.380 ;
        RECT 2799.020 2804.370 2802.020 2804.380 ;
        RECT 2931.300 2804.370 2934.300 2804.380 ;
        RECT -14.680 2627.380 -11.680 2627.390 ;
        RECT 99.020 2627.380 102.020 2627.390 ;
        RECT 279.020 2627.380 282.020 2627.390 ;
        RECT 459.020 2627.380 462.020 2627.390 ;
        RECT 639.020 2627.380 642.020 2627.390 ;
        RECT 819.020 2627.380 822.020 2627.390 ;
        RECT 999.020 2627.380 1002.020 2627.390 ;
        RECT 1179.020 2627.380 1182.020 2627.390 ;
        RECT 1359.020 2627.380 1362.020 2627.390 ;
        RECT 1539.020 2627.380 1542.020 2627.390 ;
        RECT 1719.020 2627.380 1722.020 2627.390 ;
        RECT 1899.020 2627.380 1902.020 2627.390 ;
        RECT 2079.020 2627.380 2082.020 2627.390 ;
        RECT 2259.020 2627.380 2262.020 2627.390 ;
        RECT 2439.020 2627.380 2442.020 2627.390 ;
        RECT 2619.020 2627.380 2622.020 2627.390 ;
        RECT 2799.020 2627.380 2802.020 2627.390 ;
        RECT 2931.300 2627.380 2934.300 2627.390 ;
        RECT -14.680 2624.380 2934.300 2627.380 ;
        RECT -14.680 2624.370 -11.680 2624.380 ;
        RECT 99.020 2624.370 102.020 2624.380 ;
        RECT 279.020 2624.370 282.020 2624.380 ;
        RECT 459.020 2624.370 462.020 2624.380 ;
        RECT 639.020 2624.370 642.020 2624.380 ;
        RECT 819.020 2624.370 822.020 2624.380 ;
        RECT 999.020 2624.370 1002.020 2624.380 ;
        RECT 1179.020 2624.370 1182.020 2624.380 ;
        RECT 1359.020 2624.370 1362.020 2624.380 ;
        RECT 1539.020 2624.370 1542.020 2624.380 ;
        RECT 1719.020 2624.370 1722.020 2624.380 ;
        RECT 1899.020 2624.370 1902.020 2624.380 ;
        RECT 2079.020 2624.370 2082.020 2624.380 ;
        RECT 2259.020 2624.370 2262.020 2624.380 ;
        RECT 2439.020 2624.370 2442.020 2624.380 ;
        RECT 2619.020 2624.370 2622.020 2624.380 ;
        RECT 2799.020 2624.370 2802.020 2624.380 ;
        RECT 2931.300 2624.370 2934.300 2624.380 ;
        RECT -14.680 2447.380 -11.680 2447.390 ;
        RECT 99.020 2447.380 102.020 2447.390 ;
        RECT 279.020 2447.380 282.020 2447.390 ;
        RECT 459.020 2447.380 462.020 2447.390 ;
        RECT 639.020 2447.380 642.020 2447.390 ;
        RECT 819.020 2447.380 822.020 2447.390 ;
        RECT 999.020 2447.380 1002.020 2447.390 ;
        RECT 1179.020 2447.380 1182.020 2447.390 ;
        RECT 1359.020 2447.380 1362.020 2447.390 ;
        RECT 1539.020 2447.380 1542.020 2447.390 ;
        RECT 1719.020 2447.380 1722.020 2447.390 ;
        RECT 1899.020 2447.380 1902.020 2447.390 ;
        RECT 2079.020 2447.380 2082.020 2447.390 ;
        RECT 2259.020 2447.380 2262.020 2447.390 ;
        RECT 2439.020 2447.380 2442.020 2447.390 ;
        RECT 2619.020 2447.380 2622.020 2447.390 ;
        RECT 2799.020 2447.380 2802.020 2447.390 ;
        RECT 2931.300 2447.380 2934.300 2447.390 ;
        RECT -14.680 2444.380 2934.300 2447.380 ;
        RECT -14.680 2444.370 -11.680 2444.380 ;
        RECT 99.020 2444.370 102.020 2444.380 ;
        RECT 279.020 2444.370 282.020 2444.380 ;
        RECT 459.020 2444.370 462.020 2444.380 ;
        RECT 639.020 2444.370 642.020 2444.380 ;
        RECT 819.020 2444.370 822.020 2444.380 ;
        RECT 999.020 2444.370 1002.020 2444.380 ;
        RECT 1179.020 2444.370 1182.020 2444.380 ;
        RECT 1359.020 2444.370 1362.020 2444.380 ;
        RECT 1539.020 2444.370 1542.020 2444.380 ;
        RECT 1719.020 2444.370 1722.020 2444.380 ;
        RECT 1899.020 2444.370 1902.020 2444.380 ;
        RECT 2079.020 2444.370 2082.020 2444.380 ;
        RECT 2259.020 2444.370 2262.020 2444.380 ;
        RECT 2439.020 2444.370 2442.020 2444.380 ;
        RECT 2619.020 2444.370 2622.020 2444.380 ;
        RECT 2799.020 2444.370 2802.020 2444.380 ;
        RECT 2931.300 2444.370 2934.300 2444.380 ;
        RECT -14.680 2267.380 -11.680 2267.390 ;
        RECT 99.020 2267.380 102.020 2267.390 ;
        RECT 279.020 2267.380 282.020 2267.390 ;
        RECT 459.020 2267.380 462.020 2267.390 ;
        RECT 639.020 2267.380 642.020 2267.390 ;
        RECT 819.020 2267.380 822.020 2267.390 ;
        RECT 999.020 2267.380 1002.020 2267.390 ;
        RECT 1179.020 2267.380 1182.020 2267.390 ;
        RECT 1359.020 2267.380 1362.020 2267.390 ;
        RECT 1539.020 2267.380 1542.020 2267.390 ;
        RECT 1719.020 2267.380 1722.020 2267.390 ;
        RECT 1899.020 2267.380 1902.020 2267.390 ;
        RECT 2079.020 2267.380 2082.020 2267.390 ;
        RECT 2259.020 2267.380 2262.020 2267.390 ;
        RECT 2439.020 2267.380 2442.020 2267.390 ;
        RECT 2619.020 2267.380 2622.020 2267.390 ;
        RECT 2799.020 2267.380 2802.020 2267.390 ;
        RECT 2931.300 2267.380 2934.300 2267.390 ;
        RECT -14.680 2264.380 2934.300 2267.380 ;
        RECT -14.680 2264.370 -11.680 2264.380 ;
        RECT 99.020 2264.370 102.020 2264.380 ;
        RECT 279.020 2264.370 282.020 2264.380 ;
        RECT 459.020 2264.370 462.020 2264.380 ;
        RECT 639.020 2264.370 642.020 2264.380 ;
        RECT 819.020 2264.370 822.020 2264.380 ;
        RECT 999.020 2264.370 1002.020 2264.380 ;
        RECT 1179.020 2264.370 1182.020 2264.380 ;
        RECT 1359.020 2264.370 1362.020 2264.380 ;
        RECT 1539.020 2264.370 1542.020 2264.380 ;
        RECT 1719.020 2264.370 1722.020 2264.380 ;
        RECT 1899.020 2264.370 1902.020 2264.380 ;
        RECT 2079.020 2264.370 2082.020 2264.380 ;
        RECT 2259.020 2264.370 2262.020 2264.380 ;
        RECT 2439.020 2264.370 2442.020 2264.380 ;
        RECT 2619.020 2264.370 2622.020 2264.380 ;
        RECT 2799.020 2264.370 2802.020 2264.380 ;
        RECT 2931.300 2264.370 2934.300 2264.380 ;
        RECT -14.680 2087.380 -11.680 2087.390 ;
        RECT 99.020 2087.380 102.020 2087.390 ;
        RECT 279.020 2087.380 282.020 2087.390 ;
        RECT 459.020 2087.380 462.020 2087.390 ;
        RECT 639.020 2087.380 642.020 2087.390 ;
        RECT 819.020 2087.380 822.020 2087.390 ;
        RECT 999.020 2087.380 1002.020 2087.390 ;
        RECT 1179.020 2087.380 1182.020 2087.390 ;
        RECT 1359.020 2087.380 1362.020 2087.390 ;
        RECT 1539.020 2087.380 1542.020 2087.390 ;
        RECT 1719.020 2087.380 1722.020 2087.390 ;
        RECT 1899.020 2087.380 1902.020 2087.390 ;
        RECT 2079.020 2087.380 2082.020 2087.390 ;
        RECT 2259.020 2087.380 2262.020 2087.390 ;
        RECT 2439.020 2087.380 2442.020 2087.390 ;
        RECT 2619.020 2087.380 2622.020 2087.390 ;
        RECT 2799.020 2087.380 2802.020 2087.390 ;
        RECT 2931.300 2087.380 2934.300 2087.390 ;
        RECT -14.680 2084.380 2934.300 2087.380 ;
        RECT -14.680 2084.370 -11.680 2084.380 ;
        RECT 99.020 2084.370 102.020 2084.380 ;
        RECT 279.020 2084.370 282.020 2084.380 ;
        RECT 459.020 2084.370 462.020 2084.380 ;
        RECT 639.020 2084.370 642.020 2084.380 ;
        RECT 819.020 2084.370 822.020 2084.380 ;
        RECT 999.020 2084.370 1002.020 2084.380 ;
        RECT 1179.020 2084.370 1182.020 2084.380 ;
        RECT 1359.020 2084.370 1362.020 2084.380 ;
        RECT 1539.020 2084.370 1542.020 2084.380 ;
        RECT 1719.020 2084.370 1722.020 2084.380 ;
        RECT 1899.020 2084.370 1902.020 2084.380 ;
        RECT 2079.020 2084.370 2082.020 2084.380 ;
        RECT 2259.020 2084.370 2262.020 2084.380 ;
        RECT 2439.020 2084.370 2442.020 2084.380 ;
        RECT 2619.020 2084.370 2622.020 2084.380 ;
        RECT 2799.020 2084.370 2802.020 2084.380 ;
        RECT 2931.300 2084.370 2934.300 2084.380 ;
        RECT -14.680 1907.380 -11.680 1907.390 ;
        RECT 99.020 1907.380 102.020 1907.390 ;
        RECT 279.020 1907.380 282.020 1907.390 ;
        RECT 459.020 1907.380 462.020 1907.390 ;
        RECT 639.020 1907.380 642.020 1907.390 ;
        RECT 819.020 1907.380 822.020 1907.390 ;
        RECT 999.020 1907.380 1002.020 1907.390 ;
        RECT 1179.020 1907.380 1182.020 1907.390 ;
        RECT 1359.020 1907.380 1362.020 1907.390 ;
        RECT 1539.020 1907.380 1542.020 1907.390 ;
        RECT 1719.020 1907.380 1722.020 1907.390 ;
        RECT 1899.020 1907.380 1902.020 1907.390 ;
        RECT 2079.020 1907.380 2082.020 1907.390 ;
        RECT 2259.020 1907.380 2262.020 1907.390 ;
        RECT 2439.020 1907.380 2442.020 1907.390 ;
        RECT 2619.020 1907.380 2622.020 1907.390 ;
        RECT 2799.020 1907.380 2802.020 1907.390 ;
        RECT 2931.300 1907.380 2934.300 1907.390 ;
        RECT -14.680 1904.380 2934.300 1907.380 ;
        RECT -14.680 1904.370 -11.680 1904.380 ;
        RECT 99.020 1904.370 102.020 1904.380 ;
        RECT 279.020 1904.370 282.020 1904.380 ;
        RECT 459.020 1904.370 462.020 1904.380 ;
        RECT 639.020 1904.370 642.020 1904.380 ;
        RECT 819.020 1904.370 822.020 1904.380 ;
        RECT 999.020 1904.370 1002.020 1904.380 ;
        RECT 1179.020 1904.370 1182.020 1904.380 ;
        RECT 1359.020 1904.370 1362.020 1904.380 ;
        RECT 1539.020 1904.370 1542.020 1904.380 ;
        RECT 1719.020 1904.370 1722.020 1904.380 ;
        RECT 1899.020 1904.370 1902.020 1904.380 ;
        RECT 2079.020 1904.370 2082.020 1904.380 ;
        RECT 2259.020 1904.370 2262.020 1904.380 ;
        RECT 2439.020 1904.370 2442.020 1904.380 ;
        RECT 2619.020 1904.370 2622.020 1904.380 ;
        RECT 2799.020 1904.370 2802.020 1904.380 ;
        RECT 2931.300 1904.370 2934.300 1904.380 ;
        RECT -14.680 1727.380 -11.680 1727.390 ;
        RECT 99.020 1727.380 102.020 1727.390 ;
        RECT 279.020 1727.380 282.020 1727.390 ;
        RECT 459.020 1727.380 462.020 1727.390 ;
        RECT 639.020 1727.380 642.020 1727.390 ;
        RECT 819.020 1727.380 822.020 1727.390 ;
        RECT 999.020 1727.380 1002.020 1727.390 ;
        RECT 1179.020 1727.380 1182.020 1727.390 ;
        RECT 1359.020 1727.380 1362.020 1727.390 ;
        RECT 1539.020 1727.380 1542.020 1727.390 ;
        RECT 1719.020 1727.380 1722.020 1727.390 ;
        RECT 1899.020 1727.380 1902.020 1727.390 ;
        RECT 2079.020 1727.380 2082.020 1727.390 ;
        RECT 2259.020 1727.380 2262.020 1727.390 ;
        RECT 2439.020 1727.380 2442.020 1727.390 ;
        RECT 2619.020 1727.380 2622.020 1727.390 ;
        RECT 2799.020 1727.380 2802.020 1727.390 ;
        RECT 2931.300 1727.380 2934.300 1727.390 ;
        RECT -14.680 1724.380 2934.300 1727.380 ;
        RECT -14.680 1724.370 -11.680 1724.380 ;
        RECT 99.020 1724.370 102.020 1724.380 ;
        RECT 279.020 1724.370 282.020 1724.380 ;
        RECT 459.020 1724.370 462.020 1724.380 ;
        RECT 639.020 1724.370 642.020 1724.380 ;
        RECT 819.020 1724.370 822.020 1724.380 ;
        RECT 999.020 1724.370 1002.020 1724.380 ;
        RECT 1179.020 1724.370 1182.020 1724.380 ;
        RECT 1359.020 1724.370 1362.020 1724.380 ;
        RECT 1539.020 1724.370 1542.020 1724.380 ;
        RECT 1719.020 1724.370 1722.020 1724.380 ;
        RECT 1899.020 1724.370 1902.020 1724.380 ;
        RECT 2079.020 1724.370 2082.020 1724.380 ;
        RECT 2259.020 1724.370 2262.020 1724.380 ;
        RECT 2439.020 1724.370 2442.020 1724.380 ;
        RECT 2619.020 1724.370 2622.020 1724.380 ;
        RECT 2799.020 1724.370 2802.020 1724.380 ;
        RECT 2931.300 1724.370 2934.300 1724.380 ;
        RECT -14.680 1547.380 -11.680 1547.390 ;
        RECT 99.020 1547.380 102.020 1547.390 ;
        RECT 279.020 1547.380 282.020 1547.390 ;
        RECT 459.020 1547.380 462.020 1547.390 ;
        RECT 639.020 1547.380 642.020 1547.390 ;
        RECT 819.020 1547.380 822.020 1547.390 ;
        RECT 999.020 1547.380 1002.020 1547.390 ;
        RECT 1179.020 1547.380 1182.020 1547.390 ;
        RECT 1359.020 1547.380 1362.020 1547.390 ;
        RECT 1539.020 1547.380 1542.020 1547.390 ;
        RECT 1719.020 1547.380 1722.020 1547.390 ;
        RECT 1899.020 1547.380 1902.020 1547.390 ;
        RECT 2079.020 1547.380 2082.020 1547.390 ;
        RECT 2259.020 1547.380 2262.020 1547.390 ;
        RECT 2439.020 1547.380 2442.020 1547.390 ;
        RECT 2619.020 1547.380 2622.020 1547.390 ;
        RECT 2799.020 1547.380 2802.020 1547.390 ;
        RECT 2931.300 1547.380 2934.300 1547.390 ;
        RECT -14.680 1544.380 2934.300 1547.380 ;
        RECT -14.680 1544.370 -11.680 1544.380 ;
        RECT 99.020 1544.370 102.020 1544.380 ;
        RECT 279.020 1544.370 282.020 1544.380 ;
        RECT 459.020 1544.370 462.020 1544.380 ;
        RECT 639.020 1544.370 642.020 1544.380 ;
        RECT 819.020 1544.370 822.020 1544.380 ;
        RECT 999.020 1544.370 1002.020 1544.380 ;
        RECT 1179.020 1544.370 1182.020 1544.380 ;
        RECT 1359.020 1544.370 1362.020 1544.380 ;
        RECT 1539.020 1544.370 1542.020 1544.380 ;
        RECT 1719.020 1544.370 1722.020 1544.380 ;
        RECT 1899.020 1544.370 1902.020 1544.380 ;
        RECT 2079.020 1544.370 2082.020 1544.380 ;
        RECT 2259.020 1544.370 2262.020 1544.380 ;
        RECT 2439.020 1544.370 2442.020 1544.380 ;
        RECT 2619.020 1544.370 2622.020 1544.380 ;
        RECT 2799.020 1544.370 2802.020 1544.380 ;
        RECT 2931.300 1544.370 2934.300 1544.380 ;
        RECT -14.680 1367.380 -11.680 1367.390 ;
        RECT 99.020 1367.380 102.020 1367.390 ;
        RECT 279.020 1367.380 282.020 1367.390 ;
        RECT 459.020 1367.380 462.020 1367.390 ;
        RECT 639.020 1367.380 642.020 1367.390 ;
        RECT 819.020 1367.380 822.020 1367.390 ;
        RECT 999.020 1367.380 1002.020 1367.390 ;
        RECT 1179.020 1367.380 1182.020 1367.390 ;
        RECT 1359.020 1367.380 1362.020 1367.390 ;
        RECT 1539.020 1367.380 1542.020 1367.390 ;
        RECT 1719.020 1367.380 1722.020 1367.390 ;
        RECT 1899.020 1367.380 1902.020 1367.390 ;
        RECT 2079.020 1367.380 2082.020 1367.390 ;
        RECT 2259.020 1367.380 2262.020 1367.390 ;
        RECT 2439.020 1367.380 2442.020 1367.390 ;
        RECT 2619.020 1367.380 2622.020 1367.390 ;
        RECT 2799.020 1367.380 2802.020 1367.390 ;
        RECT 2931.300 1367.380 2934.300 1367.390 ;
        RECT -14.680 1364.380 2934.300 1367.380 ;
        RECT -14.680 1364.370 -11.680 1364.380 ;
        RECT 99.020 1364.370 102.020 1364.380 ;
        RECT 279.020 1364.370 282.020 1364.380 ;
        RECT 459.020 1364.370 462.020 1364.380 ;
        RECT 639.020 1364.370 642.020 1364.380 ;
        RECT 819.020 1364.370 822.020 1364.380 ;
        RECT 999.020 1364.370 1002.020 1364.380 ;
        RECT 1179.020 1364.370 1182.020 1364.380 ;
        RECT 1359.020 1364.370 1362.020 1364.380 ;
        RECT 1539.020 1364.370 1542.020 1364.380 ;
        RECT 1719.020 1364.370 1722.020 1364.380 ;
        RECT 1899.020 1364.370 1902.020 1364.380 ;
        RECT 2079.020 1364.370 2082.020 1364.380 ;
        RECT 2259.020 1364.370 2262.020 1364.380 ;
        RECT 2439.020 1364.370 2442.020 1364.380 ;
        RECT 2619.020 1364.370 2622.020 1364.380 ;
        RECT 2799.020 1364.370 2802.020 1364.380 ;
        RECT 2931.300 1364.370 2934.300 1364.380 ;
        RECT -14.680 1187.380 -11.680 1187.390 ;
        RECT 99.020 1187.380 102.020 1187.390 ;
        RECT 279.020 1187.380 282.020 1187.390 ;
        RECT 459.020 1187.380 462.020 1187.390 ;
        RECT 639.020 1187.380 642.020 1187.390 ;
        RECT 819.020 1187.380 822.020 1187.390 ;
        RECT 999.020 1187.380 1002.020 1187.390 ;
        RECT 1179.020 1187.380 1182.020 1187.390 ;
        RECT 1359.020 1187.380 1362.020 1187.390 ;
        RECT 1539.020 1187.380 1542.020 1187.390 ;
        RECT 1719.020 1187.380 1722.020 1187.390 ;
        RECT 1899.020 1187.380 1902.020 1187.390 ;
        RECT 2079.020 1187.380 2082.020 1187.390 ;
        RECT 2259.020 1187.380 2262.020 1187.390 ;
        RECT 2439.020 1187.380 2442.020 1187.390 ;
        RECT 2619.020 1187.380 2622.020 1187.390 ;
        RECT 2799.020 1187.380 2802.020 1187.390 ;
        RECT 2931.300 1187.380 2934.300 1187.390 ;
        RECT -14.680 1184.380 2934.300 1187.380 ;
        RECT -14.680 1184.370 -11.680 1184.380 ;
        RECT 99.020 1184.370 102.020 1184.380 ;
        RECT 279.020 1184.370 282.020 1184.380 ;
        RECT 459.020 1184.370 462.020 1184.380 ;
        RECT 639.020 1184.370 642.020 1184.380 ;
        RECT 819.020 1184.370 822.020 1184.380 ;
        RECT 999.020 1184.370 1002.020 1184.380 ;
        RECT 1179.020 1184.370 1182.020 1184.380 ;
        RECT 1359.020 1184.370 1362.020 1184.380 ;
        RECT 1539.020 1184.370 1542.020 1184.380 ;
        RECT 1719.020 1184.370 1722.020 1184.380 ;
        RECT 1899.020 1184.370 1902.020 1184.380 ;
        RECT 2079.020 1184.370 2082.020 1184.380 ;
        RECT 2259.020 1184.370 2262.020 1184.380 ;
        RECT 2439.020 1184.370 2442.020 1184.380 ;
        RECT 2619.020 1184.370 2622.020 1184.380 ;
        RECT 2799.020 1184.370 2802.020 1184.380 ;
        RECT 2931.300 1184.370 2934.300 1184.380 ;
        RECT -14.680 1007.380 -11.680 1007.390 ;
        RECT 99.020 1007.380 102.020 1007.390 ;
        RECT 279.020 1007.380 282.020 1007.390 ;
        RECT 459.020 1007.380 462.020 1007.390 ;
        RECT 639.020 1007.380 642.020 1007.390 ;
        RECT 819.020 1007.380 822.020 1007.390 ;
        RECT 999.020 1007.380 1002.020 1007.390 ;
        RECT 1179.020 1007.380 1182.020 1007.390 ;
        RECT 1359.020 1007.380 1362.020 1007.390 ;
        RECT 1539.020 1007.380 1542.020 1007.390 ;
        RECT 1719.020 1007.380 1722.020 1007.390 ;
        RECT 1899.020 1007.380 1902.020 1007.390 ;
        RECT 2079.020 1007.380 2082.020 1007.390 ;
        RECT 2259.020 1007.380 2262.020 1007.390 ;
        RECT 2439.020 1007.380 2442.020 1007.390 ;
        RECT 2619.020 1007.380 2622.020 1007.390 ;
        RECT 2799.020 1007.380 2802.020 1007.390 ;
        RECT 2931.300 1007.380 2934.300 1007.390 ;
        RECT -14.680 1004.380 2934.300 1007.380 ;
        RECT -14.680 1004.370 -11.680 1004.380 ;
        RECT 99.020 1004.370 102.020 1004.380 ;
        RECT 279.020 1004.370 282.020 1004.380 ;
        RECT 459.020 1004.370 462.020 1004.380 ;
        RECT 639.020 1004.370 642.020 1004.380 ;
        RECT 819.020 1004.370 822.020 1004.380 ;
        RECT 999.020 1004.370 1002.020 1004.380 ;
        RECT 1179.020 1004.370 1182.020 1004.380 ;
        RECT 1359.020 1004.370 1362.020 1004.380 ;
        RECT 1539.020 1004.370 1542.020 1004.380 ;
        RECT 1719.020 1004.370 1722.020 1004.380 ;
        RECT 1899.020 1004.370 1902.020 1004.380 ;
        RECT 2079.020 1004.370 2082.020 1004.380 ;
        RECT 2259.020 1004.370 2262.020 1004.380 ;
        RECT 2439.020 1004.370 2442.020 1004.380 ;
        RECT 2619.020 1004.370 2622.020 1004.380 ;
        RECT 2799.020 1004.370 2802.020 1004.380 ;
        RECT 2931.300 1004.370 2934.300 1004.380 ;
        RECT -14.680 827.380 -11.680 827.390 ;
        RECT 99.020 827.380 102.020 827.390 ;
        RECT 279.020 827.380 282.020 827.390 ;
        RECT 459.020 827.380 462.020 827.390 ;
        RECT 639.020 827.380 642.020 827.390 ;
        RECT 819.020 827.380 822.020 827.390 ;
        RECT 999.020 827.380 1002.020 827.390 ;
        RECT 1179.020 827.380 1182.020 827.390 ;
        RECT 1359.020 827.380 1362.020 827.390 ;
        RECT 1539.020 827.380 1542.020 827.390 ;
        RECT 1719.020 827.380 1722.020 827.390 ;
        RECT 1899.020 827.380 1902.020 827.390 ;
        RECT 2079.020 827.380 2082.020 827.390 ;
        RECT 2259.020 827.380 2262.020 827.390 ;
        RECT 2439.020 827.380 2442.020 827.390 ;
        RECT 2619.020 827.380 2622.020 827.390 ;
        RECT 2799.020 827.380 2802.020 827.390 ;
        RECT 2931.300 827.380 2934.300 827.390 ;
        RECT -14.680 824.380 2934.300 827.380 ;
        RECT -14.680 824.370 -11.680 824.380 ;
        RECT 99.020 824.370 102.020 824.380 ;
        RECT 279.020 824.370 282.020 824.380 ;
        RECT 459.020 824.370 462.020 824.380 ;
        RECT 639.020 824.370 642.020 824.380 ;
        RECT 819.020 824.370 822.020 824.380 ;
        RECT 999.020 824.370 1002.020 824.380 ;
        RECT 1179.020 824.370 1182.020 824.380 ;
        RECT 1359.020 824.370 1362.020 824.380 ;
        RECT 1539.020 824.370 1542.020 824.380 ;
        RECT 1719.020 824.370 1722.020 824.380 ;
        RECT 1899.020 824.370 1902.020 824.380 ;
        RECT 2079.020 824.370 2082.020 824.380 ;
        RECT 2259.020 824.370 2262.020 824.380 ;
        RECT 2439.020 824.370 2442.020 824.380 ;
        RECT 2619.020 824.370 2622.020 824.380 ;
        RECT 2799.020 824.370 2802.020 824.380 ;
        RECT 2931.300 824.370 2934.300 824.380 ;
        RECT -14.680 647.380 -11.680 647.390 ;
        RECT 99.020 647.380 102.020 647.390 ;
        RECT 279.020 647.380 282.020 647.390 ;
        RECT 459.020 647.380 462.020 647.390 ;
        RECT 639.020 647.380 642.020 647.390 ;
        RECT 819.020 647.380 822.020 647.390 ;
        RECT 999.020 647.380 1002.020 647.390 ;
        RECT 1179.020 647.380 1182.020 647.390 ;
        RECT 1359.020 647.380 1362.020 647.390 ;
        RECT 1539.020 647.380 1542.020 647.390 ;
        RECT 1719.020 647.380 1722.020 647.390 ;
        RECT 1899.020 647.380 1902.020 647.390 ;
        RECT 2079.020 647.380 2082.020 647.390 ;
        RECT 2259.020 647.380 2262.020 647.390 ;
        RECT 2439.020 647.380 2442.020 647.390 ;
        RECT 2619.020 647.380 2622.020 647.390 ;
        RECT 2799.020 647.380 2802.020 647.390 ;
        RECT 2931.300 647.380 2934.300 647.390 ;
        RECT -14.680 644.380 2934.300 647.380 ;
        RECT -14.680 644.370 -11.680 644.380 ;
        RECT 99.020 644.370 102.020 644.380 ;
        RECT 279.020 644.370 282.020 644.380 ;
        RECT 459.020 644.370 462.020 644.380 ;
        RECT 639.020 644.370 642.020 644.380 ;
        RECT 819.020 644.370 822.020 644.380 ;
        RECT 999.020 644.370 1002.020 644.380 ;
        RECT 1179.020 644.370 1182.020 644.380 ;
        RECT 1359.020 644.370 1362.020 644.380 ;
        RECT 1539.020 644.370 1542.020 644.380 ;
        RECT 1719.020 644.370 1722.020 644.380 ;
        RECT 1899.020 644.370 1902.020 644.380 ;
        RECT 2079.020 644.370 2082.020 644.380 ;
        RECT 2259.020 644.370 2262.020 644.380 ;
        RECT 2439.020 644.370 2442.020 644.380 ;
        RECT 2619.020 644.370 2622.020 644.380 ;
        RECT 2799.020 644.370 2802.020 644.380 ;
        RECT 2931.300 644.370 2934.300 644.380 ;
        RECT -14.680 467.380 -11.680 467.390 ;
        RECT 99.020 467.380 102.020 467.390 ;
        RECT 279.020 467.380 282.020 467.390 ;
        RECT 459.020 467.380 462.020 467.390 ;
        RECT 639.020 467.380 642.020 467.390 ;
        RECT 819.020 467.380 822.020 467.390 ;
        RECT 999.020 467.380 1002.020 467.390 ;
        RECT 1179.020 467.380 1182.020 467.390 ;
        RECT 1359.020 467.380 1362.020 467.390 ;
        RECT 1539.020 467.380 1542.020 467.390 ;
        RECT 1719.020 467.380 1722.020 467.390 ;
        RECT 1899.020 467.380 1902.020 467.390 ;
        RECT 2079.020 467.380 2082.020 467.390 ;
        RECT 2259.020 467.380 2262.020 467.390 ;
        RECT 2439.020 467.380 2442.020 467.390 ;
        RECT 2619.020 467.380 2622.020 467.390 ;
        RECT 2799.020 467.380 2802.020 467.390 ;
        RECT 2931.300 467.380 2934.300 467.390 ;
        RECT -14.680 464.380 2934.300 467.380 ;
        RECT -14.680 464.370 -11.680 464.380 ;
        RECT 99.020 464.370 102.020 464.380 ;
        RECT 279.020 464.370 282.020 464.380 ;
        RECT 459.020 464.370 462.020 464.380 ;
        RECT 639.020 464.370 642.020 464.380 ;
        RECT 819.020 464.370 822.020 464.380 ;
        RECT 999.020 464.370 1002.020 464.380 ;
        RECT 1179.020 464.370 1182.020 464.380 ;
        RECT 1359.020 464.370 1362.020 464.380 ;
        RECT 1539.020 464.370 1542.020 464.380 ;
        RECT 1719.020 464.370 1722.020 464.380 ;
        RECT 1899.020 464.370 1902.020 464.380 ;
        RECT 2079.020 464.370 2082.020 464.380 ;
        RECT 2259.020 464.370 2262.020 464.380 ;
        RECT 2439.020 464.370 2442.020 464.380 ;
        RECT 2619.020 464.370 2622.020 464.380 ;
        RECT 2799.020 464.370 2802.020 464.380 ;
        RECT 2931.300 464.370 2934.300 464.380 ;
        RECT -14.680 287.380 -11.680 287.390 ;
        RECT 99.020 287.380 102.020 287.390 ;
        RECT 279.020 287.380 282.020 287.390 ;
        RECT 459.020 287.380 462.020 287.390 ;
        RECT 639.020 287.380 642.020 287.390 ;
        RECT 819.020 287.380 822.020 287.390 ;
        RECT 999.020 287.380 1002.020 287.390 ;
        RECT 1179.020 287.380 1182.020 287.390 ;
        RECT 1359.020 287.380 1362.020 287.390 ;
        RECT 1539.020 287.380 1542.020 287.390 ;
        RECT 1719.020 287.380 1722.020 287.390 ;
        RECT 1899.020 287.380 1902.020 287.390 ;
        RECT 2079.020 287.380 2082.020 287.390 ;
        RECT 2259.020 287.380 2262.020 287.390 ;
        RECT 2439.020 287.380 2442.020 287.390 ;
        RECT 2619.020 287.380 2622.020 287.390 ;
        RECT 2799.020 287.380 2802.020 287.390 ;
        RECT 2931.300 287.380 2934.300 287.390 ;
        RECT -14.680 284.380 2934.300 287.380 ;
        RECT -14.680 284.370 -11.680 284.380 ;
        RECT 99.020 284.370 102.020 284.380 ;
        RECT 279.020 284.370 282.020 284.380 ;
        RECT 459.020 284.370 462.020 284.380 ;
        RECT 639.020 284.370 642.020 284.380 ;
        RECT 819.020 284.370 822.020 284.380 ;
        RECT 999.020 284.370 1002.020 284.380 ;
        RECT 1179.020 284.370 1182.020 284.380 ;
        RECT 1359.020 284.370 1362.020 284.380 ;
        RECT 1539.020 284.370 1542.020 284.380 ;
        RECT 1719.020 284.370 1722.020 284.380 ;
        RECT 1899.020 284.370 1902.020 284.380 ;
        RECT 2079.020 284.370 2082.020 284.380 ;
        RECT 2259.020 284.370 2262.020 284.380 ;
        RECT 2439.020 284.370 2442.020 284.380 ;
        RECT 2619.020 284.370 2622.020 284.380 ;
        RECT 2799.020 284.370 2802.020 284.380 ;
        RECT 2931.300 284.370 2934.300 284.380 ;
        RECT -14.680 107.380 -11.680 107.390 ;
        RECT 99.020 107.380 102.020 107.390 ;
        RECT 279.020 107.380 282.020 107.390 ;
        RECT 459.020 107.380 462.020 107.390 ;
        RECT 639.020 107.380 642.020 107.390 ;
        RECT 819.020 107.380 822.020 107.390 ;
        RECT 999.020 107.380 1002.020 107.390 ;
        RECT 1179.020 107.380 1182.020 107.390 ;
        RECT 1359.020 107.380 1362.020 107.390 ;
        RECT 1539.020 107.380 1542.020 107.390 ;
        RECT 1719.020 107.380 1722.020 107.390 ;
        RECT 1899.020 107.380 1902.020 107.390 ;
        RECT 2079.020 107.380 2082.020 107.390 ;
        RECT 2259.020 107.380 2262.020 107.390 ;
        RECT 2439.020 107.380 2442.020 107.390 ;
        RECT 2619.020 107.380 2622.020 107.390 ;
        RECT 2799.020 107.380 2802.020 107.390 ;
        RECT 2931.300 107.380 2934.300 107.390 ;
        RECT -14.680 104.380 2934.300 107.380 ;
        RECT -14.680 104.370 -11.680 104.380 ;
        RECT 99.020 104.370 102.020 104.380 ;
        RECT 279.020 104.370 282.020 104.380 ;
        RECT 459.020 104.370 462.020 104.380 ;
        RECT 639.020 104.370 642.020 104.380 ;
        RECT 819.020 104.370 822.020 104.380 ;
        RECT 999.020 104.370 1002.020 104.380 ;
        RECT 1179.020 104.370 1182.020 104.380 ;
        RECT 1359.020 104.370 1362.020 104.380 ;
        RECT 1539.020 104.370 1542.020 104.380 ;
        RECT 1719.020 104.370 1722.020 104.380 ;
        RECT 1899.020 104.370 1902.020 104.380 ;
        RECT 2079.020 104.370 2082.020 104.380 ;
        RECT 2259.020 104.370 2262.020 104.380 ;
        RECT 2439.020 104.370 2442.020 104.380 ;
        RECT 2619.020 104.370 2622.020 104.380 ;
        RECT 2799.020 104.370 2802.020 104.380 ;
        RECT 2931.300 104.370 2934.300 104.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 99.020 -6.320 102.020 -6.310 ;
        RECT 279.020 -6.320 282.020 -6.310 ;
        RECT 459.020 -6.320 462.020 -6.310 ;
        RECT 639.020 -6.320 642.020 -6.310 ;
        RECT 819.020 -6.320 822.020 -6.310 ;
        RECT 999.020 -6.320 1002.020 -6.310 ;
        RECT 1179.020 -6.320 1182.020 -6.310 ;
        RECT 1359.020 -6.320 1362.020 -6.310 ;
        RECT 1539.020 -6.320 1542.020 -6.310 ;
        RECT 1719.020 -6.320 1722.020 -6.310 ;
        RECT 1899.020 -6.320 1902.020 -6.310 ;
        RECT 2079.020 -6.320 2082.020 -6.310 ;
        RECT 2259.020 -6.320 2262.020 -6.310 ;
        RECT 2439.020 -6.320 2442.020 -6.310 ;
        RECT 2619.020 -6.320 2622.020 -6.310 ;
        RECT 2799.020 -6.320 2802.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 99.020 -9.330 102.020 -9.320 ;
        RECT 279.020 -9.330 282.020 -9.320 ;
        RECT 459.020 -9.330 462.020 -9.320 ;
        RECT 639.020 -9.330 642.020 -9.320 ;
        RECT 819.020 -9.330 822.020 -9.320 ;
        RECT 999.020 -9.330 1002.020 -9.320 ;
        RECT 1179.020 -9.330 1182.020 -9.320 ;
        RECT 1359.020 -9.330 1362.020 -9.320 ;
        RECT 1539.020 -9.330 1542.020 -9.320 ;
        RECT 1719.020 -9.330 1722.020 -9.320 ;
        RECT 1899.020 -9.330 1902.020 -9.320 ;
        RECT 2079.020 -9.330 2082.020 -9.320 ;
        RECT 2259.020 -9.330 2262.020 -9.320 ;
        RECT 2439.020 -9.330 2442.020 -9.320 ;
        RECT 2619.020 -9.330 2622.020 -9.320 ;
        RECT 2799.020 -9.330 2802.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 27.020 -18.720 30.020 3538.400 ;
        RECT 207.020 -18.720 210.020 3538.400 ;
        RECT 387.020 -18.720 390.020 3538.400 ;
        RECT 567.020 -18.720 570.020 3538.400 ;
        RECT 747.020 -18.720 750.020 3538.400 ;
        RECT 927.020 -18.720 930.020 3538.400 ;
        RECT 1107.020 -18.720 1110.020 3538.400 ;
        RECT 1287.020 -18.720 1290.020 3538.400 ;
        RECT 1467.020 -18.720 1470.020 3538.400 ;
        RECT 1647.020 -18.720 1650.020 3538.400 ;
        RECT 1827.020 -18.720 1830.020 3538.400 ;
        RECT 2007.020 -18.720 2010.020 3538.400 ;
        RECT 2187.020 -18.720 2190.020 3538.400 ;
        RECT 2367.020 -18.720 2370.020 3538.400 ;
        RECT 2547.020 -18.720 2550.020 3538.400 ;
        RECT 2727.020 -18.720 2730.020 3538.400 ;
        RECT 2907.020 -18.720 2910.020 3538.400 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 3454.090 -17.290 3455.270 ;
        RECT -18.470 3452.490 -17.290 3453.670 ;
        RECT -18.470 3274.090 -17.290 3275.270 ;
        RECT -18.470 3272.490 -17.290 3273.670 ;
        RECT -18.470 3094.090 -17.290 3095.270 ;
        RECT -18.470 3092.490 -17.290 3093.670 ;
        RECT -18.470 2914.090 -17.290 2915.270 ;
        RECT -18.470 2912.490 -17.290 2913.670 ;
        RECT -18.470 2734.090 -17.290 2735.270 ;
        RECT -18.470 2732.490 -17.290 2733.670 ;
        RECT -18.470 2554.090 -17.290 2555.270 ;
        RECT -18.470 2552.490 -17.290 2553.670 ;
        RECT -18.470 2374.090 -17.290 2375.270 ;
        RECT -18.470 2372.490 -17.290 2373.670 ;
        RECT -18.470 2194.090 -17.290 2195.270 ;
        RECT -18.470 2192.490 -17.290 2193.670 ;
        RECT -18.470 2014.090 -17.290 2015.270 ;
        RECT -18.470 2012.490 -17.290 2013.670 ;
        RECT -18.470 1834.090 -17.290 1835.270 ;
        RECT -18.470 1832.490 -17.290 1833.670 ;
        RECT -18.470 1654.090 -17.290 1655.270 ;
        RECT -18.470 1652.490 -17.290 1653.670 ;
        RECT -18.470 1474.090 -17.290 1475.270 ;
        RECT -18.470 1472.490 -17.290 1473.670 ;
        RECT -18.470 1294.090 -17.290 1295.270 ;
        RECT -18.470 1292.490 -17.290 1293.670 ;
        RECT -18.470 1114.090 -17.290 1115.270 ;
        RECT -18.470 1112.490 -17.290 1113.670 ;
        RECT -18.470 934.090 -17.290 935.270 ;
        RECT -18.470 932.490 -17.290 933.670 ;
        RECT -18.470 754.090 -17.290 755.270 ;
        RECT -18.470 752.490 -17.290 753.670 ;
        RECT -18.470 574.090 -17.290 575.270 ;
        RECT -18.470 572.490 -17.290 573.670 ;
        RECT -18.470 394.090 -17.290 395.270 ;
        RECT -18.470 392.490 -17.290 393.670 ;
        RECT -18.470 214.090 -17.290 215.270 ;
        RECT -18.470 212.490 -17.290 213.670 ;
        RECT -18.470 34.090 -17.290 35.270 ;
        RECT -18.470 32.490 -17.290 33.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 27.930 3532.410 29.110 3533.590 ;
        RECT 27.930 3530.810 29.110 3531.990 ;
        RECT 27.930 3454.090 29.110 3455.270 ;
        RECT 27.930 3452.490 29.110 3453.670 ;
        RECT 27.930 3274.090 29.110 3275.270 ;
        RECT 27.930 3272.490 29.110 3273.670 ;
        RECT 27.930 3094.090 29.110 3095.270 ;
        RECT 27.930 3092.490 29.110 3093.670 ;
        RECT 27.930 2914.090 29.110 2915.270 ;
        RECT 27.930 2912.490 29.110 2913.670 ;
        RECT 27.930 2734.090 29.110 2735.270 ;
        RECT 27.930 2732.490 29.110 2733.670 ;
        RECT 27.930 2554.090 29.110 2555.270 ;
        RECT 27.930 2552.490 29.110 2553.670 ;
        RECT 27.930 2374.090 29.110 2375.270 ;
        RECT 27.930 2372.490 29.110 2373.670 ;
        RECT 27.930 2194.090 29.110 2195.270 ;
        RECT 27.930 2192.490 29.110 2193.670 ;
        RECT 27.930 2014.090 29.110 2015.270 ;
        RECT 27.930 2012.490 29.110 2013.670 ;
        RECT 27.930 1834.090 29.110 1835.270 ;
        RECT 27.930 1832.490 29.110 1833.670 ;
        RECT 27.930 1654.090 29.110 1655.270 ;
        RECT 27.930 1652.490 29.110 1653.670 ;
        RECT 27.930 1474.090 29.110 1475.270 ;
        RECT 27.930 1472.490 29.110 1473.670 ;
        RECT 27.930 1294.090 29.110 1295.270 ;
        RECT 27.930 1292.490 29.110 1293.670 ;
        RECT 27.930 1114.090 29.110 1115.270 ;
        RECT 27.930 1112.490 29.110 1113.670 ;
        RECT 27.930 934.090 29.110 935.270 ;
        RECT 27.930 932.490 29.110 933.670 ;
        RECT 27.930 754.090 29.110 755.270 ;
        RECT 27.930 752.490 29.110 753.670 ;
        RECT 27.930 574.090 29.110 575.270 ;
        RECT 27.930 572.490 29.110 573.670 ;
        RECT 27.930 394.090 29.110 395.270 ;
        RECT 27.930 392.490 29.110 393.670 ;
        RECT 27.930 214.090 29.110 215.270 ;
        RECT 27.930 212.490 29.110 213.670 ;
        RECT 27.930 34.090 29.110 35.270 ;
        RECT 27.930 32.490 29.110 33.670 ;
        RECT 27.930 -12.310 29.110 -11.130 ;
        RECT 27.930 -13.910 29.110 -12.730 ;
        RECT 207.930 3532.410 209.110 3533.590 ;
        RECT 207.930 3530.810 209.110 3531.990 ;
        RECT 207.930 3454.090 209.110 3455.270 ;
        RECT 207.930 3452.490 209.110 3453.670 ;
        RECT 207.930 3274.090 209.110 3275.270 ;
        RECT 207.930 3272.490 209.110 3273.670 ;
        RECT 207.930 3094.090 209.110 3095.270 ;
        RECT 207.930 3092.490 209.110 3093.670 ;
        RECT 207.930 2914.090 209.110 2915.270 ;
        RECT 207.930 2912.490 209.110 2913.670 ;
        RECT 207.930 2734.090 209.110 2735.270 ;
        RECT 207.930 2732.490 209.110 2733.670 ;
        RECT 207.930 2554.090 209.110 2555.270 ;
        RECT 207.930 2552.490 209.110 2553.670 ;
        RECT 207.930 2374.090 209.110 2375.270 ;
        RECT 207.930 2372.490 209.110 2373.670 ;
        RECT 207.930 2194.090 209.110 2195.270 ;
        RECT 207.930 2192.490 209.110 2193.670 ;
        RECT 207.930 2014.090 209.110 2015.270 ;
        RECT 207.930 2012.490 209.110 2013.670 ;
        RECT 207.930 1834.090 209.110 1835.270 ;
        RECT 207.930 1832.490 209.110 1833.670 ;
        RECT 207.930 1654.090 209.110 1655.270 ;
        RECT 207.930 1652.490 209.110 1653.670 ;
        RECT 207.930 1474.090 209.110 1475.270 ;
        RECT 207.930 1472.490 209.110 1473.670 ;
        RECT 207.930 1294.090 209.110 1295.270 ;
        RECT 207.930 1292.490 209.110 1293.670 ;
        RECT 207.930 1114.090 209.110 1115.270 ;
        RECT 207.930 1112.490 209.110 1113.670 ;
        RECT 207.930 934.090 209.110 935.270 ;
        RECT 207.930 932.490 209.110 933.670 ;
        RECT 207.930 754.090 209.110 755.270 ;
        RECT 207.930 752.490 209.110 753.670 ;
        RECT 207.930 574.090 209.110 575.270 ;
        RECT 207.930 572.490 209.110 573.670 ;
        RECT 207.930 394.090 209.110 395.270 ;
        RECT 207.930 392.490 209.110 393.670 ;
        RECT 207.930 214.090 209.110 215.270 ;
        RECT 207.930 212.490 209.110 213.670 ;
        RECT 207.930 34.090 209.110 35.270 ;
        RECT 207.930 32.490 209.110 33.670 ;
        RECT 207.930 -12.310 209.110 -11.130 ;
        RECT 207.930 -13.910 209.110 -12.730 ;
        RECT 387.930 3532.410 389.110 3533.590 ;
        RECT 387.930 3530.810 389.110 3531.990 ;
        RECT 387.930 3454.090 389.110 3455.270 ;
        RECT 387.930 3452.490 389.110 3453.670 ;
        RECT 387.930 3274.090 389.110 3275.270 ;
        RECT 387.930 3272.490 389.110 3273.670 ;
        RECT 387.930 3094.090 389.110 3095.270 ;
        RECT 387.930 3092.490 389.110 3093.670 ;
        RECT 387.930 2914.090 389.110 2915.270 ;
        RECT 387.930 2912.490 389.110 2913.670 ;
        RECT 387.930 2734.090 389.110 2735.270 ;
        RECT 387.930 2732.490 389.110 2733.670 ;
        RECT 387.930 2554.090 389.110 2555.270 ;
        RECT 387.930 2552.490 389.110 2553.670 ;
        RECT 387.930 2374.090 389.110 2375.270 ;
        RECT 387.930 2372.490 389.110 2373.670 ;
        RECT 387.930 2194.090 389.110 2195.270 ;
        RECT 387.930 2192.490 389.110 2193.670 ;
        RECT 387.930 2014.090 389.110 2015.270 ;
        RECT 387.930 2012.490 389.110 2013.670 ;
        RECT 387.930 1834.090 389.110 1835.270 ;
        RECT 387.930 1832.490 389.110 1833.670 ;
        RECT 387.930 1654.090 389.110 1655.270 ;
        RECT 387.930 1652.490 389.110 1653.670 ;
        RECT 387.930 1474.090 389.110 1475.270 ;
        RECT 387.930 1472.490 389.110 1473.670 ;
        RECT 387.930 1294.090 389.110 1295.270 ;
        RECT 387.930 1292.490 389.110 1293.670 ;
        RECT 387.930 1114.090 389.110 1115.270 ;
        RECT 387.930 1112.490 389.110 1113.670 ;
        RECT 387.930 934.090 389.110 935.270 ;
        RECT 387.930 932.490 389.110 933.670 ;
        RECT 387.930 754.090 389.110 755.270 ;
        RECT 387.930 752.490 389.110 753.670 ;
        RECT 387.930 574.090 389.110 575.270 ;
        RECT 387.930 572.490 389.110 573.670 ;
        RECT 387.930 394.090 389.110 395.270 ;
        RECT 387.930 392.490 389.110 393.670 ;
        RECT 387.930 214.090 389.110 215.270 ;
        RECT 387.930 212.490 389.110 213.670 ;
        RECT 387.930 34.090 389.110 35.270 ;
        RECT 387.930 32.490 389.110 33.670 ;
        RECT 387.930 -12.310 389.110 -11.130 ;
        RECT 387.930 -13.910 389.110 -12.730 ;
        RECT 567.930 3532.410 569.110 3533.590 ;
        RECT 567.930 3530.810 569.110 3531.990 ;
        RECT 567.930 3454.090 569.110 3455.270 ;
        RECT 567.930 3452.490 569.110 3453.670 ;
        RECT 567.930 3274.090 569.110 3275.270 ;
        RECT 567.930 3272.490 569.110 3273.670 ;
        RECT 567.930 3094.090 569.110 3095.270 ;
        RECT 567.930 3092.490 569.110 3093.670 ;
        RECT 567.930 2914.090 569.110 2915.270 ;
        RECT 567.930 2912.490 569.110 2913.670 ;
        RECT 567.930 2734.090 569.110 2735.270 ;
        RECT 567.930 2732.490 569.110 2733.670 ;
        RECT 567.930 2554.090 569.110 2555.270 ;
        RECT 567.930 2552.490 569.110 2553.670 ;
        RECT 567.930 2374.090 569.110 2375.270 ;
        RECT 567.930 2372.490 569.110 2373.670 ;
        RECT 567.930 2194.090 569.110 2195.270 ;
        RECT 567.930 2192.490 569.110 2193.670 ;
        RECT 567.930 2014.090 569.110 2015.270 ;
        RECT 567.930 2012.490 569.110 2013.670 ;
        RECT 567.930 1834.090 569.110 1835.270 ;
        RECT 567.930 1832.490 569.110 1833.670 ;
        RECT 567.930 1654.090 569.110 1655.270 ;
        RECT 567.930 1652.490 569.110 1653.670 ;
        RECT 567.930 1474.090 569.110 1475.270 ;
        RECT 567.930 1472.490 569.110 1473.670 ;
        RECT 567.930 1294.090 569.110 1295.270 ;
        RECT 567.930 1292.490 569.110 1293.670 ;
        RECT 567.930 1114.090 569.110 1115.270 ;
        RECT 567.930 1112.490 569.110 1113.670 ;
        RECT 567.930 934.090 569.110 935.270 ;
        RECT 567.930 932.490 569.110 933.670 ;
        RECT 567.930 754.090 569.110 755.270 ;
        RECT 567.930 752.490 569.110 753.670 ;
        RECT 567.930 574.090 569.110 575.270 ;
        RECT 567.930 572.490 569.110 573.670 ;
        RECT 567.930 394.090 569.110 395.270 ;
        RECT 567.930 392.490 569.110 393.670 ;
        RECT 567.930 214.090 569.110 215.270 ;
        RECT 567.930 212.490 569.110 213.670 ;
        RECT 567.930 34.090 569.110 35.270 ;
        RECT 567.930 32.490 569.110 33.670 ;
        RECT 567.930 -12.310 569.110 -11.130 ;
        RECT 567.930 -13.910 569.110 -12.730 ;
        RECT 747.930 3532.410 749.110 3533.590 ;
        RECT 747.930 3530.810 749.110 3531.990 ;
        RECT 747.930 3454.090 749.110 3455.270 ;
        RECT 747.930 3452.490 749.110 3453.670 ;
        RECT 747.930 3274.090 749.110 3275.270 ;
        RECT 747.930 3272.490 749.110 3273.670 ;
        RECT 747.930 3094.090 749.110 3095.270 ;
        RECT 747.930 3092.490 749.110 3093.670 ;
        RECT 747.930 2914.090 749.110 2915.270 ;
        RECT 747.930 2912.490 749.110 2913.670 ;
        RECT 747.930 2734.090 749.110 2735.270 ;
        RECT 747.930 2732.490 749.110 2733.670 ;
        RECT 747.930 2554.090 749.110 2555.270 ;
        RECT 747.930 2552.490 749.110 2553.670 ;
        RECT 747.930 2374.090 749.110 2375.270 ;
        RECT 747.930 2372.490 749.110 2373.670 ;
        RECT 747.930 2194.090 749.110 2195.270 ;
        RECT 747.930 2192.490 749.110 2193.670 ;
        RECT 747.930 2014.090 749.110 2015.270 ;
        RECT 747.930 2012.490 749.110 2013.670 ;
        RECT 747.930 1834.090 749.110 1835.270 ;
        RECT 747.930 1832.490 749.110 1833.670 ;
        RECT 747.930 1654.090 749.110 1655.270 ;
        RECT 747.930 1652.490 749.110 1653.670 ;
        RECT 747.930 1474.090 749.110 1475.270 ;
        RECT 747.930 1472.490 749.110 1473.670 ;
        RECT 747.930 1294.090 749.110 1295.270 ;
        RECT 747.930 1292.490 749.110 1293.670 ;
        RECT 747.930 1114.090 749.110 1115.270 ;
        RECT 747.930 1112.490 749.110 1113.670 ;
        RECT 747.930 934.090 749.110 935.270 ;
        RECT 747.930 932.490 749.110 933.670 ;
        RECT 747.930 754.090 749.110 755.270 ;
        RECT 747.930 752.490 749.110 753.670 ;
        RECT 747.930 574.090 749.110 575.270 ;
        RECT 747.930 572.490 749.110 573.670 ;
        RECT 747.930 394.090 749.110 395.270 ;
        RECT 747.930 392.490 749.110 393.670 ;
        RECT 747.930 214.090 749.110 215.270 ;
        RECT 747.930 212.490 749.110 213.670 ;
        RECT 747.930 34.090 749.110 35.270 ;
        RECT 747.930 32.490 749.110 33.670 ;
        RECT 747.930 -12.310 749.110 -11.130 ;
        RECT 747.930 -13.910 749.110 -12.730 ;
        RECT 927.930 3532.410 929.110 3533.590 ;
        RECT 927.930 3530.810 929.110 3531.990 ;
        RECT 927.930 3454.090 929.110 3455.270 ;
        RECT 927.930 3452.490 929.110 3453.670 ;
        RECT 927.930 3274.090 929.110 3275.270 ;
        RECT 927.930 3272.490 929.110 3273.670 ;
        RECT 927.930 3094.090 929.110 3095.270 ;
        RECT 927.930 3092.490 929.110 3093.670 ;
        RECT 927.930 2914.090 929.110 2915.270 ;
        RECT 927.930 2912.490 929.110 2913.670 ;
        RECT 927.930 2734.090 929.110 2735.270 ;
        RECT 927.930 2732.490 929.110 2733.670 ;
        RECT 927.930 2554.090 929.110 2555.270 ;
        RECT 927.930 2552.490 929.110 2553.670 ;
        RECT 927.930 2374.090 929.110 2375.270 ;
        RECT 927.930 2372.490 929.110 2373.670 ;
        RECT 927.930 2194.090 929.110 2195.270 ;
        RECT 927.930 2192.490 929.110 2193.670 ;
        RECT 927.930 2014.090 929.110 2015.270 ;
        RECT 927.930 2012.490 929.110 2013.670 ;
        RECT 927.930 1834.090 929.110 1835.270 ;
        RECT 927.930 1832.490 929.110 1833.670 ;
        RECT 927.930 1654.090 929.110 1655.270 ;
        RECT 927.930 1652.490 929.110 1653.670 ;
        RECT 927.930 1474.090 929.110 1475.270 ;
        RECT 927.930 1472.490 929.110 1473.670 ;
        RECT 927.930 1294.090 929.110 1295.270 ;
        RECT 927.930 1292.490 929.110 1293.670 ;
        RECT 927.930 1114.090 929.110 1115.270 ;
        RECT 927.930 1112.490 929.110 1113.670 ;
        RECT 927.930 934.090 929.110 935.270 ;
        RECT 927.930 932.490 929.110 933.670 ;
        RECT 927.930 754.090 929.110 755.270 ;
        RECT 927.930 752.490 929.110 753.670 ;
        RECT 927.930 574.090 929.110 575.270 ;
        RECT 927.930 572.490 929.110 573.670 ;
        RECT 927.930 394.090 929.110 395.270 ;
        RECT 927.930 392.490 929.110 393.670 ;
        RECT 927.930 214.090 929.110 215.270 ;
        RECT 927.930 212.490 929.110 213.670 ;
        RECT 927.930 34.090 929.110 35.270 ;
        RECT 927.930 32.490 929.110 33.670 ;
        RECT 927.930 -12.310 929.110 -11.130 ;
        RECT 927.930 -13.910 929.110 -12.730 ;
        RECT 1107.930 3532.410 1109.110 3533.590 ;
        RECT 1107.930 3530.810 1109.110 3531.990 ;
        RECT 1107.930 3454.090 1109.110 3455.270 ;
        RECT 1107.930 3452.490 1109.110 3453.670 ;
        RECT 1107.930 3274.090 1109.110 3275.270 ;
        RECT 1107.930 3272.490 1109.110 3273.670 ;
        RECT 1107.930 3094.090 1109.110 3095.270 ;
        RECT 1107.930 3092.490 1109.110 3093.670 ;
        RECT 1107.930 2914.090 1109.110 2915.270 ;
        RECT 1107.930 2912.490 1109.110 2913.670 ;
        RECT 1107.930 2734.090 1109.110 2735.270 ;
        RECT 1107.930 2732.490 1109.110 2733.670 ;
        RECT 1107.930 2554.090 1109.110 2555.270 ;
        RECT 1107.930 2552.490 1109.110 2553.670 ;
        RECT 1107.930 2374.090 1109.110 2375.270 ;
        RECT 1107.930 2372.490 1109.110 2373.670 ;
        RECT 1107.930 2194.090 1109.110 2195.270 ;
        RECT 1107.930 2192.490 1109.110 2193.670 ;
        RECT 1107.930 2014.090 1109.110 2015.270 ;
        RECT 1107.930 2012.490 1109.110 2013.670 ;
        RECT 1107.930 1834.090 1109.110 1835.270 ;
        RECT 1107.930 1832.490 1109.110 1833.670 ;
        RECT 1107.930 1654.090 1109.110 1655.270 ;
        RECT 1107.930 1652.490 1109.110 1653.670 ;
        RECT 1107.930 1474.090 1109.110 1475.270 ;
        RECT 1107.930 1472.490 1109.110 1473.670 ;
        RECT 1107.930 1294.090 1109.110 1295.270 ;
        RECT 1107.930 1292.490 1109.110 1293.670 ;
        RECT 1107.930 1114.090 1109.110 1115.270 ;
        RECT 1107.930 1112.490 1109.110 1113.670 ;
        RECT 1107.930 934.090 1109.110 935.270 ;
        RECT 1107.930 932.490 1109.110 933.670 ;
        RECT 1107.930 754.090 1109.110 755.270 ;
        RECT 1107.930 752.490 1109.110 753.670 ;
        RECT 1107.930 574.090 1109.110 575.270 ;
        RECT 1107.930 572.490 1109.110 573.670 ;
        RECT 1107.930 394.090 1109.110 395.270 ;
        RECT 1107.930 392.490 1109.110 393.670 ;
        RECT 1107.930 214.090 1109.110 215.270 ;
        RECT 1107.930 212.490 1109.110 213.670 ;
        RECT 1107.930 34.090 1109.110 35.270 ;
        RECT 1107.930 32.490 1109.110 33.670 ;
        RECT 1107.930 -12.310 1109.110 -11.130 ;
        RECT 1107.930 -13.910 1109.110 -12.730 ;
        RECT 1287.930 3532.410 1289.110 3533.590 ;
        RECT 1287.930 3530.810 1289.110 3531.990 ;
        RECT 1287.930 3454.090 1289.110 3455.270 ;
        RECT 1287.930 3452.490 1289.110 3453.670 ;
        RECT 1287.930 3274.090 1289.110 3275.270 ;
        RECT 1287.930 3272.490 1289.110 3273.670 ;
        RECT 1287.930 3094.090 1289.110 3095.270 ;
        RECT 1287.930 3092.490 1289.110 3093.670 ;
        RECT 1287.930 2914.090 1289.110 2915.270 ;
        RECT 1287.930 2912.490 1289.110 2913.670 ;
        RECT 1287.930 2734.090 1289.110 2735.270 ;
        RECT 1287.930 2732.490 1289.110 2733.670 ;
        RECT 1287.930 2554.090 1289.110 2555.270 ;
        RECT 1287.930 2552.490 1289.110 2553.670 ;
        RECT 1287.930 2374.090 1289.110 2375.270 ;
        RECT 1287.930 2372.490 1289.110 2373.670 ;
        RECT 1287.930 2194.090 1289.110 2195.270 ;
        RECT 1287.930 2192.490 1289.110 2193.670 ;
        RECT 1287.930 2014.090 1289.110 2015.270 ;
        RECT 1287.930 2012.490 1289.110 2013.670 ;
        RECT 1287.930 1834.090 1289.110 1835.270 ;
        RECT 1287.930 1832.490 1289.110 1833.670 ;
        RECT 1287.930 1654.090 1289.110 1655.270 ;
        RECT 1287.930 1652.490 1289.110 1653.670 ;
        RECT 1287.930 1474.090 1289.110 1475.270 ;
        RECT 1287.930 1472.490 1289.110 1473.670 ;
        RECT 1287.930 1294.090 1289.110 1295.270 ;
        RECT 1287.930 1292.490 1289.110 1293.670 ;
        RECT 1287.930 1114.090 1289.110 1115.270 ;
        RECT 1287.930 1112.490 1289.110 1113.670 ;
        RECT 1287.930 934.090 1289.110 935.270 ;
        RECT 1287.930 932.490 1289.110 933.670 ;
        RECT 1287.930 754.090 1289.110 755.270 ;
        RECT 1287.930 752.490 1289.110 753.670 ;
        RECT 1287.930 574.090 1289.110 575.270 ;
        RECT 1287.930 572.490 1289.110 573.670 ;
        RECT 1287.930 394.090 1289.110 395.270 ;
        RECT 1287.930 392.490 1289.110 393.670 ;
        RECT 1287.930 214.090 1289.110 215.270 ;
        RECT 1287.930 212.490 1289.110 213.670 ;
        RECT 1287.930 34.090 1289.110 35.270 ;
        RECT 1287.930 32.490 1289.110 33.670 ;
        RECT 1287.930 -12.310 1289.110 -11.130 ;
        RECT 1287.930 -13.910 1289.110 -12.730 ;
        RECT 1467.930 3532.410 1469.110 3533.590 ;
        RECT 1467.930 3530.810 1469.110 3531.990 ;
        RECT 1467.930 3454.090 1469.110 3455.270 ;
        RECT 1467.930 3452.490 1469.110 3453.670 ;
        RECT 1467.930 3274.090 1469.110 3275.270 ;
        RECT 1467.930 3272.490 1469.110 3273.670 ;
        RECT 1467.930 3094.090 1469.110 3095.270 ;
        RECT 1467.930 3092.490 1469.110 3093.670 ;
        RECT 1467.930 2914.090 1469.110 2915.270 ;
        RECT 1467.930 2912.490 1469.110 2913.670 ;
        RECT 1467.930 2734.090 1469.110 2735.270 ;
        RECT 1467.930 2732.490 1469.110 2733.670 ;
        RECT 1467.930 2554.090 1469.110 2555.270 ;
        RECT 1467.930 2552.490 1469.110 2553.670 ;
        RECT 1467.930 2374.090 1469.110 2375.270 ;
        RECT 1467.930 2372.490 1469.110 2373.670 ;
        RECT 1467.930 2194.090 1469.110 2195.270 ;
        RECT 1467.930 2192.490 1469.110 2193.670 ;
        RECT 1467.930 2014.090 1469.110 2015.270 ;
        RECT 1467.930 2012.490 1469.110 2013.670 ;
        RECT 1467.930 1834.090 1469.110 1835.270 ;
        RECT 1467.930 1832.490 1469.110 1833.670 ;
        RECT 1467.930 1654.090 1469.110 1655.270 ;
        RECT 1467.930 1652.490 1469.110 1653.670 ;
        RECT 1467.930 1474.090 1469.110 1475.270 ;
        RECT 1467.930 1472.490 1469.110 1473.670 ;
        RECT 1467.930 1294.090 1469.110 1295.270 ;
        RECT 1467.930 1292.490 1469.110 1293.670 ;
        RECT 1467.930 1114.090 1469.110 1115.270 ;
        RECT 1467.930 1112.490 1469.110 1113.670 ;
        RECT 1467.930 934.090 1469.110 935.270 ;
        RECT 1467.930 932.490 1469.110 933.670 ;
        RECT 1467.930 754.090 1469.110 755.270 ;
        RECT 1467.930 752.490 1469.110 753.670 ;
        RECT 1467.930 574.090 1469.110 575.270 ;
        RECT 1467.930 572.490 1469.110 573.670 ;
        RECT 1467.930 394.090 1469.110 395.270 ;
        RECT 1467.930 392.490 1469.110 393.670 ;
        RECT 1467.930 214.090 1469.110 215.270 ;
        RECT 1467.930 212.490 1469.110 213.670 ;
        RECT 1467.930 34.090 1469.110 35.270 ;
        RECT 1467.930 32.490 1469.110 33.670 ;
        RECT 1467.930 -12.310 1469.110 -11.130 ;
        RECT 1467.930 -13.910 1469.110 -12.730 ;
        RECT 1647.930 3532.410 1649.110 3533.590 ;
        RECT 1647.930 3530.810 1649.110 3531.990 ;
        RECT 1647.930 3454.090 1649.110 3455.270 ;
        RECT 1647.930 3452.490 1649.110 3453.670 ;
        RECT 1647.930 3274.090 1649.110 3275.270 ;
        RECT 1647.930 3272.490 1649.110 3273.670 ;
        RECT 1647.930 3094.090 1649.110 3095.270 ;
        RECT 1647.930 3092.490 1649.110 3093.670 ;
        RECT 1647.930 2914.090 1649.110 2915.270 ;
        RECT 1647.930 2912.490 1649.110 2913.670 ;
        RECT 1647.930 2734.090 1649.110 2735.270 ;
        RECT 1647.930 2732.490 1649.110 2733.670 ;
        RECT 1647.930 2554.090 1649.110 2555.270 ;
        RECT 1647.930 2552.490 1649.110 2553.670 ;
        RECT 1647.930 2374.090 1649.110 2375.270 ;
        RECT 1647.930 2372.490 1649.110 2373.670 ;
        RECT 1647.930 2194.090 1649.110 2195.270 ;
        RECT 1647.930 2192.490 1649.110 2193.670 ;
        RECT 1647.930 2014.090 1649.110 2015.270 ;
        RECT 1647.930 2012.490 1649.110 2013.670 ;
        RECT 1647.930 1834.090 1649.110 1835.270 ;
        RECT 1647.930 1832.490 1649.110 1833.670 ;
        RECT 1647.930 1654.090 1649.110 1655.270 ;
        RECT 1647.930 1652.490 1649.110 1653.670 ;
        RECT 1647.930 1474.090 1649.110 1475.270 ;
        RECT 1647.930 1472.490 1649.110 1473.670 ;
        RECT 1647.930 1294.090 1649.110 1295.270 ;
        RECT 1647.930 1292.490 1649.110 1293.670 ;
        RECT 1647.930 1114.090 1649.110 1115.270 ;
        RECT 1647.930 1112.490 1649.110 1113.670 ;
        RECT 1647.930 934.090 1649.110 935.270 ;
        RECT 1647.930 932.490 1649.110 933.670 ;
        RECT 1647.930 754.090 1649.110 755.270 ;
        RECT 1647.930 752.490 1649.110 753.670 ;
        RECT 1647.930 574.090 1649.110 575.270 ;
        RECT 1647.930 572.490 1649.110 573.670 ;
        RECT 1647.930 394.090 1649.110 395.270 ;
        RECT 1647.930 392.490 1649.110 393.670 ;
        RECT 1647.930 214.090 1649.110 215.270 ;
        RECT 1647.930 212.490 1649.110 213.670 ;
        RECT 1647.930 34.090 1649.110 35.270 ;
        RECT 1647.930 32.490 1649.110 33.670 ;
        RECT 1647.930 -12.310 1649.110 -11.130 ;
        RECT 1647.930 -13.910 1649.110 -12.730 ;
        RECT 1827.930 3532.410 1829.110 3533.590 ;
        RECT 1827.930 3530.810 1829.110 3531.990 ;
        RECT 1827.930 3454.090 1829.110 3455.270 ;
        RECT 1827.930 3452.490 1829.110 3453.670 ;
        RECT 1827.930 3274.090 1829.110 3275.270 ;
        RECT 1827.930 3272.490 1829.110 3273.670 ;
        RECT 1827.930 3094.090 1829.110 3095.270 ;
        RECT 1827.930 3092.490 1829.110 3093.670 ;
        RECT 1827.930 2914.090 1829.110 2915.270 ;
        RECT 1827.930 2912.490 1829.110 2913.670 ;
        RECT 1827.930 2734.090 1829.110 2735.270 ;
        RECT 1827.930 2732.490 1829.110 2733.670 ;
        RECT 1827.930 2554.090 1829.110 2555.270 ;
        RECT 1827.930 2552.490 1829.110 2553.670 ;
        RECT 1827.930 2374.090 1829.110 2375.270 ;
        RECT 1827.930 2372.490 1829.110 2373.670 ;
        RECT 1827.930 2194.090 1829.110 2195.270 ;
        RECT 1827.930 2192.490 1829.110 2193.670 ;
        RECT 1827.930 2014.090 1829.110 2015.270 ;
        RECT 1827.930 2012.490 1829.110 2013.670 ;
        RECT 1827.930 1834.090 1829.110 1835.270 ;
        RECT 1827.930 1832.490 1829.110 1833.670 ;
        RECT 1827.930 1654.090 1829.110 1655.270 ;
        RECT 1827.930 1652.490 1829.110 1653.670 ;
        RECT 1827.930 1474.090 1829.110 1475.270 ;
        RECT 1827.930 1472.490 1829.110 1473.670 ;
        RECT 1827.930 1294.090 1829.110 1295.270 ;
        RECT 1827.930 1292.490 1829.110 1293.670 ;
        RECT 1827.930 1114.090 1829.110 1115.270 ;
        RECT 1827.930 1112.490 1829.110 1113.670 ;
        RECT 1827.930 934.090 1829.110 935.270 ;
        RECT 1827.930 932.490 1829.110 933.670 ;
        RECT 1827.930 754.090 1829.110 755.270 ;
        RECT 1827.930 752.490 1829.110 753.670 ;
        RECT 1827.930 574.090 1829.110 575.270 ;
        RECT 1827.930 572.490 1829.110 573.670 ;
        RECT 1827.930 394.090 1829.110 395.270 ;
        RECT 1827.930 392.490 1829.110 393.670 ;
        RECT 1827.930 214.090 1829.110 215.270 ;
        RECT 1827.930 212.490 1829.110 213.670 ;
        RECT 1827.930 34.090 1829.110 35.270 ;
        RECT 1827.930 32.490 1829.110 33.670 ;
        RECT 1827.930 -12.310 1829.110 -11.130 ;
        RECT 1827.930 -13.910 1829.110 -12.730 ;
        RECT 2007.930 3532.410 2009.110 3533.590 ;
        RECT 2007.930 3530.810 2009.110 3531.990 ;
        RECT 2007.930 3454.090 2009.110 3455.270 ;
        RECT 2007.930 3452.490 2009.110 3453.670 ;
        RECT 2007.930 3274.090 2009.110 3275.270 ;
        RECT 2007.930 3272.490 2009.110 3273.670 ;
        RECT 2007.930 3094.090 2009.110 3095.270 ;
        RECT 2007.930 3092.490 2009.110 3093.670 ;
        RECT 2007.930 2914.090 2009.110 2915.270 ;
        RECT 2007.930 2912.490 2009.110 2913.670 ;
        RECT 2007.930 2734.090 2009.110 2735.270 ;
        RECT 2007.930 2732.490 2009.110 2733.670 ;
        RECT 2007.930 2554.090 2009.110 2555.270 ;
        RECT 2007.930 2552.490 2009.110 2553.670 ;
        RECT 2007.930 2374.090 2009.110 2375.270 ;
        RECT 2007.930 2372.490 2009.110 2373.670 ;
        RECT 2007.930 2194.090 2009.110 2195.270 ;
        RECT 2007.930 2192.490 2009.110 2193.670 ;
        RECT 2007.930 2014.090 2009.110 2015.270 ;
        RECT 2007.930 2012.490 2009.110 2013.670 ;
        RECT 2007.930 1834.090 2009.110 1835.270 ;
        RECT 2007.930 1832.490 2009.110 1833.670 ;
        RECT 2007.930 1654.090 2009.110 1655.270 ;
        RECT 2007.930 1652.490 2009.110 1653.670 ;
        RECT 2007.930 1474.090 2009.110 1475.270 ;
        RECT 2007.930 1472.490 2009.110 1473.670 ;
        RECT 2007.930 1294.090 2009.110 1295.270 ;
        RECT 2007.930 1292.490 2009.110 1293.670 ;
        RECT 2007.930 1114.090 2009.110 1115.270 ;
        RECT 2007.930 1112.490 2009.110 1113.670 ;
        RECT 2007.930 934.090 2009.110 935.270 ;
        RECT 2007.930 932.490 2009.110 933.670 ;
        RECT 2007.930 754.090 2009.110 755.270 ;
        RECT 2007.930 752.490 2009.110 753.670 ;
        RECT 2007.930 574.090 2009.110 575.270 ;
        RECT 2007.930 572.490 2009.110 573.670 ;
        RECT 2007.930 394.090 2009.110 395.270 ;
        RECT 2007.930 392.490 2009.110 393.670 ;
        RECT 2007.930 214.090 2009.110 215.270 ;
        RECT 2007.930 212.490 2009.110 213.670 ;
        RECT 2007.930 34.090 2009.110 35.270 ;
        RECT 2007.930 32.490 2009.110 33.670 ;
        RECT 2007.930 -12.310 2009.110 -11.130 ;
        RECT 2007.930 -13.910 2009.110 -12.730 ;
        RECT 2187.930 3532.410 2189.110 3533.590 ;
        RECT 2187.930 3530.810 2189.110 3531.990 ;
        RECT 2187.930 3454.090 2189.110 3455.270 ;
        RECT 2187.930 3452.490 2189.110 3453.670 ;
        RECT 2187.930 3274.090 2189.110 3275.270 ;
        RECT 2187.930 3272.490 2189.110 3273.670 ;
        RECT 2187.930 3094.090 2189.110 3095.270 ;
        RECT 2187.930 3092.490 2189.110 3093.670 ;
        RECT 2187.930 2914.090 2189.110 2915.270 ;
        RECT 2187.930 2912.490 2189.110 2913.670 ;
        RECT 2187.930 2734.090 2189.110 2735.270 ;
        RECT 2187.930 2732.490 2189.110 2733.670 ;
        RECT 2187.930 2554.090 2189.110 2555.270 ;
        RECT 2187.930 2552.490 2189.110 2553.670 ;
        RECT 2187.930 2374.090 2189.110 2375.270 ;
        RECT 2187.930 2372.490 2189.110 2373.670 ;
        RECT 2187.930 2194.090 2189.110 2195.270 ;
        RECT 2187.930 2192.490 2189.110 2193.670 ;
        RECT 2187.930 2014.090 2189.110 2015.270 ;
        RECT 2187.930 2012.490 2189.110 2013.670 ;
        RECT 2187.930 1834.090 2189.110 1835.270 ;
        RECT 2187.930 1832.490 2189.110 1833.670 ;
        RECT 2187.930 1654.090 2189.110 1655.270 ;
        RECT 2187.930 1652.490 2189.110 1653.670 ;
        RECT 2187.930 1474.090 2189.110 1475.270 ;
        RECT 2187.930 1472.490 2189.110 1473.670 ;
        RECT 2187.930 1294.090 2189.110 1295.270 ;
        RECT 2187.930 1292.490 2189.110 1293.670 ;
        RECT 2187.930 1114.090 2189.110 1115.270 ;
        RECT 2187.930 1112.490 2189.110 1113.670 ;
        RECT 2187.930 934.090 2189.110 935.270 ;
        RECT 2187.930 932.490 2189.110 933.670 ;
        RECT 2187.930 754.090 2189.110 755.270 ;
        RECT 2187.930 752.490 2189.110 753.670 ;
        RECT 2187.930 574.090 2189.110 575.270 ;
        RECT 2187.930 572.490 2189.110 573.670 ;
        RECT 2187.930 394.090 2189.110 395.270 ;
        RECT 2187.930 392.490 2189.110 393.670 ;
        RECT 2187.930 214.090 2189.110 215.270 ;
        RECT 2187.930 212.490 2189.110 213.670 ;
        RECT 2187.930 34.090 2189.110 35.270 ;
        RECT 2187.930 32.490 2189.110 33.670 ;
        RECT 2187.930 -12.310 2189.110 -11.130 ;
        RECT 2187.930 -13.910 2189.110 -12.730 ;
        RECT 2367.930 3532.410 2369.110 3533.590 ;
        RECT 2367.930 3530.810 2369.110 3531.990 ;
        RECT 2367.930 3454.090 2369.110 3455.270 ;
        RECT 2367.930 3452.490 2369.110 3453.670 ;
        RECT 2367.930 3274.090 2369.110 3275.270 ;
        RECT 2367.930 3272.490 2369.110 3273.670 ;
        RECT 2367.930 3094.090 2369.110 3095.270 ;
        RECT 2367.930 3092.490 2369.110 3093.670 ;
        RECT 2367.930 2914.090 2369.110 2915.270 ;
        RECT 2367.930 2912.490 2369.110 2913.670 ;
        RECT 2367.930 2734.090 2369.110 2735.270 ;
        RECT 2367.930 2732.490 2369.110 2733.670 ;
        RECT 2367.930 2554.090 2369.110 2555.270 ;
        RECT 2367.930 2552.490 2369.110 2553.670 ;
        RECT 2367.930 2374.090 2369.110 2375.270 ;
        RECT 2367.930 2372.490 2369.110 2373.670 ;
        RECT 2367.930 2194.090 2369.110 2195.270 ;
        RECT 2367.930 2192.490 2369.110 2193.670 ;
        RECT 2367.930 2014.090 2369.110 2015.270 ;
        RECT 2367.930 2012.490 2369.110 2013.670 ;
        RECT 2367.930 1834.090 2369.110 1835.270 ;
        RECT 2367.930 1832.490 2369.110 1833.670 ;
        RECT 2367.930 1654.090 2369.110 1655.270 ;
        RECT 2367.930 1652.490 2369.110 1653.670 ;
        RECT 2367.930 1474.090 2369.110 1475.270 ;
        RECT 2367.930 1472.490 2369.110 1473.670 ;
        RECT 2367.930 1294.090 2369.110 1295.270 ;
        RECT 2367.930 1292.490 2369.110 1293.670 ;
        RECT 2367.930 1114.090 2369.110 1115.270 ;
        RECT 2367.930 1112.490 2369.110 1113.670 ;
        RECT 2367.930 934.090 2369.110 935.270 ;
        RECT 2367.930 932.490 2369.110 933.670 ;
        RECT 2367.930 754.090 2369.110 755.270 ;
        RECT 2367.930 752.490 2369.110 753.670 ;
        RECT 2367.930 574.090 2369.110 575.270 ;
        RECT 2367.930 572.490 2369.110 573.670 ;
        RECT 2367.930 394.090 2369.110 395.270 ;
        RECT 2367.930 392.490 2369.110 393.670 ;
        RECT 2367.930 214.090 2369.110 215.270 ;
        RECT 2367.930 212.490 2369.110 213.670 ;
        RECT 2367.930 34.090 2369.110 35.270 ;
        RECT 2367.930 32.490 2369.110 33.670 ;
        RECT 2367.930 -12.310 2369.110 -11.130 ;
        RECT 2367.930 -13.910 2369.110 -12.730 ;
        RECT 2547.930 3532.410 2549.110 3533.590 ;
        RECT 2547.930 3530.810 2549.110 3531.990 ;
        RECT 2547.930 3454.090 2549.110 3455.270 ;
        RECT 2547.930 3452.490 2549.110 3453.670 ;
        RECT 2547.930 3274.090 2549.110 3275.270 ;
        RECT 2547.930 3272.490 2549.110 3273.670 ;
        RECT 2547.930 3094.090 2549.110 3095.270 ;
        RECT 2547.930 3092.490 2549.110 3093.670 ;
        RECT 2547.930 2914.090 2549.110 2915.270 ;
        RECT 2547.930 2912.490 2549.110 2913.670 ;
        RECT 2547.930 2734.090 2549.110 2735.270 ;
        RECT 2547.930 2732.490 2549.110 2733.670 ;
        RECT 2547.930 2554.090 2549.110 2555.270 ;
        RECT 2547.930 2552.490 2549.110 2553.670 ;
        RECT 2547.930 2374.090 2549.110 2375.270 ;
        RECT 2547.930 2372.490 2549.110 2373.670 ;
        RECT 2547.930 2194.090 2549.110 2195.270 ;
        RECT 2547.930 2192.490 2549.110 2193.670 ;
        RECT 2547.930 2014.090 2549.110 2015.270 ;
        RECT 2547.930 2012.490 2549.110 2013.670 ;
        RECT 2547.930 1834.090 2549.110 1835.270 ;
        RECT 2547.930 1832.490 2549.110 1833.670 ;
        RECT 2547.930 1654.090 2549.110 1655.270 ;
        RECT 2547.930 1652.490 2549.110 1653.670 ;
        RECT 2547.930 1474.090 2549.110 1475.270 ;
        RECT 2547.930 1472.490 2549.110 1473.670 ;
        RECT 2547.930 1294.090 2549.110 1295.270 ;
        RECT 2547.930 1292.490 2549.110 1293.670 ;
        RECT 2547.930 1114.090 2549.110 1115.270 ;
        RECT 2547.930 1112.490 2549.110 1113.670 ;
        RECT 2547.930 934.090 2549.110 935.270 ;
        RECT 2547.930 932.490 2549.110 933.670 ;
        RECT 2547.930 754.090 2549.110 755.270 ;
        RECT 2547.930 752.490 2549.110 753.670 ;
        RECT 2547.930 574.090 2549.110 575.270 ;
        RECT 2547.930 572.490 2549.110 573.670 ;
        RECT 2547.930 394.090 2549.110 395.270 ;
        RECT 2547.930 392.490 2549.110 393.670 ;
        RECT 2547.930 214.090 2549.110 215.270 ;
        RECT 2547.930 212.490 2549.110 213.670 ;
        RECT 2547.930 34.090 2549.110 35.270 ;
        RECT 2547.930 32.490 2549.110 33.670 ;
        RECT 2547.930 -12.310 2549.110 -11.130 ;
        RECT 2547.930 -13.910 2549.110 -12.730 ;
        RECT 2727.930 3532.410 2729.110 3533.590 ;
        RECT 2727.930 3530.810 2729.110 3531.990 ;
        RECT 2727.930 3454.090 2729.110 3455.270 ;
        RECT 2727.930 3452.490 2729.110 3453.670 ;
        RECT 2727.930 3274.090 2729.110 3275.270 ;
        RECT 2727.930 3272.490 2729.110 3273.670 ;
        RECT 2727.930 3094.090 2729.110 3095.270 ;
        RECT 2727.930 3092.490 2729.110 3093.670 ;
        RECT 2727.930 2914.090 2729.110 2915.270 ;
        RECT 2727.930 2912.490 2729.110 2913.670 ;
        RECT 2727.930 2734.090 2729.110 2735.270 ;
        RECT 2727.930 2732.490 2729.110 2733.670 ;
        RECT 2727.930 2554.090 2729.110 2555.270 ;
        RECT 2727.930 2552.490 2729.110 2553.670 ;
        RECT 2727.930 2374.090 2729.110 2375.270 ;
        RECT 2727.930 2372.490 2729.110 2373.670 ;
        RECT 2727.930 2194.090 2729.110 2195.270 ;
        RECT 2727.930 2192.490 2729.110 2193.670 ;
        RECT 2727.930 2014.090 2729.110 2015.270 ;
        RECT 2727.930 2012.490 2729.110 2013.670 ;
        RECT 2727.930 1834.090 2729.110 1835.270 ;
        RECT 2727.930 1832.490 2729.110 1833.670 ;
        RECT 2727.930 1654.090 2729.110 1655.270 ;
        RECT 2727.930 1652.490 2729.110 1653.670 ;
        RECT 2727.930 1474.090 2729.110 1475.270 ;
        RECT 2727.930 1472.490 2729.110 1473.670 ;
        RECT 2727.930 1294.090 2729.110 1295.270 ;
        RECT 2727.930 1292.490 2729.110 1293.670 ;
        RECT 2727.930 1114.090 2729.110 1115.270 ;
        RECT 2727.930 1112.490 2729.110 1113.670 ;
        RECT 2727.930 934.090 2729.110 935.270 ;
        RECT 2727.930 932.490 2729.110 933.670 ;
        RECT 2727.930 754.090 2729.110 755.270 ;
        RECT 2727.930 752.490 2729.110 753.670 ;
        RECT 2727.930 574.090 2729.110 575.270 ;
        RECT 2727.930 572.490 2729.110 573.670 ;
        RECT 2727.930 394.090 2729.110 395.270 ;
        RECT 2727.930 392.490 2729.110 393.670 ;
        RECT 2727.930 214.090 2729.110 215.270 ;
        RECT 2727.930 212.490 2729.110 213.670 ;
        RECT 2727.930 34.090 2729.110 35.270 ;
        RECT 2727.930 32.490 2729.110 33.670 ;
        RECT 2727.930 -12.310 2729.110 -11.130 ;
        RECT 2727.930 -13.910 2729.110 -12.730 ;
        RECT 2907.930 3532.410 2909.110 3533.590 ;
        RECT 2907.930 3530.810 2909.110 3531.990 ;
        RECT 2907.930 3454.090 2909.110 3455.270 ;
        RECT 2907.930 3452.490 2909.110 3453.670 ;
        RECT 2907.930 3274.090 2909.110 3275.270 ;
        RECT 2907.930 3272.490 2909.110 3273.670 ;
        RECT 2907.930 3094.090 2909.110 3095.270 ;
        RECT 2907.930 3092.490 2909.110 3093.670 ;
        RECT 2907.930 2914.090 2909.110 2915.270 ;
        RECT 2907.930 2912.490 2909.110 2913.670 ;
        RECT 2907.930 2734.090 2909.110 2735.270 ;
        RECT 2907.930 2732.490 2909.110 2733.670 ;
        RECT 2907.930 2554.090 2909.110 2555.270 ;
        RECT 2907.930 2552.490 2909.110 2553.670 ;
        RECT 2907.930 2374.090 2909.110 2375.270 ;
        RECT 2907.930 2372.490 2909.110 2373.670 ;
        RECT 2907.930 2194.090 2909.110 2195.270 ;
        RECT 2907.930 2192.490 2909.110 2193.670 ;
        RECT 2907.930 2014.090 2909.110 2015.270 ;
        RECT 2907.930 2012.490 2909.110 2013.670 ;
        RECT 2907.930 1834.090 2909.110 1835.270 ;
        RECT 2907.930 1832.490 2909.110 1833.670 ;
        RECT 2907.930 1654.090 2909.110 1655.270 ;
        RECT 2907.930 1652.490 2909.110 1653.670 ;
        RECT 2907.930 1474.090 2909.110 1475.270 ;
        RECT 2907.930 1472.490 2909.110 1473.670 ;
        RECT 2907.930 1294.090 2909.110 1295.270 ;
        RECT 2907.930 1292.490 2909.110 1293.670 ;
        RECT 2907.930 1114.090 2909.110 1115.270 ;
        RECT 2907.930 1112.490 2909.110 1113.670 ;
        RECT 2907.930 934.090 2909.110 935.270 ;
        RECT 2907.930 932.490 2909.110 933.670 ;
        RECT 2907.930 754.090 2909.110 755.270 ;
        RECT 2907.930 752.490 2909.110 753.670 ;
        RECT 2907.930 574.090 2909.110 575.270 ;
        RECT 2907.930 572.490 2909.110 573.670 ;
        RECT 2907.930 394.090 2909.110 395.270 ;
        RECT 2907.930 392.490 2909.110 393.670 ;
        RECT 2907.930 214.090 2909.110 215.270 ;
        RECT 2907.930 212.490 2909.110 213.670 ;
        RECT 2907.930 34.090 2909.110 35.270 ;
        RECT 2907.930 32.490 2909.110 33.670 ;
        RECT 2907.930 -12.310 2909.110 -11.130 ;
        RECT 2907.930 -13.910 2909.110 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 3454.090 2938.090 3455.270 ;
        RECT 2936.910 3452.490 2938.090 3453.670 ;
        RECT 2936.910 3274.090 2938.090 3275.270 ;
        RECT 2936.910 3272.490 2938.090 3273.670 ;
        RECT 2936.910 3094.090 2938.090 3095.270 ;
        RECT 2936.910 3092.490 2938.090 3093.670 ;
        RECT 2936.910 2914.090 2938.090 2915.270 ;
        RECT 2936.910 2912.490 2938.090 2913.670 ;
        RECT 2936.910 2734.090 2938.090 2735.270 ;
        RECT 2936.910 2732.490 2938.090 2733.670 ;
        RECT 2936.910 2554.090 2938.090 2555.270 ;
        RECT 2936.910 2552.490 2938.090 2553.670 ;
        RECT 2936.910 2374.090 2938.090 2375.270 ;
        RECT 2936.910 2372.490 2938.090 2373.670 ;
        RECT 2936.910 2194.090 2938.090 2195.270 ;
        RECT 2936.910 2192.490 2938.090 2193.670 ;
        RECT 2936.910 2014.090 2938.090 2015.270 ;
        RECT 2936.910 2012.490 2938.090 2013.670 ;
        RECT 2936.910 1834.090 2938.090 1835.270 ;
        RECT 2936.910 1832.490 2938.090 1833.670 ;
        RECT 2936.910 1654.090 2938.090 1655.270 ;
        RECT 2936.910 1652.490 2938.090 1653.670 ;
        RECT 2936.910 1474.090 2938.090 1475.270 ;
        RECT 2936.910 1472.490 2938.090 1473.670 ;
        RECT 2936.910 1294.090 2938.090 1295.270 ;
        RECT 2936.910 1292.490 2938.090 1293.670 ;
        RECT 2936.910 1114.090 2938.090 1115.270 ;
        RECT 2936.910 1112.490 2938.090 1113.670 ;
        RECT 2936.910 934.090 2938.090 935.270 ;
        RECT 2936.910 932.490 2938.090 933.670 ;
        RECT 2936.910 754.090 2938.090 755.270 ;
        RECT 2936.910 752.490 2938.090 753.670 ;
        RECT 2936.910 574.090 2938.090 575.270 ;
        RECT 2936.910 572.490 2938.090 573.670 ;
        RECT 2936.910 394.090 2938.090 395.270 ;
        RECT 2936.910 392.490 2938.090 393.670 ;
        RECT 2936.910 214.090 2938.090 215.270 ;
        RECT 2936.910 212.490 2938.090 213.670 ;
        RECT 2936.910 34.090 2938.090 35.270 ;
        RECT 2936.910 32.490 2938.090 33.670 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 27.020 3533.700 30.020 3533.710 ;
        RECT 207.020 3533.700 210.020 3533.710 ;
        RECT 387.020 3533.700 390.020 3533.710 ;
        RECT 567.020 3533.700 570.020 3533.710 ;
        RECT 747.020 3533.700 750.020 3533.710 ;
        RECT 927.020 3533.700 930.020 3533.710 ;
        RECT 1107.020 3533.700 1110.020 3533.710 ;
        RECT 1287.020 3533.700 1290.020 3533.710 ;
        RECT 1467.020 3533.700 1470.020 3533.710 ;
        RECT 1647.020 3533.700 1650.020 3533.710 ;
        RECT 1827.020 3533.700 1830.020 3533.710 ;
        RECT 2007.020 3533.700 2010.020 3533.710 ;
        RECT 2187.020 3533.700 2190.020 3533.710 ;
        RECT 2367.020 3533.700 2370.020 3533.710 ;
        RECT 2547.020 3533.700 2550.020 3533.710 ;
        RECT 2727.020 3533.700 2730.020 3533.710 ;
        RECT 2907.020 3533.700 2910.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 27.020 3530.690 30.020 3530.700 ;
        RECT 207.020 3530.690 210.020 3530.700 ;
        RECT 387.020 3530.690 390.020 3530.700 ;
        RECT 567.020 3530.690 570.020 3530.700 ;
        RECT 747.020 3530.690 750.020 3530.700 ;
        RECT 927.020 3530.690 930.020 3530.700 ;
        RECT 1107.020 3530.690 1110.020 3530.700 ;
        RECT 1287.020 3530.690 1290.020 3530.700 ;
        RECT 1467.020 3530.690 1470.020 3530.700 ;
        RECT 1647.020 3530.690 1650.020 3530.700 ;
        RECT 1827.020 3530.690 1830.020 3530.700 ;
        RECT 2007.020 3530.690 2010.020 3530.700 ;
        RECT 2187.020 3530.690 2190.020 3530.700 ;
        RECT 2367.020 3530.690 2370.020 3530.700 ;
        RECT 2547.020 3530.690 2550.020 3530.700 ;
        RECT 2727.020 3530.690 2730.020 3530.700 ;
        RECT 2907.020 3530.690 2910.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3455.380 -16.380 3455.390 ;
        RECT 27.020 3455.380 30.020 3455.390 ;
        RECT 207.020 3455.380 210.020 3455.390 ;
        RECT 387.020 3455.380 390.020 3455.390 ;
        RECT 567.020 3455.380 570.020 3455.390 ;
        RECT 747.020 3455.380 750.020 3455.390 ;
        RECT 927.020 3455.380 930.020 3455.390 ;
        RECT 1107.020 3455.380 1110.020 3455.390 ;
        RECT 1287.020 3455.380 1290.020 3455.390 ;
        RECT 1467.020 3455.380 1470.020 3455.390 ;
        RECT 1647.020 3455.380 1650.020 3455.390 ;
        RECT 1827.020 3455.380 1830.020 3455.390 ;
        RECT 2007.020 3455.380 2010.020 3455.390 ;
        RECT 2187.020 3455.380 2190.020 3455.390 ;
        RECT 2367.020 3455.380 2370.020 3455.390 ;
        RECT 2547.020 3455.380 2550.020 3455.390 ;
        RECT 2727.020 3455.380 2730.020 3455.390 ;
        RECT 2907.020 3455.380 2910.020 3455.390 ;
        RECT 2936.000 3455.380 2939.000 3455.390 ;
        RECT -24.080 3452.380 2943.700 3455.380 ;
        RECT -19.380 3452.370 -16.380 3452.380 ;
        RECT 27.020 3452.370 30.020 3452.380 ;
        RECT 207.020 3452.370 210.020 3452.380 ;
        RECT 387.020 3452.370 390.020 3452.380 ;
        RECT 567.020 3452.370 570.020 3452.380 ;
        RECT 747.020 3452.370 750.020 3452.380 ;
        RECT 927.020 3452.370 930.020 3452.380 ;
        RECT 1107.020 3452.370 1110.020 3452.380 ;
        RECT 1287.020 3452.370 1290.020 3452.380 ;
        RECT 1467.020 3452.370 1470.020 3452.380 ;
        RECT 1647.020 3452.370 1650.020 3452.380 ;
        RECT 1827.020 3452.370 1830.020 3452.380 ;
        RECT 2007.020 3452.370 2010.020 3452.380 ;
        RECT 2187.020 3452.370 2190.020 3452.380 ;
        RECT 2367.020 3452.370 2370.020 3452.380 ;
        RECT 2547.020 3452.370 2550.020 3452.380 ;
        RECT 2727.020 3452.370 2730.020 3452.380 ;
        RECT 2907.020 3452.370 2910.020 3452.380 ;
        RECT 2936.000 3452.370 2939.000 3452.380 ;
        RECT -19.380 3275.380 -16.380 3275.390 ;
        RECT 27.020 3275.380 30.020 3275.390 ;
        RECT 207.020 3275.380 210.020 3275.390 ;
        RECT 387.020 3275.380 390.020 3275.390 ;
        RECT 567.020 3275.380 570.020 3275.390 ;
        RECT 747.020 3275.380 750.020 3275.390 ;
        RECT 927.020 3275.380 930.020 3275.390 ;
        RECT 1107.020 3275.380 1110.020 3275.390 ;
        RECT 1287.020 3275.380 1290.020 3275.390 ;
        RECT 1467.020 3275.380 1470.020 3275.390 ;
        RECT 1647.020 3275.380 1650.020 3275.390 ;
        RECT 1827.020 3275.380 1830.020 3275.390 ;
        RECT 2007.020 3275.380 2010.020 3275.390 ;
        RECT 2187.020 3275.380 2190.020 3275.390 ;
        RECT 2367.020 3275.380 2370.020 3275.390 ;
        RECT 2547.020 3275.380 2550.020 3275.390 ;
        RECT 2727.020 3275.380 2730.020 3275.390 ;
        RECT 2907.020 3275.380 2910.020 3275.390 ;
        RECT 2936.000 3275.380 2939.000 3275.390 ;
        RECT -24.080 3272.380 2943.700 3275.380 ;
        RECT -19.380 3272.370 -16.380 3272.380 ;
        RECT 27.020 3272.370 30.020 3272.380 ;
        RECT 207.020 3272.370 210.020 3272.380 ;
        RECT 387.020 3272.370 390.020 3272.380 ;
        RECT 567.020 3272.370 570.020 3272.380 ;
        RECT 747.020 3272.370 750.020 3272.380 ;
        RECT 927.020 3272.370 930.020 3272.380 ;
        RECT 1107.020 3272.370 1110.020 3272.380 ;
        RECT 1287.020 3272.370 1290.020 3272.380 ;
        RECT 1467.020 3272.370 1470.020 3272.380 ;
        RECT 1647.020 3272.370 1650.020 3272.380 ;
        RECT 1827.020 3272.370 1830.020 3272.380 ;
        RECT 2007.020 3272.370 2010.020 3272.380 ;
        RECT 2187.020 3272.370 2190.020 3272.380 ;
        RECT 2367.020 3272.370 2370.020 3272.380 ;
        RECT 2547.020 3272.370 2550.020 3272.380 ;
        RECT 2727.020 3272.370 2730.020 3272.380 ;
        RECT 2907.020 3272.370 2910.020 3272.380 ;
        RECT 2936.000 3272.370 2939.000 3272.380 ;
        RECT -19.380 3095.380 -16.380 3095.390 ;
        RECT 27.020 3095.380 30.020 3095.390 ;
        RECT 207.020 3095.380 210.020 3095.390 ;
        RECT 387.020 3095.380 390.020 3095.390 ;
        RECT 567.020 3095.380 570.020 3095.390 ;
        RECT 747.020 3095.380 750.020 3095.390 ;
        RECT 927.020 3095.380 930.020 3095.390 ;
        RECT 1107.020 3095.380 1110.020 3095.390 ;
        RECT 1287.020 3095.380 1290.020 3095.390 ;
        RECT 1467.020 3095.380 1470.020 3095.390 ;
        RECT 1647.020 3095.380 1650.020 3095.390 ;
        RECT 1827.020 3095.380 1830.020 3095.390 ;
        RECT 2007.020 3095.380 2010.020 3095.390 ;
        RECT 2187.020 3095.380 2190.020 3095.390 ;
        RECT 2367.020 3095.380 2370.020 3095.390 ;
        RECT 2547.020 3095.380 2550.020 3095.390 ;
        RECT 2727.020 3095.380 2730.020 3095.390 ;
        RECT 2907.020 3095.380 2910.020 3095.390 ;
        RECT 2936.000 3095.380 2939.000 3095.390 ;
        RECT -24.080 3092.380 2943.700 3095.380 ;
        RECT -19.380 3092.370 -16.380 3092.380 ;
        RECT 27.020 3092.370 30.020 3092.380 ;
        RECT 207.020 3092.370 210.020 3092.380 ;
        RECT 387.020 3092.370 390.020 3092.380 ;
        RECT 567.020 3092.370 570.020 3092.380 ;
        RECT 747.020 3092.370 750.020 3092.380 ;
        RECT 927.020 3092.370 930.020 3092.380 ;
        RECT 1107.020 3092.370 1110.020 3092.380 ;
        RECT 1287.020 3092.370 1290.020 3092.380 ;
        RECT 1467.020 3092.370 1470.020 3092.380 ;
        RECT 1647.020 3092.370 1650.020 3092.380 ;
        RECT 1827.020 3092.370 1830.020 3092.380 ;
        RECT 2007.020 3092.370 2010.020 3092.380 ;
        RECT 2187.020 3092.370 2190.020 3092.380 ;
        RECT 2367.020 3092.370 2370.020 3092.380 ;
        RECT 2547.020 3092.370 2550.020 3092.380 ;
        RECT 2727.020 3092.370 2730.020 3092.380 ;
        RECT 2907.020 3092.370 2910.020 3092.380 ;
        RECT 2936.000 3092.370 2939.000 3092.380 ;
        RECT -19.380 2915.380 -16.380 2915.390 ;
        RECT 27.020 2915.380 30.020 2915.390 ;
        RECT 207.020 2915.380 210.020 2915.390 ;
        RECT 387.020 2915.380 390.020 2915.390 ;
        RECT 567.020 2915.380 570.020 2915.390 ;
        RECT 747.020 2915.380 750.020 2915.390 ;
        RECT 927.020 2915.380 930.020 2915.390 ;
        RECT 1107.020 2915.380 1110.020 2915.390 ;
        RECT 1287.020 2915.380 1290.020 2915.390 ;
        RECT 1467.020 2915.380 1470.020 2915.390 ;
        RECT 1647.020 2915.380 1650.020 2915.390 ;
        RECT 1827.020 2915.380 1830.020 2915.390 ;
        RECT 2007.020 2915.380 2010.020 2915.390 ;
        RECT 2187.020 2915.380 2190.020 2915.390 ;
        RECT 2367.020 2915.380 2370.020 2915.390 ;
        RECT 2547.020 2915.380 2550.020 2915.390 ;
        RECT 2727.020 2915.380 2730.020 2915.390 ;
        RECT 2907.020 2915.380 2910.020 2915.390 ;
        RECT 2936.000 2915.380 2939.000 2915.390 ;
        RECT -24.080 2912.380 2943.700 2915.380 ;
        RECT -19.380 2912.370 -16.380 2912.380 ;
        RECT 27.020 2912.370 30.020 2912.380 ;
        RECT 207.020 2912.370 210.020 2912.380 ;
        RECT 387.020 2912.370 390.020 2912.380 ;
        RECT 567.020 2912.370 570.020 2912.380 ;
        RECT 747.020 2912.370 750.020 2912.380 ;
        RECT 927.020 2912.370 930.020 2912.380 ;
        RECT 1107.020 2912.370 1110.020 2912.380 ;
        RECT 1287.020 2912.370 1290.020 2912.380 ;
        RECT 1467.020 2912.370 1470.020 2912.380 ;
        RECT 1647.020 2912.370 1650.020 2912.380 ;
        RECT 1827.020 2912.370 1830.020 2912.380 ;
        RECT 2007.020 2912.370 2010.020 2912.380 ;
        RECT 2187.020 2912.370 2190.020 2912.380 ;
        RECT 2367.020 2912.370 2370.020 2912.380 ;
        RECT 2547.020 2912.370 2550.020 2912.380 ;
        RECT 2727.020 2912.370 2730.020 2912.380 ;
        RECT 2907.020 2912.370 2910.020 2912.380 ;
        RECT 2936.000 2912.370 2939.000 2912.380 ;
        RECT -19.380 2735.380 -16.380 2735.390 ;
        RECT 27.020 2735.380 30.020 2735.390 ;
        RECT 207.020 2735.380 210.020 2735.390 ;
        RECT 387.020 2735.380 390.020 2735.390 ;
        RECT 567.020 2735.380 570.020 2735.390 ;
        RECT 747.020 2735.380 750.020 2735.390 ;
        RECT 927.020 2735.380 930.020 2735.390 ;
        RECT 1107.020 2735.380 1110.020 2735.390 ;
        RECT 1287.020 2735.380 1290.020 2735.390 ;
        RECT 1467.020 2735.380 1470.020 2735.390 ;
        RECT 1647.020 2735.380 1650.020 2735.390 ;
        RECT 1827.020 2735.380 1830.020 2735.390 ;
        RECT 2007.020 2735.380 2010.020 2735.390 ;
        RECT 2187.020 2735.380 2190.020 2735.390 ;
        RECT 2367.020 2735.380 2370.020 2735.390 ;
        RECT 2547.020 2735.380 2550.020 2735.390 ;
        RECT 2727.020 2735.380 2730.020 2735.390 ;
        RECT 2907.020 2735.380 2910.020 2735.390 ;
        RECT 2936.000 2735.380 2939.000 2735.390 ;
        RECT -24.080 2732.380 2943.700 2735.380 ;
        RECT -19.380 2732.370 -16.380 2732.380 ;
        RECT 27.020 2732.370 30.020 2732.380 ;
        RECT 207.020 2732.370 210.020 2732.380 ;
        RECT 387.020 2732.370 390.020 2732.380 ;
        RECT 567.020 2732.370 570.020 2732.380 ;
        RECT 747.020 2732.370 750.020 2732.380 ;
        RECT 927.020 2732.370 930.020 2732.380 ;
        RECT 1107.020 2732.370 1110.020 2732.380 ;
        RECT 1287.020 2732.370 1290.020 2732.380 ;
        RECT 1467.020 2732.370 1470.020 2732.380 ;
        RECT 1647.020 2732.370 1650.020 2732.380 ;
        RECT 1827.020 2732.370 1830.020 2732.380 ;
        RECT 2007.020 2732.370 2010.020 2732.380 ;
        RECT 2187.020 2732.370 2190.020 2732.380 ;
        RECT 2367.020 2732.370 2370.020 2732.380 ;
        RECT 2547.020 2732.370 2550.020 2732.380 ;
        RECT 2727.020 2732.370 2730.020 2732.380 ;
        RECT 2907.020 2732.370 2910.020 2732.380 ;
        RECT 2936.000 2732.370 2939.000 2732.380 ;
        RECT -19.380 2555.380 -16.380 2555.390 ;
        RECT 27.020 2555.380 30.020 2555.390 ;
        RECT 207.020 2555.380 210.020 2555.390 ;
        RECT 387.020 2555.380 390.020 2555.390 ;
        RECT 567.020 2555.380 570.020 2555.390 ;
        RECT 747.020 2555.380 750.020 2555.390 ;
        RECT 927.020 2555.380 930.020 2555.390 ;
        RECT 1107.020 2555.380 1110.020 2555.390 ;
        RECT 1287.020 2555.380 1290.020 2555.390 ;
        RECT 1467.020 2555.380 1470.020 2555.390 ;
        RECT 1647.020 2555.380 1650.020 2555.390 ;
        RECT 1827.020 2555.380 1830.020 2555.390 ;
        RECT 2007.020 2555.380 2010.020 2555.390 ;
        RECT 2187.020 2555.380 2190.020 2555.390 ;
        RECT 2367.020 2555.380 2370.020 2555.390 ;
        RECT 2547.020 2555.380 2550.020 2555.390 ;
        RECT 2727.020 2555.380 2730.020 2555.390 ;
        RECT 2907.020 2555.380 2910.020 2555.390 ;
        RECT 2936.000 2555.380 2939.000 2555.390 ;
        RECT -24.080 2552.380 2943.700 2555.380 ;
        RECT -19.380 2552.370 -16.380 2552.380 ;
        RECT 27.020 2552.370 30.020 2552.380 ;
        RECT 207.020 2552.370 210.020 2552.380 ;
        RECT 387.020 2552.370 390.020 2552.380 ;
        RECT 567.020 2552.370 570.020 2552.380 ;
        RECT 747.020 2552.370 750.020 2552.380 ;
        RECT 927.020 2552.370 930.020 2552.380 ;
        RECT 1107.020 2552.370 1110.020 2552.380 ;
        RECT 1287.020 2552.370 1290.020 2552.380 ;
        RECT 1467.020 2552.370 1470.020 2552.380 ;
        RECT 1647.020 2552.370 1650.020 2552.380 ;
        RECT 1827.020 2552.370 1830.020 2552.380 ;
        RECT 2007.020 2552.370 2010.020 2552.380 ;
        RECT 2187.020 2552.370 2190.020 2552.380 ;
        RECT 2367.020 2552.370 2370.020 2552.380 ;
        RECT 2547.020 2552.370 2550.020 2552.380 ;
        RECT 2727.020 2552.370 2730.020 2552.380 ;
        RECT 2907.020 2552.370 2910.020 2552.380 ;
        RECT 2936.000 2552.370 2939.000 2552.380 ;
        RECT -19.380 2375.380 -16.380 2375.390 ;
        RECT 27.020 2375.380 30.020 2375.390 ;
        RECT 207.020 2375.380 210.020 2375.390 ;
        RECT 387.020 2375.380 390.020 2375.390 ;
        RECT 567.020 2375.380 570.020 2375.390 ;
        RECT 747.020 2375.380 750.020 2375.390 ;
        RECT 927.020 2375.380 930.020 2375.390 ;
        RECT 1107.020 2375.380 1110.020 2375.390 ;
        RECT 1287.020 2375.380 1290.020 2375.390 ;
        RECT 1467.020 2375.380 1470.020 2375.390 ;
        RECT 1647.020 2375.380 1650.020 2375.390 ;
        RECT 1827.020 2375.380 1830.020 2375.390 ;
        RECT 2007.020 2375.380 2010.020 2375.390 ;
        RECT 2187.020 2375.380 2190.020 2375.390 ;
        RECT 2367.020 2375.380 2370.020 2375.390 ;
        RECT 2547.020 2375.380 2550.020 2375.390 ;
        RECT 2727.020 2375.380 2730.020 2375.390 ;
        RECT 2907.020 2375.380 2910.020 2375.390 ;
        RECT 2936.000 2375.380 2939.000 2375.390 ;
        RECT -24.080 2372.380 2943.700 2375.380 ;
        RECT -19.380 2372.370 -16.380 2372.380 ;
        RECT 27.020 2372.370 30.020 2372.380 ;
        RECT 207.020 2372.370 210.020 2372.380 ;
        RECT 387.020 2372.370 390.020 2372.380 ;
        RECT 567.020 2372.370 570.020 2372.380 ;
        RECT 747.020 2372.370 750.020 2372.380 ;
        RECT 927.020 2372.370 930.020 2372.380 ;
        RECT 1107.020 2372.370 1110.020 2372.380 ;
        RECT 1287.020 2372.370 1290.020 2372.380 ;
        RECT 1467.020 2372.370 1470.020 2372.380 ;
        RECT 1647.020 2372.370 1650.020 2372.380 ;
        RECT 1827.020 2372.370 1830.020 2372.380 ;
        RECT 2007.020 2372.370 2010.020 2372.380 ;
        RECT 2187.020 2372.370 2190.020 2372.380 ;
        RECT 2367.020 2372.370 2370.020 2372.380 ;
        RECT 2547.020 2372.370 2550.020 2372.380 ;
        RECT 2727.020 2372.370 2730.020 2372.380 ;
        RECT 2907.020 2372.370 2910.020 2372.380 ;
        RECT 2936.000 2372.370 2939.000 2372.380 ;
        RECT -19.380 2195.380 -16.380 2195.390 ;
        RECT 27.020 2195.380 30.020 2195.390 ;
        RECT 207.020 2195.380 210.020 2195.390 ;
        RECT 387.020 2195.380 390.020 2195.390 ;
        RECT 567.020 2195.380 570.020 2195.390 ;
        RECT 747.020 2195.380 750.020 2195.390 ;
        RECT 927.020 2195.380 930.020 2195.390 ;
        RECT 1107.020 2195.380 1110.020 2195.390 ;
        RECT 1287.020 2195.380 1290.020 2195.390 ;
        RECT 1467.020 2195.380 1470.020 2195.390 ;
        RECT 1647.020 2195.380 1650.020 2195.390 ;
        RECT 1827.020 2195.380 1830.020 2195.390 ;
        RECT 2007.020 2195.380 2010.020 2195.390 ;
        RECT 2187.020 2195.380 2190.020 2195.390 ;
        RECT 2367.020 2195.380 2370.020 2195.390 ;
        RECT 2547.020 2195.380 2550.020 2195.390 ;
        RECT 2727.020 2195.380 2730.020 2195.390 ;
        RECT 2907.020 2195.380 2910.020 2195.390 ;
        RECT 2936.000 2195.380 2939.000 2195.390 ;
        RECT -24.080 2192.380 2943.700 2195.380 ;
        RECT -19.380 2192.370 -16.380 2192.380 ;
        RECT 27.020 2192.370 30.020 2192.380 ;
        RECT 207.020 2192.370 210.020 2192.380 ;
        RECT 387.020 2192.370 390.020 2192.380 ;
        RECT 567.020 2192.370 570.020 2192.380 ;
        RECT 747.020 2192.370 750.020 2192.380 ;
        RECT 927.020 2192.370 930.020 2192.380 ;
        RECT 1107.020 2192.370 1110.020 2192.380 ;
        RECT 1287.020 2192.370 1290.020 2192.380 ;
        RECT 1467.020 2192.370 1470.020 2192.380 ;
        RECT 1647.020 2192.370 1650.020 2192.380 ;
        RECT 1827.020 2192.370 1830.020 2192.380 ;
        RECT 2007.020 2192.370 2010.020 2192.380 ;
        RECT 2187.020 2192.370 2190.020 2192.380 ;
        RECT 2367.020 2192.370 2370.020 2192.380 ;
        RECT 2547.020 2192.370 2550.020 2192.380 ;
        RECT 2727.020 2192.370 2730.020 2192.380 ;
        RECT 2907.020 2192.370 2910.020 2192.380 ;
        RECT 2936.000 2192.370 2939.000 2192.380 ;
        RECT -19.380 2015.380 -16.380 2015.390 ;
        RECT 27.020 2015.380 30.020 2015.390 ;
        RECT 207.020 2015.380 210.020 2015.390 ;
        RECT 387.020 2015.380 390.020 2015.390 ;
        RECT 567.020 2015.380 570.020 2015.390 ;
        RECT 747.020 2015.380 750.020 2015.390 ;
        RECT 927.020 2015.380 930.020 2015.390 ;
        RECT 1107.020 2015.380 1110.020 2015.390 ;
        RECT 1287.020 2015.380 1290.020 2015.390 ;
        RECT 1467.020 2015.380 1470.020 2015.390 ;
        RECT 1647.020 2015.380 1650.020 2015.390 ;
        RECT 1827.020 2015.380 1830.020 2015.390 ;
        RECT 2007.020 2015.380 2010.020 2015.390 ;
        RECT 2187.020 2015.380 2190.020 2015.390 ;
        RECT 2367.020 2015.380 2370.020 2015.390 ;
        RECT 2547.020 2015.380 2550.020 2015.390 ;
        RECT 2727.020 2015.380 2730.020 2015.390 ;
        RECT 2907.020 2015.380 2910.020 2015.390 ;
        RECT 2936.000 2015.380 2939.000 2015.390 ;
        RECT -24.080 2012.380 2943.700 2015.380 ;
        RECT -19.380 2012.370 -16.380 2012.380 ;
        RECT 27.020 2012.370 30.020 2012.380 ;
        RECT 207.020 2012.370 210.020 2012.380 ;
        RECT 387.020 2012.370 390.020 2012.380 ;
        RECT 567.020 2012.370 570.020 2012.380 ;
        RECT 747.020 2012.370 750.020 2012.380 ;
        RECT 927.020 2012.370 930.020 2012.380 ;
        RECT 1107.020 2012.370 1110.020 2012.380 ;
        RECT 1287.020 2012.370 1290.020 2012.380 ;
        RECT 1467.020 2012.370 1470.020 2012.380 ;
        RECT 1647.020 2012.370 1650.020 2012.380 ;
        RECT 1827.020 2012.370 1830.020 2012.380 ;
        RECT 2007.020 2012.370 2010.020 2012.380 ;
        RECT 2187.020 2012.370 2190.020 2012.380 ;
        RECT 2367.020 2012.370 2370.020 2012.380 ;
        RECT 2547.020 2012.370 2550.020 2012.380 ;
        RECT 2727.020 2012.370 2730.020 2012.380 ;
        RECT 2907.020 2012.370 2910.020 2012.380 ;
        RECT 2936.000 2012.370 2939.000 2012.380 ;
        RECT -19.380 1835.380 -16.380 1835.390 ;
        RECT 27.020 1835.380 30.020 1835.390 ;
        RECT 207.020 1835.380 210.020 1835.390 ;
        RECT 387.020 1835.380 390.020 1835.390 ;
        RECT 567.020 1835.380 570.020 1835.390 ;
        RECT 747.020 1835.380 750.020 1835.390 ;
        RECT 927.020 1835.380 930.020 1835.390 ;
        RECT 1107.020 1835.380 1110.020 1835.390 ;
        RECT 1287.020 1835.380 1290.020 1835.390 ;
        RECT 1467.020 1835.380 1470.020 1835.390 ;
        RECT 1647.020 1835.380 1650.020 1835.390 ;
        RECT 1827.020 1835.380 1830.020 1835.390 ;
        RECT 2007.020 1835.380 2010.020 1835.390 ;
        RECT 2187.020 1835.380 2190.020 1835.390 ;
        RECT 2367.020 1835.380 2370.020 1835.390 ;
        RECT 2547.020 1835.380 2550.020 1835.390 ;
        RECT 2727.020 1835.380 2730.020 1835.390 ;
        RECT 2907.020 1835.380 2910.020 1835.390 ;
        RECT 2936.000 1835.380 2939.000 1835.390 ;
        RECT -24.080 1832.380 2943.700 1835.380 ;
        RECT -19.380 1832.370 -16.380 1832.380 ;
        RECT 27.020 1832.370 30.020 1832.380 ;
        RECT 207.020 1832.370 210.020 1832.380 ;
        RECT 387.020 1832.370 390.020 1832.380 ;
        RECT 567.020 1832.370 570.020 1832.380 ;
        RECT 747.020 1832.370 750.020 1832.380 ;
        RECT 927.020 1832.370 930.020 1832.380 ;
        RECT 1107.020 1832.370 1110.020 1832.380 ;
        RECT 1287.020 1832.370 1290.020 1832.380 ;
        RECT 1467.020 1832.370 1470.020 1832.380 ;
        RECT 1647.020 1832.370 1650.020 1832.380 ;
        RECT 1827.020 1832.370 1830.020 1832.380 ;
        RECT 2007.020 1832.370 2010.020 1832.380 ;
        RECT 2187.020 1832.370 2190.020 1832.380 ;
        RECT 2367.020 1832.370 2370.020 1832.380 ;
        RECT 2547.020 1832.370 2550.020 1832.380 ;
        RECT 2727.020 1832.370 2730.020 1832.380 ;
        RECT 2907.020 1832.370 2910.020 1832.380 ;
        RECT 2936.000 1832.370 2939.000 1832.380 ;
        RECT -19.380 1655.380 -16.380 1655.390 ;
        RECT 27.020 1655.380 30.020 1655.390 ;
        RECT 207.020 1655.380 210.020 1655.390 ;
        RECT 387.020 1655.380 390.020 1655.390 ;
        RECT 567.020 1655.380 570.020 1655.390 ;
        RECT 747.020 1655.380 750.020 1655.390 ;
        RECT 927.020 1655.380 930.020 1655.390 ;
        RECT 1107.020 1655.380 1110.020 1655.390 ;
        RECT 1287.020 1655.380 1290.020 1655.390 ;
        RECT 1467.020 1655.380 1470.020 1655.390 ;
        RECT 1647.020 1655.380 1650.020 1655.390 ;
        RECT 1827.020 1655.380 1830.020 1655.390 ;
        RECT 2007.020 1655.380 2010.020 1655.390 ;
        RECT 2187.020 1655.380 2190.020 1655.390 ;
        RECT 2367.020 1655.380 2370.020 1655.390 ;
        RECT 2547.020 1655.380 2550.020 1655.390 ;
        RECT 2727.020 1655.380 2730.020 1655.390 ;
        RECT 2907.020 1655.380 2910.020 1655.390 ;
        RECT 2936.000 1655.380 2939.000 1655.390 ;
        RECT -24.080 1652.380 2943.700 1655.380 ;
        RECT -19.380 1652.370 -16.380 1652.380 ;
        RECT 27.020 1652.370 30.020 1652.380 ;
        RECT 207.020 1652.370 210.020 1652.380 ;
        RECT 387.020 1652.370 390.020 1652.380 ;
        RECT 567.020 1652.370 570.020 1652.380 ;
        RECT 747.020 1652.370 750.020 1652.380 ;
        RECT 927.020 1652.370 930.020 1652.380 ;
        RECT 1107.020 1652.370 1110.020 1652.380 ;
        RECT 1287.020 1652.370 1290.020 1652.380 ;
        RECT 1467.020 1652.370 1470.020 1652.380 ;
        RECT 1647.020 1652.370 1650.020 1652.380 ;
        RECT 1827.020 1652.370 1830.020 1652.380 ;
        RECT 2007.020 1652.370 2010.020 1652.380 ;
        RECT 2187.020 1652.370 2190.020 1652.380 ;
        RECT 2367.020 1652.370 2370.020 1652.380 ;
        RECT 2547.020 1652.370 2550.020 1652.380 ;
        RECT 2727.020 1652.370 2730.020 1652.380 ;
        RECT 2907.020 1652.370 2910.020 1652.380 ;
        RECT 2936.000 1652.370 2939.000 1652.380 ;
        RECT -19.380 1475.380 -16.380 1475.390 ;
        RECT 27.020 1475.380 30.020 1475.390 ;
        RECT 207.020 1475.380 210.020 1475.390 ;
        RECT 387.020 1475.380 390.020 1475.390 ;
        RECT 567.020 1475.380 570.020 1475.390 ;
        RECT 747.020 1475.380 750.020 1475.390 ;
        RECT 927.020 1475.380 930.020 1475.390 ;
        RECT 1107.020 1475.380 1110.020 1475.390 ;
        RECT 1287.020 1475.380 1290.020 1475.390 ;
        RECT 1467.020 1475.380 1470.020 1475.390 ;
        RECT 1647.020 1475.380 1650.020 1475.390 ;
        RECT 1827.020 1475.380 1830.020 1475.390 ;
        RECT 2007.020 1475.380 2010.020 1475.390 ;
        RECT 2187.020 1475.380 2190.020 1475.390 ;
        RECT 2367.020 1475.380 2370.020 1475.390 ;
        RECT 2547.020 1475.380 2550.020 1475.390 ;
        RECT 2727.020 1475.380 2730.020 1475.390 ;
        RECT 2907.020 1475.380 2910.020 1475.390 ;
        RECT 2936.000 1475.380 2939.000 1475.390 ;
        RECT -24.080 1472.380 2943.700 1475.380 ;
        RECT -19.380 1472.370 -16.380 1472.380 ;
        RECT 27.020 1472.370 30.020 1472.380 ;
        RECT 207.020 1472.370 210.020 1472.380 ;
        RECT 387.020 1472.370 390.020 1472.380 ;
        RECT 567.020 1472.370 570.020 1472.380 ;
        RECT 747.020 1472.370 750.020 1472.380 ;
        RECT 927.020 1472.370 930.020 1472.380 ;
        RECT 1107.020 1472.370 1110.020 1472.380 ;
        RECT 1287.020 1472.370 1290.020 1472.380 ;
        RECT 1467.020 1472.370 1470.020 1472.380 ;
        RECT 1647.020 1472.370 1650.020 1472.380 ;
        RECT 1827.020 1472.370 1830.020 1472.380 ;
        RECT 2007.020 1472.370 2010.020 1472.380 ;
        RECT 2187.020 1472.370 2190.020 1472.380 ;
        RECT 2367.020 1472.370 2370.020 1472.380 ;
        RECT 2547.020 1472.370 2550.020 1472.380 ;
        RECT 2727.020 1472.370 2730.020 1472.380 ;
        RECT 2907.020 1472.370 2910.020 1472.380 ;
        RECT 2936.000 1472.370 2939.000 1472.380 ;
        RECT -19.380 1295.380 -16.380 1295.390 ;
        RECT 27.020 1295.380 30.020 1295.390 ;
        RECT 207.020 1295.380 210.020 1295.390 ;
        RECT 387.020 1295.380 390.020 1295.390 ;
        RECT 567.020 1295.380 570.020 1295.390 ;
        RECT 747.020 1295.380 750.020 1295.390 ;
        RECT 927.020 1295.380 930.020 1295.390 ;
        RECT 1107.020 1295.380 1110.020 1295.390 ;
        RECT 1287.020 1295.380 1290.020 1295.390 ;
        RECT 1467.020 1295.380 1470.020 1295.390 ;
        RECT 1647.020 1295.380 1650.020 1295.390 ;
        RECT 1827.020 1295.380 1830.020 1295.390 ;
        RECT 2007.020 1295.380 2010.020 1295.390 ;
        RECT 2187.020 1295.380 2190.020 1295.390 ;
        RECT 2367.020 1295.380 2370.020 1295.390 ;
        RECT 2547.020 1295.380 2550.020 1295.390 ;
        RECT 2727.020 1295.380 2730.020 1295.390 ;
        RECT 2907.020 1295.380 2910.020 1295.390 ;
        RECT 2936.000 1295.380 2939.000 1295.390 ;
        RECT -24.080 1292.380 2943.700 1295.380 ;
        RECT -19.380 1292.370 -16.380 1292.380 ;
        RECT 27.020 1292.370 30.020 1292.380 ;
        RECT 207.020 1292.370 210.020 1292.380 ;
        RECT 387.020 1292.370 390.020 1292.380 ;
        RECT 567.020 1292.370 570.020 1292.380 ;
        RECT 747.020 1292.370 750.020 1292.380 ;
        RECT 927.020 1292.370 930.020 1292.380 ;
        RECT 1107.020 1292.370 1110.020 1292.380 ;
        RECT 1287.020 1292.370 1290.020 1292.380 ;
        RECT 1467.020 1292.370 1470.020 1292.380 ;
        RECT 1647.020 1292.370 1650.020 1292.380 ;
        RECT 1827.020 1292.370 1830.020 1292.380 ;
        RECT 2007.020 1292.370 2010.020 1292.380 ;
        RECT 2187.020 1292.370 2190.020 1292.380 ;
        RECT 2367.020 1292.370 2370.020 1292.380 ;
        RECT 2547.020 1292.370 2550.020 1292.380 ;
        RECT 2727.020 1292.370 2730.020 1292.380 ;
        RECT 2907.020 1292.370 2910.020 1292.380 ;
        RECT 2936.000 1292.370 2939.000 1292.380 ;
        RECT -19.380 1115.380 -16.380 1115.390 ;
        RECT 27.020 1115.380 30.020 1115.390 ;
        RECT 207.020 1115.380 210.020 1115.390 ;
        RECT 387.020 1115.380 390.020 1115.390 ;
        RECT 567.020 1115.380 570.020 1115.390 ;
        RECT 747.020 1115.380 750.020 1115.390 ;
        RECT 927.020 1115.380 930.020 1115.390 ;
        RECT 1107.020 1115.380 1110.020 1115.390 ;
        RECT 1287.020 1115.380 1290.020 1115.390 ;
        RECT 1467.020 1115.380 1470.020 1115.390 ;
        RECT 1647.020 1115.380 1650.020 1115.390 ;
        RECT 1827.020 1115.380 1830.020 1115.390 ;
        RECT 2007.020 1115.380 2010.020 1115.390 ;
        RECT 2187.020 1115.380 2190.020 1115.390 ;
        RECT 2367.020 1115.380 2370.020 1115.390 ;
        RECT 2547.020 1115.380 2550.020 1115.390 ;
        RECT 2727.020 1115.380 2730.020 1115.390 ;
        RECT 2907.020 1115.380 2910.020 1115.390 ;
        RECT 2936.000 1115.380 2939.000 1115.390 ;
        RECT -24.080 1112.380 2943.700 1115.380 ;
        RECT -19.380 1112.370 -16.380 1112.380 ;
        RECT 27.020 1112.370 30.020 1112.380 ;
        RECT 207.020 1112.370 210.020 1112.380 ;
        RECT 387.020 1112.370 390.020 1112.380 ;
        RECT 567.020 1112.370 570.020 1112.380 ;
        RECT 747.020 1112.370 750.020 1112.380 ;
        RECT 927.020 1112.370 930.020 1112.380 ;
        RECT 1107.020 1112.370 1110.020 1112.380 ;
        RECT 1287.020 1112.370 1290.020 1112.380 ;
        RECT 1467.020 1112.370 1470.020 1112.380 ;
        RECT 1647.020 1112.370 1650.020 1112.380 ;
        RECT 1827.020 1112.370 1830.020 1112.380 ;
        RECT 2007.020 1112.370 2010.020 1112.380 ;
        RECT 2187.020 1112.370 2190.020 1112.380 ;
        RECT 2367.020 1112.370 2370.020 1112.380 ;
        RECT 2547.020 1112.370 2550.020 1112.380 ;
        RECT 2727.020 1112.370 2730.020 1112.380 ;
        RECT 2907.020 1112.370 2910.020 1112.380 ;
        RECT 2936.000 1112.370 2939.000 1112.380 ;
        RECT -19.380 935.380 -16.380 935.390 ;
        RECT 27.020 935.380 30.020 935.390 ;
        RECT 207.020 935.380 210.020 935.390 ;
        RECT 387.020 935.380 390.020 935.390 ;
        RECT 567.020 935.380 570.020 935.390 ;
        RECT 747.020 935.380 750.020 935.390 ;
        RECT 927.020 935.380 930.020 935.390 ;
        RECT 1107.020 935.380 1110.020 935.390 ;
        RECT 1287.020 935.380 1290.020 935.390 ;
        RECT 1467.020 935.380 1470.020 935.390 ;
        RECT 1647.020 935.380 1650.020 935.390 ;
        RECT 1827.020 935.380 1830.020 935.390 ;
        RECT 2007.020 935.380 2010.020 935.390 ;
        RECT 2187.020 935.380 2190.020 935.390 ;
        RECT 2367.020 935.380 2370.020 935.390 ;
        RECT 2547.020 935.380 2550.020 935.390 ;
        RECT 2727.020 935.380 2730.020 935.390 ;
        RECT 2907.020 935.380 2910.020 935.390 ;
        RECT 2936.000 935.380 2939.000 935.390 ;
        RECT -24.080 932.380 2943.700 935.380 ;
        RECT -19.380 932.370 -16.380 932.380 ;
        RECT 27.020 932.370 30.020 932.380 ;
        RECT 207.020 932.370 210.020 932.380 ;
        RECT 387.020 932.370 390.020 932.380 ;
        RECT 567.020 932.370 570.020 932.380 ;
        RECT 747.020 932.370 750.020 932.380 ;
        RECT 927.020 932.370 930.020 932.380 ;
        RECT 1107.020 932.370 1110.020 932.380 ;
        RECT 1287.020 932.370 1290.020 932.380 ;
        RECT 1467.020 932.370 1470.020 932.380 ;
        RECT 1647.020 932.370 1650.020 932.380 ;
        RECT 1827.020 932.370 1830.020 932.380 ;
        RECT 2007.020 932.370 2010.020 932.380 ;
        RECT 2187.020 932.370 2190.020 932.380 ;
        RECT 2367.020 932.370 2370.020 932.380 ;
        RECT 2547.020 932.370 2550.020 932.380 ;
        RECT 2727.020 932.370 2730.020 932.380 ;
        RECT 2907.020 932.370 2910.020 932.380 ;
        RECT 2936.000 932.370 2939.000 932.380 ;
        RECT -19.380 755.380 -16.380 755.390 ;
        RECT 27.020 755.380 30.020 755.390 ;
        RECT 207.020 755.380 210.020 755.390 ;
        RECT 387.020 755.380 390.020 755.390 ;
        RECT 567.020 755.380 570.020 755.390 ;
        RECT 747.020 755.380 750.020 755.390 ;
        RECT 927.020 755.380 930.020 755.390 ;
        RECT 1107.020 755.380 1110.020 755.390 ;
        RECT 1287.020 755.380 1290.020 755.390 ;
        RECT 1467.020 755.380 1470.020 755.390 ;
        RECT 1647.020 755.380 1650.020 755.390 ;
        RECT 1827.020 755.380 1830.020 755.390 ;
        RECT 2007.020 755.380 2010.020 755.390 ;
        RECT 2187.020 755.380 2190.020 755.390 ;
        RECT 2367.020 755.380 2370.020 755.390 ;
        RECT 2547.020 755.380 2550.020 755.390 ;
        RECT 2727.020 755.380 2730.020 755.390 ;
        RECT 2907.020 755.380 2910.020 755.390 ;
        RECT 2936.000 755.380 2939.000 755.390 ;
        RECT -24.080 752.380 2943.700 755.380 ;
        RECT -19.380 752.370 -16.380 752.380 ;
        RECT 27.020 752.370 30.020 752.380 ;
        RECT 207.020 752.370 210.020 752.380 ;
        RECT 387.020 752.370 390.020 752.380 ;
        RECT 567.020 752.370 570.020 752.380 ;
        RECT 747.020 752.370 750.020 752.380 ;
        RECT 927.020 752.370 930.020 752.380 ;
        RECT 1107.020 752.370 1110.020 752.380 ;
        RECT 1287.020 752.370 1290.020 752.380 ;
        RECT 1467.020 752.370 1470.020 752.380 ;
        RECT 1647.020 752.370 1650.020 752.380 ;
        RECT 1827.020 752.370 1830.020 752.380 ;
        RECT 2007.020 752.370 2010.020 752.380 ;
        RECT 2187.020 752.370 2190.020 752.380 ;
        RECT 2367.020 752.370 2370.020 752.380 ;
        RECT 2547.020 752.370 2550.020 752.380 ;
        RECT 2727.020 752.370 2730.020 752.380 ;
        RECT 2907.020 752.370 2910.020 752.380 ;
        RECT 2936.000 752.370 2939.000 752.380 ;
        RECT -19.380 575.380 -16.380 575.390 ;
        RECT 27.020 575.380 30.020 575.390 ;
        RECT 207.020 575.380 210.020 575.390 ;
        RECT 387.020 575.380 390.020 575.390 ;
        RECT 567.020 575.380 570.020 575.390 ;
        RECT 747.020 575.380 750.020 575.390 ;
        RECT 927.020 575.380 930.020 575.390 ;
        RECT 1107.020 575.380 1110.020 575.390 ;
        RECT 1287.020 575.380 1290.020 575.390 ;
        RECT 1467.020 575.380 1470.020 575.390 ;
        RECT 1647.020 575.380 1650.020 575.390 ;
        RECT 1827.020 575.380 1830.020 575.390 ;
        RECT 2007.020 575.380 2010.020 575.390 ;
        RECT 2187.020 575.380 2190.020 575.390 ;
        RECT 2367.020 575.380 2370.020 575.390 ;
        RECT 2547.020 575.380 2550.020 575.390 ;
        RECT 2727.020 575.380 2730.020 575.390 ;
        RECT 2907.020 575.380 2910.020 575.390 ;
        RECT 2936.000 575.380 2939.000 575.390 ;
        RECT -24.080 572.380 2943.700 575.380 ;
        RECT -19.380 572.370 -16.380 572.380 ;
        RECT 27.020 572.370 30.020 572.380 ;
        RECT 207.020 572.370 210.020 572.380 ;
        RECT 387.020 572.370 390.020 572.380 ;
        RECT 567.020 572.370 570.020 572.380 ;
        RECT 747.020 572.370 750.020 572.380 ;
        RECT 927.020 572.370 930.020 572.380 ;
        RECT 1107.020 572.370 1110.020 572.380 ;
        RECT 1287.020 572.370 1290.020 572.380 ;
        RECT 1467.020 572.370 1470.020 572.380 ;
        RECT 1647.020 572.370 1650.020 572.380 ;
        RECT 1827.020 572.370 1830.020 572.380 ;
        RECT 2007.020 572.370 2010.020 572.380 ;
        RECT 2187.020 572.370 2190.020 572.380 ;
        RECT 2367.020 572.370 2370.020 572.380 ;
        RECT 2547.020 572.370 2550.020 572.380 ;
        RECT 2727.020 572.370 2730.020 572.380 ;
        RECT 2907.020 572.370 2910.020 572.380 ;
        RECT 2936.000 572.370 2939.000 572.380 ;
        RECT -19.380 395.380 -16.380 395.390 ;
        RECT 27.020 395.380 30.020 395.390 ;
        RECT 207.020 395.380 210.020 395.390 ;
        RECT 387.020 395.380 390.020 395.390 ;
        RECT 567.020 395.380 570.020 395.390 ;
        RECT 747.020 395.380 750.020 395.390 ;
        RECT 927.020 395.380 930.020 395.390 ;
        RECT 1107.020 395.380 1110.020 395.390 ;
        RECT 1287.020 395.380 1290.020 395.390 ;
        RECT 1467.020 395.380 1470.020 395.390 ;
        RECT 1647.020 395.380 1650.020 395.390 ;
        RECT 1827.020 395.380 1830.020 395.390 ;
        RECT 2007.020 395.380 2010.020 395.390 ;
        RECT 2187.020 395.380 2190.020 395.390 ;
        RECT 2367.020 395.380 2370.020 395.390 ;
        RECT 2547.020 395.380 2550.020 395.390 ;
        RECT 2727.020 395.380 2730.020 395.390 ;
        RECT 2907.020 395.380 2910.020 395.390 ;
        RECT 2936.000 395.380 2939.000 395.390 ;
        RECT -24.080 392.380 2943.700 395.380 ;
        RECT -19.380 392.370 -16.380 392.380 ;
        RECT 27.020 392.370 30.020 392.380 ;
        RECT 207.020 392.370 210.020 392.380 ;
        RECT 387.020 392.370 390.020 392.380 ;
        RECT 567.020 392.370 570.020 392.380 ;
        RECT 747.020 392.370 750.020 392.380 ;
        RECT 927.020 392.370 930.020 392.380 ;
        RECT 1107.020 392.370 1110.020 392.380 ;
        RECT 1287.020 392.370 1290.020 392.380 ;
        RECT 1467.020 392.370 1470.020 392.380 ;
        RECT 1647.020 392.370 1650.020 392.380 ;
        RECT 1827.020 392.370 1830.020 392.380 ;
        RECT 2007.020 392.370 2010.020 392.380 ;
        RECT 2187.020 392.370 2190.020 392.380 ;
        RECT 2367.020 392.370 2370.020 392.380 ;
        RECT 2547.020 392.370 2550.020 392.380 ;
        RECT 2727.020 392.370 2730.020 392.380 ;
        RECT 2907.020 392.370 2910.020 392.380 ;
        RECT 2936.000 392.370 2939.000 392.380 ;
        RECT -19.380 215.380 -16.380 215.390 ;
        RECT 27.020 215.380 30.020 215.390 ;
        RECT 207.020 215.380 210.020 215.390 ;
        RECT 387.020 215.380 390.020 215.390 ;
        RECT 567.020 215.380 570.020 215.390 ;
        RECT 747.020 215.380 750.020 215.390 ;
        RECT 927.020 215.380 930.020 215.390 ;
        RECT 1107.020 215.380 1110.020 215.390 ;
        RECT 1287.020 215.380 1290.020 215.390 ;
        RECT 1467.020 215.380 1470.020 215.390 ;
        RECT 1647.020 215.380 1650.020 215.390 ;
        RECT 1827.020 215.380 1830.020 215.390 ;
        RECT 2007.020 215.380 2010.020 215.390 ;
        RECT 2187.020 215.380 2190.020 215.390 ;
        RECT 2367.020 215.380 2370.020 215.390 ;
        RECT 2547.020 215.380 2550.020 215.390 ;
        RECT 2727.020 215.380 2730.020 215.390 ;
        RECT 2907.020 215.380 2910.020 215.390 ;
        RECT 2936.000 215.380 2939.000 215.390 ;
        RECT -24.080 212.380 2943.700 215.380 ;
        RECT -19.380 212.370 -16.380 212.380 ;
        RECT 27.020 212.370 30.020 212.380 ;
        RECT 207.020 212.370 210.020 212.380 ;
        RECT 387.020 212.370 390.020 212.380 ;
        RECT 567.020 212.370 570.020 212.380 ;
        RECT 747.020 212.370 750.020 212.380 ;
        RECT 927.020 212.370 930.020 212.380 ;
        RECT 1107.020 212.370 1110.020 212.380 ;
        RECT 1287.020 212.370 1290.020 212.380 ;
        RECT 1467.020 212.370 1470.020 212.380 ;
        RECT 1647.020 212.370 1650.020 212.380 ;
        RECT 1827.020 212.370 1830.020 212.380 ;
        RECT 2007.020 212.370 2010.020 212.380 ;
        RECT 2187.020 212.370 2190.020 212.380 ;
        RECT 2367.020 212.370 2370.020 212.380 ;
        RECT 2547.020 212.370 2550.020 212.380 ;
        RECT 2727.020 212.370 2730.020 212.380 ;
        RECT 2907.020 212.370 2910.020 212.380 ;
        RECT 2936.000 212.370 2939.000 212.380 ;
        RECT -19.380 35.380 -16.380 35.390 ;
        RECT 27.020 35.380 30.020 35.390 ;
        RECT 207.020 35.380 210.020 35.390 ;
        RECT 387.020 35.380 390.020 35.390 ;
        RECT 567.020 35.380 570.020 35.390 ;
        RECT 747.020 35.380 750.020 35.390 ;
        RECT 927.020 35.380 930.020 35.390 ;
        RECT 1107.020 35.380 1110.020 35.390 ;
        RECT 1287.020 35.380 1290.020 35.390 ;
        RECT 1467.020 35.380 1470.020 35.390 ;
        RECT 1647.020 35.380 1650.020 35.390 ;
        RECT 1827.020 35.380 1830.020 35.390 ;
        RECT 2007.020 35.380 2010.020 35.390 ;
        RECT 2187.020 35.380 2190.020 35.390 ;
        RECT 2367.020 35.380 2370.020 35.390 ;
        RECT 2547.020 35.380 2550.020 35.390 ;
        RECT 2727.020 35.380 2730.020 35.390 ;
        RECT 2907.020 35.380 2910.020 35.390 ;
        RECT 2936.000 35.380 2939.000 35.390 ;
        RECT -24.080 32.380 2943.700 35.380 ;
        RECT -19.380 32.370 -16.380 32.380 ;
        RECT 27.020 32.370 30.020 32.380 ;
        RECT 207.020 32.370 210.020 32.380 ;
        RECT 387.020 32.370 390.020 32.380 ;
        RECT 567.020 32.370 570.020 32.380 ;
        RECT 747.020 32.370 750.020 32.380 ;
        RECT 927.020 32.370 930.020 32.380 ;
        RECT 1107.020 32.370 1110.020 32.380 ;
        RECT 1287.020 32.370 1290.020 32.380 ;
        RECT 1467.020 32.370 1470.020 32.380 ;
        RECT 1647.020 32.370 1650.020 32.380 ;
        RECT 1827.020 32.370 1830.020 32.380 ;
        RECT 2007.020 32.370 2010.020 32.380 ;
        RECT 2187.020 32.370 2190.020 32.380 ;
        RECT 2367.020 32.370 2370.020 32.380 ;
        RECT 2547.020 32.370 2550.020 32.380 ;
        RECT 2727.020 32.370 2730.020 32.380 ;
        RECT 2907.020 32.370 2910.020 32.380 ;
        RECT 2936.000 32.370 2939.000 32.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 27.020 -11.020 30.020 -11.010 ;
        RECT 207.020 -11.020 210.020 -11.010 ;
        RECT 387.020 -11.020 390.020 -11.010 ;
        RECT 567.020 -11.020 570.020 -11.010 ;
        RECT 747.020 -11.020 750.020 -11.010 ;
        RECT 927.020 -11.020 930.020 -11.010 ;
        RECT 1107.020 -11.020 1110.020 -11.010 ;
        RECT 1287.020 -11.020 1290.020 -11.010 ;
        RECT 1467.020 -11.020 1470.020 -11.010 ;
        RECT 1647.020 -11.020 1650.020 -11.010 ;
        RECT 1827.020 -11.020 1830.020 -11.010 ;
        RECT 2007.020 -11.020 2010.020 -11.010 ;
        RECT 2187.020 -11.020 2190.020 -11.010 ;
        RECT 2367.020 -11.020 2370.020 -11.010 ;
        RECT 2547.020 -11.020 2550.020 -11.010 ;
        RECT 2727.020 -11.020 2730.020 -11.010 ;
        RECT 2907.020 -11.020 2910.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 27.020 -14.030 30.020 -14.020 ;
        RECT 207.020 -14.030 210.020 -14.020 ;
        RECT 387.020 -14.030 390.020 -14.020 ;
        RECT 567.020 -14.030 570.020 -14.020 ;
        RECT 747.020 -14.030 750.020 -14.020 ;
        RECT 927.020 -14.030 930.020 -14.020 ;
        RECT 1107.020 -14.030 1110.020 -14.020 ;
        RECT 1287.020 -14.030 1290.020 -14.020 ;
        RECT 1467.020 -14.030 1470.020 -14.020 ;
        RECT 1647.020 -14.030 1650.020 -14.020 ;
        RECT 1827.020 -14.030 1830.020 -14.020 ;
        RECT 2007.020 -14.030 2010.020 -14.020 ;
        RECT 2187.020 -14.030 2190.020 -14.020 ;
        RECT 2367.020 -14.030 2370.020 -14.020 ;
        RECT 2547.020 -14.030 2550.020 -14.020 ;
        RECT 2727.020 -14.030 2730.020 -14.020 ;
        RECT 2907.020 -14.030 2910.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 117.020 -18.720 120.020 3538.400 ;
        RECT 297.020 -18.720 300.020 3538.400 ;
        RECT 477.020 -18.720 480.020 3538.400 ;
        RECT 657.020 -18.720 660.020 3538.400 ;
        RECT 837.020 -18.720 840.020 3538.400 ;
        RECT 1017.020 -18.720 1020.020 3538.400 ;
        RECT 1197.020 -18.720 1200.020 3538.400 ;
        RECT 1377.020 -18.720 1380.020 3538.400 ;
        RECT 1557.020 -18.720 1560.020 3538.400 ;
        RECT 1737.020 -18.720 1740.020 3538.400 ;
        RECT 1917.020 -18.720 1920.020 3538.400 ;
        RECT 2097.020 -18.720 2100.020 3538.400 ;
        RECT 2277.020 -18.720 2280.020 3538.400 ;
        RECT 2457.020 -18.720 2460.020 3538.400 ;
        RECT 2637.020 -18.720 2640.020 3538.400 ;
        RECT 2817.020 -18.720 2820.020 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 3364.090 -21.990 3365.270 ;
        RECT -23.170 3362.490 -21.990 3363.670 ;
        RECT -23.170 3184.090 -21.990 3185.270 ;
        RECT -23.170 3182.490 -21.990 3183.670 ;
        RECT -23.170 3004.090 -21.990 3005.270 ;
        RECT -23.170 3002.490 -21.990 3003.670 ;
        RECT -23.170 2824.090 -21.990 2825.270 ;
        RECT -23.170 2822.490 -21.990 2823.670 ;
        RECT -23.170 2644.090 -21.990 2645.270 ;
        RECT -23.170 2642.490 -21.990 2643.670 ;
        RECT -23.170 2464.090 -21.990 2465.270 ;
        RECT -23.170 2462.490 -21.990 2463.670 ;
        RECT -23.170 2284.090 -21.990 2285.270 ;
        RECT -23.170 2282.490 -21.990 2283.670 ;
        RECT -23.170 2104.090 -21.990 2105.270 ;
        RECT -23.170 2102.490 -21.990 2103.670 ;
        RECT -23.170 1924.090 -21.990 1925.270 ;
        RECT -23.170 1922.490 -21.990 1923.670 ;
        RECT -23.170 1744.090 -21.990 1745.270 ;
        RECT -23.170 1742.490 -21.990 1743.670 ;
        RECT -23.170 1564.090 -21.990 1565.270 ;
        RECT -23.170 1562.490 -21.990 1563.670 ;
        RECT -23.170 1384.090 -21.990 1385.270 ;
        RECT -23.170 1382.490 -21.990 1383.670 ;
        RECT -23.170 1204.090 -21.990 1205.270 ;
        RECT -23.170 1202.490 -21.990 1203.670 ;
        RECT -23.170 1024.090 -21.990 1025.270 ;
        RECT -23.170 1022.490 -21.990 1023.670 ;
        RECT -23.170 844.090 -21.990 845.270 ;
        RECT -23.170 842.490 -21.990 843.670 ;
        RECT -23.170 664.090 -21.990 665.270 ;
        RECT -23.170 662.490 -21.990 663.670 ;
        RECT -23.170 484.090 -21.990 485.270 ;
        RECT -23.170 482.490 -21.990 483.670 ;
        RECT -23.170 304.090 -21.990 305.270 ;
        RECT -23.170 302.490 -21.990 303.670 ;
        RECT -23.170 124.090 -21.990 125.270 ;
        RECT -23.170 122.490 -21.990 123.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 117.930 3537.110 119.110 3538.290 ;
        RECT 117.930 3535.510 119.110 3536.690 ;
        RECT 117.930 3364.090 119.110 3365.270 ;
        RECT 117.930 3362.490 119.110 3363.670 ;
        RECT 117.930 3184.090 119.110 3185.270 ;
        RECT 117.930 3182.490 119.110 3183.670 ;
        RECT 117.930 3004.090 119.110 3005.270 ;
        RECT 117.930 3002.490 119.110 3003.670 ;
        RECT 117.930 2824.090 119.110 2825.270 ;
        RECT 117.930 2822.490 119.110 2823.670 ;
        RECT 117.930 2644.090 119.110 2645.270 ;
        RECT 117.930 2642.490 119.110 2643.670 ;
        RECT 117.930 2464.090 119.110 2465.270 ;
        RECT 117.930 2462.490 119.110 2463.670 ;
        RECT 117.930 2284.090 119.110 2285.270 ;
        RECT 117.930 2282.490 119.110 2283.670 ;
        RECT 117.930 2104.090 119.110 2105.270 ;
        RECT 117.930 2102.490 119.110 2103.670 ;
        RECT 117.930 1924.090 119.110 1925.270 ;
        RECT 117.930 1922.490 119.110 1923.670 ;
        RECT 117.930 1744.090 119.110 1745.270 ;
        RECT 117.930 1742.490 119.110 1743.670 ;
        RECT 117.930 1564.090 119.110 1565.270 ;
        RECT 117.930 1562.490 119.110 1563.670 ;
        RECT 117.930 1384.090 119.110 1385.270 ;
        RECT 117.930 1382.490 119.110 1383.670 ;
        RECT 117.930 1204.090 119.110 1205.270 ;
        RECT 117.930 1202.490 119.110 1203.670 ;
        RECT 117.930 1024.090 119.110 1025.270 ;
        RECT 117.930 1022.490 119.110 1023.670 ;
        RECT 117.930 844.090 119.110 845.270 ;
        RECT 117.930 842.490 119.110 843.670 ;
        RECT 117.930 664.090 119.110 665.270 ;
        RECT 117.930 662.490 119.110 663.670 ;
        RECT 117.930 484.090 119.110 485.270 ;
        RECT 117.930 482.490 119.110 483.670 ;
        RECT 117.930 304.090 119.110 305.270 ;
        RECT 117.930 302.490 119.110 303.670 ;
        RECT 117.930 124.090 119.110 125.270 ;
        RECT 117.930 122.490 119.110 123.670 ;
        RECT 117.930 -17.010 119.110 -15.830 ;
        RECT 117.930 -18.610 119.110 -17.430 ;
        RECT 297.930 3537.110 299.110 3538.290 ;
        RECT 297.930 3535.510 299.110 3536.690 ;
        RECT 297.930 3364.090 299.110 3365.270 ;
        RECT 297.930 3362.490 299.110 3363.670 ;
        RECT 297.930 3184.090 299.110 3185.270 ;
        RECT 297.930 3182.490 299.110 3183.670 ;
        RECT 297.930 3004.090 299.110 3005.270 ;
        RECT 297.930 3002.490 299.110 3003.670 ;
        RECT 297.930 2824.090 299.110 2825.270 ;
        RECT 297.930 2822.490 299.110 2823.670 ;
        RECT 297.930 2644.090 299.110 2645.270 ;
        RECT 297.930 2642.490 299.110 2643.670 ;
        RECT 297.930 2464.090 299.110 2465.270 ;
        RECT 297.930 2462.490 299.110 2463.670 ;
        RECT 297.930 2284.090 299.110 2285.270 ;
        RECT 297.930 2282.490 299.110 2283.670 ;
        RECT 297.930 2104.090 299.110 2105.270 ;
        RECT 297.930 2102.490 299.110 2103.670 ;
        RECT 297.930 1924.090 299.110 1925.270 ;
        RECT 297.930 1922.490 299.110 1923.670 ;
        RECT 297.930 1744.090 299.110 1745.270 ;
        RECT 297.930 1742.490 299.110 1743.670 ;
        RECT 297.930 1564.090 299.110 1565.270 ;
        RECT 297.930 1562.490 299.110 1563.670 ;
        RECT 297.930 1384.090 299.110 1385.270 ;
        RECT 297.930 1382.490 299.110 1383.670 ;
        RECT 297.930 1204.090 299.110 1205.270 ;
        RECT 297.930 1202.490 299.110 1203.670 ;
        RECT 297.930 1024.090 299.110 1025.270 ;
        RECT 297.930 1022.490 299.110 1023.670 ;
        RECT 297.930 844.090 299.110 845.270 ;
        RECT 297.930 842.490 299.110 843.670 ;
        RECT 297.930 664.090 299.110 665.270 ;
        RECT 297.930 662.490 299.110 663.670 ;
        RECT 297.930 484.090 299.110 485.270 ;
        RECT 297.930 482.490 299.110 483.670 ;
        RECT 297.930 304.090 299.110 305.270 ;
        RECT 297.930 302.490 299.110 303.670 ;
        RECT 297.930 124.090 299.110 125.270 ;
        RECT 297.930 122.490 299.110 123.670 ;
        RECT 297.930 -17.010 299.110 -15.830 ;
        RECT 297.930 -18.610 299.110 -17.430 ;
        RECT 477.930 3537.110 479.110 3538.290 ;
        RECT 477.930 3535.510 479.110 3536.690 ;
        RECT 477.930 3364.090 479.110 3365.270 ;
        RECT 477.930 3362.490 479.110 3363.670 ;
        RECT 477.930 3184.090 479.110 3185.270 ;
        RECT 477.930 3182.490 479.110 3183.670 ;
        RECT 477.930 3004.090 479.110 3005.270 ;
        RECT 477.930 3002.490 479.110 3003.670 ;
        RECT 477.930 2824.090 479.110 2825.270 ;
        RECT 477.930 2822.490 479.110 2823.670 ;
        RECT 477.930 2644.090 479.110 2645.270 ;
        RECT 477.930 2642.490 479.110 2643.670 ;
        RECT 477.930 2464.090 479.110 2465.270 ;
        RECT 477.930 2462.490 479.110 2463.670 ;
        RECT 477.930 2284.090 479.110 2285.270 ;
        RECT 477.930 2282.490 479.110 2283.670 ;
        RECT 477.930 2104.090 479.110 2105.270 ;
        RECT 477.930 2102.490 479.110 2103.670 ;
        RECT 477.930 1924.090 479.110 1925.270 ;
        RECT 477.930 1922.490 479.110 1923.670 ;
        RECT 477.930 1744.090 479.110 1745.270 ;
        RECT 477.930 1742.490 479.110 1743.670 ;
        RECT 477.930 1564.090 479.110 1565.270 ;
        RECT 477.930 1562.490 479.110 1563.670 ;
        RECT 477.930 1384.090 479.110 1385.270 ;
        RECT 477.930 1382.490 479.110 1383.670 ;
        RECT 477.930 1204.090 479.110 1205.270 ;
        RECT 477.930 1202.490 479.110 1203.670 ;
        RECT 477.930 1024.090 479.110 1025.270 ;
        RECT 477.930 1022.490 479.110 1023.670 ;
        RECT 477.930 844.090 479.110 845.270 ;
        RECT 477.930 842.490 479.110 843.670 ;
        RECT 477.930 664.090 479.110 665.270 ;
        RECT 477.930 662.490 479.110 663.670 ;
        RECT 477.930 484.090 479.110 485.270 ;
        RECT 477.930 482.490 479.110 483.670 ;
        RECT 477.930 304.090 479.110 305.270 ;
        RECT 477.930 302.490 479.110 303.670 ;
        RECT 477.930 124.090 479.110 125.270 ;
        RECT 477.930 122.490 479.110 123.670 ;
        RECT 477.930 -17.010 479.110 -15.830 ;
        RECT 477.930 -18.610 479.110 -17.430 ;
        RECT 657.930 3537.110 659.110 3538.290 ;
        RECT 657.930 3535.510 659.110 3536.690 ;
        RECT 657.930 3364.090 659.110 3365.270 ;
        RECT 657.930 3362.490 659.110 3363.670 ;
        RECT 657.930 3184.090 659.110 3185.270 ;
        RECT 657.930 3182.490 659.110 3183.670 ;
        RECT 657.930 3004.090 659.110 3005.270 ;
        RECT 657.930 3002.490 659.110 3003.670 ;
        RECT 657.930 2824.090 659.110 2825.270 ;
        RECT 657.930 2822.490 659.110 2823.670 ;
        RECT 657.930 2644.090 659.110 2645.270 ;
        RECT 657.930 2642.490 659.110 2643.670 ;
        RECT 657.930 2464.090 659.110 2465.270 ;
        RECT 657.930 2462.490 659.110 2463.670 ;
        RECT 657.930 2284.090 659.110 2285.270 ;
        RECT 657.930 2282.490 659.110 2283.670 ;
        RECT 657.930 2104.090 659.110 2105.270 ;
        RECT 657.930 2102.490 659.110 2103.670 ;
        RECT 657.930 1924.090 659.110 1925.270 ;
        RECT 657.930 1922.490 659.110 1923.670 ;
        RECT 657.930 1744.090 659.110 1745.270 ;
        RECT 657.930 1742.490 659.110 1743.670 ;
        RECT 657.930 1564.090 659.110 1565.270 ;
        RECT 657.930 1562.490 659.110 1563.670 ;
        RECT 657.930 1384.090 659.110 1385.270 ;
        RECT 657.930 1382.490 659.110 1383.670 ;
        RECT 657.930 1204.090 659.110 1205.270 ;
        RECT 657.930 1202.490 659.110 1203.670 ;
        RECT 657.930 1024.090 659.110 1025.270 ;
        RECT 657.930 1022.490 659.110 1023.670 ;
        RECT 657.930 844.090 659.110 845.270 ;
        RECT 657.930 842.490 659.110 843.670 ;
        RECT 657.930 664.090 659.110 665.270 ;
        RECT 657.930 662.490 659.110 663.670 ;
        RECT 657.930 484.090 659.110 485.270 ;
        RECT 657.930 482.490 659.110 483.670 ;
        RECT 657.930 304.090 659.110 305.270 ;
        RECT 657.930 302.490 659.110 303.670 ;
        RECT 657.930 124.090 659.110 125.270 ;
        RECT 657.930 122.490 659.110 123.670 ;
        RECT 657.930 -17.010 659.110 -15.830 ;
        RECT 657.930 -18.610 659.110 -17.430 ;
        RECT 837.930 3537.110 839.110 3538.290 ;
        RECT 837.930 3535.510 839.110 3536.690 ;
        RECT 837.930 3364.090 839.110 3365.270 ;
        RECT 837.930 3362.490 839.110 3363.670 ;
        RECT 837.930 3184.090 839.110 3185.270 ;
        RECT 837.930 3182.490 839.110 3183.670 ;
        RECT 837.930 3004.090 839.110 3005.270 ;
        RECT 837.930 3002.490 839.110 3003.670 ;
        RECT 837.930 2824.090 839.110 2825.270 ;
        RECT 837.930 2822.490 839.110 2823.670 ;
        RECT 837.930 2644.090 839.110 2645.270 ;
        RECT 837.930 2642.490 839.110 2643.670 ;
        RECT 837.930 2464.090 839.110 2465.270 ;
        RECT 837.930 2462.490 839.110 2463.670 ;
        RECT 837.930 2284.090 839.110 2285.270 ;
        RECT 837.930 2282.490 839.110 2283.670 ;
        RECT 837.930 2104.090 839.110 2105.270 ;
        RECT 837.930 2102.490 839.110 2103.670 ;
        RECT 837.930 1924.090 839.110 1925.270 ;
        RECT 837.930 1922.490 839.110 1923.670 ;
        RECT 837.930 1744.090 839.110 1745.270 ;
        RECT 837.930 1742.490 839.110 1743.670 ;
        RECT 837.930 1564.090 839.110 1565.270 ;
        RECT 837.930 1562.490 839.110 1563.670 ;
        RECT 837.930 1384.090 839.110 1385.270 ;
        RECT 837.930 1382.490 839.110 1383.670 ;
        RECT 837.930 1204.090 839.110 1205.270 ;
        RECT 837.930 1202.490 839.110 1203.670 ;
        RECT 837.930 1024.090 839.110 1025.270 ;
        RECT 837.930 1022.490 839.110 1023.670 ;
        RECT 837.930 844.090 839.110 845.270 ;
        RECT 837.930 842.490 839.110 843.670 ;
        RECT 837.930 664.090 839.110 665.270 ;
        RECT 837.930 662.490 839.110 663.670 ;
        RECT 837.930 484.090 839.110 485.270 ;
        RECT 837.930 482.490 839.110 483.670 ;
        RECT 837.930 304.090 839.110 305.270 ;
        RECT 837.930 302.490 839.110 303.670 ;
        RECT 837.930 124.090 839.110 125.270 ;
        RECT 837.930 122.490 839.110 123.670 ;
        RECT 837.930 -17.010 839.110 -15.830 ;
        RECT 837.930 -18.610 839.110 -17.430 ;
        RECT 1017.930 3537.110 1019.110 3538.290 ;
        RECT 1017.930 3535.510 1019.110 3536.690 ;
        RECT 1017.930 3364.090 1019.110 3365.270 ;
        RECT 1017.930 3362.490 1019.110 3363.670 ;
        RECT 1017.930 3184.090 1019.110 3185.270 ;
        RECT 1017.930 3182.490 1019.110 3183.670 ;
        RECT 1017.930 3004.090 1019.110 3005.270 ;
        RECT 1017.930 3002.490 1019.110 3003.670 ;
        RECT 1017.930 2824.090 1019.110 2825.270 ;
        RECT 1017.930 2822.490 1019.110 2823.670 ;
        RECT 1017.930 2644.090 1019.110 2645.270 ;
        RECT 1017.930 2642.490 1019.110 2643.670 ;
        RECT 1017.930 2464.090 1019.110 2465.270 ;
        RECT 1017.930 2462.490 1019.110 2463.670 ;
        RECT 1017.930 2284.090 1019.110 2285.270 ;
        RECT 1017.930 2282.490 1019.110 2283.670 ;
        RECT 1017.930 2104.090 1019.110 2105.270 ;
        RECT 1017.930 2102.490 1019.110 2103.670 ;
        RECT 1017.930 1924.090 1019.110 1925.270 ;
        RECT 1017.930 1922.490 1019.110 1923.670 ;
        RECT 1017.930 1744.090 1019.110 1745.270 ;
        RECT 1017.930 1742.490 1019.110 1743.670 ;
        RECT 1017.930 1564.090 1019.110 1565.270 ;
        RECT 1017.930 1562.490 1019.110 1563.670 ;
        RECT 1017.930 1384.090 1019.110 1385.270 ;
        RECT 1017.930 1382.490 1019.110 1383.670 ;
        RECT 1017.930 1204.090 1019.110 1205.270 ;
        RECT 1017.930 1202.490 1019.110 1203.670 ;
        RECT 1017.930 1024.090 1019.110 1025.270 ;
        RECT 1017.930 1022.490 1019.110 1023.670 ;
        RECT 1017.930 844.090 1019.110 845.270 ;
        RECT 1017.930 842.490 1019.110 843.670 ;
        RECT 1017.930 664.090 1019.110 665.270 ;
        RECT 1017.930 662.490 1019.110 663.670 ;
        RECT 1017.930 484.090 1019.110 485.270 ;
        RECT 1017.930 482.490 1019.110 483.670 ;
        RECT 1017.930 304.090 1019.110 305.270 ;
        RECT 1017.930 302.490 1019.110 303.670 ;
        RECT 1017.930 124.090 1019.110 125.270 ;
        RECT 1017.930 122.490 1019.110 123.670 ;
        RECT 1017.930 -17.010 1019.110 -15.830 ;
        RECT 1017.930 -18.610 1019.110 -17.430 ;
        RECT 1197.930 3537.110 1199.110 3538.290 ;
        RECT 1197.930 3535.510 1199.110 3536.690 ;
        RECT 1197.930 3364.090 1199.110 3365.270 ;
        RECT 1197.930 3362.490 1199.110 3363.670 ;
        RECT 1197.930 3184.090 1199.110 3185.270 ;
        RECT 1197.930 3182.490 1199.110 3183.670 ;
        RECT 1197.930 3004.090 1199.110 3005.270 ;
        RECT 1197.930 3002.490 1199.110 3003.670 ;
        RECT 1197.930 2824.090 1199.110 2825.270 ;
        RECT 1197.930 2822.490 1199.110 2823.670 ;
        RECT 1197.930 2644.090 1199.110 2645.270 ;
        RECT 1197.930 2642.490 1199.110 2643.670 ;
        RECT 1197.930 2464.090 1199.110 2465.270 ;
        RECT 1197.930 2462.490 1199.110 2463.670 ;
        RECT 1197.930 2284.090 1199.110 2285.270 ;
        RECT 1197.930 2282.490 1199.110 2283.670 ;
        RECT 1197.930 2104.090 1199.110 2105.270 ;
        RECT 1197.930 2102.490 1199.110 2103.670 ;
        RECT 1197.930 1924.090 1199.110 1925.270 ;
        RECT 1197.930 1922.490 1199.110 1923.670 ;
        RECT 1197.930 1744.090 1199.110 1745.270 ;
        RECT 1197.930 1742.490 1199.110 1743.670 ;
        RECT 1197.930 1564.090 1199.110 1565.270 ;
        RECT 1197.930 1562.490 1199.110 1563.670 ;
        RECT 1197.930 1384.090 1199.110 1385.270 ;
        RECT 1197.930 1382.490 1199.110 1383.670 ;
        RECT 1197.930 1204.090 1199.110 1205.270 ;
        RECT 1197.930 1202.490 1199.110 1203.670 ;
        RECT 1197.930 1024.090 1199.110 1025.270 ;
        RECT 1197.930 1022.490 1199.110 1023.670 ;
        RECT 1197.930 844.090 1199.110 845.270 ;
        RECT 1197.930 842.490 1199.110 843.670 ;
        RECT 1197.930 664.090 1199.110 665.270 ;
        RECT 1197.930 662.490 1199.110 663.670 ;
        RECT 1197.930 484.090 1199.110 485.270 ;
        RECT 1197.930 482.490 1199.110 483.670 ;
        RECT 1197.930 304.090 1199.110 305.270 ;
        RECT 1197.930 302.490 1199.110 303.670 ;
        RECT 1197.930 124.090 1199.110 125.270 ;
        RECT 1197.930 122.490 1199.110 123.670 ;
        RECT 1197.930 -17.010 1199.110 -15.830 ;
        RECT 1197.930 -18.610 1199.110 -17.430 ;
        RECT 1377.930 3537.110 1379.110 3538.290 ;
        RECT 1377.930 3535.510 1379.110 3536.690 ;
        RECT 1377.930 3364.090 1379.110 3365.270 ;
        RECT 1377.930 3362.490 1379.110 3363.670 ;
        RECT 1377.930 3184.090 1379.110 3185.270 ;
        RECT 1377.930 3182.490 1379.110 3183.670 ;
        RECT 1377.930 3004.090 1379.110 3005.270 ;
        RECT 1377.930 3002.490 1379.110 3003.670 ;
        RECT 1377.930 2824.090 1379.110 2825.270 ;
        RECT 1377.930 2822.490 1379.110 2823.670 ;
        RECT 1377.930 2644.090 1379.110 2645.270 ;
        RECT 1377.930 2642.490 1379.110 2643.670 ;
        RECT 1377.930 2464.090 1379.110 2465.270 ;
        RECT 1377.930 2462.490 1379.110 2463.670 ;
        RECT 1377.930 2284.090 1379.110 2285.270 ;
        RECT 1377.930 2282.490 1379.110 2283.670 ;
        RECT 1377.930 2104.090 1379.110 2105.270 ;
        RECT 1377.930 2102.490 1379.110 2103.670 ;
        RECT 1377.930 1924.090 1379.110 1925.270 ;
        RECT 1377.930 1922.490 1379.110 1923.670 ;
        RECT 1377.930 1744.090 1379.110 1745.270 ;
        RECT 1377.930 1742.490 1379.110 1743.670 ;
        RECT 1377.930 1564.090 1379.110 1565.270 ;
        RECT 1377.930 1562.490 1379.110 1563.670 ;
        RECT 1377.930 1384.090 1379.110 1385.270 ;
        RECT 1377.930 1382.490 1379.110 1383.670 ;
        RECT 1377.930 1204.090 1379.110 1205.270 ;
        RECT 1377.930 1202.490 1379.110 1203.670 ;
        RECT 1377.930 1024.090 1379.110 1025.270 ;
        RECT 1377.930 1022.490 1379.110 1023.670 ;
        RECT 1377.930 844.090 1379.110 845.270 ;
        RECT 1377.930 842.490 1379.110 843.670 ;
        RECT 1377.930 664.090 1379.110 665.270 ;
        RECT 1377.930 662.490 1379.110 663.670 ;
        RECT 1377.930 484.090 1379.110 485.270 ;
        RECT 1377.930 482.490 1379.110 483.670 ;
        RECT 1377.930 304.090 1379.110 305.270 ;
        RECT 1377.930 302.490 1379.110 303.670 ;
        RECT 1377.930 124.090 1379.110 125.270 ;
        RECT 1377.930 122.490 1379.110 123.670 ;
        RECT 1377.930 -17.010 1379.110 -15.830 ;
        RECT 1377.930 -18.610 1379.110 -17.430 ;
        RECT 1557.930 3537.110 1559.110 3538.290 ;
        RECT 1557.930 3535.510 1559.110 3536.690 ;
        RECT 1557.930 3364.090 1559.110 3365.270 ;
        RECT 1557.930 3362.490 1559.110 3363.670 ;
        RECT 1557.930 3184.090 1559.110 3185.270 ;
        RECT 1557.930 3182.490 1559.110 3183.670 ;
        RECT 1557.930 3004.090 1559.110 3005.270 ;
        RECT 1557.930 3002.490 1559.110 3003.670 ;
        RECT 1557.930 2824.090 1559.110 2825.270 ;
        RECT 1557.930 2822.490 1559.110 2823.670 ;
        RECT 1557.930 2644.090 1559.110 2645.270 ;
        RECT 1557.930 2642.490 1559.110 2643.670 ;
        RECT 1557.930 2464.090 1559.110 2465.270 ;
        RECT 1557.930 2462.490 1559.110 2463.670 ;
        RECT 1557.930 2284.090 1559.110 2285.270 ;
        RECT 1557.930 2282.490 1559.110 2283.670 ;
        RECT 1557.930 2104.090 1559.110 2105.270 ;
        RECT 1557.930 2102.490 1559.110 2103.670 ;
        RECT 1557.930 1924.090 1559.110 1925.270 ;
        RECT 1557.930 1922.490 1559.110 1923.670 ;
        RECT 1557.930 1744.090 1559.110 1745.270 ;
        RECT 1557.930 1742.490 1559.110 1743.670 ;
        RECT 1557.930 1564.090 1559.110 1565.270 ;
        RECT 1557.930 1562.490 1559.110 1563.670 ;
        RECT 1557.930 1384.090 1559.110 1385.270 ;
        RECT 1557.930 1382.490 1559.110 1383.670 ;
        RECT 1557.930 1204.090 1559.110 1205.270 ;
        RECT 1557.930 1202.490 1559.110 1203.670 ;
        RECT 1557.930 1024.090 1559.110 1025.270 ;
        RECT 1557.930 1022.490 1559.110 1023.670 ;
        RECT 1557.930 844.090 1559.110 845.270 ;
        RECT 1557.930 842.490 1559.110 843.670 ;
        RECT 1557.930 664.090 1559.110 665.270 ;
        RECT 1557.930 662.490 1559.110 663.670 ;
        RECT 1557.930 484.090 1559.110 485.270 ;
        RECT 1557.930 482.490 1559.110 483.670 ;
        RECT 1557.930 304.090 1559.110 305.270 ;
        RECT 1557.930 302.490 1559.110 303.670 ;
        RECT 1557.930 124.090 1559.110 125.270 ;
        RECT 1557.930 122.490 1559.110 123.670 ;
        RECT 1557.930 -17.010 1559.110 -15.830 ;
        RECT 1557.930 -18.610 1559.110 -17.430 ;
        RECT 1737.930 3537.110 1739.110 3538.290 ;
        RECT 1737.930 3535.510 1739.110 3536.690 ;
        RECT 1737.930 3364.090 1739.110 3365.270 ;
        RECT 1737.930 3362.490 1739.110 3363.670 ;
        RECT 1737.930 3184.090 1739.110 3185.270 ;
        RECT 1737.930 3182.490 1739.110 3183.670 ;
        RECT 1737.930 3004.090 1739.110 3005.270 ;
        RECT 1737.930 3002.490 1739.110 3003.670 ;
        RECT 1737.930 2824.090 1739.110 2825.270 ;
        RECT 1737.930 2822.490 1739.110 2823.670 ;
        RECT 1737.930 2644.090 1739.110 2645.270 ;
        RECT 1737.930 2642.490 1739.110 2643.670 ;
        RECT 1737.930 2464.090 1739.110 2465.270 ;
        RECT 1737.930 2462.490 1739.110 2463.670 ;
        RECT 1737.930 2284.090 1739.110 2285.270 ;
        RECT 1737.930 2282.490 1739.110 2283.670 ;
        RECT 1737.930 2104.090 1739.110 2105.270 ;
        RECT 1737.930 2102.490 1739.110 2103.670 ;
        RECT 1737.930 1924.090 1739.110 1925.270 ;
        RECT 1737.930 1922.490 1739.110 1923.670 ;
        RECT 1737.930 1744.090 1739.110 1745.270 ;
        RECT 1737.930 1742.490 1739.110 1743.670 ;
        RECT 1737.930 1564.090 1739.110 1565.270 ;
        RECT 1737.930 1562.490 1739.110 1563.670 ;
        RECT 1737.930 1384.090 1739.110 1385.270 ;
        RECT 1737.930 1382.490 1739.110 1383.670 ;
        RECT 1737.930 1204.090 1739.110 1205.270 ;
        RECT 1737.930 1202.490 1739.110 1203.670 ;
        RECT 1737.930 1024.090 1739.110 1025.270 ;
        RECT 1737.930 1022.490 1739.110 1023.670 ;
        RECT 1737.930 844.090 1739.110 845.270 ;
        RECT 1737.930 842.490 1739.110 843.670 ;
        RECT 1737.930 664.090 1739.110 665.270 ;
        RECT 1737.930 662.490 1739.110 663.670 ;
        RECT 1737.930 484.090 1739.110 485.270 ;
        RECT 1737.930 482.490 1739.110 483.670 ;
        RECT 1737.930 304.090 1739.110 305.270 ;
        RECT 1737.930 302.490 1739.110 303.670 ;
        RECT 1737.930 124.090 1739.110 125.270 ;
        RECT 1737.930 122.490 1739.110 123.670 ;
        RECT 1737.930 -17.010 1739.110 -15.830 ;
        RECT 1737.930 -18.610 1739.110 -17.430 ;
        RECT 1917.930 3537.110 1919.110 3538.290 ;
        RECT 1917.930 3535.510 1919.110 3536.690 ;
        RECT 1917.930 3364.090 1919.110 3365.270 ;
        RECT 1917.930 3362.490 1919.110 3363.670 ;
        RECT 1917.930 3184.090 1919.110 3185.270 ;
        RECT 1917.930 3182.490 1919.110 3183.670 ;
        RECT 1917.930 3004.090 1919.110 3005.270 ;
        RECT 1917.930 3002.490 1919.110 3003.670 ;
        RECT 1917.930 2824.090 1919.110 2825.270 ;
        RECT 1917.930 2822.490 1919.110 2823.670 ;
        RECT 1917.930 2644.090 1919.110 2645.270 ;
        RECT 1917.930 2642.490 1919.110 2643.670 ;
        RECT 1917.930 2464.090 1919.110 2465.270 ;
        RECT 1917.930 2462.490 1919.110 2463.670 ;
        RECT 1917.930 2284.090 1919.110 2285.270 ;
        RECT 1917.930 2282.490 1919.110 2283.670 ;
        RECT 1917.930 2104.090 1919.110 2105.270 ;
        RECT 1917.930 2102.490 1919.110 2103.670 ;
        RECT 1917.930 1924.090 1919.110 1925.270 ;
        RECT 1917.930 1922.490 1919.110 1923.670 ;
        RECT 1917.930 1744.090 1919.110 1745.270 ;
        RECT 1917.930 1742.490 1919.110 1743.670 ;
        RECT 1917.930 1564.090 1919.110 1565.270 ;
        RECT 1917.930 1562.490 1919.110 1563.670 ;
        RECT 1917.930 1384.090 1919.110 1385.270 ;
        RECT 1917.930 1382.490 1919.110 1383.670 ;
        RECT 1917.930 1204.090 1919.110 1205.270 ;
        RECT 1917.930 1202.490 1919.110 1203.670 ;
        RECT 1917.930 1024.090 1919.110 1025.270 ;
        RECT 1917.930 1022.490 1919.110 1023.670 ;
        RECT 1917.930 844.090 1919.110 845.270 ;
        RECT 1917.930 842.490 1919.110 843.670 ;
        RECT 1917.930 664.090 1919.110 665.270 ;
        RECT 1917.930 662.490 1919.110 663.670 ;
        RECT 1917.930 484.090 1919.110 485.270 ;
        RECT 1917.930 482.490 1919.110 483.670 ;
        RECT 1917.930 304.090 1919.110 305.270 ;
        RECT 1917.930 302.490 1919.110 303.670 ;
        RECT 1917.930 124.090 1919.110 125.270 ;
        RECT 1917.930 122.490 1919.110 123.670 ;
        RECT 1917.930 -17.010 1919.110 -15.830 ;
        RECT 1917.930 -18.610 1919.110 -17.430 ;
        RECT 2097.930 3537.110 2099.110 3538.290 ;
        RECT 2097.930 3535.510 2099.110 3536.690 ;
        RECT 2097.930 3364.090 2099.110 3365.270 ;
        RECT 2097.930 3362.490 2099.110 3363.670 ;
        RECT 2097.930 3184.090 2099.110 3185.270 ;
        RECT 2097.930 3182.490 2099.110 3183.670 ;
        RECT 2097.930 3004.090 2099.110 3005.270 ;
        RECT 2097.930 3002.490 2099.110 3003.670 ;
        RECT 2097.930 2824.090 2099.110 2825.270 ;
        RECT 2097.930 2822.490 2099.110 2823.670 ;
        RECT 2097.930 2644.090 2099.110 2645.270 ;
        RECT 2097.930 2642.490 2099.110 2643.670 ;
        RECT 2097.930 2464.090 2099.110 2465.270 ;
        RECT 2097.930 2462.490 2099.110 2463.670 ;
        RECT 2097.930 2284.090 2099.110 2285.270 ;
        RECT 2097.930 2282.490 2099.110 2283.670 ;
        RECT 2097.930 2104.090 2099.110 2105.270 ;
        RECT 2097.930 2102.490 2099.110 2103.670 ;
        RECT 2097.930 1924.090 2099.110 1925.270 ;
        RECT 2097.930 1922.490 2099.110 1923.670 ;
        RECT 2097.930 1744.090 2099.110 1745.270 ;
        RECT 2097.930 1742.490 2099.110 1743.670 ;
        RECT 2097.930 1564.090 2099.110 1565.270 ;
        RECT 2097.930 1562.490 2099.110 1563.670 ;
        RECT 2097.930 1384.090 2099.110 1385.270 ;
        RECT 2097.930 1382.490 2099.110 1383.670 ;
        RECT 2097.930 1204.090 2099.110 1205.270 ;
        RECT 2097.930 1202.490 2099.110 1203.670 ;
        RECT 2097.930 1024.090 2099.110 1025.270 ;
        RECT 2097.930 1022.490 2099.110 1023.670 ;
        RECT 2097.930 844.090 2099.110 845.270 ;
        RECT 2097.930 842.490 2099.110 843.670 ;
        RECT 2097.930 664.090 2099.110 665.270 ;
        RECT 2097.930 662.490 2099.110 663.670 ;
        RECT 2097.930 484.090 2099.110 485.270 ;
        RECT 2097.930 482.490 2099.110 483.670 ;
        RECT 2097.930 304.090 2099.110 305.270 ;
        RECT 2097.930 302.490 2099.110 303.670 ;
        RECT 2097.930 124.090 2099.110 125.270 ;
        RECT 2097.930 122.490 2099.110 123.670 ;
        RECT 2097.930 -17.010 2099.110 -15.830 ;
        RECT 2097.930 -18.610 2099.110 -17.430 ;
        RECT 2277.930 3537.110 2279.110 3538.290 ;
        RECT 2277.930 3535.510 2279.110 3536.690 ;
        RECT 2277.930 3364.090 2279.110 3365.270 ;
        RECT 2277.930 3362.490 2279.110 3363.670 ;
        RECT 2277.930 3184.090 2279.110 3185.270 ;
        RECT 2277.930 3182.490 2279.110 3183.670 ;
        RECT 2277.930 3004.090 2279.110 3005.270 ;
        RECT 2277.930 3002.490 2279.110 3003.670 ;
        RECT 2277.930 2824.090 2279.110 2825.270 ;
        RECT 2277.930 2822.490 2279.110 2823.670 ;
        RECT 2277.930 2644.090 2279.110 2645.270 ;
        RECT 2277.930 2642.490 2279.110 2643.670 ;
        RECT 2277.930 2464.090 2279.110 2465.270 ;
        RECT 2277.930 2462.490 2279.110 2463.670 ;
        RECT 2277.930 2284.090 2279.110 2285.270 ;
        RECT 2277.930 2282.490 2279.110 2283.670 ;
        RECT 2277.930 2104.090 2279.110 2105.270 ;
        RECT 2277.930 2102.490 2279.110 2103.670 ;
        RECT 2277.930 1924.090 2279.110 1925.270 ;
        RECT 2277.930 1922.490 2279.110 1923.670 ;
        RECT 2277.930 1744.090 2279.110 1745.270 ;
        RECT 2277.930 1742.490 2279.110 1743.670 ;
        RECT 2277.930 1564.090 2279.110 1565.270 ;
        RECT 2277.930 1562.490 2279.110 1563.670 ;
        RECT 2277.930 1384.090 2279.110 1385.270 ;
        RECT 2277.930 1382.490 2279.110 1383.670 ;
        RECT 2277.930 1204.090 2279.110 1205.270 ;
        RECT 2277.930 1202.490 2279.110 1203.670 ;
        RECT 2277.930 1024.090 2279.110 1025.270 ;
        RECT 2277.930 1022.490 2279.110 1023.670 ;
        RECT 2277.930 844.090 2279.110 845.270 ;
        RECT 2277.930 842.490 2279.110 843.670 ;
        RECT 2277.930 664.090 2279.110 665.270 ;
        RECT 2277.930 662.490 2279.110 663.670 ;
        RECT 2277.930 484.090 2279.110 485.270 ;
        RECT 2277.930 482.490 2279.110 483.670 ;
        RECT 2277.930 304.090 2279.110 305.270 ;
        RECT 2277.930 302.490 2279.110 303.670 ;
        RECT 2277.930 124.090 2279.110 125.270 ;
        RECT 2277.930 122.490 2279.110 123.670 ;
        RECT 2277.930 -17.010 2279.110 -15.830 ;
        RECT 2277.930 -18.610 2279.110 -17.430 ;
        RECT 2457.930 3537.110 2459.110 3538.290 ;
        RECT 2457.930 3535.510 2459.110 3536.690 ;
        RECT 2457.930 3364.090 2459.110 3365.270 ;
        RECT 2457.930 3362.490 2459.110 3363.670 ;
        RECT 2457.930 3184.090 2459.110 3185.270 ;
        RECT 2457.930 3182.490 2459.110 3183.670 ;
        RECT 2457.930 3004.090 2459.110 3005.270 ;
        RECT 2457.930 3002.490 2459.110 3003.670 ;
        RECT 2457.930 2824.090 2459.110 2825.270 ;
        RECT 2457.930 2822.490 2459.110 2823.670 ;
        RECT 2457.930 2644.090 2459.110 2645.270 ;
        RECT 2457.930 2642.490 2459.110 2643.670 ;
        RECT 2457.930 2464.090 2459.110 2465.270 ;
        RECT 2457.930 2462.490 2459.110 2463.670 ;
        RECT 2457.930 2284.090 2459.110 2285.270 ;
        RECT 2457.930 2282.490 2459.110 2283.670 ;
        RECT 2457.930 2104.090 2459.110 2105.270 ;
        RECT 2457.930 2102.490 2459.110 2103.670 ;
        RECT 2457.930 1924.090 2459.110 1925.270 ;
        RECT 2457.930 1922.490 2459.110 1923.670 ;
        RECT 2457.930 1744.090 2459.110 1745.270 ;
        RECT 2457.930 1742.490 2459.110 1743.670 ;
        RECT 2457.930 1564.090 2459.110 1565.270 ;
        RECT 2457.930 1562.490 2459.110 1563.670 ;
        RECT 2457.930 1384.090 2459.110 1385.270 ;
        RECT 2457.930 1382.490 2459.110 1383.670 ;
        RECT 2457.930 1204.090 2459.110 1205.270 ;
        RECT 2457.930 1202.490 2459.110 1203.670 ;
        RECT 2457.930 1024.090 2459.110 1025.270 ;
        RECT 2457.930 1022.490 2459.110 1023.670 ;
        RECT 2457.930 844.090 2459.110 845.270 ;
        RECT 2457.930 842.490 2459.110 843.670 ;
        RECT 2457.930 664.090 2459.110 665.270 ;
        RECT 2457.930 662.490 2459.110 663.670 ;
        RECT 2457.930 484.090 2459.110 485.270 ;
        RECT 2457.930 482.490 2459.110 483.670 ;
        RECT 2457.930 304.090 2459.110 305.270 ;
        RECT 2457.930 302.490 2459.110 303.670 ;
        RECT 2457.930 124.090 2459.110 125.270 ;
        RECT 2457.930 122.490 2459.110 123.670 ;
        RECT 2457.930 -17.010 2459.110 -15.830 ;
        RECT 2457.930 -18.610 2459.110 -17.430 ;
        RECT 2637.930 3537.110 2639.110 3538.290 ;
        RECT 2637.930 3535.510 2639.110 3536.690 ;
        RECT 2637.930 3364.090 2639.110 3365.270 ;
        RECT 2637.930 3362.490 2639.110 3363.670 ;
        RECT 2637.930 3184.090 2639.110 3185.270 ;
        RECT 2637.930 3182.490 2639.110 3183.670 ;
        RECT 2637.930 3004.090 2639.110 3005.270 ;
        RECT 2637.930 3002.490 2639.110 3003.670 ;
        RECT 2637.930 2824.090 2639.110 2825.270 ;
        RECT 2637.930 2822.490 2639.110 2823.670 ;
        RECT 2637.930 2644.090 2639.110 2645.270 ;
        RECT 2637.930 2642.490 2639.110 2643.670 ;
        RECT 2637.930 2464.090 2639.110 2465.270 ;
        RECT 2637.930 2462.490 2639.110 2463.670 ;
        RECT 2637.930 2284.090 2639.110 2285.270 ;
        RECT 2637.930 2282.490 2639.110 2283.670 ;
        RECT 2637.930 2104.090 2639.110 2105.270 ;
        RECT 2637.930 2102.490 2639.110 2103.670 ;
        RECT 2637.930 1924.090 2639.110 1925.270 ;
        RECT 2637.930 1922.490 2639.110 1923.670 ;
        RECT 2637.930 1744.090 2639.110 1745.270 ;
        RECT 2637.930 1742.490 2639.110 1743.670 ;
        RECT 2637.930 1564.090 2639.110 1565.270 ;
        RECT 2637.930 1562.490 2639.110 1563.670 ;
        RECT 2637.930 1384.090 2639.110 1385.270 ;
        RECT 2637.930 1382.490 2639.110 1383.670 ;
        RECT 2637.930 1204.090 2639.110 1205.270 ;
        RECT 2637.930 1202.490 2639.110 1203.670 ;
        RECT 2637.930 1024.090 2639.110 1025.270 ;
        RECT 2637.930 1022.490 2639.110 1023.670 ;
        RECT 2637.930 844.090 2639.110 845.270 ;
        RECT 2637.930 842.490 2639.110 843.670 ;
        RECT 2637.930 664.090 2639.110 665.270 ;
        RECT 2637.930 662.490 2639.110 663.670 ;
        RECT 2637.930 484.090 2639.110 485.270 ;
        RECT 2637.930 482.490 2639.110 483.670 ;
        RECT 2637.930 304.090 2639.110 305.270 ;
        RECT 2637.930 302.490 2639.110 303.670 ;
        RECT 2637.930 124.090 2639.110 125.270 ;
        RECT 2637.930 122.490 2639.110 123.670 ;
        RECT 2637.930 -17.010 2639.110 -15.830 ;
        RECT 2637.930 -18.610 2639.110 -17.430 ;
        RECT 2817.930 3537.110 2819.110 3538.290 ;
        RECT 2817.930 3535.510 2819.110 3536.690 ;
        RECT 2817.930 3364.090 2819.110 3365.270 ;
        RECT 2817.930 3362.490 2819.110 3363.670 ;
        RECT 2817.930 3184.090 2819.110 3185.270 ;
        RECT 2817.930 3182.490 2819.110 3183.670 ;
        RECT 2817.930 3004.090 2819.110 3005.270 ;
        RECT 2817.930 3002.490 2819.110 3003.670 ;
        RECT 2817.930 2824.090 2819.110 2825.270 ;
        RECT 2817.930 2822.490 2819.110 2823.670 ;
        RECT 2817.930 2644.090 2819.110 2645.270 ;
        RECT 2817.930 2642.490 2819.110 2643.670 ;
        RECT 2817.930 2464.090 2819.110 2465.270 ;
        RECT 2817.930 2462.490 2819.110 2463.670 ;
        RECT 2817.930 2284.090 2819.110 2285.270 ;
        RECT 2817.930 2282.490 2819.110 2283.670 ;
        RECT 2817.930 2104.090 2819.110 2105.270 ;
        RECT 2817.930 2102.490 2819.110 2103.670 ;
        RECT 2817.930 1924.090 2819.110 1925.270 ;
        RECT 2817.930 1922.490 2819.110 1923.670 ;
        RECT 2817.930 1744.090 2819.110 1745.270 ;
        RECT 2817.930 1742.490 2819.110 1743.670 ;
        RECT 2817.930 1564.090 2819.110 1565.270 ;
        RECT 2817.930 1562.490 2819.110 1563.670 ;
        RECT 2817.930 1384.090 2819.110 1385.270 ;
        RECT 2817.930 1382.490 2819.110 1383.670 ;
        RECT 2817.930 1204.090 2819.110 1205.270 ;
        RECT 2817.930 1202.490 2819.110 1203.670 ;
        RECT 2817.930 1024.090 2819.110 1025.270 ;
        RECT 2817.930 1022.490 2819.110 1023.670 ;
        RECT 2817.930 844.090 2819.110 845.270 ;
        RECT 2817.930 842.490 2819.110 843.670 ;
        RECT 2817.930 664.090 2819.110 665.270 ;
        RECT 2817.930 662.490 2819.110 663.670 ;
        RECT 2817.930 484.090 2819.110 485.270 ;
        RECT 2817.930 482.490 2819.110 483.670 ;
        RECT 2817.930 304.090 2819.110 305.270 ;
        RECT 2817.930 302.490 2819.110 303.670 ;
        RECT 2817.930 124.090 2819.110 125.270 ;
        RECT 2817.930 122.490 2819.110 123.670 ;
        RECT 2817.930 -17.010 2819.110 -15.830 ;
        RECT 2817.930 -18.610 2819.110 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 3364.090 2942.790 3365.270 ;
        RECT 2941.610 3362.490 2942.790 3363.670 ;
        RECT 2941.610 3184.090 2942.790 3185.270 ;
        RECT 2941.610 3182.490 2942.790 3183.670 ;
        RECT 2941.610 3004.090 2942.790 3005.270 ;
        RECT 2941.610 3002.490 2942.790 3003.670 ;
        RECT 2941.610 2824.090 2942.790 2825.270 ;
        RECT 2941.610 2822.490 2942.790 2823.670 ;
        RECT 2941.610 2644.090 2942.790 2645.270 ;
        RECT 2941.610 2642.490 2942.790 2643.670 ;
        RECT 2941.610 2464.090 2942.790 2465.270 ;
        RECT 2941.610 2462.490 2942.790 2463.670 ;
        RECT 2941.610 2284.090 2942.790 2285.270 ;
        RECT 2941.610 2282.490 2942.790 2283.670 ;
        RECT 2941.610 2104.090 2942.790 2105.270 ;
        RECT 2941.610 2102.490 2942.790 2103.670 ;
        RECT 2941.610 1924.090 2942.790 1925.270 ;
        RECT 2941.610 1922.490 2942.790 1923.670 ;
        RECT 2941.610 1744.090 2942.790 1745.270 ;
        RECT 2941.610 1742.490 2942.790 1743.670 ;
        RECT 2941.610 1564.090 2942.790 1565.270 ;
        RECT 2941.610 1562.490 2942.790 1563.670 ;
        RECT 2941.610 1384.090 2942.790 1385.270 ;
        RECT 2941.610 1382.490 2942.790 1383.670 ;
        RECT 2941.610 1204.090 2942.790 1205.270 ;
        RECT 2941.610 1202.490 2942.790 1203.670 ;
        RECT 2941.610 1024.090 2942.790 1025.270 ;
        RECT 2941.610 1022.490 2942.790 1023.670 ;
        RECT 2941.610 844.090 2942.790 845.270 ;
        RECT 2941.610 842.490 2942.790 843.670 ;
        RECT 2941.610 664.090 2942.790 665.270 ;
        RECT 2941.610 662.490 2942.790 663.670 ;
        RECT 2941.610 484.090 2942.790 485.270 ;
        RECT 2941.610 482.490 2942.790 483.670 ;
        RECT 2941.610 304.090 2942.790 305.270 ;
        RECT 2941.610 302.490 2942.790 303.670 ;
        RECT 2941.610 124.090 2942.790 125.270 ;
        RECT 2941.610 122.490 2942.790 123.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 117.020 3538.400 120.020 3538.410 ;
        RECT 297.020 3538.400 300.020 3538.410 ;
        RECT 477.020 3538.400 480.020 3538.410 ;
        RECT 657.020 3538.400 660.020 3538.410 ;
        RECT 837.020 3538.400 840.020 3538.410 ;
        RECT 1017.020 3538.400 1020.020 3538.410 ;
        RECT 1197.020 3538.400 1200.020 3538.410 ;
        RECT 1377.020 3538.400 1380.020 3538.410 ;
        RECT 1557.020 3538.400 1560.020 3538.410 ;
        RECT 1737.020 3538.400 1740.020 3538.410 ;
        RECT 1917.020 3538.400 1920.020 3538.410 ;
        RECT 2097.020 3538.400 2100.020 3538.410 ;
        RECT 2277.020 3538.400 2280.020 3538.410 ;
        RECT 2457.020 3538.400 2460.020 3538.410 ;
        RECT 2637.020 3538.400 2640.020 3538.410 ;
        RECT 2817.020 3538.400 2820.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 117.020 3535.390 120.020 3535.400 ;
        RECT 297.020 3535.390 300.020 3535.400 ;
        RECT 477.020 3535.390 480.020 3535.400 ;
        RECT 657.020 3535.390 660.020 3535.400 ;
        RECT 837.020 3535.390 840.020 3535.400 ;
        RECT 1017.020 3535.390 1020.020 3535.400 ;
        RECT 1197.020 3535.390 1200.020 3535.400 ;
        RECT 1377.020 3535.390 1380.020 3535.400 ;
        RECT 1557.020 3535.390 1560.020 3535.400 ;
        RECT 1737.020 3535.390 1740.020 3535.400 ;
        RECT 1917.020 3535.390 1920.020 3535.400 ;
        RECT 2097.020 3535.390 2100.020 3535.400 ;
        RECT 2277.020 3535.390 2280.020 3535.400 ;
        RECT 2457.020 3535.390 2460.020 3535.400 ;
        RECT 2637.020 3535.390 2640.020 3535.400 ;
        RECT 2817.020 3535.390 2820.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3365.380 -21.080 3365.390 ;
        RECT 117.020 3365.380 120.020 3365.390 ;
        RECT 297.020 3365.380 300.020 3365.390 ;
        RECT 477.020 3365.380 480.020 3365.390 ;
        RECT 657.020 3365.380 660.020 3365.390 ;
        RECT 837.020 3365.380 840.020 3365.390 ;
        RECT 1017.020 3365.380 1020.020 3365.390 ;
        RECT 1197.020 3365.380 1200.020 3365.390 ;
        RECT 1377.020 3365.380 1380.020 3365.390 ;
        RECT 1557.020 3365.380 1560.020 3365.390 ;
        RECT 1737.020 3365.380 1740.020 3365.390 ;
        RECT 1917.020 3365.380 1920.020 3365.390 ;
        RECT 2097.020 3365.380 2100.020 3365.390 ;
        RECT 2277.020 3365.380 2280.020 3365.390 ;
        RECT 2457.020 3365.380 2460.020 3365.390 ;
        RECT 2637.020 3365.380 2640.020 3365.390 ;
        RECT 2817.020 3365.380 2820.020 3365.390 ;
        RECT 2940.700 3365.380 2943.700 3365.390 ;
        RECT -24.080 3362.380 2943.700 3365.380 ;
        RECT -24.080 3362.370 -21.080 3362.380 ;
        RECT 117.020 3362.370 120.020 3362.380 ;
        RECT 297.020 3362.370 300.020 3362.380 ;
        RECT 477.020 3362.370 480.020 3362.380 ;
        RECT 657.020 3362.370 660.020 3362.380 ;
        RECT 837.020 3362.370 840.020 3362.380 ;
        RECT 1017.020 3362.370 1020.020 3362.380 ;
        RECT 1197.020 3362.370 1200.020 3362.380 ;
        RECT 1377.020 3362.370 1380.020 3362.380 ;
        RECT 1557.020 3362.370 1560.020 3362.380 ;
        RECT 1737.020 3362.370 1740.020 3362.380 ;
        RECT 1917.020 3362.370 1920.020 3362.380 ;
        RECT 2097.020 3362.370 2100.020 3362.380 ;
        RECT 2277.020 3362.370 2280.020 3362.380 ;
        RECT 2457.020 3362.370 2460.020 3362.380 ;
        RECT 2637.020 3362.370 2640.020 3362.380 ;
        RECT 2817.020 3362.370 2820.020 3362.380 ;
        RECT 2940.700 3362.370 2943.700 3362.380 ;
        RECT -24.080 3185.380 -21.080 3185.390 ;
        RECT 117.020 3185.380 120.020 3185.390 ;
        RECT 297.020 3185.380 300.020 3185.390 ;
        RECT 477.020 3185.380 480.020 3185.390 ;
        RECT 657.020 3185.380 660.020 3185.390 ;
        RECT 837.020 3185.380 840.020 3185.390 ;
        RECT 1017.020 3185.380 1020.020 3185.390 ;
        RECT 1197.020 3185.380 1200.020 3185.390 ;
        RECT 1377.020 3185.380 1380.020 3185.390 ;
        RECT 1557.020 3185.380 1560.020 3185.390 ;
        RECT 1737.020 3185.380 1740.020 3185.390 ;
        RECT 1917.020 3185.380 1920.020 3185.390 ;
        RECT 2097.020 3185.380 2100.020 3185.390 ;
        RECT 2277.020 3185.380 2280.020 3185.390 ;
        RECT 2457.020 3185.380 2460.020 3185.390 ;
        RECT 2637.020 3185.380 2640.020 3185.390 ;
        RECT 2817.020 3185.380 2820.020 3185.390 ;
        RECT 2940.700 3185.380 2943.700 3185.390 ;
        RECT -24.080 3182.380 2943.700 3185.380 ;
        RECT -24.080 3182.370 -21.080 3182.380 ;
        RECT 117.020 3182.370 120.020 3182.380 ;
        RECT 297.020 3182.370 300.020 3182.380 ;
        RECT 477.020 3182.370 480.020 3182.380 ;
        RECT 657.020 3182.370 660.020 3182.380 ;
        RECT 837.020 3182.370 840.020 3182.380 ;
        RECT 1017.020 3182.370 1020.020 3182.380 ;
        RECT 1197.020 3182.370 1200.020 3182.380 ;
        RECT 1377.020 3182.370 1380.020 3182.380 ;
        RECT 1557.020 3182.370 1560.020 3182.380 ;
        RECT 1737.020 3182.370 1740.020 3182.380 ;
        RECT 1917.020 3182.370 1920.020 3182.380 ;
        RECT 2097.020 3182.370 2100.020 3182.380 ;
        RECT 2277.020 3182.370 2280.020 3182.380 ;
        RECT 2457.020 3182.370 2460.020 3182.380 ;
        RECT 2637.020 3182.370 2640.020 3182.380 ;
        RECT 2817.020 3182.370 2820.020 3182.380 ;
        RECT 2940.700 3182.370 2943.700 3182.380 ;
        RECT -24.080 3005.380 -21.080 3005.390 ;
        RECT 117.020 3005.380 120.020 3005.390 ;
        RECT 297.020 3005.380 300.020 3005.390 ;
        RECT 477.020 3005.380 480.020 3005.390 ;
        RECT 657.020 3005.380 660.020 3005.390 ;
        RECT 837.020 3005.380 840.020 3005.390 ;
        RECT 1017.020 3005.380 1020.020 3005.390 ;
        RECT 1197.020 3005.380 1200.020 3005.390 ;
        RECT 1377.020 3005.380 1380.020 3005.390 ;
        RECT 1557.020 3005.380 1560.020 3005.390 ;
        RECT 1737.020 3005.380 1740.020 3005.390 ;
        RECT 1917.020 3005.380 1920.020 3005.390 ;
        RECT 2097.020 3005.380 2100.020 3005.390 ;
        RECT 2277.020 3005.380 2280.020 3005.390 ;
        RECT 2457.020 3005.380 2460.020 3005.390 ;
        RECT 2637.020 3005.380 2640.020 3005.390 ;
        RECT 2817.020 3005.380 2820.020 3005.390 ;
        RECT 2940.700 3005.380 2943.700 3005.390 ;
        RECT -24.080 3002.380 2943.700 3005.380 ;
        RECT -24.080 3002.370 -21.080 3002.380 ;
        RECT 117.020 3002.370 120.020 3002.380 ;
        RECT 297.020 3002.370 300.020 3002.380 ;
        RECT 477.020 3002.370 480.020 3002.380 ;
        RECT 657.020 3002.370 660.020 3002.380 ;
        RECT 837.020 3002.370 840.020 3002.380 ;
        RECT 1017.020 3002.370 1020.020 3002.380 ;
        RECT 1197.020 3002.370 1200.020 3002.380 ;
        RECT 1377.020 3002.370 1380.020 3002.380 ;
        RECT 1557.020 3002.370 1560.020 3002.380 ;
        RECT 1737.020 3002.370 1740.020 3002.380 ;
        RECT 1917.020 3002.370 1920.020 3002.380 ;
        RECT 2097.020 3002.370 2100.020 3002.380 ;
        RECT 2277.020 3002.370 2280.020 3002.380 ;
        RECT 2457.020 3002.370 2460.020 3002.380 ;
        RECT 2637.020 3002.370 2640.020 3002.380 ;
        RECT 2817.020 3002.370 2820.020 3002.380 ;
        RECT 2940.700 3002.370 2943.700 3002.380 ;
        RECT -24.080 2825.380 -21.080 2825.390 ;
        RECT 117.020 2825.380 120.020 2825.390 ;
        RECT 297.020 2825.380 300.020 2825.390 ;
        RECT 477.020 2825.380 480.020 2825.390 ;
        RECT 657.020 2825.380 660.020 2825.390 ;
        RECT 837.020 2825.380 840.020 2825.390 ;
        RECT 1017.020 2825.380 1020.020 2825.390 ;
        RECT 1197.020 2825.380 1200.020 2825.390 ;
        RECT 1377.020 2825.380 1380.020 2825.390 ;
        RECT 1557.020 2825.380 1560.020 2825.390 ;
        RECT 1737.020 2825.380 1740.020 2825.390 ;
        RECT 1917.020 2825.380 1920.020 2825.390 ;
        RECT 2097.020 2825.380 2100.020 2825.390 ;
        RECT 2277.020 2825.380 2280.020 2825.390 ;
        RECT 2457.020 2825.380 2460.020 2825.390 ;
        RECT 2637.020 2825.380 2640.020 2825.390 ;
        RECT 2817.020 2825.380 2820.020 2825.390 ;
        RECT 2940.700 2825.380 2943.700 2825.390 ;
        RECT -24.080 2822.380 2943.700 2825.380 ;
        RECT -24.080 2822.370 -21.080 2822.380 ;
        RECT 117.020 2822.370 120.020 2822.380 ;
        RECT 297.020 2822.370 300.020 2822.380 ;
        RECT 477.020 2822.370 480.020 2822.380 ;
        RECT 657.020 2822.370 660.020 2822.380 ;
        RECT 837.020 2822.370 840.020 2822.380 ;
        RECT 1017.020 2822.370 1020.020 2822.380 ;
        RECT 1197.020 2822.370 1200.020 2822.380 ;
        RECT 1377.020 2822.370 1380.020 2822.380 ;
        RECT 1557.020 2822.370 1560.020 2822.380 ;
        RECT 1737.020 2822.370 1740.020 2822.380 ;
        RECT 1917.020 2822.370 1920.020 2822.380 ;
        RECT 2097.020 2822.370 2100.020 2822.380 ;
        RECT 2277.020 2822.370 2280.020 2822.380 ;
        RECT 2457.020 2822.370 2460.020 2822.380 ;
        RECT 2637.020 2822.370 2640.020 2822.380 ;
        RECT 2817.020 2822.370 2820.020 2822.380 ;
        RECT 2940.700 2822.370 2943.700 2822.380 ;
        RECT -24.080 2645.380 -21.080 2645.390 ;
        RECT 117.020 2645.380 120.020 2645.390 ;
        RECT 297.020 2645.380 300.020 2645.390 ;
        RECT 477.020 2645.380 480.020 2645.390 ;
        RECT 657.020 2645.380 660.020 2645.390 ;
        RECT 837.020 2645.380 840.020 2645.390 ;
        RECT 1017.020 2645.380 1020.020 2645.390 ;
        RECT 1197.020 2645.380 1200.020 2645.390 ;
        RECT 1377.020 2645.380 1380.020 2645.390 ;
        RECT 1557.020 2645.380 1560.020 2645.390 ;
        RECT 1737.020 2645.380 1740.020 2645.390 ;
        RECT 1917.020 2645.380 1920.020 2645.390 ;
        RECT 2097.020 2645.380 2100.020 2645.390 ;
        RECT 2277.020 2645.380 2280.020 2645.390 ;
        RECT 2457.020 2645.380 2460.020 2645.390 ;
        RECT 2637.020 2645.380 2640.020 2645.390 ;
        RECT 2817.020 2645.380 2820.020 2645.390 ;
        RECT 2940.700 2645.380 2943.700 2645.390 ;
        RECT -24.080 2642.380 2943.700 2645.380 ;
        RECT -24.080 2642.370 -21.080 2642.380 ;
        RECT 117.020 2642.370 120.020 2642.380 ;
        RECT 297.020 2642.370 300.020 2642.380 ;
        RECT 477.020 2642.370 480.020 2642.380 ;
        RECT 657.020 2642.370 660.020 2642.380 ;
        RECT 837.020 2642.370 840.020 2642.380 ;
        RECT 1017.020 2642.370 1020.020 2642.380 ;
        RECT 1197.020 2642.370 1200.020 2642.380 ;
        RECT 1377.020 2642.370 1380.020 2642.380 ;
        RECT 1557.020 2642.370 1560.020 2642.380 ;
        RECT 1737.020 2642.370 1740.020 2642.380 ;
        RECT 1917.020 2642.370 1920.020 2642.380 ;
        RECT 2097.020 2642.370 2100.020 2642.380 ;
        RECT 2277.020 2642.370 2280.020 2642.380 ;
        RECT 2457.020 2642.370 2460.020 2642.380 ;
        RECT 2637.020 2642.370 2640.020 2642.380 ;
        RECT 2817.020 2642.370 2820.020 2642.380 ;
        RECT 2940.700 2642.370 2943.700 2642.380 ;
        RECT -24.080 2465.380 -21.080 2465.390 ;
        RECT 117.020 2465.380 120.020 2465.390 ;
        RECT 297.020 2465.380 300.020 2465.390 ;
        RECT 477.020 2465.380 480.020 2465.390 ;
        RECT 657.020 2465.380 660.020 2465.390 ;
        RECT 837.020 2465.380 840.020 2465.390 ;
        RECT 1017.020 2465.380 1020.020 2465.390 ;
        RECT 1197.020 2465.380 1200.020 2465.390 ;
        RECT 1377.020 2465.380 1380.020 2465.390 ;
        RECT 1557.020 2465.380 1560.020 2465.390 ;
        RECT 1737.020 2465.380 1740.020 2465.390 ;
        RECT 1917.020 2465.380 1920.020 2465.390 ;
        RECT 2097.020 2465.380 2100.020 2465.390 ;
        RECT 2277.020 2465.380 2280.020 2465.390 ;
        RECT 2457.020 2465.380 2460.020 2465.390 ;
        RECT 2637.020 2465.380 2640.020 2465.390 ;
        RECT 2817.020 2465.380 2820.020 2465.390 ;
        RECT 2940.700 2465.380 2943.700 2465.390 ;
        RECT -24.080 2462.380 2943.700 2465.380 ;
        RECT -24.080 2462.370 -21.080 2462.380 ;
        RECT 117.020 2462.370 120.020 2462.380 ;
        RECT 297.020 2462.370 300.020 2462.380 ;
        RECT 477.020 2462.370 480.020 2462.380 ;
        RECT 657.020 2462.370 660.020 2462.380 ;
        RECT 837.020 2462.370 840.020 2462.380 ;
        RECT 1017.020 2462.370 1020.020 2462.380 ;
        RECT 1197.020 2462.370 1200.020 2462.380 ;
        RECT 1377.020 2462.370 1380.020 2462.380 ;
        RECT 1557.020 2462.370 1560.020 2462.380 ;
        RECT 1737.020 2462.370 1740.020 2462.380 ;
        RECT 1917.020 2462.370 1920.020 2462.380 ;
        RECT 2097.020 2462.370 2100.020 2462.380 ;
        RECT 2277.020 2462.370 2280.020 2462.380 ;
        RECT 2457.020 2462.370 2460.020 2462.380 ;
        RECT 2637.020 2462.370 2640.020 2462.380 ;
        RECT 2817.020 2462.370 2820.020 2462.380 ;
        RECT 2940.700 2462.370 2943.700 2462.380 ;
        RECT -24.080 2285.380 -21.080 2285.390 ;
        RECT 117.020 2285.380 120.020 2285.390 ;
        RECT 297.020 2285.380 300.020 2285.390 ;
        RECT 477.020 2285.380 480.020 2285.390 ;
        RECT 657.020 2285.380 660.020 2285.390 ;
        RECT 837.020 2285.380 840.020 2285.390 ;
        RECT 1017.020 2285.380 1020.020 2285.390 ;
        RECT 1197.020 2285.380 1200.020 2285.390 ;
        RECT 1377.020 2285.380 1380.020 2285.390 ;
        RECT 1557.020 2285.380 1560.020 2285.390 ;
        RECT 1737.020 2285.380 1740.020 2285.390 ;
        RECT 1917.020 2285.380 1920.020 2285.390 ;
        RECT 2097.020 2285.380 2100.020 2285.390 ;
        RECT 2277.020 2285.380 2280.020 2285.390 ;
        RECT 2457.020 2285.380 2460.020 2285.390 ;
        RECT 2637.020 2285.380 2640.020 2285.390 ;
        RECT 2817.020 2285.380 2820.020 2285.390 ;
        RECT 2940.700 2285.380 2943.700 2285.390 ;
        RECT -24.080 2282.380 2943.700 2285.380 ;
        RECT -24.080 2282.370 -21.080 2282.380 ;
        RECT 117.020 2282.370 120.020 2282.380 ;
        RECT 297.020 2282.370 300.020 2282.380 ;
        RECT 477.020 2282.370 480.020 2282.380 ;
        RECT 657.020 2282.370 660.020 2282.380 ;
        RECT 837.020 2282.370 840.020 2282.380 ;
        RECT 1017.020 2282.370 1020.020 2282.380 ;
        RECT 1197.020 2282.370 1200.020 2282.380 ;
        RECT 1377.020 2282.370 1380.020 2282.380 ;
        RECT 1557.020 2282.370 1560.020 2282.380 ;
        RECT 1737.020 2282.370 1740.020 2282.380 ;
        RECT 1917.020 2282.370 1920.020 2282.380 ;
        RECT 2097.020 2282.370 2100.020 2282.380 ;
        RECT 2277.020 2282.370 2280.020 2282.380 ;
        RECT 2457.020 2282.370 2460.020 2282.380 ;
        RECT 2637.020 2282.370 2640.020 2282.380 ;
        RECT 2817.020 2282.370 2820.020 2282.380 ;
        RECT 2940.700 2282.370 2943.700 2282.380 ;
        RECT -24.080 2105.380 -21.080 2105.390 ;
        RECT 117.020 2105.380 120.020 2105.390 ;
        RECT 297.020 2105.380 300.020 2105.390 ;
        RECT 477.020 2105.380 480.020 2105.390 ;
        RECT 657.020 2105.380 660.020 2105.390 ;
        RECT 837.020 2105.380 840.020 2105.390 ;
        RECT 1017.020 2105.380 1020.020 2105.390 ;
        RECT 1197.020 2105.380 1200.020 2105.390 ;
        RECT 1377.020 2105.380 1380.020 2105.390 ;
        RECT 1557.020 2105.380 1560.020 2105.390 ;
        RECT 1737.020 2105.380 1740.020 2105.390 ;
        RECT 1917.020 2105.380 1920.020 2105.390 ;
        RECT 2097.020 2105.380 2100.020 2105.390 ;
        RECT 2277.020 2105.380 2280.020 2105.390 ;
        RECT 2457.020 2105.380 2460.020 2105.390 ;
        RECT 2637.020 2105.380 2640.020 2105.390 ;
        RECT 2817.020 2105.380 2820.020 2105.390 ;
        RECT 2940.700 2105.380 2943.700 2105.390 ;
        RECT -24.080 2102.380 2943.700 2105.380 ;
        RECT -24.080 2102.370 -21.080 2102.380 ;
        RECT 117.020 2102.370 120.020 2102.380 ;
        RECT 297.020 2102.370 300.020 2102.380 ;
        RECT 477.020 2102.370 480.020 2102.380 ;
        RECT 657.020 2102.370 660.020 2102.380 ;
        RECT 837.020 2102.370 840.020 2102.380 ;
        RECT 1017.020 2102.370 1020.020 2102.380 ;
        RECT 1197.020 2102.370 1200.020 2102.380 ;
        RECT 1377.020 2102.370 1380.020 2102.380 ;
        RECT 1557.020 2102.370 1560.020 2102.380 ;
        RECT 1737.020 2102.370 1740.020 2102.380 ;
        RECT 1917.020 2102.370 1920.020 2102.380 ;
        RECT 2097.020 2102.370 2100.020 2102.380 ;
        RECT 2277.020 2102.370 2280.020 2102.380 ;
        RECT 2457.020 2102.370 2460.020 2102.380 ;
        RECT 2637.020 2102.370 2640.020 2102.380 ;
        RECT 2817.020 2102.370 2820.020 2102.380 ;
        RECT 2940.700 2102.370 2943.700 2102.380 ;
        RECT -24.080 1925.380 -21.080 1925.390 ;
        RECT 117.020 1925.380 120.020 1925.390 ;
        RECT 297.020 1925.380 300.020 1925.390 ;
        RECT 477.020 1925.380 480.020 1925.390 ;
        RECT 657.020 1925.380 660.020 1925.390 ;
        RECT 837.020 1925.380 840.020 1925.390 ;
        RECT 1017.020 1925.380 1020.020 1925.390 ;
        RECT 1197.020 1925.380 1200.020 1925.390 ;
        RECT 1377.020 1925.380 1380.020 1925.390 ;
        RECT 1557.020 1925.380 1560.020 1925.390 ;
        RECT 1737.020 1925.380 1740.020 1925.390 ;
        RECT 1917.020 1925.380 1920.020 1925.390 ;
        RECT 2097.020 1925.380 2100.020 1925.390 ;
        RECT 2277.020 1925.380 2280.020 1925.390 ;
        RECT 2457.020 1925.380 2460.020 1925.390 ;
        RECT 2637.020 1925.380 2640.020 1925.390 ;
        RECT 2817.020 1925.380 2820.020 1925.390 ;
        RECT 2940.700 1925.380 2943.700 1925.390 ;
        RECT -24.080 1922.380 2943.700 1925.380 ;
        RECT -24.080 1922.370 -21.080 1922.380 ;
        RECT 117.020 1922.370 120.020 1922.380 ;
        RECT 297.020 1922.370 300.020 1922.380 ;
        RECT 477.020 1922.370 480.020 1922.380 ;
        RECT 657.020 1922.370 660.020 1922.380 ;
        RECT 837.020 1922.370 840.020 1922.380 ;
        RECT 1017.020 1922.370 1020.020 1922.380 ;
        RECT 1197.020 1922.370 1200.020 1922.380 ;
        RECT 1377.020 1922.370 1380.020 1922.380 ;
        RECT 1557.020 1922.370 1560.020 1922.380 ;
        RECT 1737.020 1922.370 1740.020 1922.380 ;
        RECT 1917.020 1922.370 1920.020 1922.380 ;
        RECT 2097.020 1922.370 2100.020 1922.380 ;
        RECT 2277.020 1922.370 2280.020 1922.380 ;
        RECT 2457.020 1922.370 2460.020 1922.380 ;
        RECT 2637.020 1922.370 2640.020 1922.380 ;
        RECT 2817.020 1922.370 2820.020 1922.380 ;
        RECT 2940.700 1922.370 2943.700 1922.380 ;
        RECT -24.080 1745.380 -21.080 1745.390 ;
        RECT 117.020 1745.380 120.020 1745.390 ;
        RECT 297.020 1745.380 300.020 1745.390 ;
        RECT 477.020 1745.380 480.020 1745.390 ;
        RECT 657.020 1745.380 660.020 1745.390 ;
        RECT 837.020 1745.380 840.020 1745.390 ;
        RECT 1017.020 1745.380 1020.020 1745.390 ;
        RECT 1197.020 1745.380 1200.020 1745.390 ;
        RECT 1377.020 1745.380 1380.020 1745.390 ;
        RECT 1557.020 1745.380 1560.020 1745.390 ;
        RECT 1737.020 1745.380 1740.020 1745.390 ;
        RECT 1917.020 1745.380 1920.020 1745.390 ;
        RECT 2097.020 1745.380 2100.020 1745.390 ;
        RECT 2277.020 1745.380 2280.020 1745.390 ;
        RECT 2457.020 1745.380 2460.020 1745.390 ;
        RECT 2637.020 1745.380 2640.020 1745.390 ;
        RECT 2817.020 1745.380 2820.020 1745.390 ;
        RECT 2940.700 1745.380 2943.700 1745.390 ;
        RECT -24.080 1742.380 2943.700 1745.380 ;
        RECT -24.080 1742.370 -21.080 1742.380 ;
        RECT 117.020 1742.370 120.020 1742.380 ;
        RECT 297.020 1742.370 300.020 1742.380 ;
        RECT 477.020 1742.370 480.020 1742.380 ;
        RECT 657.020 1742.370 660.020 1742.380 ;
        RECT 837.020 1742.370 840.020 1742.380 ;
        RECT 1017.020 1742.370 1020.020 1742.380 ;
        RECT 1197.020 1742.370 1200.020 1742.380 ;
        RECT 1377.020 1742.370 1380.020 1742.380 ;
        RECT 1557.020 1742.370 1560.020 1742.380 ;
        RECT 1737.020 1742.370 1740.020 1742.380 ;
        RECT 1917.020 1742.370 1920.020 1742.380 ;
        RECT 2097.020 1742.370 2100.020 1742.380 ;
        RECT 2277.020 1742.370 2280.020 1742.380 ;
        RECT 2457.020 1742.370 2460.020 1742.380 ;
        RECT 2637.020 1742.370 2640.020 1742.380 ;
        RECT 2817.020 1742.370 2820.020 1742.380 ;
        RECT 2940.700 1742.370 2943.700 1742.380 ;
        RECT -24.080 1565.380 -21.080 1565.390 ;
        RECT 117.020 1565.380 120.020 1565.390 ;
        RECT 297.020 1565.380 300.020 1565.390 ;
        RECT 477.020 1565.380 480.020 1565.390 ;
        RECT 657.020 1565.380 660.020 1565.390 ;
        RECT 837.020 1565.380 840.020 1565.390 ;
        RECT 1017.020 1565.380 1020.020 1565.390 ;
        RECT 1197.020 1565.380 1200.020 1565.390 ;
        RECT 1377.020 1565.380 1380.020 1565.390 ;
        RECT 1557.020 1565.380 1560.020 1565.390 ;
        RECT 1737.020 1565.380 1740.020 1565.390 ;
        RECT 1917.020 1565.380 1920.020 1565.390 ;
        RECT 2097.020 1565.380 2100.020 1565.390 ;
        RECT 2277.020 1565.380 2280.020 1565.390 ;
        RECT 2457.020 1565.380 2460.020 1565.390 ;
        RECT 2637.020 1565.380 2640.020 1565.390 ;
        RECT 2817.020 1565.380 2820.020 1565.390 ;
        RECT 2940.700 1565.380 2943.700 1565.390 ;
        RECT -24.080 1562.380 2943.700 1565.380 ;
        RECT -24.080 1562.370 -21.080 1562.380 ;
        RECT 117.020 1562.370 120.020 1562.380 ;
        RECT 297.020 1562.370 300.020 1562.380 ;
        RECT 477.020 1562.370 480.020 1562.380 ;
        RECT 657.020 1562.370 660.020 1562.380 ;
        RECT 837.020 1562.370 840.020 1562.380 ;
        RECT 1017.020 1562.370 1020.020 1562.380 ;
        RECT 1197.020 1562.370 1200.020 1562.380 ;
        RECT 1377.020 1562.370 1380.020 1562.380 ;
        RECT 1557.020 1562.370 1560.020 1562.380 ;
        RECT 1737.020 1562.370 1740.020 1562.380 ;
        RECT 1917.020 1562.370 1920.020 1562.380 ;
        RECT 2097.020 1562.370 2100.020 1562.380 ;
        RECT 2277.020 1562.370 2280.020 1562.380 ;
        RECT 2457.020 1562.370 2460.020 1562.380 ;
        RECT 2637.020 1562.370 2640.020 1562.380 ;
        RECT 2817.020 1562.370 2820.020 1562.380 ;
        RECT 2940.700 1562.370 2943.700 1562.380 ;
        RECT -24.080 1385.380 -21.080 1385.390 ;
        RECT 117.020 1385.380 120.020 1385.390 ;
        RECT 297.020 1385.380 300.020 1385.390 ;
        RECT 477.020 1385.380 480.020 1385.390 ;
        RECT 657.020 1385.380 660.020 1385.390 ;
        RECT 837.020 1385.380 840.020 1385.390 ;
        RECT 1017.020 1385.380 1020.020 1385.390 ;
        RECT 1197.020 1385.380 1200.020 1385.390 ;
        RECT 1377.020 1385.380 1380.020 1385.390 ;
        RECT 1557.020 1385.380 1560.020 1385.390 ;
        RECT 1737.020 1385.380 1740.020 1385.390 ;
        RECT 1917.020 1385.380 1920.020 1385.390 ;
        RECT 2097.020 1385.380 2100.020 1385.390 ;
        RECT 2277.020 1385.380 2280.020 1385.390 ;
        RECT 2457.020 1385.380 2460.020 1385.390 ;
        RECT 2637.020 1385.380 2640.020 1385.390 ;
        RECT 2817.020 1385.380 2820.020 1385.390 ;
        RECT 2940.700 1385.380 2943.700 1385.390 ;
        RECT -24.080 1382.380 2943.700 1385.380 ;
        RECT -24.080 1382.370 -21.080 1382.380 ;
        RECT 117.020 1382.370 120.020 1382.380 ;
        RECT 297.020 1382.370 300.020 1382.380 ;
        RECT 477.020 1382.370 480.020 1382.380 ;
        RECT 657.020 1382.370 660.020 1382.380 ;
        RECT 837.020 1382.370 840.020 1382.380 ;
        RECT 1017.020 1382.370 1020.020 1382.380 ;
        RECT 1197.020 1382.370 1200.020 1382.380 ;
        RECT 1377.020 1382.370 1380.020 1382.380 ;
        RECT 1557.020 1382.370 1560.020 1382.380 ;
        RECT 1737.020 1382.370 1740.020 1382.380 ;
        RECT 1917.020 1382.370 1920.020 1382.380 ;
        RECT 2097.020 1382.370 2100.020 1382.380 ;
        RECT 2277.020 1382.370 2280.020 1382.380 ;
        RECT 2457.020 1382.370 2460.020 1382.380 ;
        RECT 2637.020 1382.370 2640.020 1382.380 ;
        RECT 2817.020 1382.370 2820.020 1382.380 ;
        RECT 2940.700 1382.370 2943.700 1382.380 ;
        RECT -24.080 1205.380 -21.080 1205.390 ;
        RECT 117.020 1205.380 120.020 1205.390 ;
        RECT 297.020 1205.380 300.020 1205.390 ;
        RECT 477.020 1205.380 480.020 1205.390 ;
        RECT 657.020 1205.380 660.020 1205.390 ;
        RECT 837.020 1205.380 840.020 1205.390 ;
        RECT 1017.020 1205.380 1020.020 1205.390 ;
        RECT 1197.020 1205.380 1200.020 1205.390 ;
        RECT 1377.020 1205.380 1380.020 1205.390 ;
        RECT 1557.020 1205.380 1560.020 1205.390 ;
        RECT 1737.020 1205.380 1740.020 1205.390 ;
        RECT 1917.020 1205.380 1920.020 1205.390 ;
        RECT 2097.020 1205.380 2100.020 1205.390 ;
        RECT 2277.020 1205.380 2280.020 1205.390 ;
        RECT 2457.020 1205.380 2460.020 1205.390 ;
        RECT 2637.020 1205.380 2640.020 1205.390 ;
        RECT 2817.020 1205.380 2820.020 1205.390 ;
        RECT 2940.700 1205.380 2943.700 1205.390 ;
        RECT -24.080 1202.380 2943.700 1205.380 ;
        RECT -24.080 1202.370 -21.080 1202.380 ;
        RECT 117.020 1202.370 120.020 1202.380 ;
        RECT 297.020 1202.370 300.020 1202.380 ;
        RECT 477.020 1202.370 480.020 1202.380 ;
        RECT 657.020 1202.370 660.020 1202.380 ;
        RECT 837.020 1202.370 840.020 1202.380 ;
        RECT 1017.020 1202.370 1020.020 1202.380 ;
        RECT 1197.020 1202.370 1200.020 1202.380 ;
        RECT 1377.020 1202.370 1380.020 1202.380 ;
        RECT 1557.020 1202.370 1560.020 1202.380 ;
        RECT 1737.020 1202.370 1740.020 1202.380 ;
        RECT 1917.020 1202.370 1920.020 1202.380 ;
        RECT 2097.020 1202.370 2100.020 1202.380 ;
        RECT 2277.020 1202.370 2280.020 1202.380 ;
        RECT 2457.020 1202.370 2460.020 1202.380 ;
        RECT 2637.020 1202.370 2640.020 1202.380 ;
        RECT 2817.020 1202.370 2820.020 1202.380 ;
        RECT 2940.700 1202.370 2943.700 1202.380 ;
        RECT -24.080 1025.380 -21.080 1025.390 ;
        RECT 117.020 1025.380 120.020 1025.390 ;
        RECT 297.020 1025.380 300.020 1025.390 ;
        RECT 477.020 1025.380 480.020 1025.390 ;
        RECT 657.020 1025.380 660.020 1025.390 ;
        RECT 837.020 1025.380 840.020 1025.390 ;
        RECT 1017.020 1025.380 1020.020 1025.390 ;
        RECT 1197.020 1025.380 1200.020 1025.390 ;
        RECT 1377.020 1025.380 1380.020 1025.390 ;
        RECT 1557.020 1025.380 1560.020 1025.390 ;
        RECT 1737.020 1025.380 1740.020 1025.390 ;
        RECT 1917.020 1025.380 1920.020 1025.390 ;
        RECT 2097.020 1025.380 2100.020 1025.390 ;
        RECT 2277.020 1025.380 2280.020 1025.390 ;
        RECT 2457.020 1025.380 2460.020 1025.390 ;
        RECT 2637.020 1025.380 2640.020 1025.390 ;
        RECT 2817.020 1025.380 2820.020 1025.390 ;
        RECT 2940.700 1025.380 2943.700 1025.390 ;
        RECT -24.080 1022.380 2943.700 1025.380 ;
        RECT -24.080 1022.370 -21.080 1022.380 ;
        RECT 117.020 1022.370 120.020 1022.380 ;
        RECT 297.020 1022.370 300.020 1022.380 ;
        RECT 477.020 1022.370 480.020 1022.380 ;
        RECT 657.020 1022.370 660.020 1022.380 ;
        RECT 837.020 1022.370 840.020 1022.380 ;
        RECT 1017.020 1022.370 1020.020 1022.380 ;
        RECT 1197.020 1022.370 1200.020 1022.380 ;
        RECT 1377.020 1022.370 1380.020 1022.380 ;
        RECT 1557.020 1022.370 1560.020 1022.380 ;
        RECT 1737.020 1022.370 1740.020 1022.380 ;
        RECT 1917.020 1022.370 1920.020 1022.380 ;
        RECT 2097.020 1022.370 2100.020 1022.380 ;
        RECT 2277.020 1022.370 2280.020 1022.380 ;
        RECT 2457.020 1022.370 2460.020 1022.380 ;
        RECT 2637.020 1022.370 2640.020 1022.380 ;
        RECT 2817.020 1022.370 2820.020 1022.380 ;
        RECT 2940.700 1022.370 2943.700 1022.380 ;
        RECT -24.080 845.380 -21.080 845.390 ;
        RECT 117.020 845.380 120.020 845.390 ;
        RECT 297.020 845.380 300.020 845.390 ;
        RECT 477.020 845.380 480.020 845.390 ;
        RECT 657.020 845.380 660.020 845.390 ;
        RECT 837.020 845.380 840.020 845.390 ;
        RECT 1017.020 845.380 1020.020 845.390 ;
        RECT 1197.020 845.380 1200.020 845.390 ;
        RECT 1377.020 845.380 1380.020 845.390 ;
        RECT 1557.020 845.380 1560.020 845.390 ;
        RECT 1737.020 845.380 1740.020 845.390 ;
        RECT 1917.020 845.380 1920.020 845.390 ;
        RECT 2097.020 845.380 2100.020 845.390 ;
        RECT 2277.020 845.380 2280.020 845.390 ;
        RECT 2457.020 845.380 2460.020 845.390 ;
        RECT 2637.020 845.380 2640.020 845.390 ;
        RECT 2817.020 845.380 2820.020 845.390 ;
        RECT 2940.700 845.380 2943.700 845.390 ;
        RECT -24.080 842.380 2943.700 845.380 ;
        RECT -24.080 842.370 -21.080 842.380 ;
        RECT 117.020 842.370 120.020 842.380 ;
        RECT 297.020 842.370 300.020 842.380 ;
        RECT 477.020 842.370 480.020 842.380 ;
        RECT 657.020 842.370 660.020 842.380 ;
        RECT 837.020 842.370 840.020 842.380 ;
        RECT 1017.020 842.370 1020.020 842.380 ;
        RECT 1197.020 842.370 1200.020 842.380 ;
        RECT 1377.020 842.370 1380.020 842.380 ;
        RECT 1557.020 842.370 1560.020 842.380 ;
        RECT 1737.020 842.370 1740.020 842.380 ;
        RECT 1917.020 842.370 1920.020 842.380 ;
        RECT 2097.020 842.370 2100.020 842.380 ;
        RECT 2277.020 842.370 2280.020 842.380 ;
        RECT 2457.020 842.370 2460.020 842.380 ;
        RECT 2637.020 842.370 2640.020 842.380 ;
        RECT 2817.020 842.370 2820.020 842.380 ;
        RECT 2940.700 842.370 2943.700 842.380 ;
        RECT -24.080 665.380 -21.080 665.390 ;
        RECT 117.020 665.380 120.020 665.390 ;
        RECT 297.020 665.380 300.020 665.390 ;
        RECT 477.020 665.380 480.020 665.390 ;
        RECT 657.020 665.380 660.020 665.390 ;
        RECT 837.020 665.380 840.020 665.390 ;
        RECT 1017.020 665.380 1020.020 665.390 ;
        RECT 1197.020 665.380 1200.020 665.390 ;
        RECT 1377.020 665.380 1380.020 665.390 ;
        RECT 1557.020 665.380 1560.020 665.390 ;
        RECT 1737.020 665.380 1740.020 665.390 ;
        RECT 1917.020 665.380 1920.020 665.390 ;
        RECT 2097.020 665.380 2100.020 665.390 ;
        RECT 2277.020 665.380 2280.020 665.390 ;
        RECT 2457.020 665.380 2460.020 665.390 ;
        RECT 2637.020 665.380 2640.020 665.390 ;
        RECT 2817.020 665.380 2820.020 665.390 ;
        RECT 2940.700 665.380 2943.700 665.390 ;
        RECT -24.080 662.380 2943.700 665.380 ;
        RECT -24.080 662.370 -21.080 662.380 ;
        RECT 117.020 662.370 120.020 662.380 ;
        RECT 297.020 662.370 300.020 662.380 ;
        RECT 477.020 662.370 480.020 662.380 ;
        RECT 657.020 662.370 660.020 662.380 ;
        RECT 837.020 662.370 840.020 662.380 ;
        RECT 1017.020 662.370 1020.020 662.380 ;
        RECT 1197.020 662.370 1200.020 662.380 ;
        RECT 1377.020 662.370 1380.020 662.380 ;
        RECT 1557.020 662.370 1560.020 662.380 ;
        RECT 1737.020 662.370 1740.020 662.380 ;
        RECT 1917.020 662.370 1920.020 662.380 ;
        RECT 2097.020 662.370 2100.020 662.380 ;
        RECT 2277.020 662.370 2280.020 662.380 ;
        RECT 2457.020 662.370 2460.020 662.380 ;
        RECT 2637.020 662.370 2640.020 662.380 ;
        RECT 2817.020 662.370 2820.020 662.380 ;
        RECT 2940.700 662.370 2943.700 662.380 ;
        RECT -24.080 485.380 -21.080 485.390 ;
        RECT 117.020 485.380 120.020 485.390 ;
        RECT 297.020 485.380 300.020 485.390 ;
        RECT 477.020 485.380 480.020 485.390 ;
        RECT 657.020 485.380 660.020 485.390 ;
        RECT 837.020 485.380 840.020 485.390 ;
        RECT 1017.020 485.380 1020.020 485.390 ;
        RECT 1197.020 485.380 1200.020 485.390 ;
        RECT 1377.020 485.380 1380.020 485.390 ;
        RECT 1557.020 485.380 1560.020 485.390 ;
        RECT 1737.020 485.380 1740.020 485.390 ;
        RECT 1917.020 485.380 1920.020 485.390 ;
        RECT 2097.020 485.380 2100.020 485.390 ;
        RECT 2277.020 485.380 2280.020 485.390 ;
        RECT 2457.020 485.380 2460.020 485.390 ;
        RECT 2637.020 485.380 2640.020 485.390 ;
        RECT 2817.020 485.380 2820.020 485.390 ;
        RECT 2940.700 485.380 2943.700 485.390 ;
        RECT -24.080 482.380 2943.700 485.380 ;
        RECT -24.080 482.370 -21.080 482.380 ;
        RECT 117.020 482.370 120.020 482.380 ;
        RECT 297.020 482.370 300.020 482.380 ;
        RECT 477.020 482.370 480.020 482.380 ;
        RECT 657.020 482.370 660.020 482.380 ;
        RECT 837.020 482.370 840.020 482.380 ;
        RECT 1017.020 482.370 1020.020 482.380 ;
        RECT 1197.020 482.370 1200.020 482.380 ;
        RECT 1377.020 482.370 1380.020 482.380 ;
        RECT 1557.020 482.370 1560.020 482.380 ;
        RECT 1737.020 482.370 1740.020 482.380 ;
        RECT 1917.020 482.370 1920.020 482.380 ;
        RECT 2097.020 482.370 2100.020 482.380 ;
        RECT 2277.020 482.370 2280.020 482.380 ;
        RECT 2457.020 482.370 2460.020 482.380 ;
        RECT 2637.020 482.370 2640.020 482.380 ;
        RECT 2817.020 482.370 2820.020 482.380 ;
        RECT 2940.700 482.370 2943.700 482.380 ;
        RECT -24.080 305.380 -21.080 305.390 ;
        RECT 117.020 305.380 120.020 305.390 ;
        RECT 297.020 305.380 300.020 305.390 ;
        RECT 477.020 305.380 480.020 305.390 ;
        RECT 657.020 305.380 660.020 305.390 ;
        RECT 837.020 305.380 840.020 305.390 ;
        RECT 1017.020 305.380 1020.020 305.390 ;
        RECT 1197.020 305.380 1200.020 305.390 ;
        RECT 1377.020 305.380 1380.020 305.390 ;
        RECT 1557.020 305.380 1560.020 305.390 ;
        RECT 1737.020 305.380 1740.020 305.390 ;
        RECT 1917.020 305.380 1920.020 305.390 ;
        RECT 2097.020 305.380 2100.020 305.390 ;
        RECT 2277.020 305.380 2280.020 305.390 ;
        RECT 2457.020 305.380 2460.020 305.390 ;
        RECT 2637.020 305.380 2640.020 305.390 ;
        RECT 2817.020 305.380 2820.020 305.390 ;
        RECT 2940.700 305.380 2943.700 305.390 ;
        RECT -24.080 302.380 2943.700 305.380 ;
        RECT -24.080 302.370 -21.080 302.380 ;
        RECT 117.020 302.370 120.020 302.380 ;
        RECT 297.020 302.370 300.020 302.380 ;
        RECT 477.020 302.370 480.020 302.380 ;
        RECT 657.020 302.370 660.020 302.380 ;
        RECT 837.020 302.370 840.020 302.380 ;
        RECT 1017.020 302.370 1020.020 302.380 ;
        RECT 1197.020 302.370 1200.020 302.380 ;
        RECT 1377.020 302.370 1380.020 302.380 ;
        RECT 1557.020 302.370 1560.020 302.380 ;
        RECT 1737.020 302.370 1740.020 302.380 ;
        RECT 1917.020 302.370 1920.020 302.380 ;
        RECT 2097.020 302.370 2100.020 302.380 ;
        RECT 2277.020 302.370 2280.020 302.380 ;
        RECT 2457.020 302.370 2460.020 302.380 ;
        RECT 2637.020 302.370 2640.020 302.380 ;
        RECT 2817.020 302.370 2820.020 302.380 ;
        RECT 2940.700 302.370 2943.700 302.380 ;
        RECT -24.080 125.380 -21.080 125.390 ;
        RECT 117.020 125.380 120.020 125.390 ;
        RECT 297.020 125.380 300.020 125.390 ;
        RECT 477.020 125.380 480.020 125.390 ;
        RECT 657.020 125.380 660.020 125.390 ;
        RECT 837.020 125.380 840.020 125.390 ;
        RECT 1017.020 125.380 1020.020 125.390 ;
        RECT 1197.020 125.380 1200.020 125.390 ;
        RECT 1377.020 125.380 1380.020 125.390 ;
        RECT 1557.020 125.380 1560.020 125.390 ;
        RECT 1737.020 125.380 1740.020 125.390 ;
        RECT 1917.020 125.380 1920.020 125.390 ;
        RECT 2097.020 125.380 2100.020 125.390 ;
        RECT 2277.020 125.380 2280.020 125.390 ;
        RECT 2457.020 125.380 2460.020 125.390 ;
        RECT 2637.020 125.380 2640.020 125.390 ;
        RECT 2817.020 125.380 2820.020 125.390 ;
        RECT 2940.700 125.380 2943.700 125.390 ;
        RECT -24.080 122.380 2943.700 125.380 ;
        RECT -24.080 122.370 -21.080 122.380 ;
        RECT 117.020 122.370 120.020 122.380 ;
        RECT 297.020 122.370 300.020 122.380 ;
        RECT 477.020 122.370 480.020 122.380 ;
        RECT 657.020 122.370 660.020 122.380 ;
        RECT 837.020 122.370 840.020 122.380 ;
        RECT 1017.020 122.370 1020.020 122.380 ;
        RECT 1197.020 122.370 1200.020 122.380 ;
        RECT 1377.020 122.370 1380.020 122.380 ;
        RECT 1557.020 122.370 1560.020 122.380 ;
        RECT 1737.020 122.370 1740.020 122.380 ;
        RECT 1917.020 122.370 1920.020 122.380 ;
        RECT 2097.020 122.370 2100.020 122.380 ;
        RECT 2277.020 122.370 2280.020 122.380 ;
        RECT 2457.020 122.370 2460.020 122.380 ;
        RECT 2637.020 122.370 2640.020 122.380 ;
        RECT 2817.020 122.370 2820.020 122.380 ;
        RECT 2940.700 122.370 2943.700 122.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 117.020 -15.720 120.020 -15.710 ;
        RECT 297.020 -15.720 300.020 -15.710 ;
        RECT 477.020 -15.720 480.020 -15.710 ;
        RECT 657.020 -15.720 660.020 -15.710 ;
        RECT 837.020 -15.720 840.020 -15.710 ;
        RECT 1017.020 -15.720 1020.020 -15.710 ;
        RECT 1197.020 -15.720 1200.020 -15.710 ;
        RECT 1377.020 -15.720 1380.020 -15.710 ;
        RECT 1557.020 -15.720 1560.020 -15.710 ;
        RECT 1737.020 -15.720 1740.020 -15.710 ;
        RECT 1917.020 -15.720 1920.020 -15.710 ;
        RECT 2097.020 -15.720 2100.020 -15.710 ;
        RECT 2277.020 -15.720 2280.020 -15.710 ;
        RECT 2457.020 -15.720 2460.020 -15.710 ;
        RECT 2637.020 -15.720 2640.020 -15.710 ;
        RECT 2817.020 -15.720 2820.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 117.020 -18.730 120.020 -18.720 ;
        RECT 297.020 -18.730 300.020 -18.720 ;
        RECT 477.020 -18.730 480.020 -18.720 ;
        RECT 657.020 -18.730 660.020 -18.720 ;
        RECT 837.020 -18.730 840.020 -18.720 ;
        RECT 1017.020 -18.730 1020.020 -18.720 ;
        RECT 1197.020 -18.730 1200.020 -18.720 ;
        RECT 1377.020 -18.730 1380.020 -18.720 ;
        RECT 1557.020 -18.730 1560.020 -18.720 ;
        RECT 1737.020 -18.730 1740.020 -18.720 ;
        RECT 1917.020 -18.730 1920.020 -18.720 ;
        RECT 2097.020 -18.730 2100.020 -18.720 ;
        RECT 2277.020 -18.730 2280.020 -18.720 ;
        RECT 2457.020 -18.730 2460.020 -18.720 ;
        RECT 2637.020 -18.730 2640.020 -18.720 ;
        RECT 2817.020 -18.730 2820.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 45.020 -28.120 48.020 3547.800 ;
        RECT 225.020 -28.120 228.020 3547.800 ;
        RECT 405.020 -28.120 408.020 3547.800 ;
        RECT 585.020 -28.120 588.020 3547.800 ;
        RECT 765.020 -28.120 768.020 3547.800 ;
        RECT 945.020 -28.120 948.020 3547.800 ;
        RECT 1125.020 -28.120 1128.020 3547.800 ;
        RECT 1305.020 -28.120 1308.020 3547.800 ;
        RECT 1485.020 -28.120 1488.020 3547.800 ;
        RECT 1665.020 -28.120 1668.020 3547.800 ;
        RECT 1845.020 -28.120 1848.020 3547.800 ;
        RECT 2025.020 -28.120 2028.020 3547.800 ;
        RECT 2205.020 -28.120 2208.020 3547.800 ;
        RECT 2385.020 -28.120 2388.020 3547.800 ;
        RECT 2565.020 -28.120 2568.020 3547.800 ;
        RECT 2745.020 -28.120 2748.020 3547.800 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 3472.090 -26.690 3473.270 ;
        RECT -27.870 3470.490 -26.690 3471.670 ;
        RECT -27.870 3292.090 -26.690 3293.270 ;
        RECT -27.870 3290.490 -26.690 3291.670 ;
        RECT -27.870 3112.090 -26.690 3113.270 ;
        RECT -27.870 3110.490 -26.690 3111.670 ;
        RECT -27.870 2932.090 -26.690 2933.270 ;
        RECT -27.870 2930.490 -26.690 2931.670 ;
        RECT -27.870 2752.090 -26.690 2753.270 ;
        RECT -27.870 2750.490 -26.690 2751.670 ;
        RECT -27.870 2572.090 -26.690 2573.270 ;
        RECT -27.870 2570.490 -26.690 2571.670 ;
        RECT -27.870 2392.090 -26.690 2393.270 ;
        RECT -27.870 2390.490 -26.690 2391.670 ;
        RECT -27.870 2212.090 -26.690 2213.270 ;
        RECT -27.870 2210.490 -26.690 2211.670 ;
        RECT -27.870 2032.090 -26.690 2033.270 ;
        RECT -27.870 2030.490 -26.690 2031.670 ;
        RECT -27.870 1852.090 -26.690 1853.270 ;
        RECT -27.870 1850.490 -26.690 1851.670 ;
        RECT -27.870 1672.090 -26.690 1673.270 ;
        RECT -27.870 1670.490 -26.690 1671.670 ;
        RECT -27.870 1492.090 -26.690 1493.270 ;
        RECT -27.870 1490.490 -26.690 1491.670 ;
        RECT -27.870 1312.090 -26.690 1313.270 ;
        RECT -27.870 1310.490 -26.690 1311.670 ;
        RECT -27.870 1132.090 -26.690 1133.270 ;
        RECT -27.870 1130.490 -26.690 1131.670 ;
        RECT -27.870 952.090 -26.690 953.270 ;
        RECT -27.870 950.490 -26.690 951.670 ;
        RECT -27.870 772.090 -26.690 773.270 ;
        RECT -27.870 770.490 -26.690 771.670 ;
        RECT -27.870 592.090 -26.690 593.270 ;
        RECT -27.870 590.490 -26.690 591.670 ;
        RECT -27.870 412.090 -26.690 413.270 ;
        RECT -27.870 410.490 -26.690 411.670 ;
        RECT -27.870 232.090 -26.690 233.270 ;
        RECT -27.870 230.490 -26.690 231.670 ;
        RECT -27.870 52.090 -26.690 53.270 ;
        RECT -27.870 50.490 -26.690 51.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 45.930 3541.810 47.110 3542.990 ;
        RECT 45.930 3540.210 47.110 3541.390 ;
        RECT 45.930 3472.090 47.110 3473.270 ;
        RECT 45.930 3470.490 47.110 3471.670 ;
        RECT 45.930 3292.090 47.110 3293.270 ;
        RECT 45.930 3290.490 47.110 3291.670 ;
        RECT 45.930 3112.090 47.110 3113.270 ;
        RECT 45.930 3110.490 47.110 3111.670 ;
        RECT 45.930 2932.090 47.110 2933.270 ;
        RECT 45.930 2930.490 47.110 2931.670 ;
        RECT 45.930 2752.090 47.110 2753.270 ;
        RECT 45.930 2750.490 47.110 2751.670 ;
        RECT 45.930 2572.090 47.110 2573.270 ;
        RECT 45.930 2570.490 47.110 2571.670 ;
        RECT 45.930 2392.090 47.110 2393.270 ;
        RECT 45.930 2390.490 47.110 2391.670 ;
        RECT 45.930 2212.090 47.110 2213.270 ;
        RECT 45.930 2210.490 47.110 2211.670 ;
        RECT 45.930 2032.090 47.110 2033.270 ;
        RECT 45.930 2030.490 47.110 2031.670 ;
        RECT 45.930 1852.090 47.110 1853.270 ;
        RECT 45.930 1850.490 47.110 1851.670 ;
        RECT 45.930 1672.090 47.110 1673.270 ;
        RECT 45.930 1670.490 47.110 1671.670 ;
        RECT 45.930 1492.090 47.110 1493.270 ;
        RECT 45.930 1490.490 47.110 1491.670 ;
        RECT 45.930 1312.090 47.110 1313.270 ;
        RECT 45.930 1310.490 47.110 1311.670 ;
        RECT 45.930 1132.090 47.110 1133.270 ;
        RECT 45.930 1130.490 47.110 1131.670 ;
        RECT 45.930 952.090 47.110 953.270 ;
        RECT 45.930 950.490 47.110 951.670 ;
        RECT 45.930 772.090 47.110 773.270 ;
        RECT 45.930 770.490 47.110 771.670 ;
        RECT 45.930 592.090 47.110 593.270 ;
        RECT 45.930 590.490 47.110 591.670 ;
        RECT 45.930 412.090 47.110 413.270 ;
        RECT 45.930 410.490 47.110 411.670 ;
        RECT 45.930 232.090 47.110 233.270 ;
        RECT 45.930 230.490 47.110 231.670 ;
        RECT 45.930 52.090 47.110 53.270 ;
        RECT 45.930 50.490 47.110 51.670 ;
        RECT 45.930 -21.710 47.110 -20.530 ;
        RECT 45.930 -23.310 47.110 -22.130 ;
        RECT 225.930 3541.810 227.110 3542.990 ;
        RECT 225.930 3540.210 227.110 3541.390 ;
        RECT 225.930 3472.090 227.110 3473.270 ;
        RECT 225.930 3470.490 227.110 3471.670 ;
        RECT 225.930 3292.090 227.110 3293.270 ;
        RECT 225.930 3290.490 227.110 3291.670 ;
        RECT 225.930 3112.090 227.110 3113.270 ;
        RECT 225.930 3110.490 227.110 3111.670 ;
        RECT 225.930 2932.090 227.110 2933.270 ;
        RECT 225.930 2930.490 227.110 2931.670 ;
        RECT 225.930 2752.090 227.110 2753.270 ;
        RECT 225.930 2750.490 227.110 2751.670 ;
        RECT 225.930 2572.090 227.110 2573.270 ;
        RECT 225.930 2570.490 227.110 2571.670 ;
        RECT 225.930 2392.090 227.110 2393.270 ;
        RECT 225.930 2390.490 227.110 2391.670 ;
        RECT 225.930 2212.090 227.110 2213.270 ;
        RECT 225.930 2210.490 227.110 2211.670 ;
        RECT 225.930 2032.090 227.110 2033.270 ;
        RECT 225.930 2030.490 227.110 2031.670 ;
        RECT 225.930 1852.090 227.110 1853.270 ;
        RECT 225.930 1850.490 227.110 1851.670 ;
        RECT 225.930 1672.090 227.110 1673.270 ;
        RECT 225.930 1670.490 227.110 1671.670 ;
        RECT 225.930 1492.090 227.110 1493.270 ;
        RECT 225.930 1490.490 227.110 1491.670 ;
        RECT 225.930 1312.090 227.110 1313.270 ;
        RECT 225.930 1310.490 227.110 1311.670 ;
        RECT 225.930 1132.090 227.110 1133.270 ;
        RECT 225.930 1130.490 227.110 1131.670 ;
        RECT 225.930 952.090 227.110 953.270 ;
        RECT 225.930 950.490 227.110 951.670 ;
        RECT 225.930 772.090 227.110 773.270 ;
        RECT 225.930 770.490 227.110 771.670 ;
        RECT 225.930 592.090 227.110 593.270 ;
        RECT 225.930 590.490 227.110 591.670 ;
        RECT 225.930 412.090 227.110 413.270 ;
        RECT 225.930 410.490 227.110 411.670 ;
        RECT 225.930 232.090 227.110 233.270 ;
        RECT 225.930 230.490 227.110 231.670 ;
        RECT 225.930 52.090 227.110 53.270 ;
        RECT 225.930 50.490 227.110 51.670 ;
        RECT 225.930 -21.710 227.110 -20.530 ;
        RECT 225.930 -23.310 227.110 -22.130 ;
        RECT 405.930 3541.810 407.110 3542.990 ;
        RECT 405.930 3540.210 407.110 3541.390 ;
        RECT 405.930 3472.090 407.110 3473.270 ;
        RECT 405.930 3470.490 407.110 3471.670 ;
        RECT 405.930 3292.090 407.110 3293.270 ;
        RECT 405.930 3290.490 407.110 3291.670 ;
        RECT 405.930 3112.090 407.110 3113.270 ;
        RECT 405.930 3110.490 407.110 3111.670 ;
        RECT 405.930 2932.090 407.110 2933.270 ;
        RECT 405.930 2930.490 407.110 2931.670 ;
        RECT 405.930 2752.090 407.110 2753.270 ;
        RECT 405.930 2750.490 407.110 2751.670 ;
        RECT 405.930 2572.090 407.110 2573.270 ;
        RECT 405.930 2570.490 407.110 2571.670 ;
        RECT 405.930 2392.090 407.110 2393.270 ;
        RECT 405.930 2390.490 407.110 2391.670 ;
        RECT 405.930 2212.090 407.110 2213.270 ;
        RECT 405.930 2210.490 407.110 2211.670 ;
        RECT 405.930 2032.090 407.110 2033.270 ;
        RECT 405.930 2030.490 407.110 2031.670 ;
        RECT 405.930 1852.090 407.110 1853.270 ;
        RECT 405.930 1850.490 407.110 1851.670 ;
        RECT 405.930 1672.090 407.110 1673.270 ;
        RECT 405.930 1670.490 407.110 1671.670 ;
        RECT 405.930 1492.090 407.110 1493.270 ;
        RECT 405.930 1490.490 407.110 1491.670 ;
        RECT 405.930 1312.090 407.110 1313.270 ;
        RECT 405.930 1310.490 407.110 1311.670 ;
        RECT 405.930 1132.090 407.110 1133.270 ;
        RECT 405.930 1130.490 407.110 1131.670 ;
        RECT 405.930 952.090 407.110 953.270 ;
        RECT 405.930 950.490 407.110 951.670 ;
        RECT 405.930 772.090 407.110 773.270 ;
        RECT 405.930 770.490 407.110 771.670 ;
        RECT 405.930 592.090 407.110 593.270 ;
        RECT 405.930 590.490 407.110 591.670 ;
        RECT 405.930 412.090 407.110 413.270 ;
        RECT 405.930 410.490 407.110 411.670 ;
        RECT 405.930 232.090 407.110 233.270 ;
        RECT 405.930 230.490 407.110 231.670 ;
        RECT 405.930 52.090 407.110 53.270 ;
        RECT 405.930 50.490 407.110 51.670 ;
        RECT 405.930 -21.710 407.110 -20.530 ;
        RECT 405.930 -23.310 407.110 -22.130 ;
        RECT 585.930 3541.810 587.110 3542.990 ;
        RECT 585.930 3540.210 587.110 3541.390 ;
        RECT 585.930 3472.090 587.110 3473.270 ;
        RECT 585.930 3470.490 587.110 3471.670 ;
        RECT 585.930 3292.090 587.110 3293.270 ;
        RECT 585.930 3290.490 587.110 3291.670 ;
        RECT 585.930 3112.090 587.110 3113.270 ;
        RECT 585.930 3110.490 587.110 3111.670 ;
        RECT 585.930 2932.090 587.110 2933.270 ;
        RECT 585.930 2930.490 587.110 2931.670 ;
        RECT 585.930 2752.090 587.110 2753.270 ;
        RECT 585.930 2750.490 587.110 2751.670 ;
        RECT 585.930 2572.090 587.110 2573.270 ;
        RECT 585.930 2570.490 587.110 2571.670 ;
        RECT 585.930 2392.090 587.110 2393.270 ;
        RECT 585.930 2390.490 587.110 2391.670 ;
        RECT 585.930 2212.090 587.110 2213.270 ;
        RECT 585.930 2210.490 587.110 2211.670 ;
        RECT 585.930 2032.090 587.110 2033.270 ;
        RECT 585.930 2030.490 587.110 2031.670 ;
        RECT 585.930 1852.090 587.110 1853.270 ;
        RECT 585.930 1850.490 587.110 1851.670 ;
        RECT 585.930 1672.090 587.110 1673.270 ;
        RECT 585.930 1670.490 587.110 1671.670 ;
        RECT 585.930 1492.090 587.110 1493.270 ;
        RECT 585.930 1490.490 587.110 1491.670 ;
        RECT 585.930 1312.090 587.110 1313.270 ;
        RECT 585.930 1310.490 587.110 1311.670 ;
        RECT 585.930 1132.090 587.110 1133.270 ;
        RECT 585.930 1130.490 587.110 1131.670 ;
        RECT 585.930 952.090 587.110 953.270 ;
        RECT 585.930 950.490 587.110 951.670 ;
        RECT 585.930 772.090 587.110 773.270 ;
        RECT 585.930 770.490 587.110 771.670 ;
        RECT 585.930 592.090 587.110 593.270 ;
        RECT 585.930 590.490 587.110 591.670 ;
        RECT 585.930 412.090 587.110 413.270 ;
        RECT 585.930 410.490 587.110 411.670 ;
        RECT 585.930 232.090 587.110 233.270 ;
        RECT 585.930 230.490 587.110 231.670 ;
        RECT 585.930 52.090 587.110 53.270 ;
        RECT 585.930 50.490 587.110 51.670 ;
        RECT 585.930 -21.710 587.110 -20.530 ;
        RECT 585.930 -23.310 587.110 -22.130 ;
        RECT 765.930 3541.810 767.110 3542.990 ;
        RECT 765.930 3540.210 767.110 3541.390 ;
        RECT 765.930 3472.090 767.110 3473.270 ;
        RECT 765.930 3470.490 767.110 3471.670 ;
        RECT 765.930 3292.090 767.110 3293.270 ;
        RECT 765.930 3290.490 767.110 3291.670 ;
        RECT 765.930 3112.090 767.110 3113.270 ;
        RECT 765.930 3110.490 767.110 3111.670 ;
        RECT 765.930 2932.090 767.110 2933.270 ;
        RECT 765.930 2930.490 767.110 2931.670 ;
        RECT 765.930 2752.090 767.110 2753.270 ;
        RECT 765.930 2750.490 767.110 2751.670 ;
        RECT 765.930 2572.090 767.110 2573.270 ;
        RECT 765.930 2570.490 767.110 2571.670 ;
        RECT 765.930 2392.090 767.110 2393.270 ;
        RECT 765.930 2390.490 767.110 2391.670 ;
        RECT 765.930 2212.090 767.110 2213.270 ;
        RECT 765.930 2210.490 767.110 2211.670 ;
        RECT 765.930 2032.090 767.110 2033.270 ;
        RECT 765.930 2030.490 767.110 2031.670 ;
        RECT 765.930 1852.090 767.110 1853.270 ;
        RECT 765.930 1850.490 767.110 1851.670 ;
        RECT 765.930 1672.090 767.110 1673.270 ;
        RECT 765.930 1670.490 767.110 1671.670 ;
        RECT 765.930 1492.090 767.110 1493.270 ;
        RECT 765.930 1490.490 767.110 1491.670 ;
        RECT 765.930 1312.090 767.110 1313.270 ;
        RECT 765.930 1310.490 767.110 1311.670 ;
        RECT 765.930 1132.090 767.110 1133.270 ;
        RECT 765.930 1130.490 767.110 1131.670 ;
        RECT 765.930 952.090 767.110 953.270 ;
        RECT 765.930 950.490 767.110 951.670 ;
        RECT 765.930 772.090 767.110 773.270 ;
        RECT 765.930 770.490 767.110 771.670 ;
        RECT 765.930 592.090 767.110 593.270 ;
        RECT 765.930 590.490 767.110 591.670 ;
        RECT 765.930 412.090 767.110 413.270 ;
        RECT 765.930 410.490 767.110 411.670 ;
        RECT 765.930 232.090 767.110 233.270 ;
        RECT 765.930 230.490 767.110 231.670 ;
        RECT 765.930 52.090 767.110 53.270 ;
        RECT 765.930 50.490 767.110 51.670 ;
        RECT 765.930 -21.710 767.110 -20.530 ;
        RECT 765.930 -23.310 767.110 -22.130 ;
        RECT 945.930 3541.810 947.110 3542.990 ;
        RECT 945.930 3540.210 947.110 3541.390 ;
        RECT 945.930 3472.090 947.110 3473.270 ;
        RECT 945.930 3470.490 947.110 3471.670 ;
        RECT 945.930 3292.090 947.110 3293.270 ;
        RECT 945.930 3290.490 947.110 3291.670 ;
        RECT 945.930 3112.090 947.110 3113.270 ;
        RECT 945.930 3110.490 947.110 3111.670 ;
        RECT 945.930 2932.090 947.110 2933.270 ;
        RECT 945.930 2930.490 947.110 2931.670 ;
        RECT 945.930 2752.090 947.110 2753.270 ;
        RECT 945.930 2750.490 947.110 2751.670 ;
        RECT 945.930 2572.090 947.110 2573.270 ;
        RECT 945.930 2570.490 947.110 2571.670 ;
        RECT 945.930 2392.090 947.110 2393.270 ;
        RECT 945.930 2390.490 947.110 2391.670 ;
        RECT 945.930 2212.090 947.110 2213.270 ;
        RECT 945.930 2210.490 947.110 2211.670 ;
        RECT 945.930 2032.090 947.110 2033.270 ;
        RECT 945.930 2030.490 947.110 2031.670 ;
        RECT 945.930 1852.090 947.110 1853.270 ;
        RECT 945.930 1850.490 947.110 1851.670 ;
        RECT 945.930 1672.090 947.110 1673.270 ;
        RECT 945.930 1670.490 947.110 1671.670 ;
        RECT 945.930 1492.090 947.110 1493.270 ;
        RECT 945.930 1490.490 947.110 1491.670 ;
        RECT 945.930 1312.090 947.110 1313.270 ;
        RECT 945.930 1310.490 947.110 1311.670 ;
        RECT 945.930 1132.090 947.110 1133.270 ;
        RECT 945.930 1130.490 947.110 1131.670 ;
        RECT 945.930 952.090 947.110 953.270 ;
        RECT 945.930 950.490 947.110 951.670 ;
        RECT 945.930 772.090 947.110 773.270 ;
        RECT 945.930 770.490 947.110 771.670 ;
        RECT 945.930 592.090 947.110 593.270 ;
        RECT 945.930 590.490 947.110 591.670 ;
        RECT 945.930 412.090 947.110 413.270 ;
        RECT 945.930 410.490 947.110 411.670 ;
        RECT 945.930 232.090 947.110 233.270 ;
        RECT 945.930 230.490 947.110 231.670 ;
        RECT 945.930 52.090 947.110 53.270 ;
        RECT 945.930 50.490 947.110 51.670 ;
        RECT 945.930 -21.710 947.110 -20.530 ;
        RECT 945.930 -23.310 947.110 -22.130 ;
        RECT 1125.930 3541.810 1127.110 3542.990 ;
        RECT 1125.930 3540.210 1127.110 3541.390 ;
        RECT 1125.930 3472.090 1127.110 3473.270 ;
        RECT 1125.930 3470.490 1127.110 3471.670 ;
        RECT 1125.930 3292.090 1127.110 3293.270 ;
        RECT 1125.930 3290.490 1127.110 3291.670 ;
        RECT 1125.930 3112.090 1127.110 3113.270 ;
        RECT 1125.930 3110.490 1127.110 3111.670 ;
        RECT 1125.930 2932.090 1127.110 2933.270 ;
        RECT 1125.930 2930.490 1127.110 2931.670 ;
        RECT 1125.930 2752.090 1127.110 2753.270 ;
        RECT 1125.930 2750.490 1127.110 2751.670 ;
        RECT 1125.930 2572.090 1127.110 2573.270 ;
        RECT 1125.930 2570.490 1127.110 2571.670 ;
        RECT 1125.930 2392.090 1127.110 2393.270 ;
        RECT 1125.930 2390.490 1127.110 2391.670 ;
        RECT 1125.930 2212.090 1127.110 2213.270 ;
        RECT 1125.930 2210.490 1127.110 2211.670 ;
        RECT 1125.930 2032.090 1127.110 2033.270 ;
        RECT 1125.930 2030.490 1127.110 2031.670 ;
        RECT 1125.930 1852.090 1127.110 1853.270 ;
        RECT 1125.930 1850.490 1127.110 1851.670 ;
        RECT 1125.930 1672.090 1127.110 1673.270 ;
        RECT 1125.930 1670.490 1127.110 1671.670 ;
        RECT 1125.930 1492.090 1127.110 1493.270 ;
        RECT 1125.930 1490.490 1127.110 1491.670 ;
        RECT 1125.930 1312.090 1127.110 1313.270 ;
        RECT 1125.930 1310.490 1127.110 1311.670 ;
        RECT 1125.930 1132.090 1127.110 1133.270 ;
        RECT 1125.930 1130.490 1127.110 1131.670 ;
        RECT 1125.930 952.090 1127.110 953.270 ;
        RECT 1125.930 950.490 1127.110 951.670 ;
        RECT 1125.930 772.090 1127.110 773.270 ;
        RECT 1125.930 770.490 1127.110 771.670 ;
        RECT 1125.930 592.090 1127.110 593.270 ;
        RECT 1125.930 590.490 1127.110 591.670 ;
        RECT 1125.930 412.090 1127.110 413.270 ;
        RECT 1125.930 410.490 1127.110 411.670 ;
        RECT 1125.930 232.090 1127.110 233.270 ;
        RECT 1125.930 230.490 1127.110 231.670 ;
        RECT 1125.930 52.090 1127.110 53.270 ;
        RECT 1125.930 50.490 1127.110 51.670 ;
        RECT 1125.930 -21.710 1127.110 -20.530 ;
        RECT 1125.930 -23.310 1127.110 -22.130 ;
        RECT 1305.930 3541.810 1307.110 3542.990 ;
        RECT 1305.930 3540.210 1307.110 3541.390 ;
        RECT 1305.930 3472.090 1307.110 3473.270 ;
        RECT 1305.930 3470.490 1307.110 3471.670 ;
        RECT 1305.930 3292.090 1307.110 3293.270 ;
        RECT 1305.930 3290.490 1307.110 3291.670 ;
        RECT 1305.930 3112.090 1307.110 3113.270 ;
        RECT 1305.930 3110.490 1307.110 3111.670 ;
        RECT 1305.930 2932.090 1307.110 2933.270 ;
        RECT 1305.930 2930.490 1307.110 2931.670 ;
        RECT 1305.930 2752.090 1307.110 2753.270 ;
        RECT 1305.930 2750.490 1307.110 2751.670 ;
        RECT 1305.930 2572.090 1307.110 2573.270 ;
        RECT 1305.930 2570.490 1307.110 2571.670 ;
        RECT 1305.930 2392.090 1307.110 2393.270 ;
        RECT 1305.930 2390.490 1307.110 2391.670 ;
        RECT 1305.930 2212.090 1307.110 2213.270 ;
        RECT 1305.930 2210.490 1307.110 2211.670 ;
        RECT 1305.930 2032.090 1307.110 2033.270 ;
        RECT 1305.930 2030.490 1307.110 2031.670 ;
        RECT 1305.930 1852.090 1307.110 1853.270 ;
        RECT 1305.930 1850.490 1307.110 1851.670 ;
        RECT 1305.930 1672.090 1307.110 1673.270 ;
        RECT 1305.930 1670.490 1307.110 1671.670 ;
        RECT 1305.930 1492.090 1307.110 1493.270 ;
        RECT 1305.930 1490.490 1307.110 1491.670 ;
        RECT 1305.930 1312.090 1307.110 1313.270 ;
        RECT 1305.930 1310.490 1307.110 1311.670 ;
        RECT 1305.930 1132.090 1307.110 1133.270 ;
        RECT 1305.930 1130.490 1307.110 1131.670 ;
        RECT 1305.930 952.090 1307.110 953.270 ;
        RECT 1305.930 950.490 1307.110 951.670 ;
        RECT 1305.930 772.090 1307.110 773.270 ;
        RECT 1305.930 770.490 1307.110 771.670 ;
        RECT 1305.930 592.090 1307.110 593.270 ;
        RECT 1305.930 590.490 1307.110 591.670 ;
        RECT 1305.930 412.090 1307.110 413.270 ;
        RECT 1305.930 410.490 1307.110 411.670 ;
        RECT 1305.930 232.090 1307.110 233.270 ;
        RECT 1305.930 230.490 1307.110 231.670 ;
        RECT 1305.930 52.090 1307.110 53.270 ;
        RECT 1305.930 50.490 1307.110 51.670 ;
        RECT 1305.930 -21.710 1307.110 -20.530 ;
        RECT 1305.930 -23.310 1307.110 -22.130 ;
        RECT 1485.930 3541.810 1487.110 3542.990 ;
        RECT 1485.930 3540.210 1487.110 3541.390 ;
        RECT 1485.930 3472.090 1487.110 3473.270 ;
        RECT 1485.930 3470.490 1487.110 3471.670 ;
        RECT 1485.930 3292.090 1487.110 3293.270 ;
        RECT 1485.930 3290.490 1487.110 3291.670 ;
        RECT 1485.930 3112.090 1487.110 3113.270 ;
        RECT 1485.930 3110.490 1487.110 3111.670 ;
        RECT 1485.930 2932.090 1487.110 2933.270 ;
        RECT 1485.930 2930.490 1487.110 2931.670 ;
        RECT 1485.930 2752.090 1487.110 2753.270 ;
        RECT 1485.930 2750.490 1487.110 2751.670 ;
        RECT 1485.930 2572.090 1487.110 2573.270 ;
        RECT 1485.930 2570.490 1487.110 2571.670 ;
        RECT 1485.930 2392.090 1487.110 2393.270 ;
        RECT 1485.930 2390.490 1487.110 2391.670 ;
        RECT 1485.930 2212.090 1487.110 2213.270 ;
        RECT 1485.930 2210.490 1487.110 2211.670 ;
        RECT 1485.930 2032.090 1487.110 2033.270 ;
        RECT 1485.930 2030.490 1487.110 2031.670 ;
        RECT 1485.930 1852.090 1487.110 1853.270 ;
        RECT 1485.930 1850.490 1487.110 1851.670 ;
        RECT 1485.930 1672.090 1487.110 1673.270 ;
        RECT 1485.930 1670.490 1487.110 1671.670 ;
        RECT 1485.930 1492.090 1487.110 1493.270 ;
        RECT 1485.930 1490.490 1487.110 1491.670 ;
        RECT 1485.930 1312.090 1487.110 1313.270 ;
        RECT 1485.930 1310.490 1487.110 1311.670 ;
        RECT 1485.930 1132.090 1487.110 1133.270 ;
        RECT 1485.930 1130.490 1487.110 1131.670 ;
        RECT 1485.930 952.090 1487.110 953.270 ;
        RECT 1485.930 950.490 1487.110 951.670 ;
        RECT 1485.930 772.090 1487.110 773.270 ;
        RECT 1485.930 770.490 1487.110 771.670 ;
        RECT 1485.930 592.090 1487.110 593.270 ;
        RECT 1485.930 590.490 1487.110 591.670 ;
        RECT 1485.930 412.090 1487.110 413.270 ;
        RECT 1485.930 410.490 1487.110 411.670 ;
        RECT 1485.930 232.090 1487.110 233.270 ;
        RECT 1485.930 230.490 1487.110 231.670 ;
        RECT 1485.930 52.090 1487.110 53.270 ;
        RECT 1485.930 50.490 1487.110 51.670 ;
        RECT 1485.930 -21.710 1487.110 -20.530 ;
        RECT 1485.930 -23.310 1487.110 -22.130 ;
        RECT 1665.930 3541.810 1667.110 3542.990 ;
        RECT 1665.930 3540.210 1667.110 3541.390 ;
        RECT 1665.930 3472.090 1667.110 3473.270 ;
        RECT 1665.930 3470.490 1667.110 3471.670 ;
        RECT 1665.930 3292.090 1667.110 3293.270 ;
        RECT 1665.930 3290.490 1667.110 3291.670 ;
        RECT 1665.930 3112.090 1667.110 3113.270 ;
        RECT 1665.930 3110.490 1667.110 3111.670 ;
        RECT 1665.930 2932.090 1667.110 2933.270 ;
        RECT 1665.930 2930.490 1667.110 2931.670 ;
        RECT 1665.930 2752.090 1667.110 2753.270 ;
        RECT 1665.930 2750.490 1667.110 2751.670 ;
        RECT 1665.930 2572.090 1667.110 2573.270 ;
        RECT 1665.930 2570.490 1667.110 2571.670 ;
        RECT 1665.930 2392.090 1667.110 2393.270 ;
        RECT 1665.930 2390.490 1667.110 2391.670 ;
        RECT 1665.930 2212.090 1667.110 2213.270 ;
        RECT 1665.930 2210.490 1667.110 2211.670 ;
        RECT 1665.930 2032.090 1667.110 2033.270 ;
        RECT 1665.930 2030.490 1667.110 2031.670 ;
        RECT 1665.930 1852.090 1667.110 1853.270 ;
        RECT 1665.930 1850.490 1667.110 1851.670 ;
        RECT 1665.930 1672.090 1667.110 1673.270 ;
        RECT 1665.930 1670.490 1667.110 1671.670 ;
        RECT 1665.930 1492.090 1667.110 1493.270 ;
        RECT 1665.930 1490.490 1667.110 1491.670 ;
        RECT 1665.930 1312.090 1667.110 1313.270 ;
        RECT 1665.930 1310.490 1667.110 1311.670 ;
        RECT 1665.930 1132.090 1667.110 1133.270 ;
        RECT 1665.930 1130.490 1667.110 1131.670 ;
        RECT 1665.930 952.090 1667.110 953.270 ;
        RECT 1665.930 950.490 1667.110 951.670 ;
        RECT 1665.930 772.090 1667.110 773.270 ;
        RECT 1665.930 770.490 1667.110 771.670 ;
        RECT 1665.930 592.090 1667.110 593.270 ;
        RECT 1665.930 590.490 1667.110 591.670 ;
        RECT 1665.930 412.090 1667.110 413.270 ;
        RECT 1665.930 410.490 1667.110 411.670 ;
        RECT 1665.930 232.090 1667.110 233.270 ;
        RECT 1665.930 230.490 1667.110 231.670 ;
        RECT 1665.930 52.090 1667.110 53.270 ;
        RECT 1665.930 50.490 1667.110 51.670 ;
        RECT 1665.930 -21.710 1667.110 -20.530 ;
        RECT 1665.930 -23.310 1667.110 -22.130 ;
        RECT 1845.930 3541.810 1847.110 3542.990 ;
        RECT 1845.930 3540.210 1847.110 3541.390 ;
        RECT 1845.930 3472.090 1847.110 3473.270 ;
        RECT 1845.930 3470.490 1847.110 3471.670 ;
        RECT 1845.930 3292.090 1847.110 3293.270 ;
        RECT 1845.930 3290.490 1847.110 3291.670 ;
        RECT 1845.930 3112.090 1847.110 3113.270 ;
        RECT 1845.930 3110.490 1847.110 3111.670 ;
        RECT 1845.930 2932.090 1847.110 2933.270 ;
        RECT 1845.930 2930.490 1847.110 2931.670 ;
        RECT 1845.930 2752.090 1847.110 2753.270 ;
        RECT 1845.930 2750.490 1847.110 2751.670 ;
        RECT 1845.930 2572.090 1847.110 2573.270 ;
        RECT 1845.930 2570.490 1847.110 2571.670 ;
        RECT 1845.930 2392.090 1847.110 2393.270 ;
        RECT 1845.930 2390.490 1847.110 2391.670 ;
        RECT 1845.930 2212.090 1847.110 2213.270 ;
        RECT 1845.930 2210.490 1847.110 2211.670 ;
        RECT 1845.930 2032.090 1847.110 2033.270 ;
        RECT 1845.930 2030.490 1847.110 2031.670 ;
        RECT 1845.930 1852.090 1847.110 1853.270 ;
        RECT 1845.930 1850.490 1847.110 1851.670 ;
        RECT 1845.930 1672.090 1847.110 1673.270 ;
        RECT 1845.930 1670.490 1847.110 1671.670 ;
        RECT 1845.930 1492.090 1847.110 1493.270 ;
        RECT 1845.930 1490.490 1847.110 1491.670 ;
        RECT 1845.930 1312.090 1847.110 1313.270 ;
        RECT 1845.930 1310.490 1847.110 1311.670 ;
        RECT 1845.930 1132.090 1847.110 1133.270 ;
        RECT 1845.930 1130.490 1847.110 1131.670 ;
        RECT 1845.930 952.090 1847.110 953.270 ;
        RECT 1845.930 950.490 1847.110 951.670 ;
        RECT 1845.930 772.090 1847.110 773.270 ;
        RECT 1845.930 770.490 1847.110 771.670 ;
        RECT 1845.930 592.090 1847.110 593.270 ;
        RECT 1845.930 590.490 1847.110 591.670 ;
        RECT 1845.930 412.090 1847.110 413.270 ;
        RECT 1845.930 410.490 1847.110 411.670 ;
        RECT 1845.930 232.090 1847.110 233.270 ;
        RECT 1845.930 230.490 1847.110 231.670 ;
        RECT 1845.930 52.090 1847.110 53.270 ;
        RECT 1845.930 50.490 1847.110 51.670 ;
        RECT 1845.930 -21.710 1847.110 -20.530 ;
        RECT 1845.930 -23.310 1847.110 -22.130 ;
        RECT 2025.930 3541.810 2027.110 3542.990 ;
        RECT 2025.930 3540.210 2027.110 3541.390 ;
        RECT 2025.930 3472.090 2027.110 3473.270 ;
        RECT 2025.930 3470.490 2027.110 3471.670 ;
        RECT 2025.930 3292.090 2027.110 3293.270 ;
        RECT 2025.930 3290.490 2027.110 3291.670 ;
        RECT 2025.930 3112.090 2027.110 3113.270 ;
        RECT 2025.930 3110.490 2027.110 3111.670 ;
        RECT 2025.930 2932.090 2027.110 2933.270 ;
        RECT 2025.930 2930.490 2027.110 2931.670 ;
        RECT 2025.930 2752.090 2027.110 2753.270 ;
        RECT 2025.930 2750.490 2027.110 2751.670 ;
        RECT 2025.930 2572.090 2027.110 2573.270 ;
        RECT 2025.930 2570.490 2027.110 2571.670 ;
        RECT 2025.930 2392.090 2027.110 2393.270 ;
        RECT 2025.930 2390.490 2027.110 2391.670 ;
        RECT 2025.930 2212.090 2027.110 2213.270 ;
        RECT 2025.930 2210.490 2027.110 2211.670 ;
        RECT 2025.930 2032.090 2027.110 2033.270 ;
        RECT 2025.930 2030.490 2027.110 2031.670 ;
        RECT 2025.930 1852.090 2027.110 1853.270 ;
        RECT 2025.930 1850.490 2027.110 1851.670 ;
        RECT 2025.930 1672.090 2027.110 1673.270 ;
        RECT 2025.930 1670.490 2027.110 1671.670 ;
        RECT 2025.930 1492.090 2027.110 1493.270 ;
        RECT 2025.930 1490.490 2027.110 1491.670 ;
        RECT 2025.930 1312.090 2027.110 1313.270 ;
        RECT 2025.930 1310.490 2027.110 1311.670 ;
        RECT 2025.930 1132.090 2027.110 1133.270 ;
        RECT 2025.930 1130.490 2027.110 1131.670 ;
        RECT 2025.930 952.090 2027.110 953.270 ;
        RECT 2025.930 950.490 2027.110 951.670 ;
        RECT 2025.930 772.090 2027.110 773.270 ;
        RECT 2025.930 770.490 2027.110 771.670 ;
        RECT 2025.930 592.090 2027.110 593.270 ;
        RECT 2025.930 590.490 2027.110 591.670 ;
        RECT 2025.930 412.090 2027.110 413.270 ;
        RECT 2025.930 410.490 2027.110 411.670 ;
        RECT 2025.930 232.090 2027.110 233.270 ;
        RECT 2025.930 230.490 2027.110 231.670 ;
        RECT 2025.930 52.090 2027.110 53.270 ;
        RECT 2025.930 50.490 2027.110 51.670 ;
        RECT 2025.930 -21.710 2027.110 -20.530 ;
        RECT 2025.930 -23.310 2027.110 -22.130 ;
        RECT 2205.930 3541.810 2207.110 3542.990 ;
        RECT 2205.930 3540.210 2207.110 3541.390 ;
        RECT 2205.930 3472.090 2207.110 3473.270 ;
        RECT 2205.930 3470.490 2207.110 3471.670 ;
        RECT 2205.930 3292.090 2207.110 3293.270 ;
        RECT 2205.930 3290.490 2207.110 3291.670 ;
        RECT 2205.930 3112.090 2207.110 3113.270 ;
        RECT 2205.930 3110.490 2207.110 3111.670 ;
        RECT 2205.930 2932.090 2207.110 2933.270 ;
        RECT 2205.930 2930.490 2207.110 2931.670 ;
        RECT 2205.930 2752.090 2207.110 2753.270 ;
        RECT 2205.930 2750.490 2207.110 2751.670 ;
        RECT 2205.930 2572.090 2207.110 2573.270 ;
        RECT 2205.930 2570.490 2207.110 2571.670 ;
        RECT 2205.930 2392.090 2207.110 2393.270 ;
        RECT 2205.930 2390.490 2207.110 2391.670 ;
        RECT 2205.930 2212.090 2207.110 2213.270 ;
        RECT 2205.930 2210.490 2207.110 2211.670 ;
        RECT 2205.930 2032.090 2207.110 2033.270 ;
        RECT 2205.930 2030.490 2207.110 2031.670 ;
        RECT 2205.930 1852.090 2207.110 1853.270 ;
        RECT 2205.930 1850.490 2207.110 1851.670 ;
        RECT 2205.930 1672.090 2207.110 1673.270 ;
        RECT 2205.930 1670.490 2207.110 1671.670 ;
        RECT 2205.930 1492.090 2207.110 1493.270 ;
        RECT 2205.930 1490.490 2207.110 1491.670 ;
        RECT 2205.930 1312.090 2207.110 1313.270 ;
        RECT 2205.930 1310.490 2207.110 1311.670 ;
        RECT 2205.930 1132.090 2207.110 1133.270 ;
        RECT 2205.930 1130.490 2207.110 1131.670 ;
        RECT 2205.930 952.090 2207.110 953.270 ;
        RECT 2205.930 950.490 2207.110 951.670 ;
        RECT 2205.930 772.090 2207.110 773.270 ;
        RECT 2205.930 770.490 2207.110 771.670 ;
        RECT 2205.930 592.090 2207.110 593.270 ;
        RECT 2205.930 590.490 2207.110 591.670 ;
        RECT 2205.930 412.090 2207.110 413.270 ;
        RECT 2205.930 410.490 2207.110 411.670 ;
        RECT 2205.930 232.090 2207.110 233.270 ;
        RECT 2205.930 230.490 2207.110 231.670 ;
        RECT 2205.930 52.090 2207.110 53.270 ;
        RECT 2205.930 50.490 2207.110 51.670 ;
        RECT 2205.930 -21.710 2207.110 -20.530 ;
        RECT 2205.930 -23.310 2207.110 -22.130 ;
        RECT 2385.930 3541.810 2387.110 3542.990 ;
        RECT 2385.930 3540.210 2387.110 3541.390 ;
        RECT 2385.930 3472.090 2387.110 3473.270 ;
        RECT 2385.930 3470.490 2387.110 3471.670 ;
        RECT 2385.930 3292.090 2387.110 3293.270 ;
        RECT 2385.930 3290.490 2387.110 3291.670 ;
        RECT 2385.930 3112.090 2387.110 3113.270 ;
        RECT 2385.930 3110.490 2387.110 3111.670 ;
        RECT 2385.930 2932.090 2387.110 2933.270 ;
        RECT 2385.930 2930.490 2387.110 2931.670 ;
        RECT 2385.930 2752.090 2387.110 2753.270 ;
        RECT 2385.930 2750.490 2387.110 2751.670 ;
        RECT 2385.930 2572.090 2387.110 2573.270 ;
        RECT 2385.930 2570.490 2387.110 2571.670 ;
        RECT 2385.930 2392.090 2387.110 2393.270 ;
        RECT 2385.930 2390.490 2387.110 2391.670 ;
        RECT 2385.930 2212.090 2387.110 2213.270 ;
        RECT 2385.930 2210.490 2387.110 2211.670 ;
        RECT 2385.930 2032.090 2387.110 2033.270 ;
        RECT 2385.930 2030.490 2387.110 2031.670 ;
        RECT 2385.930 1852.090 2387.110 1853.270 ;
        RECT 2385.930 1850.490 2387.110 1851.670 ;
        RECT 2385.930 1672.090 2387.110 1673.270 ;
        RECT 2385.930 1670.490 2387.110 1671.670 ;
        RECT 2385.930 1492.090 2387.110 1493.270 ;
        RECT 2385.930 1490.490 2387.110 1491.670 ;
        RECT 2385.930 1312.090 2387.110 1313.270 ;
        RECT 2385.930 1310.490 2387.110 1311.670 ;
        RECT 2385.930 1132.090 2387.110 1133.270 ;
        RECT 2385.930 1130.490 2387.110 1131.670 ;
        RECT 2385.930 952.090 2387.110 953.270 ;
        RECT 2385.930 950.490 2387.110 951.670 ;
        RECT 2385.930 772.090 2387.110 773.270 ;
        RECT 2385.930 770.490 2387.110 771.670 ;
        RECT 2385.930 592.090 2387.110 593.270 ;
        RECT 2385.930 590.490 2387.110 591.670 ;
        RECT 2385.930 412.090 2387.110 413.270 ;
        RECT 2385.930 410.490 2387.110 411.670 ;
        RECT 2385.930 232.090 2387.110 233.270 ;
        RECT 2385.930 230.490 2387.110 231.670 ;
        RECT 2385.930 52.090 2387.110 53.270 ;
        RECT 2385.930 50.490 2387.110 51.670 ;
        RECT 2385.930 -21.710 2387.110 -20.530 ;
        RECT 2385.930 -23.310 2387.110 -22.130 ;
        RECT 2565.930 3541.810 2567.110 3542.990 ;
        RECT 2565.930 3540.210 2567.110 3541.390 ;
        RECT 2565.930 3472.090 2567.110 3473.270 ;
        RECT 2565.930 3470.490 2567.110 3471.670 ;
        RECT 2565.930 3292.090 2567.110 3293.270 ;
        RECT 2565.930 3290.490 2567.110 3291.670 ;
        RECT 2565.930 3112.090 2567.110 3113.270 ;
        RECT 2565.930 3110.490 2567.110 3111.670 ;
        RECT 2565.930 2932.090 2567.110 2933.270 ;
        RECT 2565.930 2930.490 2567.110 2931.670 ;
        RECT 2565.930 2752.090 2567.110 2753.270 ;
        RECT 2565.930 2750.490 2567.110 2751.670 ;
        RECT 2565.930 2572.090 2567.110 2573.270 ;
        RECT 2565.930 2570.490 2567.110 2571.670 ;
        RECT 2565.930 2392.090 2567.110 2393.270 ;
        RECT 2565.930 2390.490 2567.110 2391.670 ;
        RECT 2565.930 2212.090 2567.110 2213.270 ;
        RECT 2565.930 2210.490 2567.110 2211.670 ;
        RECT 2565.930 2032.090 2567.110 2033.270 ;
        RECT 2565.930 2030.490 2567.110 2031.670 ;
        RECT 2565.930 1852.090 2567.110 1853.270 ;
        RECT 2565.930 1850.490 2567.110 1851.670 ;
        RECT 2565.930 1672.090 2567.110 1673.270 ;
        RECT 2565.930 1670.490 2567.110 1671.670 ;
        RECT 2565.930 1492.090 2567.110 1493.270 ;
        RECT 2565.930 1490.490 2567.110 1491.670 ;
        RECT 2565.930 1312.090 2567.110 1313.270 ;
        RECT 2565.930 1310.490 2567.110 1311.670 ;
        RECT 2565.930 1132.090 2567.110 1133.270 ;
        RECT 2565.930 1130.490 2567.110 1131.670 ;
        RECT 2565.930 952.090 2567.110 953.270 ;
        RECT 2565.930 950.490 2567.110 951.670 ;
        RECT 2565.930 772.090 2567.110 773.270 ;
        RECT 2565.930 770.490 2567.110 771.670 ;
        RECT 2565.930 592.090 2567.110 593.270 ;
        RECT 2565.930 590.490 2567.110 591.670 ;
        RECT 2565.930 412.090 2567.110 413.270 ;
        RECT 2565.930 410.490 2567.110 411.670 ;
        RECT 2565.930 232.090 2567.110 233.270 ;
        RECT 2565.930 230.490 2567.110 231.670 ;
        RECT 2565.930 52.090 2567.110 53.270 ;
        RECT 2565.930 50.490 2567.110 51.670 ;
        RECT 2565.930 -21.710 2567.110 -20.530 ;
        RECT 2565.930 -23.310 2567.110 -22.130 ;
        RECT 2745.930 3541.810 2747.110 3542.990 ;
        RECT 2745.930 3540.210 2747.110 3541.390 ;
        RECT 2745.930 3472.090 2747.110 3473.270 ;
        RECT 2745.930 3470.490 2747.110 3471.670 ;
        RECT 2745.930 3292.090 2747.110 3293.270 ;
        RECT 2745.930 3290.490 2747.110 3291.670 ;
        RECT 2745.930 3112.090 2747.110 3113.270 ;
        RECT 2745.930 3110.490 2747.110 3111.670 ;
        RECT 2745.930 2932.090 2747.110 2933.270 ;
        RECT 2745.930 2930.490 2747.110 2931.670 ;
        RECT 2745.930 2752.090 2747.110 2753.270 ;
        RECT 2745.930 2750.490 2747.110 2751.670 ;
        RECT 2745.930 2572.090 2747.110 2573.270 ;
        RECT 2745.930 2570.490 2747.110 2571.670 ;
        RECT 2745.930 2392.090 2747.110 2393.270 ;
        RECT 2745.930 2390.490 2747.110 2391.670 ;
        RECT 2745.930 2212.090 2747.110 2213.270 ;
        RECT 2745.930 2210.490 2747.110 2211.670 ;
        RECT 2745.930 2032.090 2747.110 2033.270 ;
        RECT 2745.930 2030.490 2747.110 2031.670 ;
        RECT 2745.930 1852.090 2747.110 1853.270 ;
        RECT 2745.930 1850.490 2747.110 1851.670 ;
        RECT 2745.930 1672.090 2747.110 1673.270 ;
        RECT 2745.930 1670.490 2747.110 1671.670 ;
        RECT 2745.930 1492.090 2747.110 1493.270 ;
        RECT 2745.930 1490.490 2747.110 1491.670 ;
        RECT 2745.930 1312.090 2747.110 1313.270 ;
        RECT 2745.930 1310.490 2747.110 1311.670 ;
        RECT 2745.930 1132.090 2747.110 1133.270 ;
        RECT 2745.930 1130.490 2747.110 1131.670 ;
        RECT 2745.930 952.090 2747.110 953.270 ;
        RECT 2745.930 950.490 2747.110 951.670 ;
        RECT 2745.930 772.090 2747.110 773.270 ;
        RECT 2745.930 770.490 2747.110 771.670 ;
        RECT 2745.930 592.090 2747.110 593.270 ;
        RECT 2745.930 590.490 2747.110 591.670 ;
        RECT 2745.930 412.090 2747.110 413.270 ;
        RECT 2745.930 410.490 2747.110 411.670 ;
        RECT 2745.930 232.090 2747.110 233.270 ;
        RECT 2745.930 230.490 2747.110 231.670 ;
        RECT 2745.930 52.090 2747.110 53.270 ;
        RECT 2745.930 50.490 2747.110 51.670 ;
        RECT 2745.930 -21.710 2747.110 -20.530 ;
        RECT 2745.930 -23.310 2747.110 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 3472.090 2947.490 3473.270 ;
        RECT 2946.310 3470.490 2947.490 3471.670 ;
        RECT 2946.310 3292.090 2947.490 3293.270 ;
        RECT 2946.310 3290.490 2947.490 3291.670 ;
        RECT 2946.310 3112.090 2947.490 3113.270 ;
        RECT 2946.310 3110.490 2947.490 3111.670 ;
        RECT 2946.310 2932.090 2947.490 2933.270 ;
        RECT 2946.310 2930.490 2947.490 2931.670 ;
        RECT 2946.310 2752.090 2947.490 2753.270 ;
        RECT 2946.310 2750.490 2947.490 2751.670 ;
        RECT 2946.310 2572.090 2947.490 2573.270 ;
        RECT 2946.310 2570.490 2947.490 2571.670 ;
        RECT 2946.310 2392.090 2947.490 2393.270 ;
        RECT 2946.310 2390.490 2947.490 2391.670 ;
        RECT 2946.310 2212.090 2947.490 2213.270 ;
        RECT 2946.310 2210.490 2947.490 2211.670 ;
        RECT 2946.310 2032.090 2947.490 2033.270 ;
        RECT 2946.310 2030.490 2947.490 2031.670 ;
        RECT 2946.310 1852.090 2947.490 1853.270 ;
        RECT 2946.310 1850.490 2947.490 1851.670 ;
        RECT 2946.310 1672.090 2947.490 1673.270 ;
        RECT 2946.310 1670.490 2947.490 1671.670 ;
        RECT 2946.310 1492.090 2947.490 1493.270 ;
        RECT 2946.310 1490.490 2947.490 1491.670 ;
        RECT 2946.310 1312.090 2947.490 1313.270 ;
        RECT 2946.310 1310.490 2947.490 1311.670 ;
        RECT 2946.310 1132.090 2947.490 1133.270 ;
        RECT 2946.310 1130.490 2947.490 1131.670 ;
        RECT 2946.310 952.090 2947.490 953.270 ;
        RECT 2946.310 950.490 2947.490 951.670 ;
        RECT 2946.310 772.090 2947.490 773.270 ;
        RECT 2946.310 770.490 2947.490 771.670 ;
        RECT 2946.310 592.090 2947.490 593.270 ;
        RECT 2946.310 590.490 2947.490 591.670 ;
        RECT 2946.310 412.090 2947.490 413.270 ;
        RECT 2946.310 410.490 2947.490 411.670 ;
        RECT 2946.310 232.090 2947.490 233.270 ;
        RECT 2946.310 230.490 2947.490 231.670 ;
        RECT 2946.310 52.090 2947.490 53.270 ;
        RECT 2946.310 50.490 2947.490 51.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 45.020 3543.100 48.020 3543.110 ;
        RECT 225.020 3543.100 228.020 3543.110 ;
        RECT 405.020 3543.100 408.020 3543.110 ;
        RECT 585.020 3543.100 588.020 3543.110 ;
        RECT 765.020 3543.100 768.020 3543.110 ;
        RECT 945.020 3543.100 948.020 3543.110 ;
        RECT 1125.020 3543.100 1128.020 3543.110 ;
        RECT 1305.020 3543.100 1308.020 3543.110 ;
        RECT 1485.020 3543.100 1488.020 3543.110 ;
        RECT 1665.020 3543.100 1668.020 3543.110 ;
        RECT 1845.020 3543.100 1848.020 3543.110 ;
        RECT 2025.020 3543.100 2028.020 3543.110 ;
        RECT 2205.020 3543.100 2208.020 3543.110 ;
        RECT 2385.020 3543.100 2388.020 3543.110 ;
        RECT 2565.020 3543.100 2568.020 3543.110 ;
        RECT 2745.020 3543.100 2748.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 45.020 3540.090 48.020 3540.100 ;
        RECT 225.020 3540.090 228.020 3540.100 ;
        RECT 405.020 3540.090 408.020 3540.100 ;
        RECT 585.020 3540.090 588.020 3540.100 ;
        RECT 765.020 3540.090 768.020 3540.100 ;
        RECT 945.020 3540.090 948.020 3540.100 ;
        RECT 1125.020 3540.090 1128.020 3540.100 ;
        RECT 1305.020 3540.090 1308.020 3540.100 ;
        RECT 1485.020 3540.090 1488.020 3540.100 ;
        RECT 1665.020 3540.090 1668.020 3540.100 ;
        RECT 1845.020 3540.090 1848.020 3540.100 ;
        RECT 2025.020 3540.090 2028.020 3540.100 ;
        RECT 2205.020 3540.090 2208.020 3540.100 ;
        RECT 2385.020 3540.090 2388.020 3540.100 ;
        RECT 2565.020 3540.090 2568.020 3540.100 ;
        RECT 2745.020 3540.090 2748.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3473.380 -25.780 3473.390 ;
        RECT 45.020 3473.380 48.020 3473.390 ;
        RECT 225.020 3473.380 228.020 3473.390 ;
        RECT 405.020 3473.380 408.020 3473.390 ;
        RECT 585.020 3473.380 588.020 3473.390 ;
        RECT 765.020 3473.380 768.020 3473.390 ;
        RECT 945.020 3473.380 948.020 3473.390 ;
        RECT 1125.020 3473.380 1128.020 3473.390 ;
        RECT 1305.020 3473.380 1308.020 3473.390 ;
        RECT 1485.020 3473.380 1488.020 3473.390 ;
        RECT 1665.020 3473.380 1668.020 3473.390 ;
        RECT 1845.020 3473.380 1848.020 3473.390 ;
        RECT 2025.020 3473.380 2028.020 3473.390 ;
        RECT 2205.020 3473.380 2208.020 3473.390 ;
        RECT 2385.020 3473.380 2388.020 3473.390 ;
        RECT 2565.020 3473.380 2568.020 3473.390 ;
        RECT 2745.020 3473.380 2748.020 3473.390 ;
        RECT 2945.400 3473.380 2948.400 3473.390 ;
        RECT -33.480 3470.380 2953.100 3473.380 ;
        RECT -28.780 3470.370 -25.780 3470.380 ;
        RECT 45.020 3470.370 48.020 3470.380 ;
        RECT 225.020 3470.370 228.020 3470.380 ;
        RECT 405.020 3470.370 408.020 3470.380 ;
        RECT 585.020 3470.370 588.020 3470.380 ;
        RECT 765.020 3470.370 768.020 3470.380 ;
        RECT 945.020 3470.370 948.020 3470.380 ;
        RECT 1125.020 3470.370 1128.020 3470.380 ;
        RECT 1305.020 3470.370 1308.020 3470.380 ;
        RECT 1485.020 3470.370 1488.020 3470.380 ;
        RECT 1665.020 3470.370 1668.020 3470.380 ;
        RECT 1845.020 3470.370 1848.020 3470.380 ;
        RECT 2025.020 3470.370 2028.020 3470.380 ;
        RECT 2205.020 3470.370 2208.020 3470.380 ;
        RECT 2385.020 3470.370 2388.020 3470.380 ;
        RECT 2565.020 3470.370 2568.020 3470.380 ;
        RECT 2745.020 3470.370 2748.020 3470.380 ;
        RECT 2945.400 3470.370 2948.400 3470.380 ;
        RECT -28.780 3293.380 -25.780 3293.390 ;
        RECT 45.020 3293.380 48.020 3293.390 ;
        RECT 225.020 3293.380 228.020 3293.390 ;
        RECT 405.020 3293.380 408.020 3293.390 ;
        RECT 585.020 3293.380 588.020 3293.390 ;
        RECT 765.020 3293.380 768.020 3293.390 ;
        RECT 945.020 3293.380 948.020 3293.390 ;
        RECT 1125.020 3293.380 1128.020 3293.390 ;
        RECT 1305.020 3293.380 1308.020 3293.390 ;
        RECT 1485.020 3293.380 1488.020 3293.390 ;
        RECT 1665.020 3293.380 1668.020 3293.390 ;
        RECT 1845.020 3293.380 1848.020 3293.390 ;
        RECT 2025.020 3293.380 2028.020 3293.390 ;
        RECT 2205.020 3293.380 2208.020 3293.390 ;
        RECT 2385.020 3293.380 2388.020 3293.390 ;
        RECT 2565.020 3293.380 2568.020 3293.390 ;
        RECT 2745.020 3293.380 2748.020 3293.390 ;
        RECT 2945.400 3293.380 2948.400 3293.390 ;
        RECT -33.480 3290.380 2953.100 3293.380 ;
        RECT -28.780 3290.370 -25.780 3290.380 ;
        RECT 45.020 3290.370 48.020 3290.380 ;
        RECT 225.020 3290.370 228.020 3290.380 ;
        RECT 405.020 3290.370 408.020 3290.380 ;
        RECT 585.020 3290.370 588.020 3290.380 ;
        RECT 765.020 3290.370 768.020 3290.380 ;
        RECT 945.020 3290.370 948.020 3290.380 ;
        RECT 1125.020 3290.370 1128.020 3290.380 ;
        RECT 1305.020 3290.370 1308.020 3290.380 ;
        RECT 1485.020 3290.370 1488.020 3290.380 ;
        RECT 1665.020 3290.370 1668.020 3290.380 ;
        RECT 1845.020 3290.370 1848.020 3290.380 ;
        RECT 2025.020 3290.370 2028.020 3290.380 ;
        RECT 2205.020 3290.370 2208.020 3290.380 ;
        RECT 2385.020 3290.370 2388.020 3290.380 ;
        RECT 2565.020 3290.370 2568.020 3290.380 ;
        RECT 2745.020 3290.370 2748.020 3290.380 ;
        RECT 2945.400 3290.370 2948.400 3290.380 ;
        RECT -28.780 3113.380 -25.780 3113.390 ;
        RECT 45.020 3113.380 48.020 3113.390 ;
        RECT 225.020 3113.380 228.020 3113.390 ;
        RECT 405.020 3113.380 408.020 3113.390 ;
        RECT 585.020 3113.380 588.020 3113.390 ;
        RECT 765.020 3113.380 768.020 3113.390 ;
        RECT 945.020 3113.380 948.020 3113.390 ;
        RECT 1125.020 3113.380 1128.020 3113.390 ;
        RECT 1305.020 3113.380 1308.020 3113.390 ;
        RECT 1485.020 3113.380 1488.020 3113.390 ;
        RECT 1665.020 3113.380 1668.020 3113.390 ;
        RECT 1845.020 3113.380 1848.020 3113.390 ;
        RECT 2025.020 3113.380 2028.020 3113.390 ;
        RECT 2205.020 3113.380 2208.020 3113.390 ;
        RECT 2385.020 3113.380 2388.020 3113.390 ;
        RECT 2565.020 3113.380 2568.020 3113.390 ;
        RECT 2745.020 3113.380 2748.020 3113.390 ;
        RECT 2945.400 3113.380 2948.400 3113.390 ;
        RECT -33.480 3110.380 2953.100 3113.380 ;
        RECT -28.780 3110.370 -25.780 3110.380 ;
        RECT 45.020 3110.370 48.020 3110.380 ;
        RECT 225.020 3110.370 228.020 3110.380 ;
        RECT 405.020 3110.370 408.020 3110.380 ;
        RECT 585.020 3110.370 588.020 3110.380 ;
        RECT 765.020 3110.370 768.020 3110.380 ;
        RECT 945.020 3110.370 948.020 3110.380 ;
        RECT 1125.020 3110.370 1128.020 3110.380 ;
        RECT 1305.020 3110.370 1308.020 3110.380 ;
        RECT 1485.020 3110.370 1488.020 3110.380 ;
        RECT 1665.020 3110.370 1668.020 3110.380 ;
        RECT 1845.020 3110.370 1848.020 3110.380 ;
        RECT 2025.020 3110.370 2028.020 3110.380 ;
        RECT 2205.020 3110.370 2208.020 3110.380 ;
        RECT 2385.020 3110.370 2388.020 3110.380 ;
        RECT 2565.020 3110.370 2568.020 3110.380 ;
        RECT 2745.020 3110.370 2748.020 3110.380 ;
        RECT 2945.400 3110.370 2948.400 3110.380 ;
        RECT -28.780 2933.380 -25.780 2933.390 ;
        RECT 45.020 2933.380 48.020 2933.390 ;
        RECT 225.020 2933.380 228.020 2933.390 ;
        RECT 405.020 2933.380 408.020 2933.390 ;
        RECT 585.020 2933.380 588.020 2933.390 ;
        RECT 765.020 2933.380 768.020 2933.390 ;
        RECT 945.020 2933.380 948.020 2933.390 ;
        RECT 1125.020 2933.380 1128.020 2933.390 ;
        RECT 1305.020 2933.380 1308.020 2933.390 ;
        RECT 1485.020 2933.380 1488.020 2933.390 ;
        RECT 1665.020 2933.380 1668.020 2933.390 ;
        RECT 1845.020 2933.380 1848.020 2933.390 ;
        RECT 2025.020 2933.380 2028.020 2933.390 ;
        RECT 2205.020 2933.380 2208.020 2933.390 ;
        RECT 2385.020 2933.380 2388.020 2933.390 ;
        RECT 2565.020 2933.380 2568.020 2933.390 ;
        RECT 2745.020 2933.380 2748.020 2933.390 ;
        RECT 2945.400 2933.380 2948.400 2933.390 ;
        RECT -33.480 2930.380 2953.100 2933.380 ;
        RECT -28.780 2930.370 -25.780 2930.380 ;
        RECT 45.020 2930.370 48.020 2930.380 ;
        RECT 225.020 2930.370 228.020 2930.380 ;
        RECT 405.020 2930.370 408.020 2930.380 ;
        RECT 585.020 2930.370 588.020 2930.380 ;
        RECT 765.020 2930.370 768.020 2930.380 ;
        RECT 945.020 2930.370 948.020 2930.380 ;
        RECT 1125.020 2930.370 1128.020 2930.380 ;
        RECT 1305.020 2930.370 1308.020 2930.380 ;
        RECT 1485.020 2930.370 1488.020 2930.380 ;
        RECT 1665.020 2930.370 1668.020 2930.380 ;
        RECT 1845.020 2930.370 1848.020 2930.380 ;
        RECT 2025.020 2930.370 2028.020 2930.380 ;
        RECT 2205.020 2930.370 2208.020 2930.380 ;
        RECT 2385.020 2930.370 2388.020 2930.380 ;
        RECT 2565.020 2930.370 2568.020 2930.380 ;
        RECT 2745.020 2930.370 2748.020 2930.380 ;
        RECT 2945.400 2930.370 2948.400 2930.380 ;
        RECT -28.780 2753.380 -25.780 2753.390 ;
        RECT 45.020 2753.380 48.020 2753.390 ;
        RECT 225.020 2753.380 228.020 2753.390 ;
        RECT 405.020 2753.380 408.020 2753.390 ;
        RECT 585.020 2753.380 588.020 2753.390 ;
        RECT 765.020 2753.380 768.020 2753.390 ;
        RECT 945.020 2753.380 948.020 2753.390 ;
        RECT 1125.020 2753.380 1128.020 2753.390 ;
        RECT 1305.020 2753.380 1308.020 2753.390 ;
        RECT 1485.020 2753.380 1488.020 2753.390 ;
        RECT 1665.020 2753.380 1668.020 2753.390 ;
        RECT 1845.020 2753.380 1848.020 2753.390 ;
        RECT 2025.020 2753.380 2028.020 2753.390 ;
        RECT 2205.020 2753.380 2208.020 2753.390 ;
        RECT 2385.020 2753.380 2388.020 2753.390 ;
        RECT 2565.020 2753.380 2568.020 2753.390 ;
        RECT 2745.020 2753.380 2748.020 2753.390 ;
        RECT 2945.400 2753.380 2948.400 2753.390 ;
        RECT -33.480 2750.380 2953.100 2753.380 ;
        RECT -28.780 2750.370 -25.780 2750.380 ;
        RECT 45.020 2750.370 48.020 2750.380 ;
        RECT 225.020 2750.370 228.020 2750.380 ;
        RECT 405.020 2750.370 408.020 2750.380 ;
        RECT 585.020 2750.370 588.020 2750.380 ;
        RECT 765.020 2750.370 768.020 2750.380 ;
        RECT 945.020 2750.370 948.020 2750.380 ;
        RECT 1125.020 2750.370 1128.020 2750.380 ;
        RECT 1305.020 2750.370 1308.020 2750.380 ;
        RECT 1485.020 2750.370 1488.020 2750.380 ;
        RECT 1665.020 2750.370 1668.020 2750.380 ;
        RECT 1845.020 2750.370 1848.020 2750.380 ;
        RECT 2025.020 2750.370 2028.020 2750.380 ;
        RECT 2205.020 2750.370 2208.020 2750.380 ;
        RECT 2385.020 2750.370 2388.020 2750.380 ;
        RECT 2565.020 2750.370 2568.020 2750.380 ;
        RECT 2745.020 2750.370 2748.020 2750.380 ;
        RECT 2945.400 2750.370 2948.400 2750.380 ;
        RECT -28.780 2573.380 -25.780 2573.390 ;
        RECT 45.020 2573.380 48.020 2573.390 ;
        RECT 225.020 2573.380 228.020 2573.390 ;
        RECT 405.020 2573.380 408.020 2573.390 ;
        RECT 585.020 2573.380 588.020 2573.390 ;
        RECT 765.020 2573.380 768.020 2573.390 ;
        RECT 945.020 2573.380 948.020 2573.390 ;
        RECT 1125.020 2573.380 1128.020 2573.390 ;
        RECT 1305.020 2573.380 1308.020 2573.390 ;
        RECT 1485.020 2573.380 1488.020 2573.390 ;
        RECT 1665.020 2573.380 1668.020 2573.390 ;
        RECT 1845.020 2573.380 1848.020 2573.390 ;
        RECT 2025.020 2573.380 2028.020 2573.390 ;
        RECT 2205.020 2573.380 2208.020 2573.390 ;
        RECT 2385.020 2573.380 2388.020 2573.390 ;
        RECT 2565.020 2573.380 2568.020 2573.390 ;
        RECT 2745.020 2573.380 2748.020 2573.390 ;
        RECT 2945.400 2573.380 2948.400 2573.390 ;
        RECT -33.480 2570.380 2953.100 2573.380 ;
        RECT -28.780 2570.370 -25.780 2570.380 ;
        RECT 45.020 2570.370 48.020 2570.380 ;
        RECT 225.020 2570.370 228.020 2570.380 ;
        RECT 405.020 2570.370 408.020 2570.380 ;
        RECT 585.020 2570.370 588.020 2570.380 ;
        RECT 765.020 2570.370 768.020 2570.380 ;
        RECT 945.020 2570.370 948.020 2570.380 ;
        RECT 1125.020 2570.370 1128.020 2570.380 ;
        RECT 1305.020 2570.370 1308.020 2570.380 ;
        RECT 1485.020 2570.370 1488.020 2570.380 ;
        RECT 1665.020 2570.370 1668.020 2570.380 ;
        RECT 1845.020 2570.370 1848.020 2570.380 ;
        RECT 2025.020 2570.370 2028.020 2570.380 ;
        RECT 2205.020 2570.370 2208.020 2570.380 ;
        RECT 2385.020 2570.370 2388.020 2570.380 ;
        RECT 2565.020 2570.370 2568.020 2570.380 ;
        RECT 2745.020 2570.370 2748.020 2570.380 ;
        RECT 2945.400 2570.370 2948.400 2570.380 ;
        RECT -28.780 2393.380 -25.780 2393.390 ;
        RECT 45.020 2393.380 48.020 2393.390 ;
        RECT 225.020 2393.380 228.020 2393.390 ;
        RECT 405.020 2393.380 408.020 2393.390 ;
        RECT 585.020 2393.380 588.020 2393.390 ;
        RECT 765.020 2393.380 768.020 2393.390 ;
        RECT 945.020 2393.380 948.020 2393.390 ;
        RECT 1125.020 2393.380 1128.020 2393.390 ;
        RECT 1305.020 2393.380 1308.020 2393.390 ;
        RECT 1485.020 2393.380 1488.020 2393.390 ;
        RECT 1665.020 2393.380 1668.020 2393.390 ;
        RECT 1845.020 2393.380 1848.020 2393.390 ;
        RECT 2025.020 2393.380 2028.020 2393.390 ;
        RECT 2205.020 2393.380 2208.020 2393.390 ;
        RECT 2385.020 2393.380 2388.020 2393.390 ;
        RECT 2565.020 2393.380 2568.020 2393.390 ;
        RECT 2745.020 2393.380 2748.020 2393.390 ;
        RECT 2945.400 2393.380 2948.400 2393.390 ;
        RECT -33.480 2390.380 2953.100 2393.380 ;
        RECT -28.780 2390.370 -25.780 2390.380 ;
        RECT 45.020 2390.370 48.020 2390.380 ;
        RECT 225.020 2390.370 228.020 2390.380 ;
        RECT 405.020 2390.370 408.020 2390.380 ;
        RECT 585.020 2390.370 588.020 2390.380 ;
        RECT 765.020 2390.370 768.020 2390.380 ;
        RECT 945.020 2390.370 948.020 2390.380 ;
        RECT 1125.020 2390.370 1128.020 2390.380 ;
        RECT 1305.020 2390.370 1308.020 2390.380 ;
        RECT 1485.020 2390.370 1488.020 2390.380 ;
        RECT 1665.020 2390.370 1668.020 2390.380 ;
        RECT 1845.020 2390.370 1848.020 2390.380 ;
        RECT 2025.020 2390.370 2028.020 2390.380 ;
        RECT 2205.020 2390.370 2208.020 2390.380 ;
        RECT 2385.020 2390.370 2388.020 2390.380 ;
        RECT 2565.020 2390.370 2568.020 2390.380 ;
        RECT 2745.020 2390.370 2748.020 2390.380 ;
        RECT 2945.400 2390.370 2948.400 2390.380 ;
        RECT -28.780 2213.380 -25.780 2213.390 ;
        RECT 45.020 2213.380 48.020 2213.390 ;
        RECT 225.020 2213.380 228.020 2213.390 ;
        RECT 405.020 2213.380 408.020 2213.390 ;
        RECT 585.020 2213.380 588.020 2213.390 ;
        RECT 765.020 2213.380 768.020 2213.390 ;
        RECT 945.020 2213.380 948.020 2213.390 ;
        RECT 1125.020 2213.380 1128.020 2213.390 ;
        RECT 1305.020 2213.380 1308.020 2213.390 ;
        RECT 1485.020 2213.380 1488.020 2213.390 ;
        RECT 1665.020 2213.380 1668.020 2213.390 ;
        RECT 1845.020 2213.380 1848.020 2213.390 ;
        RECT 2025.020 2213.380 2028.020 2213.390 ;
        RECT 2205.020 2213.380 2208.020 2213.390 ;
        RECT 2385.020 2213.380 2388.020 2213.390 ;
        RECT 2565.020 2213.380 2568.020 2213.390 ;
        RECT 2745.020 2213.380 2748.020 2213.390 ;
        RECT 2945.400 2213.380 2948.400 2213.390 ;
        RECT -33.480 2210.380 2953.100 2213.380 ;
        RECT -28.780 2210.370 -25.780 2210.380 ;
        RECT 45.020 2210.370 48.020 2210.380 ;
        RECT 225.020 2210.370 228.020 2210.380 ;
        RECT 405.020 2210.370 408.020 2210.380 ;
        RECT 585.020 2210.370 588.020 2210.380 ;
        RECT 765.020 2210.370 768.020 2210.380 ;
        RECT 945.020 2210.370 948.020 2210.380 ;
        RECT 1125.020 2210.370 1128.020 2210.380 ;
        RECT 1305.020 2210.370 1308.020 2210.380 ;
        RECT 1485.020 2210.370 1488.020 2210.380 ;
        RECT 1665.020 2210.370 1668.020 2210.380 ;
        RECT 1845.020 2210.370 1848.020 2210.380 ;
        RECT 2025.020 2210.370 2028.020 2210.380 ;
        RECT 2205.020 2210.370 2208.020 2210.380 ;
        RECT 2385.020 2210.370 2388.020 2210.380 ;
        RECT 2565.020 2210.370 2568.020 2210.380 ;
        RECT 2745.020 2210.370 2748.020 2210.380 ;
        RECT 2945.400 2210.370 2948.400 2210.380 ;
        RECT -28.780 2033.380 -25.780 2033.390 ;
        RECT 45.020 2033.380 48.020 2033.390 ;
        RECT 225.020 2033.380 228.020 2033.390 ;
        RECT 405.020 2033.380 408.020 2033.390 ;
        RECT 585.020 2033.380 588.020 2033.390 ;
        RECT 765.020 2033.380 768.020 2033.390 ;
        RECT 945.020 2033.380 948.020 2033.390 ;
        RECT 1125.020 2033.380 1128.020 2033.390 ;
        RECT 1305.020 2033.380 1308.020 2033.390 ;
        RECT 1485.020 2033.380 1488.020 2033.390 ;
        RECT 1665.020 2033.380 1668.020 2033.390 ;
        RECT 1845.020 2033.380 1848.020 2033.390 ;
        RECT 2025.020 2033.380 2028.020 2033.390 ;
        RECT 2205.020 2033.380 2208.020 2033.390 ;
        RECT 2385.020 2033.380 2388.020 2033.390 ;
        RECT 2565.020 2033.380 2568.020 2033.390 ;
        RECT 2745.020 2033.380 2748.020 2033.390 ;
        RECT 2945.400 2033.380 2948.400 2033.390 ;
        RECT -33.480 2030.380 2953.100 2033.380 ;
        RECT -28.780 2030.370 -25.780 2030.380 ;
        RECT 45.020 2030.370 48.020 2030.380 ;
        RECT 225.020 2030.370 228.020 2030.380 ;
        RECT 405.020 2030.370 408.020 2030.380 ;
        RECT 585.020 2030.370 588.020 2030.380 ;
        RECT 765.020 2030.370 768.020 2030.380 ;
        RECT 945.020 2030.370 948.020 2030.380 ;
        RECT 1125.020 2030.370 1128.020 2030.380 ;
        RECT 1305.020 2030.370 1308.020 2030.380 ;
        RECT 1485.020 2030.370 1488.020 2030.380 ;
        RECT 1665.020 2030.370 1668.020 2030.380 ;
        RECT 1845.020 2030.370 1848.020 2030.380 ;
        RECT 2025.020 2030.370 2028.020 2030.380 ;
        RECT 2205.020 2030.370 2208.020 2030.380 ;
        RECT 2385.020 2030.370 2388.020 2030.380 ;
        RECT 2565.020 2030.370 2568.020 2030.380 ;
        RECT 2745.020 2030.370 2748.020 2030.380 ;
        RECT 2945.400 2030.370 2948.400 2030.380 ;
        RECT -28.780 1853.380 -25.780 1853.390 ;
        RECT 45.020 1853.380 48.020 1853.390 ;
        RECT 225.020 1853.380 228.020 1853.390 ;
        RECT 405.020 1853.380 408.020 1853.390 ;
        RECT 585.020 1853.380 588.020 1853.390 ;
        RECT 765.020 1853.380 768.020 1853.390 ;
        RECT 945.020 1853.380 948.020 1853.390 ;
        RECT 1125.020 1853.380 1128.020 1853.390 ;
        RECT 1305.020 1853.380 1308.020 1853.390 ;
        RECT 1485.020 1853.380 1488.020 1853.390 ;
        RECT 1665.020 1853.380 1668.020 1853.390 ;
        RECT 1845.020 1853.380 1848.020 1853.390 ;
        RECT 2025.020 1853.380 2028.020 1853.390 ;
        RECT 2205.020 1853.380 2208.020 1853.390 ;
        RECT 2385.020 1853.380 2388.020 1853.390 ;
        RECT 2565.020 1853.380 2568.020 1853.390 ;
        RECT 2745.020 1853.380 2748.020 1853.390 ;
        RECT 2945.400 1853.380 2948.400 1853.390 ;
        RECT -33.480 1850.380 2953.100 1853.380 ;
        RECT -28.780 1850.370 -25.780 1850.380 ;
        RECT 45.020 1850.370 48.020 1850.380 ;
        RECT 225.020 1850.370 228.020 1850.380 ;
        RECT 405.020 1850.370 408.020 1850.380 ;
        RECT 585.020 1850.370 588.020 1850.380 ;
        RECT 765.020 1850.370 768.020 1850.380 ;
        RECT 945.020 1850.370 948.020 1850.380 ;
        RECT 1125.020 1850.370 1128.020 1850.380 ;
        RECT 1305.020 1850.370 1308.020 1850.380 ;
        RECT 1485.020 1850.370 1488.020 1850.380 ;
        RECT 1665.020 1850.370 1668.020 1850.380 ;
        RECT 1845.020 1850.370 1848.020 1850.380 ;
        RECT 2025.020 1850.370 2028.020 1850.380 ;
        RECT 2205.020 1850.370 2208.020 1850.380 ;
        RECT 2385.020 1850.370 2388.020 1850.380 ;
        RECT 2565.020 1850.370 2568.020 1850.380 ;
        RECT 2745.020 1850.370 2748.020 1850.380 ;
        RECT 2945.400 1850.370 2948.400 1850.380 ;
        RECT -28.780 1673.380 -25.780 1673.390 ;
        RECT 45.020 1673.380 48.020 1673.390 ;
        RECT 225.020 1673.380 228.020 1673.390 ;
        RECT 405.020 1673.380 408.020 1673.390 ;
        RECT 585.020 1673.380 588.020 1673.390 ;
        RECT 765.020 1673.380 768.020 1673.390 ;
        RECT 945.020 1673.380 948.020 1673.390 ;
        RECT 1125.020 1673.380 1128.020 1673.390 ;
        RECT 1305.020 1673.380 1308.020 1673.390 ;
        RECT 1485.020 1673.380 1488.020 1673.390 ;
        RECT 1665.020 1673.380 1668.020 1673.390 ;
        RECT 1845.020 1673.380 1848.020 1673.390 ;
        RECT 2025.020 1673.380 2028.020 1673.390 ;
        RECT 2205.020 1673.380 2208.020 1673.390 ;
        RECT 2385.020 1673.380 2388.020 1673.390 ;
        RECT 2565.020 1673.380 2568.020 1673.390 ;
        RECT 2745.020 1673.380 2748.020 1673.390 ;
        RECT 2945.400 1673.380 2948.400 1673.390 ;
        RECT -33.480 1670.380 2953.100 1673.380 ;
        RECT -28.780 1670.370 -25.780 1670.380 ;
        RECT 45.020 1670.370 48.020 1670.380 ;
        RECT 225.020 1670.370 228.020 1670.380 ;
        RECT 405.020 1670.370 408.020 1670.380 ;
        RECT 585.020 1670.370 588.020 1670.380 ;
        RECT 765.020 1670.370 768.020 1670.380 ;
        RECT 945.020 1670.370 948.020 1670.380 ;
        RECT 1125.020 1670.370 1128.020 1670.380 ;
        RECT 1305.020 1670.370 1308.020 1670.380 ;
        RECT 1485.020 1670.370 1488.020 1670.380 ;
        RECT 1665.020 1670.370 1668.020 1670.380 ;
        RECT 1845.020 1670.370 1848.020 1670.380 ;
        RECT 2025.020 1670.370 2028.020 1670.380 ;
        RECT 2205.020 1670.370 2208.020 1670.380 ;
        RECT 2385.020 1670.370 2388.020 1670.380 ;
        RECT 2565.020 1670.370 2568.020 1670.380 ;
        RECT 2745.020 1670.370 2748.020 1670.380 ;
        RECT 2945.400 1670.370 2948.400 1670.380 ;
        RECT -28.780 1493.380 -25.780 1493.390 ;
        RECT 45.020 1493.380 48.020 1493.390 ;
        RECT 225.020 1493.380 228.020 1493.390 ;
        RECT 405.020 1493.380 408.020 1493.390 ;
        RECT 585.020 1493.380 588.020 1493.390 ;
        RECT 765.020 1493.380 768.020 1493.390 ;
        RECT 945.020 1493.380 948.020 1493.390 ;
        RECT 1125.020 1493.380 1128.020 1493.390 ;
        RECT 1305.020 1493.380 1308.020 1493.390 ;
        RECT 1485.020 1493.380 1488.020 1493.390 ;
        RECT 1665.020 1493.380 1668.020 1493.390 ;
        RECT 1845.020 1493.380 1848.020 1493.390 ;
        RECT 2025.020 1493.380 2028.020 1493.390 ;
        RECT 2205.020 1493.380 2208.020 1493.390 ;
        RECT 2385.020 1493.380 2388.020 1493.390 ;
        RECT 2565.020 1493.380 2568.020 1493.390 ;
        RECT 2745.020 1493.380 2748.020 1493.390 ;
        RECT 2945.400 1493.380 2948.400 1493.390 ;
        RECT -33.480 1490.380 2953.100 1493.380 ;
        RECT -28.780 1490.370 -25.780 1490.380 ;
        RECT 45.020 1490.370 48.020 1490.380 ;
        RECT 225.020 1490.370 228.020 1490.380 ;
        RECT 405.020 1490.370 408.020 1490.380 ;
        RECT 585.020 1490.370 588.020 1490.380 ;
        RECT 765.020 1490.370 768.020 1490.380 ;
        RECT 945.020 1490.370 948.020 1490.380 ;
        RECT 1125.020 1490.370 1128.020 1490.380 ;
        RECT 1305.020 1490.370 1308.020 1490.380 ;
        RECT 1485.020 1490.370 1488.020 1490.380 ;
        RECT 1665.020 1490.370 1668.020 1490.380 ;
        RECT 1845.020 1490.370 1848.020 1490.380 ;
        RECT 2025.020 1490.370 2028.020 1490.380 ;
        RECT 2205.020 1490.370 2208.020 1490.380 ;
        RECT 2385.020 1490.370 2388.020 1490.380 ;
        RECT 2565.020 1490.370 2568.020 1490.380 ;
        RECT 2745.020 1490.370 2748.020 1490.380 ;
        RECT 2945.400 1490.370 2948.400 1490.380 ;
        RECT -28.780 1313.380 -25.780 1313.390 ;
        RECT 45.020 1313.380 48.020 1313.390 ;
        RECT 225.020 1313.380 228.020 1313.390 ;
        RECT 405.020 1313.380 408.020 1313.390 ;
        RECT 585.020 1313.380 588.020 1313.390 ;
        RECT 765.020 1313.380 768.020 1313.390 ;
        RECT 945.020 1313.380 948.020 1313.390 ;
        RECT 1125.020 1313.380 1128.020 1313.390 ;
        RECT 1305.020 1313.380 1308.020 1313.390 ;
        RECT 1485.020 1313.380 1488.020 1313.390 ;
        RECT 1665.020 1313.380 1668.020 1313.390 ;
        RECT 1845.020 1313.380 1848.020 1313.390 ;
        RECT 2025.020 1313.380 2028.020 1313.390 ;
        RECT 2205.020 1313.380 2208.020 1313.390 ;
        RECT 2385.020 1313.380 2388.020 1313.390 ;
        RECT 2565.020 1313.380 2568.020 1313.390 ;
        RECT 2745.020 1313.380 2748.020 1313.390 ;
        RECT 2945.400 1313.380 2948.400 1313.390 ;
        RECT -33.480 1310.380 2953.100 1313.380 ;
        RECT -28.780 1310.370 -25.780 1310.380 ;
        RECT 45.020 1310.370 48.020 1310.380 ;
        RECT 225.020 1310.370 228.020 1310.380 ;
        RECT 405.020 1310.370 408.020 1310.380 ;
        RECT 585.020 1310.370 588.020 1310.380 ;
        RECT 765.020 1310.370 768.020 1310.380 ;
        RECT 945.020 1310.370 948.020 1310.380 ;
        RECT 1125.020 1310.370 1128.020 1310.380 ;
        RECT 1305.020 1310.370 1308.020 1310.380 ;
        RECT 1485.020 1310.370 1488.020 1310.380 ;
        RECT 1665.020 1310.370 1668.020 1310.380 ;
        RECT 1845.020 1310.370 1848.020 1310.380 ;
        RECT 2025.020 1310.370 2028.020 1310.380 ;
        RECT 2205.020 1310.370 2208.020 1310.380 ;
        RECT 2385.020 1310.370 2388.020 1310.380 ;
        RECT 2565.020 1310.370 2568.020 1310.380 ;
        RECT 2745.020 1310.370 2748.020 1310.380 ;
        RECT 2945.400 1310.370 2948.400 1310.380 ;
        RECT -28.780 1133.380 -25.780 1133.390 ;
        RECT 45.020 1133.380 48.020 1133.390 ;
        RECT 225.020 1133.380 228.020 1133.390 ;
        RECT 405.020 1133.380 408.020 1133.390 ;
        RECT 585.020 1133.380 588.020 1133.390 ;
        RECT 765.020 1133.380 768.020 1133.390 ;
        RECT 945.020 1133.380 948.020 1133.390 ;
        RECT 1125.020 1133.380 1128.020 1133.390 ;
        RECT 1305.020 1133.380 1308.020 1133.390 ;
        RECT 1485.020 1133.380 1488.020 1133.390 ;
        RECT 1665.020 1133.380 1668.020 1133.390 ;
        RECT 1845.020 1133.380 1848.020 1133.390 ;
        RECT 2025.020 1133.380 2028.020 1133.390 ;
        RECT 2205.020 1133.380 2208.020 1133.390 ;
        RECT 2385.020 1133.380 2388.020 1133.390 ;
        RECT 2565.020 1133.380 2568.020 1133.390 ;
        RECT 2745.020 1133.380 2748.020 1133.390 ;
        RECT 2945.400 1133.380 2948.400 1133.390 ;
        RECT -33.480 1130.380 2953.100 1133.380 ;
        RECT -28.780 1130.370 -25.780 1130.380 ;
        RECT 45.020 1130.370 48.020 1130.380 ;
        RECT 225.020 1130.370 228.020 1130.380 ;
        RECT 405.020 1130.370 408.020 1130.380 ;
        RECT 585.020 1130.370 588.020 1130.380 ;
        RECT 765.020 1130.370 768.020 1130.380 ;
        RECT 945.020 1130.370 948.020 1130.380 ;
        RECT 1125.020 1130.370 1128.020 1130.380 ;
        RECT 1305.020 1130.370 1308.020 1130.380 ;
        RECT 1485.020 1130.370 1488.020 1130.380 ;
        RECT 1665.020 1130.370 1668.020 1130.380 ;
        RECT 1845.020 1130.370 1848.020 1130.380 ;
        RECT 2025.020 1130.370 2028.020 1130.380 ;
        RECT 2205.020 1130.370 2208.020 1130.380 ;
        RECT 2385.020 1130.370 2388.020 1130.380 ;
        RECT 2565.020 1130.370 2568.020 1130.380 ;
        RECT 2745.020 1130.370 2748.020 1130.380 ;
        RECT 2945.400 1130.370 2948.400 1130.380 ;
        RECT -28.780 953.380 -25.780 953.390 ;
        RECT 45.020 953.380 48.020 953.390 ;
        RECT 225.020 953.380 228.020 953.390 ;
        RECT 405.020 953.380 408.020 953.390 ;
        RECT 585.020 953.380 588.020 953.390 ;
        RECT 765.020 953.380 768.020 953.390 ;
        RECT 945.020 953.380 948.020 953.390 ;
        RECT 1125.020 953.380 1128.020 953.390 ;
        RECT 1305.020 953.380 1308.020 953.390 ;
        RECT 1485.020 953.380 1488.020 953.390 ;
        RECT 1665.020 953.380 1668.020 953.390 ;
        RECT 1845.020 953.380 1848.020 953.390 ;
        RECT 2025.020 953.380 2028.020 953.390 ;
        RECT 2205.020 953.380 2208.020 953.390 ;
        RECT 2385.020 953.380 2388.020 953.390 ;
        RECT 2565.020 953.380 2568.020 953.390 ;
        RECT 2745.020 953.380 2748.020 953.390 ;
        RECT 2945.400 953.380 2948.400 953.390 ;
        RECT -33.480 950.380 2953.100 953.380 ;
        RECT -28.780 950.370 -25.780 950.380 ;
        RECT 45.020 950.370 48.020 950.380 ;
        RECT 225.020 950.370 228.020 950.380 ;
        RECT 405.020 950.370 408.020 950.380 ;
        RECT 585.020 950.370 588.020 950.380 ;
        RECT 765.020 950.370 768.020 950.380 ;
        RECT 945.020 950.370 948.020 950.380 ;
        RECT 1125.020 950.370 1128.020 950.380 ;
        RECT 1305.020 950.370 1308.020 950.380 ;
        RECT 1485.020 950.370 1488.020 950.380 ;
        RECT 1665.020 950.370 1668.020 950.380 ;
        RECT 1845.020 950.370 1848.020 950.380 ;
        RECT 2025.020 950.370 2028.020 950.380 ;
        RECT 2205.020 950.370 2208.020 950.380 ;
        RECT 2385.020 950.370 2388.020 950.380 ;
        RECT 2565.020 950.370 2568.020 950.380 ;
        RECT 2745.020 950.370 2748.020 950.380 ;
        RECT 2945.400 950.370 2948.400 950.380 ;
        RECT -28.780 773.380 -25.780 773.390 ;
        RECT 45.020 773.380 48.020 773.390 ;
        RECT 225.020 773.380 228.020 773.390 ;
        RECT 405.020 773.380 408.020 773.390 ;
        RECT 585.020 773.380 588.020 773.390 ;
        RECT 765.020 773.380 768.020 773.390 ;
        RECT 945.020 773.380 948.020 773.390 ;
        RECT 1125.020 773.380 1128.020 773.390 ;
        RECT 1305.020 773.380 1308.020 773.390 ;
        RECT 1485.020 773.380 1488.020 773.390 ;
        RECT 1665.020 773.380 1668.020 773.390 ;
        RECT 1845.020 773.380 1848.020 773.390 ;
        RECT 2025.020 773.380 2028.020 773.390 ;
        RECT 2205.020 773.380 2208.020 773.390 ;
        RECT 2385.020 773.380 2388.020 773.390 ;
        RECT 2565.020 773.380 2568.020 773.390 ;
        RECT 2745.020 773.380 2748.020 773.390 ;
        RECT 2945.400 773.380 2948.400 773.390 ;
        RECT -33.480 770.380 2953.100 773.380 ;
        RECT -28.780 770.370 -25.780 770.380 ;
        RECT 45.020 770.370 48.020 770.380 ;
        RECT 225.020 770.370 228.020 770.380 ;
        RECT 405.020 770.370 408.020 770.380 ;
        RECT 585.020 770.370 588.020 770.380 ;
        RECT 765.020 770.370 768.020 770.380 ;
        RECT 945.020 770.370 948.020 770.380 ;
        RECT 1125.020 770.370 1128.020 770.380 ;
        RECT 1305.020 770.370 1308.020 770.380 ;
        RECT 1485.020 770.370 1488.020 770.380 ;
        RECT 1665.020 770.370 1668.020 770.380 ;
        RECT 1845.020 770.370 1848.020 770.380 ;
        RECT 2025.020 770.370 2028.020 770.380 ;
        RECT 2205.020 770.370 2208.020 770.380 ;
        RECT 2385.020 770.370 2388.020 770.380 ;
        RECT 2565.020 770.370 2568.020 770.380 ;
        RECT 2745.020 770.370 2748.020 770.380 ;
        RECT 2945.400 770.370 2948.400 770.380 ;
        RECT -28.780 593.380 -25.780 593.390 ;
        RECT 45.020 593.380 48.020 593.390 ;
        RECT 225.020 593.380 228.020 593.390 ;
        RECT 405.020 593.380 408.020 593.390 ;
        RECT 585.020 593.380 588.020 593.390 ;
        RECT 765.020 593.380 768.020 593.390 ;
        RECT 945.020 593.380 948.020 593.390 ;
        RECT 1125.020 593.380 1128.020 593.390 ;
        RECT 1305.020 593.380 1308.020 593.390 ;
        RECT 1485.020 593.380 1488.020 593.390 ;
        RECT 1665.020 593.380 1668.020 593.390 ;
        RECT 1845.020 593.380 1848.020 593.390 ;
        RECT 2025.020 593.380 2028.020 593.390 ;
        RECT 2205.020 593.380 2208.020 593.390 ;
        RECT 2385.020 593.380 2388.020 593.390 ;
        RECT 2565.020 593.380 2568.020 593.390 ;
        RECT 2745.020 593.380 2748.020 593.390 ;
        RECT 2945.400 593.380 2948.400 593.390 ;
        RECT -33.480 590.380 2953.100 593.380 ;
        RECT -28.780 590.370 -25.780 590.380 ;
        RECT 45.020 590.370 48.020 590.380 ;
        RECT 225.020 590.370 228.020 590.380 ;
        RECT 405.020 590.370 408.020 590.380 ;
        RECT 585.020 590.370 588.020 590.380 ;
        RECT 765.020 590.370 768.020 590.380 ;
        RECT 945.020 590.370 948.020 590.380 ;
        RECT 1125.020 590.370 1128.020 590.380 ;
        RECT 1305.020 590.370 1308.020 590.380 ;
        RECT 1485.020 590.370 1488.020 590.380 ;
        RECT 1665.020 590.370 1668.020 590.380 ;
        RECT 1845.020 590.370 1848.020 590.380 ;
        RECT 2025.020 590.370 2028.020 590.380 ;
        RECT 2205.020 590.370 2208.020 590.380 ;
        RECT 2385.020 590.370 2388.020 590.380 ;
        RECT 2565.020 590.370 2568.020 590.380 ;
        RECT 2745.020 590.370 2748.020 590.380 ;
        RECT 2945.400 590.370 2948.400 590.380 ;
        RECT -28.780 413.380 -25.780 413.390 ;
        RECT 45.020 413.380 48.020 413.390 ;
        RECT 225.020 413.380 228.020 413.390 ;
        RECT 405.020 413.380 408.020 413.390 ;
        RECT 585.020 413.380 588.020 413.390 ;
        RECT 765.020 413.380 768.020 413.390 ;
        RECT 945.020 413.380 948.020 413.390 ;
        RECT 1125.020 413.380 1128.020 413.390 ;
        RECT 1305.020 413.380 1308.020 413.390 ;
        RECT 1485.020 413.380 1488.020 413.390 ;
        RECT 1665.020 413.380 1668.020 413.390 ;
        RECT 1845.020 413.380 1848.020 413.390 ;
        RECT 2025.020 413.380 2028.020 413.390 ;
        RECT 2205.020 413.380 2208.020 413.390 ;
        RECT 2385.020 413.380 2388.020 413.390 ;
        RECT 2565.020 413.380 2568.020 413.390 ;
        RECT 2745.020 413.380 2748.020 413.390 ;
        RECT 2945.400 413.380 2948.400 413.390 ;
        RECT -33.480 410.380 2953.100 413.380 ;
        RECT -28.780 410.370 -25.780 410.380 ;
        RECT 45.020 410.370 48.020 410.380 ;
        RECT 225.020 410.370 228.020 410.380 ;
        RECT 405.020 410.370 408.020 410.380 ;
        RECT 585.020 410.370 588.020 410.380 ;
        RECT 765.020 410.370 768.020 410.380 ;
        RECT 945.020 410.370 948.020 410.380 ;
        RECT 1125.020 410.370 1128.020 410.380 ;
        RECT 1305.020 410.370 1308.020 410.380 ;
        RECT 1485.020 410.370 1488.020 410.380 ;
        RECT 1665.020 410.370 1668.020 410.380 ;
        RECT 1845.020 410.370 1848.020 410.380 ;
        RECT 2025.020 410.370 2028.020 410.380 ;
        RECT 2205.020 410.370 2208.020 410.380 ;
        RECT 2385.020 410.370 2388.020 410.380 ;
        RECT 2565.020 410.370 2568.020 410.380 ;
        RECT 2745.020 410.370 2748.020 410.380 ;
        RECT 2945.400 410.370 2948.400 410.380 ;
        RECT -28.780 233.380 -25.780 233.390 ;
        RECT 45.020 233.380 48.020 233.390 ;
        RECT 225.020 233.380 228.020 233.390 ;
        RECT 405.020 233.380 408.020 233.390 ;
        RECT 585.020 233.380 588.020 233.390 ;
        RECT 765.020 233.380 768.020 233.390 ;
        RECT 945.020 233.380 948.020 233.390 ;
        RECT 1125.020 233.380 1128.020 233.390 ;
        RECT 1305.020 233.380 1308.020 233.390 ;
        RECT 1485.020 233.380 1488.020 233.390 ;
        RECT 1665.020 233.380 1668.020 233.390 ;
        RECT 1845.020 233.380 1848.020 233.390 ;
        RECT 2025.020 233.380 2028.020 233.390 ;
        RECT 2205.020 233.380 2208.020 233.390 ;
        RECT 2385.020 233.380 2388.020 233.390 ;
        RECT 2565.020 233.380 2568.020 233.390 ;
        RECT 2745.020 233.380 2748.020 233.390 ;
        RECT 2945.400 233.380 2948.400 233.390 ;
        RECT -33.480 230.380 2953.100 233.380 ;
        RECT -28.780 230.370 -25.780 230.380 ;
        RECT 45.020 230.370 48.020 230.380 ;
        RECT 225.020 230.370 228.020 230.380 ;
        RECT 405.020 230.370 408.020 230.380 ;
        RECT 585.020 230.370 588.020 230.380 ;
        RECT 765.020 230.370 768.020 230.380 ;
        RECT 945.020 230.370 948.020 230.380 ;
        RECT 1125.020 230.370 1128.020 230.380 ;
        RECT 1305.020 230.370 1308.020 230.380 ;
        RECT 1485.020 230.370 1488.020 230.380 ;
        RECT 1665.020 230.370 1668.020 230.380 ;
        RECT 1845.020 230.370 1848.020 230.380 ;
        RECT 2025.020 230.370 2028.020 230.380 ;
        RECT 2205.020 230.370 2208.020 230.380 ;
        RECT 2385.020 230.370 2388.020 230.380 ;
        RECT 2565.020 230.370 2568.020 230.380 ;
        RECT 2745.020 230.370 2748.020 230.380 ;
        RECT 2945.400 230.370 2948.400 230.380 ;
        RECT -28.780 53.380 -25.780 53.390 ;
        RECT 45.020 53.380 48.020 53.390 ;
        RECT 225.020 53.380 228.020 53.390 ;
        RECT 405.020 53.380 408.020 53.390 ;
        RECT 585.020 53.380 588.020 53.390 ;
        RECT 765.020 53.380 768.020 53.390 ;
        RECT 945.020 53.380 948.020 53.390 ;
        RECT 1125.020 53.380 1128.020 53.390 ;
        RECT 1305.020 53.380 1308.020 53.390 ;
        RECT 1485.020 53.380 1488.020 53.390 ;
        RECT 1665.020 53.380 1668.020 53.390 ;
        RECT 1845.020 53.380 1848.020 53.390 ;
        RECT 2025.020 53.380 2028.020 53.390 ;
        RECT 2205.020 53.380 2208.020 53.390 ;
        RECT 2385.020 53.380 2388.020 53.390 ;
        RECT 2565.020 53.380 2568.020 53.390 ;
        RECT 2745.020 53.380 2748.020 53.390 ;
        RECT 2945.400 53.380 2948.400 53.390 ;
        RECT -33.480 50.380 2953.100 53.380 ;
        RECT -28.780 50.370 -25.780 50.380 ;
        RECT 45.020 50.370 48.020 50.380 ;
        RECT 225.020 50.370 228.020 50.380 ;
        RECT 405.020 50.370 408.020 50.380 ;
        RECT 585.020 50.370 588.020 50.380 ;
        RECT 765.020 50.370 768.020 50.380 ;
        RECT 945.020 50.370 948.020 50.380 ;
        RECT 1125.020 50.370 1128.020 50.380 ;
        RECT 1305.020 50.370 1308.020 50.380 ;
        RECT 1485.020 50.370 1488.020 50.380 ;
        RECT 1665.020 50.370 1668.020 50.380 ;
        RECT 1845.020 50.370 1848.020 50.380 ;
        RECT 2025.020 50.370 2028.020 50.380 ;
        RECT 2205.020 50.370 2208.020 50.380 ;
        RECT 2385.020 50.370 2388.020 50.380 ;
        RECT 2565.020 50.370 2568.020 50.380 ;
        RECT 2745.020 50.370 2748.020 50.380 ;
        RECT 2945.400 50.370 2948.400 50.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 45.020 -20.420 48.020 -20.410 ;
        RECT 225.020 -20.420 228.020 -20.410 ;
        RECT 405.020 -20.420 408.020 -20.410 ;
        RECT 585.020 -20.420 588.020 -20.410 ;
        RECT 765.020 -20.420 768.020 -20.410 ;
        RECT 945.020 -20.420 948.020 -20.410 ;
        RECT 1125.020 -20.420 1128.020 -20.410 ;
        RECT 1305.020 -20.420 1308.020 -20.410 ;
        RECT 1485.020 -20.420 1488.020 -20.410 ;
        RECT 1665.020 -20.420 1668.020 -20.410 ;
        RECT 1845.020 -20.420 1848.020 -20.410 ;
        RECT 2025.020 -20.420 2028.020 -20.410 ;
        RECT 2205.020 -20.420 2208.020 -20.410 ;
        RECT 2385.020 -20.420 2388.020 -20.410 ;
        RECT 2565.020 -20.420 2568.020 -20.410 ;
        RECT 2745.020 -20.420 2748.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 45.020 -23.430 48.020 -23.420 ;
        RECT 225.020 -23.430 228.020 -23.420 ;
        RECT 405.020 -23.430 408.020 -23.420 ;
        RECT 585.020 -23.430 588.020 -23.420 ;
        RECT 765.020 -23.430 768.020 -23.420 ;
        RECT 945.020 -23.430 948.020 -23.420 ;
        RECT 1125.020 -23.430 1128.020 -23.420 ;
        RECT 1305.020 -23.430 1308.020 -23.420 ;
        RECT 1485.020 -23.430 1488.020 -23.420 ;
        RECT 1665.020 -23.430 1668.020 -23.420 ;
        RECT 1845.020 -23.430 1848.020 -23.420 ;
        RECT 2025.020 -23.430 2028.020 -23.420 ;
        RECT 2205.020 -23.430 2208.020 -23.420 ;
        RECT 2385.020 -23.430 2388.020 -23.420 ;
        RECT 2565.020 -23.430 2568.020 -23.420 ;
        RECT 2745.020 -23.430 2748.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 135.020 -28.120 138.020 3547.800 ;
        RECT 315.020 -28.120 318.020 3547.800 ;
        RECT 495.020 -28.120 498.020 3547.800 ;
        RECT 675.020 -28.120 678.020 3547.800 ;
        RECT 855.020 -28.120 858.020 3547.800 ;
        RECT 1035.020 -28.120 1038.020 3547.800 ;
        RECT 1215.020 -28.120 1218.020 3547.800 ;
        RECT 1395.020 -28.120 1398.020 3547.800 ;
        RECT 1575.020 -28.120 1578.020 3547.800 ;
        RECT 1755.020 -28.120 1758.020 3547.800 ;
        RECT 1935.020 -28.120 1938.020 3547.800 ;
        RECT 2115.020 -28.120 2118.020 3547.800 ;
        RECT 2295.020 -28.120 2298.020 3547.800 ;
        RECT 2475.020 -28.120 2478.020 3547.800 ;
        RECT 2655.020 -28.120 2658.020 3547.800 ;
        RECT 2835.020 -28.120 2838.020 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 3382.090 -31.390 3383.270 ;
        RECT -32.570 3380.490 -31.390 3381.670 ;
        RECT -32.570 3202.090 -31.390 3203.270 ;
        RECT -32.570 3200.490 -31.390 3201.670 ;
        RECT -32.570 3022.090 -31.390 3023.270 ;
        RECT -32.570 3020.490 -31.390 3021.670 ;
        RECT -32.570 2842.090 -31.390 2843.270 ;
        RECT -32.570 2840.490 -31.390 2841.670 ;
        RECT -32.570 2662.090 -31.390 2663.270 ;
        RECT -32.570 2660.490 -31.390 2661.670 ;
        RECT -32.570 2482.090 -31.390 2483.270 ;
        RECT -32.570 2480.490 -31.390 2481.670 ;
        RECT -32.570 2302.090 -31.390 2303.270 ;
        RECT -32.570 2300.490 -31.390 2301.670 ;
        RECT -32.570 2122.090 -31.390 2123.270 ;
        RECT -32.570 2120.490 -31.390 2121.670 ;
        RECT -32.570 1942.090 -31.390 1943.270 ;
        RECT -32.570 1940.490 -31.390 1941.670 ;
        RECT -32.570 1762.090 -31.390 1763.270 ;
        RECT -32.570 1760.490 -31.390 1761.670 ;
        RECT -32.570 1582.090 -31.390 1583.270 ;
        RECT -32.570 1580.490 -31.390 1581.670 ;
        RECT -32.570 1402.090 -31.390 1403.270 ;
        RECT -32.570 1400.490 -31.390 1401.670 ;
        RECT -32.570 1222.090 -31.390 1223.270 ;
        RECT -32.570 1220.490 -31.390 1221.670 ;
        RECT -32.570 1042.090 -31.390 1043.270 ;
        RECT -32.570 1040.490 -31.390 1041.670 ;
        RECT -32.570 862.090 -31.390 863.270 ;
        RECT -32.570 860.490 -31.390 861.670 ;
        RECT -32.570 682.090 -31.390 683.270 ;
        RECT -32.570 680.490 -31.390 681.670 ;
        RECT -32.570 502.090 -31.390 503.270 ;
        RECT -32.570 500.490 -31.390 501.670 ;
        RECT -32.570 322.090 -31.390 323.270 ;
        RECT -32.570 320.490 -31.390 321.670 ;
        RECT -32.570 142.090 -31.390 143.270 ;
        RECT -32.570 140.490 -31.390 141.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 135.930 3546.510 137.110 3547.690 ;
        RECT 135.930 3544.910 137.110 3546.090 ;
        RECT 135.930 3382.090 137.110 3383.270 ;
        RECT 135.930 3380.490 137.110 3381.670 ;
        RECT 135.930 3202.090 137.110 3203.270 ;
        RECT 135.930 3200.490 137.110 3201.670 ;
        RECT 135.930 3022.090 137.110 3023.270 ;
        RECT 135.930 3020.490 137.110 3021.670 ;
        RECT 135.930 2842.090 137.110 2843.270 ;
        RECT 135.930 2840.490 137.110 2841.670 ;
        RECT 135.930 2662.090 137.110 2663.270 ;
        RECT 135.930 2660.490 137.110 2661.670 ;
        RECT 135.930 2482.090 137.110 2483.270 ;
        RECT 135.930 2480.490 137.110 2481.670 ;
        RECT 135.930 2302.090 137.110 2303.270 ;
        RECT 135.930 2300.490 137.110 2301.670 ;
        RECT 135.930 2122.090 137.110 2123.270 ;
        RECT 135.930 2120.490 137.110 2121.670 ;
        RECT 135.930 1942.090 137.110 1943.270 ;
        RECT 135.930 1940.490 137.110 1941.670 ;
        RECT 135.930 1762.090 137.110 1763.270 ;
        RECT 135.930 1760.490 137.110 1761.670 ;
        RECT 135.930 1582.090 137.110 1583.270 ;
        RECT 135.930 1580.490 137.110 1581.670 ;
        RECT 135.930 1402.090 137.110 1403.270 ;
        RECT 135.930 1400.490 137.110 1401.670 ;
        RECT 135.930 1222.090 137.110 1223.270 ;
        RECT 135.930 1220.490 137.110 1221.670 ;
        RECT 135.930 1042.090 137.110 1043.270 ;
        RECT 135.930 1040.490 137.110 1041.670 ;
        RECT 135.930 862.090 137.110 863.270 ;
        RECT 135.930 860.490 137.110 861.670 ;
        RECT 135.930 682.090 137.110 683.270 ;
        RECT 135.930 680.490 137.110 681.670 ;
        RECT 135.930 502.090 137.110 503.270 ;
        RECT 135.930 500.490 137.110 501.670 ;
        RECT 135.930 322.090 137.110 323.270 ;
        RECT 135.930 320.490 137.110 321.670 ;
        RECT 135.930 142.090 137.110 143.270 ;
        RECT 135.930 140.490 137.110 141.670 ;
        RECT 135.930 -26.410 137.110 -25.230 ;
        RECT 135.930 -28.010 137.110 -26.830 ;
        RECT 315.930 3546.510 317.110 3547.690 ;
        RECT 315.930 3544.910 317.110 3546.090 ;
        RECT 315.930 3382.090 317.110 3383.270 ;
        RECT 315.930 3380.490 317.110 3381.670 ;
        RECT 315.930 3202.090 317.110 3203.270 ;
        RECT 315.930 3200.490 317.110 3201.670 ;
        RECT 315.930 3022.090 317.110 3023.270 ;
        RECT 315.930 3020.490 317.110 3021.670 ;
        RECT 315.930 2842.090 317.110 2843.270 ;
        RECT 315.930 2840.490 317.110 2841.670 ;
        RECT 315.930 2662.090 317.110 2663.270 ;
        RECT 315.930 2660.490 317.110 2661.670 ;
        RECT 315.930 2482.090 317.110 2483.270 ;
        RECT 315.930 2480.490 317.110 2481.670 ;
        RECT 315.930 2302.090 317.110 2303.270 ;
        RECT 315.930 2300.490 317.110 2301.670 ;
        RECT 315.930 2122.090 317.110 2123.270 ;
        RECT 315.930 2120.490 317.110 2121.670 ;
        RECT 315.930 1942.090 317.110 1943.270 ;
        RECT 315.930 1940.490 317.110 1941.670 ;
        RECT 315.930 1762.090 317.110 1763.270 ;
        RECT 315.930 1760.490 317.110 1761.670 ;
        RECT 315.930 1582.090 317.110 1583.270 ;
        RECT 315.930 1580.490 317.110 1581.670 ;
        RECT 315.930 1402.090 317.110 1403.270 ;
        RECT 315.930 1400.490 317.110 1401.670 ;
        RECT 315.930 1222.090 317.110 1223.270 ;
        RECT 315.930 1220.490 317.110 1221.670 ;
        RECT 315.930 1042.090 317.110 1043.270 ;
        RECT 315.930 1040.490 317.110 1041.670 ;
        RECT 315.930 862.090 317.110 863.270 ;
        RECT 315.930 860.490 317.110 861.670 ;
        RECT 315.930 682.090 317.110 683.270 ;
        RECT 315.930 680.490 317.110 681.670 ;
        RECT 315.930 502.090 317.110 503.270 ;
        RECT 315.930 500.490 317.110 501.670 ;
        RECT 315.930 322.090 317.110 323.270 ;
        RECT 315.930 320.490 317.110 321.670 ;
        RECT 315.930 142.090 317.110 143.270 ;
        RECT 315.930 140.490 317.110 141.670 ;
        RECT 315.930 -26.410 317.110 -25.230 ;
        RECT 315.930 -28.010 317.110 -26.830 ;
        RECT 495.930 3546.510 497.110 3547.690 ;
        RECT 495.930 3544.910 497.110 3546.090 ;
        RECT 495.930 3382.090 497.110 3383.270 ;
        RECT 495.930 3380.490 497.110 3381.670 ;
        RECT 495.930 3202.090 497.110 3203.270 ;
        RECT 495.930 3200.490 497.110 3201.670 ;
        RECT 495.930 3022.090 497.110 3023.270 ;
        RECT 495.930 3020.490 497.110 3021.670 ;
        RECT 495.930 2842.090 497.110 2843.270 ;
        RECT 495.930 2840.490 497.110 2841.670 ;
        RECT 495.930 2662.090 497.110 2663.270 ;
        RECT 495.930 2660.490 497.110 2661.670 ;
        RECT 495.930 2482.090 497.110 2483.270 ;
        RECT 495.930 2480.490 497.110 2481.670 ;
        RECT 495.930 2302.090 497.110 2303.270 ;
        RECT 495.930 2300.490 497.110 2301.670 ;
        RECT 495.930 2122.090 497.110 2123.270 ;
        RECT 495.930 2120.490 497.110 2121.670 ;
        RECT 495.930 1942.090 497.110 1943.270 ;
        RECT 495.930 1940.490 497.110 1941.670 ;
        RECT 495.930 1762.090 497.110 1763.270 ;
        RECT 495.930 1760.490 497.110 1761.670 ;
        RECT 495.930 1582.090 497.110 1583.270 ;
        RECT 495.930 1580.490 497.110 1581.670 ;
        RECT 495.930 1402.090 497.110 1403.270 ;
        RECT 495.930 1400.490 497.110 1401.670 ;
        RECT 495.930 1222.090 497.110 1223.270 ;
        RECT 495.930 1220.490 497.110 1221.670 ;
        RECT 495.930 1042.090 497.110 1043.270 ;
        RECT 495.930 1040.490 497.110 1041.670 ;
        RECT 495.930 862.090 497.110 863.270 ;
        RECT 495.930 860.490 497.110 861.670 ;
        RECT 495.930 682.090 497.110 683.270 ;
        RECT 495.930 680.490 497.110 681.670 ;
        RECT 495.930 502.090 497.110 503.270 ;
        RECT 495.930 500.490 497.110 501.670 ;
        RECT 495.930 322.090 497.110 323.270 ;
        RECT 495.930 320.490 497.110 321.670 ;
        RECT 495.930 142.090 497.110 143.270 ;
        RECT 495.930 140.490 497.110 141.670 ;
        RECT 495.930 -26.410 497.110 -25.230 ;
        RECT 495.930 -28.010 497.110 -26.830 ;
        RECT 675.930 3546.510 677.110 3547.690 ;
        RECT 675.930 3544.910 677.110 3546.090 ;
        RECT 675.930 3382.090 677.110 3383.270 ;
        RECT 675.930 3380.490 677.110 3381.670 ;
        RECT 675.930 3202.090 677.110 3203.270 ;
        RECT 675.930 3200.490 677.110 3201.670 ;
        RECT 675.930 3022.090 677.110 3023.270 ;
        RECT 675.930 3020.490 677.110 3021.670 ;
        RECT 675.930 2842.090 677.110 2843.270 ;
        RECT 675.930 2840.490 677.110 2841.670 ;
        RECT 675.930 2662.090 677.110 2663.270 ;
        RECT 675.930 2660.490 677.110 2661.670 ;
        RECT 675.930 2482.090 677.110 2483.270 ;
        RECT 675.930 2480.490 677.110 2481.670 ;
        RECT 675.930 2302.090 677.110 2303.270 ;
        RECT 675.930 2300.490 677.110 2301.670 ;
        RECT 675.930 2122.090 677.110 2123.270 ;
        RECT 675.930 2120.490 677.110 2121.670 ;
        RECT 675.930 1942.090 677.110 1943.270 ;
        RECT 675.930 1940.490 677.110 1941.670 ;
        RECT 675.930 1762.090 677.110 1763.270 ;
        RECT 675.930 1760.490 677.110 1761.670 ;
        RECT 675.930 1582.090 677.110 1583.270 ;
        RECT 675.930 1580.490 677.110 1581.670 ;
        RECT 675.930 1402.090 677.110 1403.270 ;
        RECT 675.930 1400.490 677.110 1401.670 ;
        RECT 675.930 1222.090 677.110 1223.270 ;
        RECT 675.930 1220.490 677.110 1221.670 ;
        RECT 675.930 1042.090 677.110 1043.270 ;
        RECT 675.930 1040.490 677.110 1041.670 ;
        RECT 675.930 862.090 677.110 863.270 ;
        RECT 675.930 860.490 677.110 861.670 ;
        RECT 675.930 682.090 677.110 683.270 ;
        RECT 675.930 680.490 677.110 681.670 ;
        RECT 675.930 502.090 677.110 503.270 ;
        RECT 675.930 500.490 677.110 501.670 ;
        RECT 675.930 322.090 677.110 323.270 ;
        RECT 675.930 320.490 677.110 321.670 ;
        RECT 675.930 142.090 677.110 143.270 ;
        RECT 675.930 140.490 677.110 141.670 ;
        RECT 675.930 -26.410 677.110 -25.230 ;
        RECT 675.930 -28.010 677.110 -26.830 ;
        RECT 855.930 3546.510 857.110 3547.690 ;
        RECT 855.930 3544.910 857.110 3546.090 ;
        RECT 855.930 3382.090 857.110 3383.270 ;
        RECT 855.930 3380.490 857.110 3381.670 ;
        RECT 855.930 3202.090 857.110 3203.270 ;
        RECT 855.930 3200.490 857.110 3201.670 ;
        RECT 855.930 3022.090 857.110 3023.270 ;
        RECT 855.930 3020.490 857.110 3021.670 ;
        RECT 855.930 2842.090 857.110 2843.270 ;
        RECT 855.930 2840.490 857.110 2841.670 ;
        RECT 855.930 2662.090 857.110 2663.270 ;
        RECT 855.930 2660.490 857.110 2661.670 ;
        RECT 855.930 2482.090 857.110 2483.270 ;
        RECT 855.930 2480.490 857.110 2481.670 ;
        RECT 855.930 2302.090 857.110 2303.270 ;
        RECT 855.930 2300.490 857.110 2301.670 ;
        RECT 855.930 2122.090 857.110 2123.270 ;
        RECT 855.930 2120.490 857.110 2121.670 ;
        RECT 855.930 1942.090 857.110 1943.270 ;
        RECT 855.930 1940.490 857.110 1941.670 ;
        RECT 855.930 1762.090 857.110 1763.270 ;
        RECT 855.930 1760.490 857.110 1761.670 ;
        RECT 855.930 1582.090 857.110 1583.270 ;
        RECT 855.930 1580.490 857.110 1581.670 ;
        RECT 855.930 1402.090 857.110 1403.270 ;
        RECT 855.930 1400.490 857.110 1401.670 ;
        RECT 855.930 1222.090 857.110 1223.270 ;
        RECT 855.930 1220.490 857.110 1221.670 ;
        RECT 855.930 1042.090 857.110 1043.270 ;
        RECT 855.930 1040.490 857.110 1041.670 ;
        RECT 855.930 862.090 857.110 863.270 ;
        RECT 855.930 860.490 857.110 861.670 ;
        RECT 855.930 682.090 857.110 683.270 ;
        RECT 855.930 680.490 857.110 681.670 ;
        RECT 855.930 502.090 857.110 503.270 ;
        RECT 855.930 500.490 857.110 501.670 ;
        RECT 855.930 322.090 857.110 323.270 ;
        RECT 855.930 320.490 857.110 321.670 ;
        RECT 855.930 142.090 857.110 143.270 ;
        RECT 855.930 140.490 857.110 141.670 ;
        RECT 855.930 -26.410 857.110 -25.230 ;
        RECT 855.930 -28.010 857.110 -26.830 ;
        RECT 1035.930 3546.510 1037.110 3547.690 ;
        RECT 1035.930 3544.910 1037.110 3546.090 ;
        RECT 1035.930 3382.090 1037.110 3383.270 ;
        RECT 1035.930 3380.490 1037.110 3381.670 ;
        RECT 1035.930 3202.090 1037.110 3203.270 ;
        RECT 1035.930 3200.490 1037.110 3201.670 ;
        RECT 1035.930 3022.090 1037.110 3023.270 ;
        RECT 1035.930 3020.490 1037.110 3021.670 ;
        RECT 1035.930 2842.090 1037.110 2843.270 ;
        RECT 1035.930 2840.490 1037.110 2841.670 ;
        RECT 1035.930 2662.090 1037.110 2663.270 ;
        RECT 1035.930 2660.490 1037.110 2661.670 ;
        RECT 1035.930 2482.090 1037.110 2483.270 ;
        RECT 1035.930 2480.490 1037.110 2481.670 ;
        RECT 1035.930 2302.090 1037.110 2303.270 ;
        RECT 1035.930 2300.490 1037.110 2301.670 ;
        RECT 1035.930 2122.090 1037.110 2123.270 ;
        RECT 1035.930 2120.490 1037.110 2121.670 ;
        RECT 1035.930 1942.090 1037.110 1943.270 ;
        RECT 1035.930 1940.490 1037.110 1941.670 ;
        RECT 1035.930 1762.090 1037.110 1763.270 ;
        RECT 1035.930 1760.490 1037.110 1761.670 ;
        RECT 1035.930 1582.090 1037.110 1583.270 ;
        RECT 1035.930 1580.490 1037.110 1581.670 ;
        RECT 1035.930 1402.090 1037.110 1403.270 ;
        RECT 1035.930 1400.490 1037.110 1401.670 ;
        RECT 1035.930 1222.090 1037.110 1223.270 ;
        RECT 1035.930 1220.490 1037.110 1221.670 ;
        RECT 1035.930 1042.090 1037.110 1043.270 ;
        RECT 1035.930 1040.490 1037.110 1041.670 ;
        RECT 1035.930 862.090 1037.110 863.270 ;
        RECT 1035.930 860.490 1037.110 861.670 ;
        RECT 1035.930 682.090 1037.110 683.270 ;
        RECT 1035.930 680.490 1037.110 681.670 ;
        RECT 1035.930 502.090 1037.110 503.270 ;
        RECT 1035.930 500.490 1037.110 501.670 ;
        RECT 1035.930 322.090 1037.110 323.270 ;
        RECT 1035.930 320.490 1037.110 321.670 ;
        RECT 1035.930 142.090 1037.110 143.270 ;
        RECT 1035.930 140.490 1037.110 141.670 ;
        RECT 1035.930 -26.410 1037.110 -25.230 ;
        RECT 1035.930 -28.010 1037.110 -26.830 ;
        RECT 1215.930 3546.510 1217.110 3547.690 ;
        RECT 1215.930 3544.910 1217.110 3546.090 ;
        RECT 1215.930 3382.090 1217.110 3383.270 ;
        RECT 1215.930 3380.490 1217.110 3381.670 ;
        RECT 1215.930 3202.090 1217.110 3203.270 ;
        RECT 1215.930 3200.490 1217.110 3201.670 ;
        RECT 1215.930 3022.090 1217.110 3023.270 ;
        RECT 1215.930 3020.490 1217.110 3021.670 ;
        RECT 1215.930 2842.090 1217.110 2843.270 ;
        RECT 1215.930 2840.490 1217.110 2841.670 ;
        RECT 1215.930 2662.090 1217.110 2663.270 ;
        RECT 1215.930 2660.490 1217.110 2661.670 ;
        RECT 1215.930 2482.090 1217.110 2483.270 ;
        RECT 1215.930 2480.490 1217.110 2481.670 ;
        RECT 1215.930 2302.090 1217.110 2303.270 ;
        RECT 1215.930 2300.490 1217.110 2301.670 ;
        RECT 1215.930 2122.090 1217.110 2123.270 ;
        RECT 1215.930 2120.490 1217.110 2121.670 ;
        RECT 1215.930 1942.090 1217.110 1943.270 ;
        RECT 1215.930 1940.490 1217.110 1941.670 ;
        RECT 1215.930 1762.090 1217.110 1763.270 ;
        RECT 1215.930 1760.490 1217.110 1761.670 ;
        RECT 1215.930 1582.090 1217.110 1583.270 ;
        RECT 1215.930 1580.490 1217.110 1581.670 ;
        RECT 1215.930 1402.090 1217.110 1403.270 ;
        RECT 1215.930 1400.490 1217.110 1401.670 ;
        RECT 1215.930 1222.090 1217.110 1223.270 ;
        RECT 1215.930 1220.490 1217.110 1221.670 ;
        RECT 1215.930 1042.090 1217.110 1043.270 ;
        RECT 1215.930 1040.490 1217.110 1041.670 ;
        RECT 1215.930 862.090 1217.110 863.270 ;
        RECT 1215.930 860.490 1217.110 861.670 ;
        RECT 1215.930 682.090 1217.110 683.270 ;
        RECT 1215.930 680.490 1217.110 681.670 ;
        RECT 1215.930 502.090 1217.110 503.270 ;
        RECT 1215.930 500.490 1217.110 501.670 ;
        RECT 1215.930 322.090 1217.110 323.270 ;
        RECT 1215.930 320.490 1217.110 321.670 ;
        RECT 1215.930 142.090 1217.110 143.270 ;
        RECT 1215.930 140.490 1217.110 141.670 ;
        RECT 1215.930 -26.410 1217.110 -25.230 ;
        RECT 1215.930 -28.010 1217.110 -26.830 ;
        RECT 1395.930 3546.510 1397.110 3547.690 ;
        RECT 1395.930 3544.910 1397.110 3546.090 ;
        RECT 1395.930 3382.090 1397.110 3383.270 ;
        RECT 1395.930 3380.490 1397.110 3381.670 ;
        RECT 1395.930 3202.090 1397.110 3203.270 ;
        RECT 1395.930 3200.490 1397.110 3201.670 ;
        RECT 1395.930 3022.090 1397.110 3023.270 ;
        RECT 1395.930 3020.490 1397.110 3021.670 ;
        RECT 1395.930 2842.090 1397.110 2843.270 ;
        RECT 1395.930 2840.490 1397.110 2841.670 ;
        RECT 1395.930 2662.090 1397.110 2663.270 ;
        RECT 1395.930 2660.490 1397.110 2661.670 ;
        RECT 1395.930 2482.090 1397.110 2483.270 ;
        RECT 1395.930 2480.490 1397.110 2481.670 ;
        RECT 1395.930 2302.090 1397.110 2303.270 ;
        RECT 1395.930 2300.490 1397.110 2301.670 ;
        RECT 1395.930 2122.090 1397.110 2123.270 ;
        RECT 1395.930 2120.490 1397.110 2121.670 ;
        RECT 1395.930 1942.090 1397.110 1943.270 ;
        RECT 1395.930 1940.490 1397.110 1941.670 ;
        RECT 1395.930 1762.090 1397.110 1763.270 ;
        RECT 1395.930 1760.490 1397.110 1761.670 ;
        RECT 1395.930 1582.090 1397.110 1583.270 ;
        RECT 1395.930 1580.490 1397.110 1581.670 ;
        RECT 1395.930 1402.090 1397.110 1403.270 ;
        RECT 1395.930 1400.490 1397.110 1401.670 ;
        RECT 1395.930 1222.090 1397.110 1223.270 ;
        RECT 1395.930 1220.490 1397.110 1221.670 ;
        RECT 1395.930 1042.090 1397.110 1043.270 ;
        RECT 1395.930 1040.490 1397.110 1041.670 ;
        RECT 1395.930 862.090 1397.110 863.270 ;
        RECT 1395.930 860.490 1397.110 861.670 ;
        RECT 1395.930 682.090 1397.110 683.270 ;
        RECT 1395.930 680.490 1397.110 681.670 ;
        RECT 1395.930 502.090 1397.110 503.270 ;
        RECT 1395.930 500.490 1397.110 501.670 ;
        RECT 1395.930 322.090 1397.110 323.270 ;
        RECT 1395.930 320.490 1397.110 321.670 ;
        RECT 1395.930 142.090 1397.110 143.270 ;
        RECT 1395.930 140.490 1397.110 141.670 ;
        RECT 1395.930 -26.410 1397.110 -25.230 ;
        RECT 1395.930 -28.010 1397.110 -26.830 ;
        RECT 1575.930 3546.510 1577.110 3547.690 ;
        RECT 1575.930 3544.910 1577.110 3546.090 ;
        RECT 1575.930 3382.090 1577.110 3383.270 ;
        RECT 1575.930 3380.490 1577.110 3381.670 ;
        RECT 1575.930 3202.090 1577.110 3203.270 ;
        RECT 1575.930 3200.490 1577.110 3201.670 ;
        RECT 1575.930 3022.090 1577.110 3023.270 ;
        RECT 1575.930 3020.490 1577.110 3021.670 ;
        RECT 1575.930 2842.090 1577.110 2843.270 ;
        RECT 1575.930 2840.490 1577.110 2841.670 ;
        RECT 1575.930 2662.090 1577.110 2663.270 ;
        RECT 1575.930 2660.490 1577.110 2661.670 ;
        RECT 1575.930 2482.090 1577.110 2483.270 ;
        RECT 1575.930 2480.490 1577.110 2481.670 ;
        RECT 1575.930 2302.090 1577.110 2303.270 ;
        RECT 1575.930 2300.490 1577.110 2301.670 ;
        RECT 1575.930 2122.090 1577.110 2123.270 ;
        RECT 1575.930 2120.490 1577.110 2121.670 ;
        RECT 1575.930 1942.090 1577.110 1943.270 ;
        RECT 1575.930 1940.490 1577.110 1941.670 ;
        RECT 1575.930 1762.090 1577.110 1763.270 ;
        RECT 1575.930 1760.490 1577.110 1761.670 ;
        RECT 1575.930 1582.090 1577.110 1583.270 ;
        RECT 1575.930 1580.490 1577.110 1581.670 ;
        RECT 1575.930 1402.090 1577.110 1403.270 ;
        RECT 1575.930 1400.490 1577.110 1401.670 ;
        RECT 1575.930 1222.090 1577.110 1223.270 ;
        RECT 1575.930 1220.490 1577.110 1221.670 ;
        RECT 1575.930 1042.090 1577.110 1043.270 ;
        RECT 1575.930 1040.490 1577.110 1041.670 ;
        RECT 1575.930 862.090 1577.110 863.270 ;
        RECT 1575.930 860.490 1577.110 861.670 ;
        RECT 1575.930 682.090 1577.110 683.270 ;
        RECT 1575.930 680.490 1577.110 681.670 ;
        RECT 1575.930 502.090 1577.110 503.270 ;
        RECT 1575.930 500.490 1577.110 501.670 ;
        RECT 1575.930 322.090 1577.110 323.270 ;
        RECT 1575.930 320.490 1577.110 321.670 ;
        RECT 1575.930 142.090 1577.110 143.270 ;
        RECT 1575.930 140.490 1577.110 141.670 ;
        RECT 1575.930 -26.410 1577.110 -25.230 ;
        RECT 1575.930 -28.010 1577.110 -26.830 ;
        RECT 1755.930 3546.510 1757.110 3547.690 ;
        RECT 1755.930 3544.910 1757.110 3546.090 ;
        RECT 1755.930 3382.090 1757.110 3383.270 ;
        RECT 1755.930 3380.490 1757.110 3381.670 ;
        RECT 1755.930 3202.090 1757.110 3203.270 ;
        RECT 1755.930 3200.490 1757.110 3201.670 ;
        RECT 1755.930 3022.090 1757.110 3023.270 ;
        RECT 1755.930 3020.490 1757.110 3021.670 ;
        RECT 1755.930 2842.090 1757.110 2843.270 ;
        RECT 1755.930 2840.490 1757.110 2841.670 ;
        RECT 1755.930 2662.090 1757.110 2663.270 ;
        RECT 1755.930 2660.490 1757.110 2661.670 ;
        RECT 1755.930 2482.090 1757.110 2483.270 ;
        RECT 1755.930 2480.490 1757.110 2481.670 ;
        RECT 1755.930 2302.090 1757.110 2303.270 ;
        RECT 1755.930 2300.490 1757.110 2301.670 ;
        RECT 1755.930 2122.090 1757.110 2123.270 ;
        RECT 1755.930 2120.490 1757.110 2121.670 ;
        RECT 1755.930 1942.090 1757.110 1943.270 ;
        RECT 1755.930 1940.490 1757.110 1941.670 ;
        RECT 1755.930 1762.090 1757.110 1763.270 ;
        RECT 1755.930 1760.490 1757.110 1761.670 ;
        RECT 1755.930 1582.090 1757.110 1583.270 ;
        RECT 1755.930 1580.490 1757.110 1581.670 ;
        RECT 1755.930 1402.090 1757.110 1403.270 ;
        RECT 1755.930 1400.490 1757.110 1401.670 ;
        RECT 1755.930 1222.090 1757.110 1223.270 ;
        RECT 1755.930 1220.490 1757.110 1221.670 ;
        RECT 1755.930 1042.090 1757.110 1043.270 ;
        RECT 1755.930 1040.490 1757.110 1041.670 ;
        RECT 1755.930 862.090 1757.110 863.270 ;
        RECT 1755.930 860.490 1757.110 861.670 ;
        RECT 1755.930 682.090 1757.110 683.270 ;
        RECT 1755.930 680.490 1757.110 681.670 ;
        RECT 1755.930 502.090 1757.110 503.270 ;
        RECT 1755.930 500.490 1757.110 501.670 ;
        RECT 1755.930 322.090 1757.110 323.270 ;
        RECT 1755.930 320.490 1757.110 321.670 ;
        RECT 1755.930 142.090 1757.110 143.270 ;
        RECT 1755.930 140.490 1757.110 141.670 ;
        RECT 1755.930 -26.410 1757.110 -25.230 ;
        RECT 1755.930 -28.010 1757.110 -26.830 ;
        RECT 1935.930 3546.510 1937.110 3547.690 ;
        RECT 1935.930 3544.910 1937.110 3546.090 ;
        RECT 1935.930 3382.090 1937.110 3383.270 ;
        RECT 1935.930 3380.490 1937.110 3381.670 ;
        RECT 1935.930 3202.090 1937.110 3203.270 ;
        RECT 1935.930 3200.490 1937.110 3201.670 ;
        RECT 1935.930 3022.090 1937.110 3023.270 ;
        RECT 1935.930 3020.490 1937.110 3021.670 ;
        RECT 1935.930 2842.090 1937.110 2843.270 ;
        RECT 1935.930 2840.490 1937.110 2841.670 ;
        RECT 1935.930 2662.090 1937.110 2663.270 ;
        RECT 1935.930 2660.490 1937.110 2661.670 ;
        RECT 1935.930 2482.090 1937.110 2483.270 ;
        RECT 1935.930 2480.490 1937.110 2481.670 ;
        RECT 1935.930 2302.090 1937.110 2303.270 ;
        RECT 1935.930 2300.490 1937.110 2301.670 ;
        RECT 1935.930 2122.090 1937.110 2123.270 ;
        RECT 1935.930 2120.490 1937.110 2121.670 ;
        RECT 1935.930 1942.090 1937.110 1943.270 ;
        RECT 1935.930 1940.490 1937.110 1941.670 ;
        RECT 1935.930 1762.090 1937.110 1763.270 ;
        RECT 1935.930 1760.490 1937.110 1761.670 ;
        RECT 1935.930 1582.090 1937.110 1583.270 ;
        RECT 1935.930 1580.490 1937.110 1581.670 ;
        RECT 1935.930 1402.090 1937.110 1403.270 ;
        RECT 1935.930 1400.490 1937.110 1401.670 ;
        RECT 1935.930 1222.090 1937.110 1223.270 ;
        RECT 1935.930 1220.490 1937.110 1221.670 ;
        RECT 1935.930 1042.090 1937.110 1043.270 ;
        RECT 1935.930 1040.490 1937.110 1041.670 ;
        RECT 1935.930 862.090 1937.110 863.270 ;
        RECT 1935.930 860.490 1937.110 861.670 ;
        RECT 1935.930 682.090 1937.110 683.270 ;
        RECT 1935.930 680.490 1937.110 681.670 ;
        RECT 1935.930 502.090 1937.110 503.270 ;
        RECT 1935.930 500.490 1937.110 501.670 ;
        RECT 1935.930 322.090 1937.110 323.270 ;
        RECT 1935.930 320.490 1937.110 321.670 ;
        RECT 1935.930 142.090 1937.110 143.270 ;
        RECT 1935.930 140.490 1937.110 141.670 ;
        RECT 1935.930 -26.410 1937.110 -25.230 ;
        RECT 1935.930 -28.010 1937.110 -26.830 ;
        RECT 2115.930 3546.510 2117.110 3547.690 ;
        RECT 2115.930 3544.910 2117.110 3546.090 ;
        RECT 2115.930 3382.090 2117.110 3383.270 ;
        RECT 2115.930 3380.490 2117.110 3381.670 ;
        RECT 2115.930 3202.090 2117.110 3203.270 ;
        RECT 2115.930 3200.490 2117.110 3201.670 ;
        RECT 2115.930 3022.090 2117.110 3023.270 ;
        RECT 2115.930 3020.490 2117.110 3021.670 ;
        RECT 2115.930 2842.090 2117.110 2843.270 ;
        RECT 2115.930 2840.490 2117.110 2841.670 ;
        RECT 2115.930 2662.090 2117.110 2663.270 ;
        RECT 2115.930 2660.490 2117.110 2661.670 ;
        RECT 2115.930 2482.090 2117.110 2483.270 ;
        RECT 2115.930 2480.490 2117.110 2481.670 ;
        RECT 2115.930 2302.090 2117.110 2303.270 ;
        RECT 2115.930 2300.490 2117.110 2301.670 ;
        RECT 2115.930 2122.090 2117.110 2123.270 ;
        RECT 2115.930 2120.490 2117.110 2121.670 ;
        RECT 2115.930 1942.090 2117.110 1943.270 ;
        RECT 2115.930 1940.490 2117.110 1941.670 ;
        RECT 2115.930 1762.090 2117.110 1763.270 ;
        RECT 2115.930 1760.490 2117.110 1761.670 ;
        RECT 2115.930 1582.090 2117.110 1583.270 ;
        RECT 2115.930 1580.490 2117.110 1581.670 ;
        RECT 2115.930 1402.090 2117.110 1403.270 ;
        RECT 2115.930 1400.490 2117.110 1401.670 ;
        RECT 2115.930 1222.090 2117.110 1223.270 ;
        RECT 2115.930 1220.490 2117.110 1221.670 ;
        RECT 2115.930 1042.090 2117.110 1043.270 ;
        RECT 2115.930 1040.490 2117.110 1041.670 ;
        RECT 2115.930 862.090 2117.110 863.270 ;
        RECT 2115.930 860.490 2117.110 861.670 ;
        RECT 2115.930 682.090 2117.110 683.270 ;
        RECT 2115.930 680.490 2117.110 681.670 ;
        RECT 2115.930 502.090 2117.110 503.270 ;
        RECT 2115.930 500.490 2117.110 501.670 ;
        RECT 2115.930 322.090 2117.110 323.270 ;
        RECT 2115.930 320.490 2117.110 321.670 ;
        RECT 2115.930 142.090 2117.110 143.270 ;
        RECT 2115.930 140.490 2117.110 141.670 ;
        RECT 2115.930 -26.410 2117.110 -25.230 ;
        RECT 2115.930 -28.010 2117.110 -26.830 ;
        RECT 2295.930 3546.510 2297.110 3547.690 ;
        RECT 2295.930 3544.910 2297.110 3546.090 ;
        RECT 2295.930 3382.090 2297.110 3383.270 ;
        RECT 2295.930 3380.490 2297.110 3381.670 ;
        RECT 2295.930 3202.090 2297.110 3203.270 ;
        RECT 2295.930 3200.490 2297.110 3201.670 ;
        RECT 2295.930 3022.090 2297.110 3023.270 ;
        RECT 2295.930 3020.490 2297.110 3021.670 ;
        RECT 2295.930 2842.090 2297.110 2843.270 ;
        RECT 2295.930 2840.490 2297.110 2841.670 ;
        RECT 2295.930 2662.090 2297.110 2663.270 ;
        RECT 2295.930 2660.490 2297.110 2661.670 ;
        RECT 2295.930 2482.090 2297.110 2483.270 ;
        RECT 2295.930 2480.490 2297.110 2481.670 ;
        RECT 2295.930 2302.090 2297.110 2303.270 ;
        RECT 2295.930 2300.490 2297.110 2301.670 ;
        RECT 2295.930 2122.090 2297.110 2123.270 ;
        RECT 2295.930 2120.490 2297.110 2121.670 ;
        RECT 2295.930 1942.090 2297.110 1943.270 ;
        RECT 2295.930 1940.490 2297.110 1941.670 ;
        RECT 2295.930 1762.090 2297.110 1763.270 ;
        RECT 2295.930 1760.490 2297.110 1761.670 ;
        RECT 2295.930 1582.090 2297.110 1583.270 ;
        RECT 2295.930 1580.490 2297.110 1581.670 ;
        RECT 2295.930 1402.090 2297.110 1403.270 ;
        RECT 2295.930 1400.490 2297.110 1401.670 ;
        RECT 2295.930 1222.090 2297.110 1223.270 ;
        RECT 2295.930 1220.490 2297.110 1221.670 ;
        RECT 2295.930 1042.090 2297.110 1043.270 ;
        RECT 2295.930 1040.490 2297.110 1041.670 ;
        RECT 2295.930 862.090 2297.110 863.270 ;
        RECT 2295.930 860.490 2297.110 861.670 ;
        RECT 2295.930 682.090 2297.110 683.270 ;
        RECT 2295.930 680.490 2297.110 681.670 ;
        RECT 2295.930 502.090 2297.110 503.270 ;
        RECT 2295.930 500.490 2297.110 501.670 ;
        RECT 2295.930 322.090 2297.110 323.270 ;
        RECT 2295.930 320.490 2297.110 321.670 ;
        RECT 2295.930 142.090 2297.110 143.270 ;
        RECT 2295.930 140.490 2297.110 141.670 ;
        RECT 2295.930 -26.410 2297.110 -25.230 ;
        RECT 2295.930 -28.010 2297.110 -26.830 ;
        RECT 2475.930 3546.510 2477.110 3547.690 ;
        RECT 2475.930 3544.910 2477.110 3546.090 ;
        RECT 2475.930 3382.090 2477.110 3383.270 ;
        RECT 2475.930 3380.490 2477.110 3381.670 ;
        RECT 2475.930 3202.090 2477.110 3203.270 ;
        RECT 2475.930 3200.490 2477.110 3201.670 ;
        RECT 2475.930 3022.090 2477.110 3023.270 ;
        RECT 2475.930 3020.490 2477.110 3021.670 ;
        RECT 2475.930 2842.090 2477.110 2843.270 ;
        RECT 2475.930 2840.490 2477.110 2841.670 ;
        RECT 2475.930 2662.090 2477.110 2663.270 ;
        RECT 2475.930 2660.490 2477.110 2661.670 ;
        RECT 2475.930 2482.090 2477.110 2483.270 ;
        RECT 2475.930 2480.490 2477.110 2481.670 ;
        RECT 2475.930 2302.090 2477.110 2303.270 ;
        RECT 2475.930 2300.490 2477.110 2301.670 ;
        RECT 2475.930 2122.090 2477.110 2123.270 ;
        RECT 2475.930 2120.490 2477.110 2121.670 ;
        RECT 2475.930 1942.090 2477.110 1943.270 ;
        RECT 2475.930 1940.490 2477.110 1941.670 ;
        RECT 2475.930 1762.090 2477.110 1763.270 ;
        RECT 2475.930 1760.490 2477.110 1761.670 ;
        RECT 2475.930 1582.090 2477.110 1583.270 ;
        RECT 2475.930 1580.490 2477.110 1581.670 ;
        RECT 2475.930 1402.090 2477.110 1403.270 ;
        RECT 2475.930 1400.490 2477.110 1401.670 ;
        RECT 2475.930 1222.090 2477.110 1223.270 ;
        RECT 2475.930 1220.490 2477.110 1221.670 ;
        RECT 2475.930 1042.090 2477.110 1043.270 ;
        RECT 2475.930 1040.490 2477.110 1041.670 ;
        RECT 2475.930 862.090 2477.110 863.270 ;
        RECT 2475.930 860.490 2477.110 861.670 ;
        RECT 2475.930 682.090 2477.110 683.270 ;
        RECT 2475.930 680.490 2477.110 681.670 ;
        RECT 2475.930 502.090 2477.110 503.270 ;
        RECT 2475.930 500.490 2477.110 501.670 ;
        RECT 2475.930 322.090 2477.110 323.270 ;
        RECT 2475.930 320.490 2477.110 321.670 ;
        RECT 2475.930 142.090 2477.110 143.270 ;
        RECT 2475.930 140.490 2477.110 141.670 ;
        RECT 2475.930 -26.410 2477.110 -25.230 ;
        RECT 2475.930 -28.010 2477.110 -26.830 ;
        RECT 2655.930 3546.510 2657.110 3547.690 ;
        RECT 2655.930 3544.910 2657.110 3546.090 ;
        RECT 2655.930 3382.090 2657.110 3383.270 ;
        RECT 2655.930 3380.490 2657.110 3381.670 ;
        RECT 2655.930 3202.090 2657.110 3203.270 ;
        RECT 2655.930 3200.490 2657.110 3201.670 ;
        RECT 2655.930 3022.090 2657.110 3023.270 ;
        RECT 2655.930 3020.490 2657.110 3021.670 ;
        RECT 2655.930 2842.090 2657.110 2843.270 ;
        RECT 2655.930 2840.490 2657.110 2841.670 ;
        RECT 2655.930 2662.090 2657.110 2663.270 ;
        RECT 2655.930 2660.490 2657.110 2661.670 ;
        RECT 2655.930 2482.090 2657.110 2483.270 ;
        RECT 2655.930 2480.490 2657.110 2481.670 ;
        RECT 2655.930 2302.090 2657.110 2303.270 ;
        RECT 2655.930 2300.490 2657.110 2301.670 ;
        RECT 2655.930 2122.090 2657.110 2123.270 ;
        RECT 2655.930 2120.490 2657.110 2121.670 ;
        RECT 2655.930 1942.090 2657.110 1943.270 ;
        RECT 2655.930 1940.490 2657.110 1941.670 ;
        RECT 2655.930 1762.090 2657.110 1763.270 ;
        RECT 2655.930 1760.490 2657.110 1761.670 ;
        RECT 2655.930 1582.090 2657.110 1583.270 ;
        RECT 2655.930 1580.490 2657.110 1581.670 ;
        RECT 2655.930 1402.090 2657.110 1403.270 ;
        RECT 2655.930 1400.490 2657.110 1401.670 ;
        RECT 2655.930 1222.090 2657.110 1223.270 ;
        RECT 2655.930 1220.490 2657.110 1221.670 ;
        RECT 2655.930 1042.090 2657.110 1043.270 ;
        RECT 2655.930 1040.490 2657.110 1041.670 ;
        RECT 2655.930 862.090 2657.110 863.270 ;
        RECT 2655.930 860.490 2657.110 861.670 ;
        RECT 2655.930 682.090 2657.110 683.270 ;
        RECT 2655.930 680.490 2657.110 681.670 ;
        RECT 2655.930 502.090 2657.110 503.270 ;
        RECT 2655.930 500.490 2657.110 501.670 ;
        RECT 2655.930 322.090 2657.110 323.270 ;
        RECT 2655.930 320.490 2657.110 321.670 ;
        RECT 2655.930 142.090 2657.110 143.270 ;
        RECT 2655.930 140.490 2657.110 141.670 ;
        RECT 2655.930 -26.410 2657.110 -25.230 ;
        RECT 2655.930 -28.010 2657.110 -26.830 ;
        RECT 2835.930 3546.510 2837.110 3547.690 ;
        RECT 2835.930 3544.910 2837.110 3546.090 ;
        RECT 2835.930 3382.090 2837.110 3383.270 ;
        RECT 2835.930 3380.490 2837.110 3381.670 ;
        RECT 2835.930 3202.090 2837.110 3203.270 ;
        RECT 2835.930 3200.490 2837.110 3201.670 ;
        RECT 2835.930 3022.090 2837.110 3023.270 ;
        RECT 2835.930 3020.490 2837.110 3021.670 ;
        RECT 2835.930 2842.090 2837.110 2843.270 ;
        RECT 2835.930 2840.490 2837.110 2841.670 ;
        RECT 2835.930 2662.090 2837.110 2663.270 ;
        RECT 2835.930 2660.490 2837.110 2661.670 ;
        RECT 2835.930 2482.090 2837.110 2483.270 ;
        RECT 2835.930 2480.490 2837.110 2481.670 ;
        RECT 2835.930 2302.090 2837.110 2303.270 ;
        RECT 2835.930 2300.490 2837.110 2301.670 ;
        RECT 2835.930 2122.090 2837.110 2123.270 ;
        RECT 2835.930 2120.490 2837.110 2121.670 ;
        RECT 2835.930 1942.090 2837.110 1943.270 ;
        RECT 2835.930 1940.490 2837.110 1941.670 ;
        RECT 2835.930 1762.090 2837.110 1763.270 ;
        RECT 2835.930 1760.490 2837.110 1761.670 ;
        RECT 2835.930 1582.090 2837.110 1583.270 ;
        RECT 2835.930 1580.490 2837.110 1581.670 ;
        RECT 2835.930 1402.090 2837.110 1403.270 ;
        RECT 2835.930 1400.490 2837.110 1401.670 ;
        RECT 2835.930 1222.090 2837.110 1223.270 ;
        RECT 2835.930 1220.490 2837.110 1221.670 ;
        RECT 2835.930 1042.090 2837.110 1043.270 ;
        RECT 2835.930 1040.490 2837.110 1041.670 ;
        RECT 2835.930 862.090 2837.110 863.270 ;
        RECT 2835.930 860.490 2837.110 861.670 ;
        RECT 2835.930 682.090 2837.110 683.270 ;
        RECT 2835.930 680.490 2837.110 681.670 ;
        RECT 2835.930 502.090 2837.110 503.270 ;
        RECT 2835.930 500.490 2837.110 501.670 ;
        RECT 2835.930 322.090 2837.110 323.270 ;
        RECT 2835.930 320.490 2837.110 321.670 ;
        RECT 2835.930 142.090 2837.110 143.270 ;
        RECT 2835.930 140.490 2837.110 141.670 ;
        RECT 2835.930 -26.410 2837.110 -25.230 ;
        RECT 2835.930 -28.010 2837.110 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 3382.090 2952.190 3383.270 ;
        RECT 2951.010 3380.490 2952.190 3381.670 ;
        RECT 2951.010 3202.090 2952.190 3203.270 ;
        RECT 2951.010 3200.490 2952.190 3201.670 ;
        RECT 2951.010 3022.090 2952.190 3023.270 ;
        RECT 2951.010 3020.490 2952.190 3021.670 ;
        RECT 2951.010 2842.090 2952.190 2843.270 ;
        RECT 2951.010 2840.490 2952.190 2841.670 ;
        RECT 2951.010 2662.090 2952.190 2663.270 ;
        RECT 2951.010 2660.490 2952.190 2661.670 ;
        RECT 2951.010 2482.090 2952.190 2483.270 ;
        RECT 2951.010 2480.490 2952.190 2481.670 ;
        RECT 2951.010 2302.090 2952.190 2303.270 ;
        RECT 2951.010 2300.490 2952.190 2301.670 ;
        RECT 2951.010 2122.090 2952.190 2123.270 ;
        RECT 2951.010 2120.490 2952.190 2121.670 ;
        RECT 2951.010 1942.090 2952.190 1943.270 ;
        RECT 2951.010 1940.490 2952.190 1941.670 ;
        RECT 2951.010 1762.090 2952.190 1763.270 ;
        RECT 2951.010 1760.490 2952.190 1761.670 ;
        RECT 2951.010 1582.090 2952.190 1583.270 ;
        RECT 2951.010 1580.490 2952.190 1581.670 ;
        RECT 2951.010 1402.090 2952.190 1403.270 ;
        RECT 2951.010 1400.490 2952.190 1401.670 ;
        RECT 2951.010 1222.090 2952.190 1223.270 ;
        RECT 2951.010 1220.490 2952.190 1221.670 ;
        RECT 2951.010 1042.090 2952.190 1043.270 ;
        RECT 2951.010 1040.490 2952.190 1041.670 ;
        RECT 2951.010 862.090 2952.190 863.270 ;
        RECT 2951.010 860.490 2952.190 861.670 ;
        RECT 2951.010 682.090 2952.190 683.270 ;
        RECT 2951.010 680.490 2952.190 681.670 ;
        RECT 2951.010 502.090 2952.190 503.270 ;
        RECT 2951.010 500.490 2952.190 501.670 ;
        RECT 2951.010 322.090 2952.190 323.270 ;
        RECT 2951.010 320.490 2952.190 321.670 ;
        RECT 2951.010 142.090 2952.190 143.270 ;
        RECT 2951.010 140.490 2952.190 141.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 135.020 3547.800 138.020 3547.810 ;
        RECT 315.020 3547.800 318.020 3547.810 ;
        RECT 495.020 3547.800 498.020 3547.810 ;
        RECT 675.020 3547.800 678.020 3547.810 ;
        RECT 855.020 3547.800 858.020 3547.810 ;
        RECT 1035.020 3547.800 1038.020 3547.810 ;
        RECT 1215.020 3547.800 1218.020 3547.810 ;
        RECT 1395.020 3547.800 1398.020 3547.810 ;
        RECT 1575.020 3547.800 1578.020 3547.810 ;
        RECT 1755.020 3547.800 1758.020 3547.810 ;
        RECT 1935.020 3547.800 1938.020 3547.810 ;
        RECT 2115.020 3547.800 2118.020 3547.810 ;
        RECT 2295.020 3547.800 2298.020 3547.810 ;
        RECT 2475.020 3547.800 2478.020 3547.810 ;
        RECT 2655.020 3547.800 2658.020 3547.810 ;
        RECT 2835.020 3547.800 2838.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 135.020 3544.790 138.020 3544.800 ;
        RECT 315.020 3544.790 318.020 3544.800 ;
        RECT 495.020 3544.790 498.020 3544.800 ;
        RECT 675.020 3544.790 678.020 3544.800 ;
        RECT 855.020 3544.790 858.020 3544.800 ;
        RECT 1035.020 3544.790 1038.020 3544.800 ;
        RECT 1215.020 3544.790 1218.020 3544.800 ;
        RECT 1395.020 3544.790 1398.020 3544.800 ;
        RECT 1575.020 3544.790 1578.020 3544.800 ;
        RECT 1755.020 3544.790 1758.020 3544.800 ;
        RECT 1935.020 3544.790 1938.020 3544.800 ;
        RECT 2115.020 3544.790 2118.020 3544.800 ;
        RECT 2295.020 3544.790 2298.020 3544.800 ;
        RECT 2475.020 3544.790 2478.020 3544.800 ;
        RECT 2655.020 3544.790 2658.020 3544.800 ;
        RECT 2835.020 3544.790 2838.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3383.380 -30.480 3383.390 ;
        RECT 135.020 3383.380 138.020 3383.390 ;
        RECT 315.020 3383.380 318.020 3383.390 ;
        RECT 495.020 3383.380 498.020 3383.390 ;
        RECT 675.020 3383.380 678.020 3383.390 ;
        RECT 855.020 3383.380 858.020 3383.390 ;
        RECT 1035.020 3383.380 1038.020 3383.390 ;
        RECT 1215.020 3383.380 1218.020 3383.390 ;
        RECT 1395.020 3383.380 1398.020 3383.390 ;
        RECT 1575.020 3383.380 1578.020 3383.390 ;
        RECT 1755.020 3383.380 1758.020 3383.390 ;
        RECT 1935.020 3383.380 1938.020 3383.390 ;
        RECT 2115.020 3383.380 2118.020 3383.390 ;
        RECT 2295.020 3383.380 2298.020 3383.390 ;
        RECT 2475.020 3383.380 2478.020 3383.390 ;
        RECT 2655.020 3383.380 2658.020 3383.390 ;
        RECT 2835.020 3383.380 2838.020 3383.390 ;
        RECT 2950.100 3383.380 2953.100 3383.390 ;
        RECT -33.480 3380.380 2953.100 3383.380 ;
        RECT -33.480 3380.370 -30.480 3380.380 ;
        RECT 135.020 3380.370 138.020 3380.380 ;
        RECT 315.020 3380.370 318.020 3380.380 ;
        RECT 495.020 3380.370 498.020 3380.380 ;
        RECT 675.020 3380.370 678.020 3380.380 ;
        RECT 855.020 3380.370 858.020 3380.380 ;
        RECT 1035.020 3380.370 1038.020 3380.380 ;
        RECT 1215.020 3380.370 1218.020 3380.380 ;
        RECT 1395.020 3380.370 1398.020 3380.380 ;
        RECT 1575.020 3380.370 1578.020 3380.380 ;
        RECT 1755.020 3380.370 1758.020 3380.380 ;
        RECT 1935.020 3380.370 1938.020 3380.380 ;
        RECT 2115.020 3380.370 2118.020 3380.380 ;
        RECT 2295.020 3380.370 2298.020 3380.380 ;
        RECT 2475.020 3380.370 2478.020 3380.380 ;
        RECT 2655.020 3380.370 2658.020 3380.380 ;
        RECT 2835.020 3380.370 2838.020 3380.380 ;
        RECT 2950.100 3380.370 2953.100 3380.380 ;
        RECT -33.480 3203.380 -30.480 3203.390 ;
        RECT 135.020 3203.380 138.020 3203.390 ;
        RECT 315.020 3203.380 318.020 3203.390 ;
        RECT 495.020 3203.380 498.020 3203.390 ;
        RECT 675.020 3203.380 678.020 3203.390 ;
        RECT 855.020 3203.380 858.020 3203.390 ;
        RECT 1035.020 3203.380 1038.020 3203.390 ;
        RECT 1215.020 3203.380 1218.020 3203.390 ;
        RECT 1395.020 3203.380 1398.020 3203.390 ;
        RECT 1575.020 3203.380 1578.020 3203.390 ;
        RECT 1755.020 3203.380 1758.020 3203.390 ;
        RECT 1935.020 3203.380 1938.020 3203.390 ;
        RECT 2115.020 3203.380 2118.020 3203.390 ;
        RECT 2295.020 3203.380 2298.020 3203.390 ;
        RECT 2475.020 3203.380 2478.020 3203.390 ;
        RECT 2655.020 3203.380 2658.020 3203.390 ;
        RECT 2835.020 3203.380 2838.020 3203.390 ;
        RECT 2950.100 3203.380 2953.100 3203.390 ;
        RECT -33.480 3200.380 2953.100 3203.380 ;
        RECT -33.480 3200.370 -30.480 3200.380 ;
        RECT 135.020 3200.370 138.020 3200.380 ;
        RECT 315.020 3200.370 318.020 3200.380 ;
        RECT 495.020 3200.370 498.020 3200.380 ;
        RECT 675.020 3200.370 678.020 3200.380 ;
        RECT 855.020 3200.370 858.020 3200.380 ;
        RECT 1035.020 3200.370 1038.020 3200.380 ;
        RECT 1215.020 3200.370 1218.020 3200.380 ;
        RECT 1395.020 3200.370 1398.020 3200.380 ;
        RECT 1575.020 3200.370 1578.020 3200.380 ;
        RECT 1755.020 3200.370 1758.020 3200.380 ;
        RECT 1935.020 3200.370 1938.020 3200.380 ;
        RECT 2115.020 3200.370 2118.020 3200.380 ;
        RECT 2295.020 3200.370 2298.020 3200.380 ;
        RECT 2475.020 3200.370 2478.020 3200.380 ;
        RECT 2655.020 3200.370 2658.020 3200.380 ;
        RECT 2835.020 3200.370 2838.020 3200.380 ;
        RECT 2950.100 3200.370 2953.100 3200.380 ;
        RECT -33.480 3023.380 -30.480 3023.390 ;
        RECT 135.020 3023.380 138.020 3023.390 ;
        RECT 315.020 3023.380 318.020 3023.390 ;
        RECT 495.020 3023.380 498.020 3023.390 ;
        RECT 675.020 3023.380 678.020 3023.390 ;
        RECT 855.020 3023.380 858.020 3023.390 ;
        RECT 1035.020 3023.380 1038.020 3023.390 ;
        RECT 1215.020 3023.380 1218.020 3023.390 ;
        RECT 1395.020 3023.380 1398.020 3023.390 ;
        RECT 1575.020 3023.380 1578.020 3023.390 ;
        RECT 1755.020 3023.380 1758.020 3023.390 ;
        RECT 1935.020 3023.380 1938.020 3023.390 ;
        RECT 2115.020 3023.380 2118.020 3023.390 ;
        RECT 2295.020 3023.380 2298.020 3023.390 ;
        RECT 2475.020 3023.380 2478.020 3023.390 ;
        RECT 2655.020 3023.380 2658.020 3023.390 ;
        RECT 2835.020 3023.380 2838.020 3023.390 ;
        RECT 2950.100 3023.380 2953.100 3023.390 ;
        RECT -33.480 3020.380 2953.100 3023.380 ;
        RECT -33.480 3020.370 -30.480 3020.380 ;
        RECT 135.020 3020.370 138.020 3020.380 ;
        RECT 315.020 3020.370 318.020 3020.380 ;
        RECT 495.020 3020.370 498.020 3020.380 ;
        RECT 675.020 3020.370 678.020 3020.380 ;
        RECT 855.020 3020.370 858.020 3020.380 ;
        RECT 1035.020 3020.370 1038.020 3020.380 ;
        RECT 1215.020 3020.370 1218.020 3020.380 ;
        RECT 1395.020 3020.370 1398.020 3020.380 ;
        RECT 1575.020 3020.370 1578.020 3020.380 ;
        RECT 1755.020 3020.370 1758.020 3020.380 ;
        RECT 1935.020 3020.370 1938.020 3020.380 ;
        RECT 2115.020 3020.370 2118.020 3020.380 ;
        RECT 2295.020 3020.370 2298.020 3020.380 ;
        RECT 2475.020 3020.370 2478.020 3020.380 ;
        RECT 2655.020 3020.370 2658.020 3020.380 ;
        RECT 2835.020 3020.370 2838.020 3020.380 ;
        RECT 2950.100 3020.370 2953.100 3020.380 ;
        RECT -33.480 2843.380 -30.480 2843.390 ;
        RECT 135.020 2843.380 138.020 2843.390 ;
        RECT 315.020 2843.380 318.020 2843.390 ;
        RECT 495.020 2843.380 498.020 2843.390 ;
        RECT 675.020 2843.380 678.020 2843.390 ;
        RECT 855.020 2843.380 858.020 2843.390 ;
        RECT 1035.020 2843.380 1038.020 2843.390 ;
        RECT 1215.020 2843.380 1218.020 2843.390 ;
        RECT 1395.020 2843.380 1398.020 2843.390 ;
        RECT 1575.020 2843.380 1578.020 2843.390 ;
        RECT 1755.020 2843.380 1758.020 2843.390 ;
        RECT 1935.020 2843.380 1938.020 2843.390 ;
        RECT 2115.020 2843.380 2118.020 2843.390 ;
        RECT 2295.020 2843.380 2298.020 2843.390 ;
        RECT 2475.020 2843.380 2478.020 2843.390 ;
        RECT 2655.020 2843.380 2658.020 2843.390 ;
        RECT 2835.020 2843.380 2838.020 2843.390 ;
        RECT 2950.100 2843.380 2953.100 2843.390 ;
        RECT -33.480 2840.380 2953.100 2843.380 ;
        RECT -33.480 2840.370 -30.480 2840.380 ;
        RECT 135.020 2840.370 138.020 2840.380 ;
        RECT 315.020 2840.370 318.020 2840.380 ;
        RECT 495.020 2840.370 498.020 2840.380 ;
        RECT 675.020 2840.370 678.020 2840.380 ;
        RECT 855.020 2840.370 858.020 2840.380 ;
        RECT 1035.020 2840.370 1038.020 2840.380 ;
        RECT 1215.020 2840.370 1218.020 2840.380 ;
        RECT 1395.020 2840.370 1398.020 2840.380 ;
        RECT 1575.020 2840.370 1578.020 2840.380 ;
        RECT 1755.020 2840.370 1758.020 2840.380 ;
        RECT 1935.020 2840.370 1938.020 2840.380 ;
        RECT 2115.020 2840.370 2118.020 2840.380 ;
        RECT 2295.020 2840.370 2298.020 2840.380 ;
        RECT 2475.020 2840.370 2478.020 2840.380 ;
        RECT 2655.020 2840.370 2658.020 2840.380 ;
        RECT 2835.020 2840.370 2838.020 2840.380 ;
        RECT 2950.100 2840.370 2953.100 2840.380 ;
        RECT -33.480 2663.380 -30.480 2663.390 ;
        RECT 135.020 2663.380 138.020 2663.390 ;
        RECT 315.020 2663.380 318.020 2663.390 ;
        RECT 495.020 2663.380 498.020 2663.390 ;
        RECT 675.020 2663.380 678.020 2663.390 ;
        RECT 855.020 2663.380 858.020 2663.390 ;
        RECT 1035.020 2663.380 1038.020 2663.390 ;
        RECT 1215.020 2663.380 1218.020 2663.390 ;
        RECT 1395.020 2663.380 1398.020 2663.390 ;
        RECT 1575.020 2663.380 1578.020 2663.390 ;
        RECT 1755.020 2663.380 1758.020 2663.390 ;
        RECT 1935.020 2663.380 1938.020 2663.390 ;
        RECT 2115.020 2663.380 2118.020 2663.390 ;
        RECT 2295.020 2663.380 2298.020 2663.390 ;
        RECT 2475.020 2663.380 2478.020 2663.390 ;
        RECT 2655.020 2663.380 2658.020 2663.390 ;
        RECT 2835.020 2663.380 2838.020 2663.390 ;
        RECT 2950.100 2663.380 2953.100 2663.390 ;
        RECT -33.480 2660.380 2953.100 2663.380 ;
        RECT -33.480 2660.370 -30.480 2660.380 ;
        RECT 135.020 2660.370 138.020 2660.380 ;
        RECT 315.020 2660.370 318.020 2660.380 ;
        RECT 495.020 2660.370 498.020 2660.380 ;
        RECT 675.020 2660.370 678.020 2660.380 ;
        RECT 855.020 2660.370 858.020 2660.380 ;
        RECT 1035.020 2660.370 1038.020 2660.380 ;
        RECT 1215.020 2660.370 1218.020 2660.380 ;
        RECT 1395.020 2660.370 1398.020 2660.380 ;
        RECT 1575.020 2660.370 1578.020 2660.380 ;
        RECT 1755.020 2660.370 1758.020 2660.380 ;
        RECT 1935.020 2660.370 1938.020 2660.380 ;
        RECT 2115.020 2660.370 2118.020 2660.380 ;
        RECT 2295.020 2660.370 2298.020 2660.380 ;
        RECT 2475.020 2660.370 2478.020 2660.380 ;
        RECT 2655.020 2660.370 2658.020 2660.380 ;
        RECT 2835.020 2660.370 2838.020 2660.380 ;
        RECT 2950.100 2660.370 2953.100 2660.380 ;
        RECT -33.480 2483.380 -30.480 2483.390 ;
        RECT 135.020 2483.380 138.020 2483.390 ;
        RECT 315.020 2483.380 318.020 2483.390 ;
        RECT 495.020 2483.380 498.020 2483.390 ;
        RECT 675.020 2483.380 678.020 2483.390 ;
        RECT 855.020 2483.380 858.020 2483.390 ;
        RECT 1035.020 2483.380 1038.020 2483.390 ;
        RECT 1215.020 2483.380 1218.020 2483.390 ;
        RECT 1395.020 2483.380 1398.020 2483.390 ;
        RECT 1575.020 2483.380 1578.020 2483.390 ;
        RECT 1755.020 2483.380 1758.020 2483.390 ;
        RECT 1935.020 2483.380 1938.020 2483.390 ;
        RECT 2115.020 2483.380 2118.020 2483.390 ;
        RECT 2295.020 2483.380 2298.020 2483.390 ;
        RECT 2475.020 2483.380 2478.020 2483.390 ;
        RECT 2655.020 2483.380 2658.020 2483.390 ;
        RECT 2835.020 2483.380 2838.020 2483.390 ;
        RECT 2950.100 2483.380 2953.100 2483.390 ;
        RECT -33.480 2480.380 2953.100 2483.380 ;
        RECT -33.480 2480.370 -30.480 2480.380 ;
        RECT 135.020 2480.370 138.020 2480.380 ;
        RECT 315.020 2480.370 318.020 2480.380 ;
        RECT 495.020 2480.370 498.020 2480.380 ;
        RECT 675.020 2480.370 678.020 2480.380 ;
        RECT 855.020 2480.370 858.020 2480.380 ;
        RECT 1035.020 2480.370 1038.020 2480.380 ;
        RECT 1215.020 2480.370 1218.020 2480.380 ;
        RECT 1395.020 2480.370 1398.020 2480.380 ;
        RECT 1575.020 2480.370 1578.020 2480.380 ;
        RECT 1755.020 2480.370 1758.020 2480.380 ;
        RECT 1935.020 2480.370 1938.020 2480.380 ;
        RECT 2115.020 2480.370 2118.020 2480.380 ;
        RECT 2295.020 2480.370 2298.020 2480.380 ;
        RECT 2475.020 2480.370 2478.020 2480.380 ;
        RECT 2655.020 2480.370 2658.020 2480.380 ;
        RECT 2835.020 2480.370 2838.020 2480.380 ;
        RECT 2950.100 2480.370 2953.100 2480.380 ;
        RECT -33.480 2303.380 -30.480 2303.390 ;
        RECT 135.020 2303.380 138.020 2303.390 ;
        RECT 315.020 2303.380 318.020 2303.390 ;
        RECT 495.020 2303.380 498.020 2303.390 ;
        RECT 675.020 2303.380 678.020 2303.390 ;
        RECT 855.020 2303.380 858.020 2303.390 ;
        RECT 1035.020 2303.380 1038.020 2303.390 ;
        RECT 1215.020 2303.380 1218.020 2303.390 ;
        RECT 1395.020 2303.380 1398.020 2303.390 ;
        RECT 1575.020 2303.380 1578.020 2303.390 ;
        RECT 1755.020 2303.380 1758.020 2303.390 ;
        RECT 1935.020 2303.380 1938.020 2303.390 ;
        RECT 2115.020 2303.380 2118.020 2303.390 ;
        RECT 2295.020 2303.380 2298.020 2303.390 ;
        RECT 2475.020 2303.380 2478.020 2303.390 ;
        RECT 2655.020 2303.380 2658.020 2303.390 ;
        RECT 2835.020 2303.380 2838.020 2303.390 ;
        RECT 2950.100 2303.380 2953.100 2303.390 ;
        RECT -33.480 2300.380 2953.100 2303.380 ;
        RECT -33.480 2300.370 -30.480 2300.380 ;
        RECT 135.020 2300.370 138.020 2300.380 ;
        RECT 315.020 2300.370 318.020 2300.380 ;
        RECT 495.020 2300.370 498.020 2300.380 ;
        RECT 675.020 2300.370 678.020 2300.380 ;
        RECT 855.020 2300.370 858.020 2300.380 ;
        RECT 1035.020 2300.370 1038.020 2300.380 ;
        RECT 1215.020 2300.370 1218.020 2300.380 ;
        RECT 1395.020 2300.370 1398.020 2300.380 ;
        RECT 1575.020 2300.370 1578.020 2300.380 ;
        RECT 1755.020 2300.370 1758.020 2300.380 ;
        RECT 1935.020 2300.370 1938.020 2300.380 ;
        RECT 2115.020 2300.370 2118.020 2300.380 ;
        RECT 2295.020 2300.370 2298.020 2300.380 ;
        RECT 2475.020 2300.370 2478.020 2300.380 ;
        RECT 2655.020 2300.370 2658.020 2300.380 ;
        RECT 2835.020 2300.370 2838.020 2300.380 ;
        RECT 2950.100 2300.370 2953.100 2300.380 ;
        RECT -33.480 2123.380 -30.480 2123.390 ;
        RECT 135.020 2123.380 138.020 2123.390 ;
        RECT 315.020 2123.380 318.020 2123.390 ;
        RECT 495.020 2123.380 498.020 2123.390 ;
        RECT 675.020 2123.380 678.020 2123.390 ;
        RECT 855.020 2123.380 858.020 2123.390 ;
        RECT 1035.020 2123.380 1038.020 2123.390 ;
        RECT 1215.020 2123.380 1218.020 2123.390 ;
        RECT 1395.020 2123.380 1398.020 2123.390 ;
        RECT 1575.020 2123.380 1578.020 2123.390 ;
        RECT 1755.020 2123.380 1758.020 2123.390 ;
        RECT 1935.020 2123.380 1938.020 2123.390 ;
        RECT 2115.020 2123.380 2118.020 2123.390 ;
        RECT 2295.020 2123.380 2298.020 2123.390 ;
        RECT 2475.020 2123.380 2478.020 2123.390 ;
        RECT 2655.020 2123.380 2658.020 2123.390 ;
        RECT 2835.020 2123.380 2838.020 2123.390 ;
        RECT 2950.100 2123.380 2953.100 2123.390 ;
        RECT -33.480 2120.380 2953.100 2123.380 ;
        RECT -33.480 2120.370 -30.480 2120.380 ;
        RECT 135.020 2120.370 138.020 2120.380 ;
        RECT 315.020 2120.370 318.020 2120.380 ;
        RECT 495.020 2120.370 498.020 2120.380 ;
        RECT 675.020 2120.370 678.020 2120.380 ;
        RECT 855.020 2120.370 858.020 2120.380 ;
        RECT 1035.020 2120.370 1038.020 2120.380 ;
        RECT 1215.020 2120.370 1218.020 2120.380 ;
        RECT 1395.020 2120.370 1398.020 2120.380 ;
        RECT 1575.020 2120.370 1578.020 2120.380 ;
        RECT 1755.020 2120.370 1758.020 2120.380 ;
        RECT 1935.020 2120.370 1938.020 2120.380 ;
        RECT 2115.020 2120.370 2118.020 2120.380 ;
        RECT 2295.020 2120.370 2298.020 2120.380 ;
        RECT 2475.020 2120.370 2478.020 2120.380 ;
        RECT 2655.020 2120.370 2658.020 2120.380 ;
        RECT 2835.020 2120.370 2838.020 2120.380 ;
        RECT 2950.100 2120.370 2953.100 2120.380 ;
        RECT -33.480 1943.380 -30.480 1943.390 ;
        RECT 135.020 1943.380 138.020 1943.390 ;
        RECT 315.020 1943.380 318.020 1943.390 ;
        RECT 495.020 1943.380 498.020 1943.390 ;
        RECT 675.020 1943.380 678.020 1943.390 ;
        RECT 855.020 1943.380 858.020 1943.390 ;
        RECT 1035.020 1943.380 1038.020 1943.390 ;
        RECT 1215.020 1943.380 1218.020 1943.390 ;
        RECT 1395.020 1943.380 1398.020 1943.390 ;
        RECT 1575.020 1943.380 1578.020 1943.390 ;
        RECT 1755.020 1943.380 1758.020 1943.390 ;
        RECT 1935.020 1943.380 1938.020 1943.390 ;
        RECT 2115.020 1943.380 2118.020 1943.390 ;
        RECT 2295.020 1943.380 2298.020 1943.390 ;
        RECT 2475.020 1943.380 2478.020 1943.390 ;
        RECT 2655.020 1943.380 2658.020 1943.390 ;
        RECT 2835.020 1943.380 2838.020 1943.390 ;
        RECT 2950.100 1943.380 2953.100 1943.390 ;
        RECT -33.480 1940.380 2953.100 1943.380 ;
        RECT -33.480 1940.370 -30.480 1940.380 ;
        RECT 135.020 1940.370 138.020 1940.380 ;
        RECT 315.020 1940.370 318.020 1940.380 ;
        RECT 495.020 1940.370 498.020 1940.380 ;
        RECT 675.020 1940.370 678.020 1940.380 ;
        RECT 855.020 1940.370 858.020 1940.380 ;
        RECT 1035.020 1940.370 1038.020 1940.380 ;
        RECT 1215.020 1940.370 1218.020 1940.380 ;
        RECT 1395.020 1940.370 1398.020 1940.380 ;
        RECT 1575.020 1940.370 1578.020 1940.380 ;
        RECT 1755.020 1940.370 1758.020 1940.380 ;
        RECT 1935.020 1940.370 1938.020 1940.380 ;
        RECT 2115.020 1940.370 2118.020 1940.380 ;
        RECT 2295.020 1940.370 2298.020 1940.380 ;
        RECT 2475.020 1940.370 2478.020 1940.380 ;
        RECT 2655.020 1940.370 2658.020 1940.380 ;
        RECT 2835.020 1940.370 2838.020 1940.380 ;
        RECT 2950.100 1940.370 2953.100 1940.380 ;
        RECT -33.480 1763.380 -30.480 1763.390 ;
        RECT 135.020 1763.380 138.020 1763.390 ;
        RECT 315.020 1763.380 318.020 1763.390 ;
        RECT 495.020 1763.380 498.020 1763.390 ;
        RECT 675.020 1763.380 678.020 1763.390 ;
        RECT 855.020 1763.380 858.020 1763.390 ;
        RECT 1035.020 1763.380 1038.020 1763.390 ;
        RECT 1215.020 1763.380 1218.020 1763.390 ;
        RECT 1395.020 1763.380 1398.020 1763.390 ;
        RECT 1575.020 1763.380 1578.020 1763.390 ;
        RECT 1755.020 1763.380 1758.020 1763.390 ;
        RECT 1935.020 1763.380 1938.020 1763.390 ;
        RECT 2115.020 1763.380 2118.020 1763.390 ;
        RECT 2295.020 1763.380 2298.020 1763.390 ;
        RECT 2475.020 1763.380 2478.020 1763.390 ;
        RECT 2655.020 1763.380 2658.020 1763.390 ;
        RECT 2835.020 1763.380 2838.020 1763.390 ;
        RECT 2950.100 1763.380 2953.100 1763.390 ;
        RECT -33.480 1760.380 2953.100 1763.380 ;
        RECT -33.480 1760.370 -30.480 1760.380 ;
        RECT 135.020 1760.370 138.020 1760.380 ;
        RECT 315.020 1760.370 318.020 1760.380 ;
        RECT 495.020 1760.370 498.020 1760.380 ;
        RECT 675.020 1760.370 678.020 1760.380 ;
        RECT 855.020 1760.370 858.020 1760.380 ;
        RECT 1035.020 1760.370 1038.020 1760.380 ;
        RECT 1215.020 1760.370 1218.020 1760.380 ;
        RECT 1395.020 1760.370 1398.020 1760.380 ;
        RECT 1575.020 1760.370 1578.020 1760.380 ;
        RECT 1755.020 1760.370 1758.020 1760.380 ;
        RECT 1935.020 1760.370 1938.020 1760.380 ;
        RECT 2115.020 1760.370 2118.020 1760.380 ;
        RECT 2295.020 1760.370 2298.020 1760.380 ;
        RECT 2475.020 1760.370 2478.020 1760.380 ;
        RECT 2655.020 1760.370 2658.020 1760.380 ;
        RECT 2835.020 1760.370 2838.020 1760.380 ;
        RECT 2950.100 1760.370 2953.100 1760.380 ;
        RECT -33.480 1583.380 -30.480 1583.390 ;
        RECT 135.020 1583.380 138.020 1583.390 ;
        RECT 315.020 1583.380 318.020 1583.390 ;
        RECT 495.020 1583.380 498.020 1583.390 ;
        RECT 675.020 1583.380 678.020 1583.390 ;
        RECT 855.020 1583.380 858.020 1583.390 ;
        RECT 1035.020 1583.380 1038.020 1583.390 ;
        RECT 1215.020 1583.380 1218.020 1583.390 ;
        RECT 1395.020 1583.380 1398.020 1583.390 ;
        RECT 1575.020 1583.380 1578.020 1583.390 ;
        RECT 1755.020 1583.380 1758.020 1583.390 ;
        RECT 1935.020 1583.380 1938.020 1583.390 ;
        RECT 2115.020 1583.380 2118.020 1583.390 ;
        RECT 2295.020 1583.380 2298.020 1583.390 ;
        RECT 2475.020 1583.380 2478.020 1583.390 ;
        RECT 2655.020 1583.380 2658.020 1583.390 ;
        RECT 2835.020 1583.380 2838.020 1583.390 ;
        RECT 2950.100 1583.380 2953.100 1583.390 ;
        RECT -33.480 1580.380 2953.100 1583.380 ;
        RECT -33.480 1580.370 -30.480 1580.380 ;
        RECT 135.020 1580.370 138.020 1580.380 ;
        RECT 315.020 1580.370 318.020 1580.380 ;
        RECT 495.020 1580.370 498.020 1580.380 ;
        RECT 675.020 1580.370 678.020 1580.380 ;
        RECT 855.020 1580.370 858.020 1580.380 ;
        RECT 1035.020 1580.370 1038.020 1580.380 ;
        RECT 1215.020 1580.370 1218.020 1580.380 ;
        RECT 1395.020 1580.370 1398.020 1580.380 ;
        RECT 1575.020 1580.370 1578.020 1580.380 ;
        RECT 1755.020 1580.370 1758.020 1580.380 ;
        RECT 1935.020 1580.370 1938.020 1580.380 ;
        RECT 2115.020 1580.370 2118.020 1580.380 ;
        RECT 2295.020 1580.370 2298.020 1580.380 ;
        RECT 2475.020 1580.370 2478.020 1580.380 ;
        RECT 2655.020 1580.370 2658.020 1580.380 ;
        RECT 2835.020 1580.370 2838.020 1580.380 ;
        RECT 2950.100 1580.370 2953.100 1580.380 ;
        RECT -33.480 1403.380 -30.480 1403.390 ;
        RECT 135.020 1403.380 138.020 1403.390 ;
        RECT 315.020 1403.380 318.020 1403.390 ;
        RECT 495.020 1403.380 498.020 1403.390 ;
        RECT 675.020 1403.380 678.020 1403.390 ;
        RECT 855.020 1403.380 858.020 1403.390 ;
        RECT 1035.020 1403.380 1038.020 1403.390 ;
        RECT 1215.020 1403.380 1218.020 1403.390 ;
        RECT 1395.020 1403.380 1398.020 1403.390 ;
        RECT 1575.020 1403.380 1578.020 1403.390 ;
        RECT 1755.020 1403.380 1758.020 1403.390 ;
        RECT 1935.020 1403.380 1938.020 1403.390 ;
        RECT 2115.020 1403.380 2118.020 1403.390 ;
        RECT 2295.020 1403.380 2298.020 1403.390 ;
        RECT 2475.020 1403.380 2478.020 1403.390 ;
        RECT 2655.020 1403.380 2658.020 1403.390 ;
        RECT 2835.020 1403.380 2838.020 1403.390 ;
        RECT 2950.100 1403.380 2953.100 1403.390 ;
        RECT -33.480 1400.380 2953.100 1403.380 ;
        RECT -33.480 1400.370 -30.480 1400.380 ;
        RECT 135.020 1400.370 138.020 1400.380 ;
        RECT 315.020 1400.370 318.020 1400.380 ;
        RECT 495.020 1400.370 498.020 1400.380 ;
        RECT 675.020 1400.370 678.020 1400.380 ;
        RECT 855.020 1400.370 858.020 1400.380 ;
        RECT 1035.020 1400.370 1038.020 1400.380 ;
        RECT 1215.020 1400.370 1218.020 1400.380 ;
        RECT 1395.020 1400.370 1398.020 1400.380 ;
        RECT 1575.020 1400.370 1578.020 1400.380 ;
        RECT 1755.020 1400.370 1758.020 1400.380 ;
        RECT 1935.020 1400.370 1938.020 1400.380 ;
        RECT 2115.020 1400.370 2118.020 1400.380 ;
        RECT 2295.020 1400.370 2298.020 1400.380 ;
        RECT 2475.020 1400.370 2478.020 1400.380 ;
        RECT 2655.020 1400.370 2658.020 1400.380 ;
        RECT 2835.020 1400.370 2838.020 1400.380 ;
        RECT 2950.100 1400.370 2953.100 1400.380 ;
        RECT -33.480 1223.380 -30.480 1223.390 ;
        RECT 135.020 1223.380 138.020 1223.390 ;
        RECT 315.020 1223.380 318.020 1223.390 ;
        RECT 495.020 1223.380 498.020 1223.390 ;
        RECT 675.020 1223.380 678.020 1223.390 ;
        RECT 855.020 1223.380 858.020 1223.390 ;
        RECT 1035.020 1223.380 1038.020 1223.390 ;
        RECT 1215.020 1223.380 1218.020 1223.390 ;
        RECT 1395.020 1223.380 1398.020 1223.390 ;
        RECT 1575.020 1223.380 1578.020 1223.390 ;
        RECT 1755.020 1223.380 1758.020 1223.390 ;
        RECT 1935.020 1223.380 1938.020 1223.390 ;
        RECT 2115.020 1223.380 2118.020 1223.390 ;
        RECT 2295.020 1223.380 2298.020 1223.390 ;
        RECT 2475.020 1223.380 2478.020 1223.390 ;
        RECT 2655.020 1223.380 2658.020 1223.390 ;
        RECT 2835.020 1223.380 2838.020 1223.390 ;
        RECT 2950.100 1223.380 2953.100 1223.390 ;
        RECT -33.480 1220.380 2953.100 1223.380 ;
        RECT -33.480 1220.370 -30.480 1220.380 ;
        RECT 135.020 1220.370 138.020 1220.380 ;
        RECT 315.020 1220.370 318.020 1220.380 ;
        RECT 495.020 1220.370 498.020 1220.380 ;
        RECT 675.020 1220.370 678.020 1220.380 ;
        RECT 855.020 1220.370 858.020 1220.380 ;
        RECT 1035.020 1220.370 1038.020 1220.380 ;
        RECT 1215.020 1220.370 1218.020 1220.380 ;
        RECT 1395.020 1220.370 1398.020 1220.380 ;
        RECT 1575.020 1220.370 1578.020 1220.380 ;
        RECT 1755.020 1220.370 1758.020 1220.380 ;
        RECT 1935.020 1220.370 1938.020 1220.380 ;
        RECT 2115.020 1220.370 2118.020 1220.380 ;
        RECT 2295.020 1220.370 2298.020 1220.380 ;
        RECT 2475.020 1220.370 2478.020 1220.380 ;
        RECT 2655.020 1220.370 2658.020 1220.380 ;
        RECT 2835.020 1220.370 2838.020 1220.380 ;
        RECT 2950.100 1220.370 2953.100 1220.380 ;
        RECT -33.480 1043.380 -30.480 1043.390 ;
        RECT 135.020 1043.380 138.020 1043.390 ;
        RECT 315.020 1043.380 318.020 1043.390 ;
        RECT 495.020 1043.380 498.020 1043.390 ;
        RECT 675.020 1043.380 678.020 1043.390 ;
        RECT 855.020 1043.380 858.020 1043.390 ;
        RECT 1035.020 1043.380 1038.020 1043.390 ;
        RECT 1215.020 1043.380 1218.020 1043.390 ;
        RECT 1395.020 1043.380 1398.020 1043.390 ;
        RECT 1575.020 1043.380 1578.020 1043.390 ;
        RECT 1755.020 1043.380 1758.020 1043.390 ;
        RECT 1935.020 1043.380 1938.020 1043.390 ;
        RECT 2115.020 1043.380 2118.020 1043.390 ;
        RECT 2295.020 1043.380 2298.020 1043.390 ;
        RECT 2475.020 1043.380 2478.020 1043.390 ;
        RECT 2655.020 1043.380 2658.020 1043.390 ;
        RECT 2835.020 1043.380 2838.020 1043.390 ;
        RECT 2950.100 1043.380 2953.100 1043.390 ;
        RECT -33.480 1040.380 2953.100 1043.380 ;
        RECT -33.480 1040.370 -30.480 1040.380 ;
        RECT 135.020 1040.370 138.020 1040.380 ;
        RECT 315.020 1040.370 318.020 1040.380 ;
        RECT 495.020 1040.370 498.020 1040.380 ;
        RECT 675.020 1040.370 678.020 1040.380 ;
        RECT 855.020 1040.370 858.020 1040.380 ;
        RECT 1035.020 1040.370 1038.020 1040.380 ;
        RECT 1215.020 1040.370 1218.020 1040.380 ;
        RECT 1395.020 1040.370 1398.020 1040.380 ;
        RECT 1575.020 1040.370 1578.020 1040.380 ;
        RECT 1755.020 1040.370 1758.020 1040.380 ;
        RECT 1935.020 1040.370 1938.020 1040.380 ;
        RECT 2115.020 1040.370 2118.020 1040.380 ;
        RECT 2295.020 1040.370 2298.020 1040.380 ;
        RECT 2475.020 1040.370 2478.020 1040.380 ;
        RECT 2655.020 1040.370 2658.020 1040.380 ;
        RECT 2835.020 1040.370 2838.020 1040.380 ;
        RECT 2950.100 1040.370 2953.100 1040.380 ;
        RECT -33.480 863.380 -30.480 863.390 ;
        RECT 135.020 863.380 138.020 863.390 ;
        RECT 315.020 863.380 318.020 863.390 ;
        RECT 495.020 863.380 498.020 863.390 ;
        RECT 675.020 863.380 678.020 863.390 ;
        RECT 855.020 863.380 858.020 863.390 ;
        RECT 1035.020 863.380 1038.020 863.390 ;
        RECT 1215.020 863.380 1218.020 863.390 ;
        RECT 1395.020 863.380 1398.020 863.390 ;
        RECT 1575.020 863.380 1578.020 863.390 ;
        RECT 1755.020 863.380 1758.020 863.390 ;
        RECT 1935.020 863.380 1938.020 863.390 ;
        RECT 2115.020 863.380 2118.020 863.390 ;
        RECT 2295.020 863.380 2298.020 863.390 ;
        RECT 2475.020 863.380 2478.020 863.390 ;
        RECT 2655.020 863.380 2658.020 863.390 ;
        RECT 2835.020 863.380 2838.020 863.390 ;
        RECT 2950.100 863.380 2953.100 863.390 ;
        RECT -33.480 860.380 2953.100 863.380 ;
        RECT -33.480 860.370 -30.480 860.380 ;
        RECT 135.020 860.370 138.020 860.380 ;
        RECT 315.020 860.370 318.020 860.380 ;
        RECT 495.020 860.370 498.020 860.380 ;
        RECT 675.020 860.370 678.020 860.380 ;
        RECT 855.020 860.370 858.020 860.380 ;
        RECT 1035.020 860.370 1038.020 860.380 ;
        RECT 1215.020 860.370 1218.020 860.380 ;
        RECT 1395.020 860.370 1398.020 860.380 ;
        RECT 1575.020 860.370 1578.020 860.380 ;
        RECT 1755.020 860.370 1758.020 860.380 ;
        RECT 1935.020 860.370 1938.020 860.380 ;
        RECT 2115.020 860.370 2118.020 860.380 ;
        RECT 2295.020 860.370 2298.020 860.380 ;
        RECT 2475.020 860.370 2478.020 860.380 ;
        RECT 2655.020 860.370 2658.020 860.380 ;
        RECT 2835.020 860.370 2838.020 860.380 ;
        RECT 2950.100 860.370 2953.100 860.380 ;
        RECT -33.480 683.380 -30.480 683.390 ;
        RECT 135.020 683.380 138.020 683.390 ;
        RECT 315.020 683.380 318.020 683.390 ;
        RECT 495.020 683.380 498.020 683.390 ;
        RECT 675.020 683.380 678.020 683.390 ;
        RECT 855.020 683.380 858.020 683.390 ;
        RECT 1035.020 683.380 1038.020 683.390 ;
        RECT 1215.020 683.380 1218.020 683.390 ;
        RECT 1395.020 683.380 1398.020 683.390 ;
        RECT 1575.020 683.380 1578.020 683.390 ;
        RECT 1755.020 683.380 1758.020 683.390 ;
        RECT 1935.020 683.380 1938.020 683.390 ;
        RECT 2115.020 683.380 2118.020 683.390 ;
        RECT 2295.020 683.380 2298.020 683.390 ;
        RECT 2475.020 683.380 2478.020 683.390 ;
        RECT 2655.020 683.380 2658.020 683.390 ;
        RECT 2835.020 683.380 2838.020 683.390 ;
        RECT 2950.100 683.380 2953.100 683.390 ;
        RECT -33.480 680.380 2953.100 683.380 ;
        RECT -33.480 680.370 -30.480 680.380 ;
        RECT 135.020 680.370 138.020 680.380 ;
        RECT 315.020 680.370 318.020 680.380 ;
        RECT 495.020 680.370 498.020 680.380 ;
        RECT 675.020 680.370 678.020 680.380 ;
        RECT 855.020 680.370 858.020 680.380 ;
        RECT 1035.020 680.370 1038.020 680.380 ;
        RECT 1215.020 680.370 1218.020 680.380 ;
        RECT 1395.020 680.370 1398.020 680.380 ;
        RECT 1575.020 680.370 1578.020 680.380 ;
        RECT 1755.020 680.370 1758.020 680.380 ;
        RECT 1935.020 680.370 1938.020 680.380 ;
        RECT 2115.020 680.370 2118.020 680.380 ;
        RECT 2295.020 680.370 2298.020 680.380 ;
        RECT 2475.020 680.370 2478.020 680.380 ;
        RECT 2655.020 680.370 2658.020 680.380 ;
        RECT 2835.020 680.370 2838.020 680.380 ;
        RECT 2950.100 680.370 2953.100 680.380 ;
        RECT -33.480 503.380 -30.480 503.390 ;
        RECT 135.020 503.380 138.020 503.390 ;
        RECT 315.020 503.380 318.020 503.390 ;
        RECT 495.020 503.380 498.020 503.390 ;
        RECT 675.020 503.380 678.020 503.390 ;
        RECT 855.020 503.380 858.020 503.390 ;
        RECT 1035.020 503.380 1038.020 503.390 ;
        RECT 1215.020 503.380 1218.020 503.390 ;
        RECT 1395.020 503.380 1398.020 503.390 ;
        RECT 1575.020 503.380 1578.020 503.390 ;
        RECT 1755.020 503.380 1758.020 503.390 ;
        RECT 1935.020 503.380 1938.020 503.390 ;
        RECT 2115.020 503.380 2118.020 503.390 ;
        RECT 2295.020 503.380 2298.020 503.390 ;
        RECT 2475.020 503.380 2478.020 503.390 ;
        RECT 2655.020 503.380 2658.020 503.390 ;
        RECT 2835.020 503.380 2838.020 503.390 ;
        RECT 2950.100 503.380 2953.100 503.390 ;
        RECT -33.480 500.380 2953.100 503.380 ;
        RECT -33.480 500.370 -30.480 500.380 ;
        RECT 135.020 500.370 138.020 500.380 ;
        RECT 315.020 500.370 318.020 500.380 ;
        RECT 495.020 500.370 498.020 500.380 ;
        RECT 675.020 500.370 678.020 500.380 ;
        RECT 855.020 500.370 858.020 500.380 ;
        RECT 1035.020 500.370 1038.020 500.380 ;
        RECT 1215.020 500.370 1218.020 500.380 ;
        RECT 1395.020 500.370 1398.020 500.380 ;
        RECT 1575.020 500.370 1578.020 500.380 ;
        RECT 1755.020 500.370 1758.020 500.380 ;
        RECT 1935.020 500.370 1938.020 500.380 ;
        RECT 2115.020 500.370 2118.020 500.380 ;
        RECT 2295.020 500.370 2298.020 500.380 ;
        RECT 2475.020 500.370 2478.020 500.380 ;
        RECT 2655.020 500.370 2658.020 500.380 ;
        RECT 2835.020 500.370 2838.020 500.380 ;
        RECT 2950.100 500.370 2953.100 500.380 ;
        RECT -33.480 323.380 -30.480 323.390 ;
        RECT 135.020 323.380 138.020 323.390 ;
        RECT 315.020 323.380 318.020 323.390 ;
        RECT 495.020 323.380 498.020 323.390 ;
        RECT 675.020 323.380 678.020 323.390 ;
        RECT 855.020 323.380 858.020 323.390 ;
        RECT 1035.020 323.380 1038.020 323.390 ;
        RECT 1215.020 323.380 1218.020 323.390 ;
        RECT 1395.020 323.380 1398.020 323.390 ;
        RECT 1575.020 323.380 1578.020 323.390 ;
        RECT 1755.020 323.380 1758.020 323.390 ;
        RECT 1935.020 323.380 1938.020 323.390 ;
        RECT 2115.020 323.380 2118.020 323.390 ;
        RECT 2295.020 323.380 2298.020 323.390 ;
        RECT 2475.020 323.380 2478.020 323.390 ;
        RECT 2655.020 323.380 2658.020 323.390 ;
        RECT 2835.020 323.380 2838.020 323.390 ;
        RECT 2950.100 323.380 2953.100 323.390 ;
        RECT -33.480 320.380 2953.100 323.380 ;
        RECT -33.480 320.370 -30.480 320.380 ;
        RECT 135.020 320.370 138.020 320.380 ;
        RECT 315.020 320.370 318.020 320.380 ;
        RECT 495.020 320.370 498.020 320.380 ;
        RECT 675.020 320.370 678.020 320.380 ;
        RECT 855.020 320.370 858.020 320.380 ;
        RECT 1035.020 320.370 1038.020 320.380 ;
        RECT 1215.020 320.370 1218.020 320.380 ;
        RECT 1395.020 320.370 1398.020 320.380 ;
        RECT 1575.020 320.370 1578.020 320.380 ;
        RECT 1755.020 320.370 1758.020 320.380 ;
        RECT 1935.020 320.370 1938.020 320.380 ;
        RECT 2115.020 320.370 2118.020 320.380 ;
        RECT 2295.020 320.370 2298.020 320.380 ;
        RECT 2475.020 320.370 2478.020 320.380 ;
        RECT 2655.020 320.370 2658.020 320.380 ;
        RECT 2835.020 320.370 2838.020 320.380 ;
        RECT 2950.100 320.370 2953.100 320.380 ;
        RECT -33.480 143.380 -30.480 143.390 ;
        RECT 135.020 143.380 138.020 143.390 ;
        RECT 315.020 143.380 318.020 143.390 ;
        RECT 495.020 143.380 498.020 143.390 ;
        RECT 675.020 143.380 678.020 143.390 ;
        RECT 855.020 143.380 858.020 143.390 ;
        RECT 1035.020 143.380 1038.020 143.390 ;
        RECT 1215.020 143.380 1218.020 143.390 ;
        RECT 1395.020 143.380 1398.020 143.390 ;
        RECT 1575.020 143.380 1578.020 143.390 ;
        RECT 1755.020 143.380 1758.020 143.390 ;
        RECT 1935.020 143.380 1938.020 143.390 ;
        RECT 2115.020 143.380 2118.020 143.390 ;
        RECT 2295.020 143.380 2298.020 143.390 ;
        RECT 2475.020 143.380 2478.020 143.390 ;
        RECT 2655.020 143.380 2658.020 143.390 ;
        RECT 2835.020 143.380 2838.020 143.390 ;
        RECT 2950.100 143.380 2953.100 143.390 ;
        RECT -33.480 140.380 2953.100 143.380 ;
        RECT -33.480 140.370 -30.480 140.380 ;
        RECT 135.020 140.370 138.020 140.380 ;
        RECT 315.020 140.370 318.020 140.380 ;
        RECT 495.020 140.370 498.020 140.380 ;
        RECT 675.020 140.370 678.020 140.380 ;
        RECT 855.020 140.370 858.020 140.380 ;
        RECT 1035.020 140.370 1038.020 140.380 ;
        RECT 1215.020 140.370 1218.020 140.380 ;
        RECT 1395.020 140.370 1398.020 140.380 ;
        RECT 1575.020 140.370 1578.020 140.380 ;
        RECT 1755.020 140.370 1758.020 140.380 ;
        RECT 1935.020 140.370 1938.020 140.380 ;
        RECT 2115.020 140.370 2118.020 140.380 ;
        RECT 2295.020 140.370 2298.020 140.380 ;
        RECT 2475.020 140.370 2478.020 140.380 ;
        RECT 2655.020 140.370 2658.020 140.380 ;
        RECT 2835.020 140.370 2838.020 140.380 ;
        RECT 2950.100 140.370 2953.100 140.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 135.020 -25.120 138.020 -25.110 ;
        RECT 315.020 -25.120 318.020 -25.110 ;
        RECT 495.020 -25.120 498.020 -25.110 ;
        RECT 675.020 -25.120 678.020 -25.110 ;
        RECT 855.020 -25.120 858.020 -25.110 ;
        RECT 1035.020 -25.120 1038.020 -25.110 ;
        RECT 1215.020 -25.120 1218.020 -25.110 ;
        RECT 1395.020 -25.120 1398.020 -25.110 ;
        RECT 1575.020 -25.120 1578.020 -25.110 ;
        RECT 1755.020 -25.120 1758.020 -25.110 ;
        RECT 1935.020 -25.120 1938.020 -25.110 ;
        RECT 2115.020 -25.120 2118.020 -25.110 ;
        RECT 2295.020 -25.120 2298.020 -25.110 ;
        RECT 2475.020 -25.120 2478.020 -25.110 ;
        RECT 2655.020 -25.120 2658.020 -25.110 ;
        RECT 2835.020 -25.120 2838.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 135.020 -28.130 138.020 -28.120 ;
        RECT 315.020 -28.130 318.020 -28.120 ;
        RECT 495.020 -28.130 498.020 -28.120 ;
        RECT 675.020 -28.130 678.020 -28.120 ;
        RECT 855.020 -28.130 858.020 -28.120 ;
        RECT 1035.020 -28.130 1038.020 -28.120 ;
        RECT 1215.020 -28.130 1218.020 -28.120 ;
        RECT 1395.020 -28.130 1398.020 -28.120 ;
        RECT 1575.020 -28.130 1578.020 -28.120 ;
        RECT 1755.020 -28.130 1758.020 -28.120 ;
        RECT 1935.020 -28.130 1938.020 -28.120 ;
        RECT 2115.020 -28.130 2118.020 -28.120 ;
        RECT 2295.020 -28.130 2298.020 -28.120 ;
        RECT 2475.020 -28.130 2478.020 -28.120 ;
        RECT 2655.020 -28.130 2658.020 -28.120 ;
        RECT 2835.020 -28.130 2838.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 63.020 -37.520 66.020 3557.200 ;
        RECT 243.020 -37.520 246.020 3557.200 ;
        RECT 423.020 -37.520 426.020 3557.200 ;
        RECT 603.020 -37.520 606.020 3557.200 ;
        RECT 783.020 -37.520 786.020 3557.200 ;
        RECT 963.020 -37.520 966.020 3557.200 ;
        RECT 1143.020 -37.520 1146.020 3557.200 ;
        RECT 1323.020 -37.520 1326.020 3557.200 ;
        RECT 1503.020 -37.520 1506.020 3557.200 ;
        RECT 1683.020 -37.520 1686.020 3557.200 ;
        RECT 1863.020 -37.520 1866.020 3557.200 ;
        RECT 2043.020 -37.520 2046.020 3557.200 ;
        RECT 2223.020 -37.520 2226.020 3557.200 ;
        RECT 2403.020 -37.520 2406.020 3557.200 ;
        RECT 2583.020 -37.520 2586.020 3557.200 ;
        RECT 2763.020 -37.520 2766.020 3557.200 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 3490.090 -36.090 3491.270 ;
        RECT -37.270 3488.490 -36.090 3489.670 ;
        RECT -37.270 3310.090 -36.090 3311.270 ;
        RECT -37.270 3308.490 -36.090 3309.670 ;
        RECT -37.270 3130.090 -36.090 3131.270 ;
        RECT -37.270 3128.490 -36.090 3129.670 ;
        RECT -37.270 2950.090 -36.090 2951.270 ;
        RECT -37.270 2948.490 -36.090 2949.670 ;
        RECT -37.270 2770.090 -36.090 2771.270 ;
        RECT -37.270 2768.490 -36.090 2769.670 ;
        RECT -37.270 2590.090 -36.090 2591.270 ;
        RECT -37.270 2588.490 -36.090 2589.670 ;
        RECT -37.270 2410.090 -36.090 2411.270 ;
        RECT -37.270 2408.490 -36.090 2409.670 ;
        RECT -37.270 2230.090 -36.090 2231.270 ;
        RECT -37.270 2228.490 -36.090 2229.670 ;
        RECT -37.270 2050.090 -36.090 2051.270 ;
        RECT -37.270 2048.490 -36.090 2049.670 ;
        RECT -37.270 1870.090 -36.090 1871.270 ;
        RECT -37.270 1868.490 -36.090 1869.670 ;
        RECT -37.270 1690.090 -36.090 1691.270 ;
        RECT -37.270 1688.490 -36.090 1689.670 ;
        RECT -37.270 1510.090 -36.090 1511.270 ;
        RECT -37.270 1508.490 -36.090 1509.670 ;
        RECT -37.270 1330.090 -36.090 1331.270 ;
        RECT -37.270 1328.490 -36.090 1329.670 ;
        RECT -37.270 1150.090 -36.090 1151.270 ;
        RECT -37.270 1148.490 -36.090 1149.670 ;
        RECT -37.270 970.090 -36.090 971.270 ;
        RECT -37.270 968.490 -36.090 969.670 ;
        RECT -37.270 790.090 -36.090 791.270 ;
        RECT -37.270 788.490 -36.090 789.670 ;
        RECT -37.270 610.090 -36.090 611.270 ;
        RECT -37.270 608.490 -36.090 609.670 ;
        RECT -37.270 430.090 -36.090 431.270 ;
        RECT -37.270 428.490 -36.090 429.670 ;
        RECT -37.270 250.090 -36.090 251.270 ;
        RECT -37.270 248.490 -36.090 249.670 ;
        RECT -37.270 70.090 -36.090 71.270 ;
        RECT -37.270 68.490 -36.090 69.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 63.930 3551.210 65.110 3552.390 ;
        RECT 63.930 3549.610 65.110 3550.790 ;
        RECT 63.930 3490.090 65.110 3491.270 ;
        RECT 63.930 3488.490 65.110 3489.670 ;
        RECT 63.930 3310.090 65.110 3311.270 ;
        RECT 63.930 3308.490 65.110 3309.670 ;
        RECT 63.930 3130.090 65.110 3131.270 ;
        RECT 63.930 3128.490 65.110 3129.670 ;
        RECT 63.930 2950.090 65.110 2951.270 ;
        RECT 63.930 2948.490 65.110 2949.670 ;
        RECT 63.930 2770.090 65.110 2771.270 ;
        RECT 63.930 2768.490 65.110 2769.670 ;
        RECT 63.930 2590.090 65.110 2591.270 ;
        RECT 63.930 2588.490 65.110 2589.670 ;
        RECT 63.930 2410.090 65.110 2411.270 ;
        RECT 63.930 2408.490 65.110 2409.670 ;
        RECT 63.930 2230.090 65.110 2231.270 ;
        RECT 63.930 2228.490 65.110 2229.670 ;
        RECT 63.930 2050.090 65.110 2051.270 ;
        RECT 63.930 2048.490 65.110 2049.670 ;
        RECT 63.930 1870.090 65.110 1871.270 ;
        RECT 63.930 1868.490 65.110 1869.670 ;
        RECT 63.930 1690.090 65.110 1691.270 ;
        RECT 63.930 1688.490 65.110 1689.670 ;
        RECT 63.930 1510.090 65.110 1511.270 ;
        RECT 63.930 1508.490 65.110 1509.670 ;
        RECT 63.930 1330.090 65.110 1331.270 ;
        RECT 63.930 1328.490 65.110 1329.670 ;
        RECT 63.930 1150.090 65.110 1151.270 ;
        RECT 63.930 1148.490 65.110 1149.670 ;
        RECT 63.930 970.090 65.110 971.270 ;
        RECT 63.930 968.490 65.110 969.670 ;
        RECT 63.930 790.090 65.110 791.270 ;
        RECT 63.930 788.490 65.110 789.670 ;
        RECT 63.930 610.090 65.110 611.270 ;
        RECT 63.930 608.490 65.110 609.670 ;
        RECT 63.930 430.090 65.110 431.270 ;
        RECT 63.930 428.490 65.110 429.670 ;
        RECT 63.930 250.090 65.110 251.270 ;
        RECT 63.930 248.490 65.110 249.670 ;
        RECT 63.930 70.090 65.110 71.270 ;
        RECT 63.930 68.490 65.110 69.670 ;
        RECT 63.930 -31.110 65.110 -29.930 ;
        RECT 63.930 -32.710 65.110 -31.530 ;
        RECT 243.930 3551.210 245.110 3552.390 ;
        RECT 243.930 3549.610 245.110 3550.790 ;
        RECT 243.930 3490.090 245.110 3491.270 ;
        RECT 243.930 3488.490 245.110 3489.670 ;
        RECT 243.930 3310.090 245.110 3311.270 ;
        RECT 243.930 3308.490 245.110 3309.670 ;
        RECT 243.930 3130.090 245.110 3131.270 ;
        RECT 243.930 3128.490 245.110 3129.670 ;
        RECT 243.930 2950.090 245.110 2951.270 ;
        RECT 243.930 2948.490 245.110 2949.670 ;
        RECT 243.930 2770.090 245.110 2771.270 ;
        RECT 243.930 2768.490 245.110 2769.670 ;
        RECT 243.930 2590.090 245.110 2591.270 ;
        RECT 243.930 2588.490 245.110 2589.670 ;
        RECT 243.930 2410.090 245.110 2411.270 ;
        RECT 243.930 2408.490 245.110 2409.670 ;
        RECT 243.930 2230.090 245.110 2231.270 ;
        RECT 243.930 2228.490 245.110 2229.670 ;
        RECT 243.930 2050.090 245.110 2051.270 ;
        RECT 243.930 2048.490 245.110 2049.670 ;
        RECT 243.930 1870.090 245.110 1871.270 ;
        RECT 243.930 1868.490 245.110 1869.670 ;
        RECT 243.930 1690.090 245.110 1691.270 ;
        RECT 243.930 1688.490 245.110 1689.670 ;
        RECT 243.930 1510.090 245.110 1511.270 ;
        RECT 243.930 1508.490 245.110 1509.670 ;
        RECT 243.930 1330.090 245.110 1331.270 ;
        RECT 243.930 1328.490 245.110 1329.670 ;
        RECT 243.930 1150.090 245.110 1151.270 ;
        RECT 243.930 1148.490 245.110 1149.670 ;
        RECT 243.930 970.090 245.110 971.270 ;
        RECT 243.930 968.490 245.110 969.670 ;
        RECT 243.930 790.090 245.110 791.270 ;
        RECT 243.930 788.490 245.110 789.670 ;
        RECT 243.930 610.090 245.110 611.270 ;
        RECT 243.930 608.490 245.110 609.670 ;
        RECT 243.930 430.090 245.110 431.270 ;
        RECT 243.930 428.490 245.110 429.670 ;
        RECT 243.930 250.090 245.110 251.270 ;
        RECT 243.930 248.490 245.110 249.670 ;
        RECT 243.930 70.090 245.110 71.270 ;
        RECT 243.930 68.490 245.110 69.670 ;
        RECT 243.930 -31.110 245.110 -29.930 ;
        RECT 243.930 -32.710 245.110 -31.530 ;
        RECT 423.930 3551.210 425.110 3552.390 ;
        RECT 423.930 3549.610 425.110 3550.790 ;
        RECT 423.930 3490.090 425.110 3491.270 ;
        RECT 423.930 3488.490 425.110 3489.670 ;
        RECT 423.930 3310.090 425.110 3311.270 ;
        RECT 423.930 3308.490 425.110 3309.670 ;
        RECT 423.930 3130.090 425.110 3131.270 ;
        RECT 423.930 3128.490 425.110 3129.670 ;
        RECT 423.930 2950.090 425.110 2951.270 ;
        RECT 423.930 2948.490 425.110 2949.670 ;
        RECT 423.930 2770.090 425.110 2771.270 ;
        RECT 423.930 2768.490 425.110 2769.670 ;
        RECT 423.930 2590.090 425.110 2591.270 ;
        RECT 423.930 2588.490 425.110 2589.670 ;
        RECT 423.930 2410.090 425.110 2411.270 ;
        RECT 423.930 2408.490 425.110 2409.670 ;
        RECT 423.930 2230.090 425.110 2231.270 ;
        RECT 423.930 2228.490 425.110 2229.670 ;
        RECT 423.930 2050.090 425.110 2051.270 ;
        RECT 423.930 2048.490 425.110 2049.670 ;
        RECT 423.930 1870.090 425.110 1871.270 ;
        RECT 423.930 1868.490 425.110 1869.670 ;
        RECT 423.930 1690.090 425.110 1691.270 ;
        RECT 423.930 1688.490 425.110 1689.670 ;
        RECT 423.930 1510.090 425.110 1511.270 ;
        RECT 423.930 1508.490 425.110 1509.670 ;
        RECT 423.930 1330.090 425.110 1331.270 ;
        RECT 423.930 1328.490 425.110 1329.670 ;
        RECT 423.930 1150.090 425.110 1151.270 ;
        RECT 423.930 1148.490 425.110 1149.670 ;
        RECT 423.930 970.090 425.110 971.270 ;
        RECT 423.930 968.490 425.110 969.670 ;
        RECT 423.930 790.090 425.110 791.270 ;
        RECT 423.930 788.490 425.110 789.670 ;
        RECT 423.930 610.090 425.110 611.270 ;
        RECT 423.930 608.490 425.110 609.670 ;
        RECT 423.930 430.090 425.110 431.270 ;
        RECT 423.930 428.490 425.110 429.670 ;
        RECT 423.930 250.090 425.110 251.270 ;
        RECT 423.930 248.490 425.110 249.670 ;
        RECT 423.930 70.090 425.110 71.270 ;
        RECT 423.930 68.490 425.110 69.670 ;
        RECT 423.930 -31.110 425.110 -29.930 ;
        RECT 423.930 -32.710 425.110 -31.530 ;
        RECT 603.930 3551.210 605.110 3552.390 ;
        RECT 603.930 3549.610 605.110 3550.790 ;
        RECT 603.930 3490.090 605.110 3491.270 ;
        RECT 603.930 3488.490 605.110 3489.670 ;
        RECT 603.930 3310.090 605.110 3311.270 ;
        RECT 603.930 3308.490 605.110 3309.670 ;
        RECT 603.930 3130.090 605.110 3131.270 ;
        RECT 603.930 3128.490 605.110 3129.670 ;
        RECT 603.930 2950.090 605.110 2951.270 ;
        RECT 603.930 2948.490 605.110 2949.670 ;
        RECT 603.930 2770.090 605.110 2771.270 ;
        RECT 603.930 2768.490 605.110 2769.670 ;
        RECT 603.930 2590.090 605.110 2591.270 ;
        RECT 603.930 2588.490 605.110 2589.670 ;
        RECT 603.930 2410.090 605.110 2411.270 ;
        RECT 603.930 2408.490 605.110 2409.670 ;
        RECT 603.930 2230.090 605.110 2231.270 ;
        RECT 603.930 2228.490 605.110 2229.670 ;
        RECT 603.930 2050.090 605.110 2051.270 ;
        RECT 603.930 2048.490 605.110 2049.670 ;
        RECT 603.930 1870.090 605.110 1871.270 ;
        RECT 603.930 1868.490 605.110 1869.670 ;
        RECT 603.930 1690.090 605.110 1691.270 ;
        RECT 603.930 1688.490 605.110 1689.670 ;
        RECT 603.930 1510.090 605.110 1511.270 ;
        RECT 603.930 1508.490 605.110 1509.670 ;
        RECT 603.930 1330.090 605.110 1331.270 ;
        RECT 603.930 1328.490 605.110 1329.670 ;
        RECT 603.930 1150.090 605.110 1151.270 ;
        RECT 603.930 1148.490 605.110 1149.670 ;
        RECT 603.930 970.090 605.110 971.270 ;
        RECT 603.930 968.490 605.110 969.670 ;
        RECT 603.930 790.090 605.110 791.270 ;
        RECT 603.930 788.490 605.110 789.670 ;
        RECT 603.930 610.090 605.110 611.270 ;
        RECT 603.930 608.490 605.110 609.670 ;
        RECT 603.930 430.090 605.110 431.270 ;
        RECT 603.930 428.490 605.110 429.670 ;
        RECT 603.930 250.090 605.110 251.270 ;
        RECT 603.930 248.490 605.110 249.670 ;
        RECT 603.930 70.090 605.110 71.270 ;
        RECT 603.930 68.490 605.110 69.670 ;
        RECT 603.930 -31.110 605.110 -29.930 ;
        RECT 603.930 -32.710 605.110 -31.530 ;
        RECT 783.930 3551.210 785.110 3552.390 ;
        RECT 783.930 3549.610 785.110 3550.790 ;
        RECT 783.930 3490.090 785.110 3491.270 ;
        RECT 783.930 3488.490 785.110 3489.670 ;
        RECT 783.930 3310.090 785.110 3311.270 ;
        RECT 783.930 3308.490 785.110 3309.670 ;
        RECT 783.930 3130.090 785.110 3131.270 ;
        RECT 783.930 3128.490 785.110 3129.670 ;
        RECT 783.930 2950.090 785.110 2951.270 ;
        RECT 783.930 2948.490 785.110 2949.670 ;
        RECT 783.930 2770.090 785.110 2771.270 ;
        RECT 783.930 2768.490 785.110 2769.670 ;
        RECT 783.930 2590.090 785.110 2591.270 ;
        RECT 783.930 2588.490 785.110 2589.670 ;
        RECT 783.930 2410.090 785.110 2411.270 ;
        RECT 783.930 2408.490 785.110 2409.670 ;
        RECT 783.930 2230.090 785.110 2231.270 ;
        RECT 783.930 2228.490 785.110 2229.670 ;
        RECT 783.930 2050.090 785.110 2051.270 ;
        RECT 783.930 2048.490 785.110 2049.670 ;
        RECT 783.930 1870.090 785.110 1871.270 ;
        RECT 783.930 1868.490 785.110 1869.670 ;
        RECT 783.930 1690.090 785.110 1691.270 ;
        RECT 783.930 1688.490 785.110 1689.670 ;
        RECT 783.930 1510.090 785.110 1511.270 ;
        RECT 783.930 1508.490 785.110 1509.670 ;
        RECT 783.930 1330.090 785.110 1331.270 ;
        RECT 783.930 1328.490 785.110 1329.670 ;
        RECT 783.930 1150.090 785.110 1151.270 ;
        RECT 783.930 1148.490 785.110 1149.670 ;
        RECT 783.930 970.090 785.110 971.270 ;
        RECT 783.930 968.490 785.110 969.670 ;
        RECT 783.930 790.090 785.110 791.270 ;
        RECT 783.930 788.490 785.110 789.670 ;
        RECT 783.930 610.090 785.110 611.270 ;
        RECT 783.930 608.490 785.110 609.670 ;
        RECT 783.930 430.090 785.110 431.270 ;
        RECT 783.930 428.490 785.110 429.670 ;
        RECT 783.930 250.090 785.110 251.270 ;
        RECT 783.930 248.490 785.110 249.670 ;
        RECT 783.930 70.090 785.110 71.270 ;
        RECT 783.930 68.490 785.110 69.670 ;
        RECT 783.930 -31.110 785.110 -29.930 ;
        RECT 783.930 -32.710 785.110 -31.530 ;
        RECT 963.930 3551.210 965.110 3552.390 ;
        RECT 963.930 3549.610 965.110 3550.790 ;
        RECT 963.930 3490.090 965.110 3491.270 ;
        RECT 963.930 3488.490 965.110 3489.670 ;
        RECT 963.930 3310.090 965.110 3311.270 ;
        RECT 963.930 3308.490 965.110 3309.670 ;
        RECT 963.930 3130.090 965.110 3131.270 ;
        RECT 963.930 3128.490 965.110 3129.670 ;
        RECT 963.930 2950.090 965.110 2951.270 ;
        RECT 963.930 2948.490 965.110 2949.670 ;
        RECT 963.930 2770.090 965.110 2771.270 ;
        RECT 963.930 2768.490 965.110 2769.670 ;
        RECT 963.930 2590.090 965.110 2591.270 ;
        RECT 963.930 2588.490 965.110 2589.670 ;
        RECT 963.930 2410.090 965.110 2411.270 ;
        RECT 963.930 2408.490 965.110 2409.670 ;
        RECT 963.930 2230.090 965.110 2231.270 ;
        RECT 963.930 2228.490 965.110 2229.670 ;
        RECT 963.930 2050.090 965.110 2051.270 ;
        RECT 963.930 2048.490 965.110 2049.670 ;
        RECT 963.930 1870.090 965.110 1871.270 ;
        RECT 963.930 1868.490 965.110 1869.670 ;
        RECT 963.930 1690.090 965.110 1691.270 ;
        RECT 963.930 1688.490 965.110 1689.670 ;
        RECT 963.930 1510.090 965.110 1511.270 ;
        RECT 963.930 1508.490 965.110 1509.670 ;
        RECT 963.930 1330.090 965.110 1331.270 ;
        RECT 963.930 1328.490 965.110 1329.670 ;
        RECT 963.930 1150.090 965.110 1151.270 ;
        RECT 963.930 1148.490 965.110 1149.670 ;
        RECT 963.930 970.090 965.110 971.270 ;
        RECT 963.930 968.490 965.110 969.670 ;
        RECT 963.930 790.090 965.110 791.270 ;
        RECT 963.930 788.490 965.110 789.670 ;
        RECT 963.930 610.090 965.110 611.270 ;
        RECT 963.930 608.490 965.110 609.670 ;
        RECT 963.930 430.090 965.110 431.270 ;
        RECT 963.930 428.490 965.110 429.670 ;
        RECT 963.930 250.090 965.110 251.270 ;
        RECT 963.930 248.490 965.110 249.670 ;
        RECT 963.930 70.090 965.110 71.270 ;
        RECT 963.930 68.490 965.110 69.670 ;
        RECT 963.930 -31.110 965.110 -29.930 ;
        RECT 963.930 -32.710 965.110 -31.530 ;
        RECT 1143.930 3551.210 1145.110 3552.390 ;
        RECT 1143.930 3549.610 1145.110 3550.790 ;
        RECT 1143.930 3490.090 1145.110 3491.270 ;
        RECT 1143.930 3488.490 1145.110 3489.670 ;
        RECT 1143.930 3310.090 1145.110 3311.270 ;
        RECT 1143.930 3308.490 1145.110 3309.670 ;
        RECT 1143.930 3130.090 1145.110 3131.270 ;
        RECT 1143.930 3128.490 1145.110 3129.670 ;
        RECT 1143.930 2950.090 1145.110 2951.270 ;
        RECT 1143.930 2948.490 1145.110 2949.670 ;
        RECT 1143.930 2770.090 1145.110 2771.270 ;
        RECT 1143.930 2768.490 1145.110 2769.670 ;
        RECT 1143.930 2590.090 1145.110 2591.270 ;
        RECT 1143.930 2588.490 1145.110 2589.670 ;
        RECT 1143.930 2410.090 1145.110 2411.270 ;
        RECT 1143.930 2408.490 1145.110 2409.670 ;
        RECT 1143.930 2230.090 1145.110 2231.270 ;
        RECT 1143.930 2228.490 1145.110 2229.670 ;
        RECT 1143.930 2050.090 1145.110 2051.270 ;
        RECT 1143.930 2048.490 1145.110 2049.670 ;
        RECT 1143.930 1870.090 1145.110 1871.270 ;
        RECT 1143.930 1868.490 1145.110 1869.670 ;
        RECT 1143.930 1690.090 1145.110 1691.270 ;
        RECT 1143.930 1688.490 1145.110 1689.670 ;
        RECT 1143.930 1510.090 1145.110 1511.270 ;
        RECT 1143.930 1508.490 1145.110 1509.670 ;
        RECT 1143.930 1330.090 1145.110 1331.270 ;
        RECT 1143.930 1328.490 1145.110 1329.670 ;
        RECT 1143.930 1150.090 1145.110 1151.270 ;
        RECT 1143.930 1148.490 1145.110 1149.670 ;
        RECT 1143.930 970.090 1145.110 971.270 ;
        RECT 1143.930 968.490 1145.110 969.670 ;
        RECT 1143.930 790.090 1145.110 791.270 ;
        RECT 1143.930 788.490 1145.110 789.670 ;
        RECT 1143.930 610.090 1145.110 611.270 ;
        RECT 1143.930 608.490 1145.110 609.670 ;
        RECT 1143.930 430.090 1145.110 431.270 ;
        RECT 1143.930 428.490 1145.110 429.670 ;
        RECT 1143.930 250.090 1145.110 251.270 ;
        RECT 1143.930 248.490 1145.110 249.670 ;
        RECT 1143.930 70.090 1145.110 71.270 ;
        RECT 1143.930 68.490 1145.110 69.670 ;
        RECT 1143.930 -31.110 1145.110 -29.930 ;
        RECT 1143.930 -32.710 1145.110 -31.530 ;
        RECT 1323.930 3551.210 1325.110 3552.390 ;
        RECT 1323.930 3549.610 1325.110 3550.790 ;
        RECT 1323.930 3490.090 1325.110 3491.270 ;
        RECT 1323.930 3488.490 1325.110 3489.670 ;
        RECT 1323.930 3310.090 1325.110 3311.270 ;
        RECT 1323.930 3308.490 1325.110 3309.670 ;
        RECT 1323.930 3130.090 1325.110 3131.270 ;
        RECT 1323.930 3128.490 1325.110 3129.670 ;
        RECT 1323.930 2950.090 1325.110 2951.270 ;
        RECT 1323.930 2948.490 1325.110 2949.670 ;
        RECT 1323.930 2770.090 1325.110 2771.270 ;
        RECT 1323.930 2768.490 1325.110 2769.670 ;
        RECT 1323.930 2590.090 1325.110 2591.270 ;
        RECT 1323.930 2588.490 1325.110 2589.670 ;
        RECT 1323.930 2410.090 1325.110 2411.270 ;
        RECT 1323.930 2408.490 1325.110 2409.670 ;
        RECT 1323.930 2230.090 1325.110 2231.270 ;
        RECT 1323.930 2228.490 1325.110 2229.670 ;
        RECT 1323.930 2050.090 1325.110 2051.270 ;
        RECT 1323.930 2048.490 1325.110 2049.670 ;
        RECT 1323.930 1870.090 1325.110 1871.270 ;
        RECT 1323.930 1868.490 1325.110 1869.670 ;
        RECT 1323.930 1690.090 1325.110 1691.270 ;
        RECT 1323.930 1688.490 1325.110 1689.670 ;
        RECT 1323.930 1510.090 1325.110 1511.270 ;
        RECT 1323.930 1508.490 1325.110 1509.670 ;
        RECT 1323.930 1330.090 1325.110 1331.270 ;
        RECT 1323.930 1328.490 1325.110 1329.670 ;
        RECT 1323.930 1150.090 1325.110 1151.270 ;
        RECT 1323.930 1148.490 1325.110 1149.670 ;
        RECT 1323.930 970.090 1325.110 971.270 ;
        RECT 1323.930 968.490 1325.110 969.670 ;
        RECT 1323.930 790.090 1325.110 791.270 ;
        RECT 1323.930 788.490 1325.110 789.670 ;
        RECT 1323.930 610.090 1325.110 611.270 ;
        RECT 1323.930 608.490 1325.110 609.670 ;
        RECT 1323.930 430.090 1325.110 431.270 ;
        RECT 1323.930 428.490 1325.110 429.670 ;
        RECT 1323.930 250.090 1325.110 251.270 ;
        RECT 1323.930 248.490 1325.110 249.670 ;
        RECT 1323.930 70.090 1325.110 71.270 ;
        RECT 1323.930 68.490 1325.110 69.670 ;
        RECT 1323.930 -31.110 1325.110 -29.930 ;
        RECT 1323.930 -32.710 1325.110 -31.530 ;
        RECT 1503.930 3551.210 1505.110 3552.390 ;
        RECT 1503.930 3549.610 1505.110 3550.790 ;
        RECT 1503.930 3490.090 1505.110 3491.270 ;
        RECT 1503.930 3488.490 1505.110 3489.670 ;
        RECT 1503.930 3310.090 1505.110 3311.270 ;
        RECT 1503.930 3308.490 1505.110 3309.670 ;
        RECT 1503.930 3130.090 1505.110 3131.270 ;
        RECT 1503.930 3128.490 1505.110 3129.670 ;
        RECT 1503.930 2950.090 1505.110 2951.270 ;
        RECT 1503.930 2948.490 1505.110 2949.670 ;
        RECT 1503.930 2770.090 1505.110 2771.270 ;
        RECT 1503.930 2768.490 1505.110 2769.670 ;
        RECT 1503.930 2590.090 1505.110 2591.270 ;
        RECT 1503.930 2588.490 1505.110 2589.670 ;
        RECT 1503.930 2410.090 1505.110 2411.270 ;
        RECT 1503.930 2408.490 1505.110 2409.670 ;
        RECT 1503.930 2230.090 1505.110 2231.270 ;
        RECT 1503.930 2228.490 1505.110 2229.670 ;
        RECT 1503.930 2050.090 1505.110 2051.270 ;
        RECT 1503.930 2048.490 1505.110 2049.670 ;
        RECT 1503.930 1870.090 1505.110 1871.270 ;
        RECT 1503.930 1868.490 1505.110 1869.670 ;
        RECT 1503.930 1690.090 1505.110 1691.270 ;
        RECT 1503.930 1688.490 1505.110 1689.670 ;
        RECT 1503.930 1510.090 1505.110 1511.270 ;
        RECT 1503.930 1508.490 1505.110 1509.670 ;
        RECT 1503.930 1330.090 1505.110 1331.270 ;
        RECT 1503.930 1328.490 1505.110 1329.670 ;
        RECT 1503.930 1150.090 1505.110 1151.270 ;
        RECT 1503.930 1148.490 1505.110 1149.670 ;
        RECT 1503.930 970.090 1505.110 971.270 ;
        RECT 1503.930 968.490 1505.110 969.670 ;
        RECT 1503.930 790.090 1505.110 791.270 ;
        RECT 1503.930 788.490 1505.110 789.670 ;
        RECT 1503.930 610.090 1505.110 611.270 ;
        RECT 1503.930 608.490 1505.110 609.670 ;
        RECT 1503.930 430.090 1505.110 431.270 ;
        RECT 1503.930 428.490 1505.110 429.670 ;
        RECT 1503.930 250.090 1505.110 251.270 ;
        RECT 1503.930 248.490 1505.110 249.670 ;
        RECT 1503.930 70.090 1505.110 71.270 ;
        RECT 1503.930 68.490 1505.110 69.670 ;
        RECT 1503.930 -31.110 1505.110 -29.930 ;
        RECT 1503.930 -32.710 1505.110 -31.530 ;
        RECT 1683.930 3551.210 1685.110 3552.390 ;
        RECT 1683.930 3549.610 1685.110 3550.790 ;
        RECT 1683.930 3490.090 1685.110 3491.270 ;
        RECT 1683.930 3488.490 1685.110 3489.670 ;
        RECT 1683.930 3310.090 1685.110 3311.270 ;
        RECT 1683.930 3308.490 1685.110 3309.670 ;
        RECT 1683.930 3130.090 1685.110 3131.270 ;
        RECT 1683.930 3128.490 1685.110 3129.670 ;
        RECT 1683.930 2950.090 1685.110 2951.270 ;
        RECT 1683.930 2948.490 1685.110 2949.670 ;
        RECT 1683.930 2770.090 1685.110 2771.270 ;
        RECT 1683.930 2768.490 1685.110 2769.670 ;
        RECT 1683.930 2590.090 1685.110 2591.270 ;
        RECT 1683.930 2588.490 1685.110 2589.670 ;
        RECT 1683.930 2410.090 1685.110 2411.270 ;
        RECT 1683.930 2408.490 1685.110 2409.670 ;
        RECT 1683.930 2230.090 1685.110 2231.270 ;
        RECT 1683.930 2228.490 1685.110 2229.670 ;
        RECT 1683.930 2050.090 1685.110 2051.270 ;
        RECT 1683.930 2048.490 1685.110 2049.670 ;
        RECT 1683.930 1870.090 1685.110 1871.270 ;
        RECT 1683.930 1868.490 1685.110 1869.670 ;
        RECT 1683.930 1690.090 1685.110 1691.270 ;
        RECT 1683.930 1688.490 1685.110 1689.670 ;
        RECT 1683.930 1510.090 1685.110 1511.270 ;
        RECT 1683.930 1508.490 1685.110 1509.670 ;
        RECT 1683.930 1330.090 1685.110 1331.270 ;
        RECT 1683.930 1328.490 1685.110 1329.670 ;
        RECT 1683.930 1150.090 1685.110 1151.270 ;
        RECT 1683.930 1148.490 1685.110 1149.670 ;
        RECT 1683.930 970.090 1685.110 971.270 ;
        RECT 1683.930 968.490 1685.110 969.670 ;
        RECT 1683.930 790.090 1685.110 791.270 ;
        RECT 1683.930 788.490 1685.110 789.670 ;
        RECT 1683.930 610.090 1685.110 611.270 ;
        RECT 1683.930 608.490 1685.110 609.670 ;
        RECT 1683.930 430.090 1685.110 431.270 ;
        RECT 1683.930 428.490 1685.110 429.670 ;
        RECT 1683.930 250.090 1685.110 251.270 ;
        RECT 1683.930 248.490 1685.110 249.670 ;
        RECT 1683.930 70.090 1685.110 71.270 ;
        RECT 1683.930 68.490 1685.110 69.670 ;
        RECT 1683.930 -31.110 1685.110 -29.930 ;
        RECT 1683.930 -32.710 1685.110 -31.530 ;
        RECT 1863.930 3551.210 1865.110 3552.390 ;
        RECT 1863.930 3549.610 1865.110 3550.790 ;
        RECT 1863.930 3490.090 1865.110 3491.270 ;
        RECT 1863.930 3488.490 1865.110 3489.670 ;
        RECT 1863.930 3310.090 1865.110 3311.270 ;
        RECT 1863.930 3308.490 1865.110 3309.670 ;
        RECT 1863.930 3130.090 1865.110 3131.270 ;
        RECT 1863.930 3128.490 1865.110 3129.670 ;
        RECT 1863.930 2950.090 1865.110 2951.270 ;
        RECT 1863.930 2948.490 1865.110 2949.670 ;
        RECT 1863.930 2770.090 1865.110 2771.270 ;
        RECT 1863.930 2768.490 1865.110 2769.670 ;
        RECT 1863.930 2590.090 1865.110 2591.270 ;
        RECT 1863.930 2588.490 1865.110 2589.670 ;
        RECT 1863.930 2410.090 1865.110 2411.270 ;
        RECT 1863.930 2408.490 1865.110 2409.670 ;
        RECT 1863.930 2230.090 1865.110 2231.270 ;
        RECT 1863.930 2228.490 1865.110 2229.670 ;
        RECT 1863.930 2050.090 1865.110 2051.270 ;
        RECT 1863.930 2048.490 1865.110 2049.670 ;
        RECT 1863.930 1870.090 1865.110 1871.270 ;
        RECT 1863.930 1868.490 1865.110 1869.670 ;
        RECT 1863.930 1690.090 1865.110 1691.270 ;
        RECT 1863.930 1688.490 1865.110 1689.670 ;
        RECT 1863.930 1510.090 1865.110 1511.270 ;
        RECT 1863.930 1508.490 1865.110 1509.670 ;
        RECT 1863.930 1330.090 1865.110 1331.270 ;
        RECT 1863.930 1328.490 1865.110 1329.670 ;
        RECT 1863.930 1150.090 1865.110 1151.270 ;
        RECT 1863.930 1148.490 1865.110 1149.670 ;
        RECT 1863.930 970.090 1865.110 971.270 ;
        RECT 1863.930 968.490 1865.110 969.670 ;
        RECT 1863.930 790.090 1865.110 791.270 ;
        RECT 1863.930 788.490 1865.110 789.670 ;
        RECT 1863.930 610.090 1865.110 611.270 ;
        RECT 1863.930 608.490 1865.110 609.670 ;
        RECT 1863.930 430.090 1865.110 431.270 ;
        RECT 1863.930 428.490 1865.110 429.670 ;
        RECT 1863.930 250.090 1865.110 251.270 ;
        RECT 1863.930 248.490 1865.110 249.670 ;
        RECT 1863.930 70.090 1865.110 71.270 ;
        RECT 1863.930 68.490 1865.110 69.670 ;
        RECT 1863.930 -31.110 1865.110 -29.930 ;
        RECT 1863.930 -32.710 1865.110 -31.530 ;
        RECT 2043.930 3551.210 2045.110 3552.390 ;
        RECT 2043.930 3549.610 2045.110 3550.790 ;
        RECT 2043.930 3490.090 2045.110 3491.270 ;
        RECT 2043.930 3488.490 2045.110 3489.670 ;
        RECT 2043.930 3310.090 2045.110 3311.270 ;
        RECT 2043.930 3308.490 2045.110 3309.670 ;
        RECT 2043.930 3130.090 2045.110 3131.270 ;
        RECT 2043.930 3128.490 2045.110 3129.670 ;
        RECT 2043.930 2950.090 2045.110 2951.270 ;
        RECT 2043.930 2948.490 2045.110 2949.670 ;
        RECT 2043.930 2770.090 2045.110 2771.270 ;
        RECT 2043.930 2768.490 2045.110 2769.670 ;
        RECT 2043.930 2590.090 2045.110 2591.270 ;
        RECT 2043.930 2588.490 2045.110 2589.670 ;
        RECT 2043.930 2410.090 2045.110 2411.270 ;
        RECT 2043.930 2408.490 2045.110 2409.670 ;
        RECT 2043.930 2230.090 2045.110 2231.270 ;
        RECT 2043.930 2228.490 2045.110 2229.670 ;
        RECT 2043.930 2050.090 2045.110 2051.270 ;
        RECT 2043.930 2048.490 2045.110 2049.670 ;
        RECT 2043.930 1870.090 2045.110 1871.270 ;
        RECT 2043.930 1868.490 2045.110 1869.670 ;
        RECT 2043.930 1690.090 2045.110 1691.270 ;
        RECT 2043.930 1688.490 2045.110 1689.670 ;
        RECT 2043.930 1510.090 2045.110 1511.270 ;
        RECT 2043.930 1508.490 2045.110 1509.670 ;
        RECT 2043.930 1330.090 2045.110 1331.270 ;
        RECT 2043.930 1328.490 2045.110 1329.670 ;
        RECT 2043.930 1150.090 2045.110 1151.270 ;
        RECT 2043.930 1148.490 2045.110 1149.670 ;
        RECT 2043.930 970.090 2045.110 971.270 ;
        RECT 2043.930 968.490 2045.110 969.670 ;
        RECT 2043.930 790.090 2045.110 791.270 ;
        RECT 2043.930 788.490 2045.110 789.670 ;
        RECT 2043.930 610.090 2045.110 611.270 ;
        RECT 2043.930 608.490 2045.110 609.670 ;
        RECT 2043.930 430.090 2045.110 431.270 ;
        RECT 2043.930 428.490 2045.110 429.670 ;
        RECT 2043.930 250.090 2045.110 251.270 ;
        RECT 2043.930 248.490 2045.110 249.670 ;
        RECT 2043.930 70.090 2045.110 71.270 ;
        RECT 2043.930 68.490 2045.110 69.670 ;
        RECT 2043.930 -31.110 2045.110 -29.930 ;
        RECT 2043.930 -32.710 2045.110 -31.530 ;
        RECT 2223.930 3551.210 2225.110 3552.390 ;
        RECT 2223.930 3549.610 2225.110 3550.790 ;
        RECT 2223.930 3490.090 2225.110 3491.270 ;
        RECT 2223.930 3488.490 2225.110 3489.670 ;
        RECT 2223.930 3310.090 2225.110 3311.270 ;
        RECT 2223.930 3308.490 2225.110 3309.670 ;
        RECT 2223.930 3130.090 2225.110 3131.270 ;
        RECT 2223.930 3128.490 2225.110 3129.670 ;
        RECT 2223.930 2950.090 2225.110 2951.270 ;
        RECT 2223.930 2948.490 2225.110 2949.670 ;
        RECT 2223.930 2770.090 2225.110 2771.270 ;
        RECT 2223.930 2768.490 2225.110 2769.670 ;
        RECT 2223.930 2590.090 2225.110 2591.270 ;
        RECT 2223.930 2588.490 2225.110 2589.670 ;
        RECT 2223.930 2410.090 2225.110 2411.270 ;
        RECT 2223.930 2408.490 2225.110 2409.670 ;
        RECT 2223.930 2230.090 2225.110 2231.270 ;
        RECT 2223.930 2228.490 2225.110 2229.670 ;
        RECT 2223.930 2050.090 2225.110 2051.270 ;
        RECT 2223.930 2048.490 2225.110 2049.670 ;
        RECT 2223.930 1870.090 2225.110 1871.270 ;
        RECT 2223.930 1868.490 2225.110 1869.670 ;
        RECT 2223.930 1690.090 2225.110 1691.270 ;
        RECT 2223.930 1688.490 2225.110 1689.670 ;
        RECT 2223.930 1510.090 2225.110 1511.270 ;
        RECT 2223.930 1508.490 2225.110 1509.670 ;
        RECT 2223.930 1330.090 2225.110 1331.270 ;
        RECT 2223.930 1328.490 2225.110 1329.670 ;
        RECT 2223.930 1150.090 2225.110 1151.270 ;
        RECT 2223.930 1148.490 2225.110 1149.670 ;
        RECT 2223.930 970.090 2225.110 971.270 ;
        RECT 2223.930 968.490 2225.110 969.670 ;
        RECT 2223.930 790.090 2225.110 791.270 ;
        RECT 2223.930 788.490 2225.110 789.670 ;
        RECT 2223.930 610.090 2225.110 611.270 ;
        RECT 2223.930 608.490 2225.110 609.670 ;
        RECT 2223.930 430.090 2225.110 431.270 ;
        RECT 2223.930 428.490 2225.110 429.670 ;
        RECT 2223.930 250.090 2225.110 251.270 ;
        RECT 2223.930 248.490 2225.110 249.670 ;
        RECT 2223.930 70.090 2225.110 71.270 ;
        RECT 2223.930 68.490 2225.110 69.670 ;
        RECT 2223.930 -31.110 2225.110 -29.930 ;
        RECT 2223.930 -32.710 2225.110 -31.530 ;
        RECT 2403.930 3551.210 2405.110 3552.390 ;
        RECT 2403.930 3549.610 2405.110 3550.790 ;
        RECT 2403.930 3490.090 2405.110 3491.270 ;
        RECT 2403.930 3488.490 2405.110 3489.670 ;
        RECT 2403.930 3310.090 2405.110 3311.270 ;
        RECT 2403.930 3308.490 2405.110 3309.670 ;
        RECT 2403.930 3130.090 2405.110 3131.270 ;
        RECT 2403.930 3128.490 2405.110 3129.670 ;
        RECT 2403.930 2950.090 2405.110 2951.270 ;
        RECT 2403.930 2948.490 2405.110 2949.670 ;
        RECT 2403.930 2770.090 2405.110 2771.270 ;
        RECT 2403.930 2768.490 2405.110 2769.670 ;
        RECT 2403.930 2590.090 2405.110 2591.270 ;
        RECT 2403.930 2588.490 2405.110 2589.670 ;
        RECT 2403.930 2410.090 2405.110 2411.270 ;
        RECT 2403.930 2408.490 2405.110 2409.670 ;
        RECT 2403.930 2230.090 2405.110 2231.270 ;
        RECT 2403.930 2228.490 2405.110 2229.670 ;
        RECT 2403.930 2050.090 2405.110 2051.270 ;
        RECT 2403.930 2048.490 2405.110 2049.670 ;
        RECT 2403.930 1870.090 2405.110 1871.270 ;
        RECT 2403.930 1868.490 2405.110 1869.670 ;
        RECT 2403.930 1690.090 2405.110 1691.270 ;
        RECT 2403.930 1688.490 2405.110 1689.670 ;
        RECT 2403.930 1510.090 2405.110 1511.270 ;
        RECT 2403.930 1508.490 2405.110 1509.670 ;
        RECT 2403.930 1330.090 2405.110 1331.270 ;
        RECT 2403.930 1328.490 2405.110 1329.670 ;
        RECT 2403.930 1150.090 2405.110 1151.270 ;
        RECT 2403.930 1148.490 2405.110 1149.670 ;
        RECT 2403.930 970.090 2405.110 971.270 ;
        RECT 2403.930 968.490 2405.110 969.670 ;
        RECT 2403.930 790.090 2405.110 791.270 ;
        RECT 2403.930 788.490 2405.110 789.670 ;
        RECT 2403.930 610.090 2405.110 611.270 ;
        RECT 2403.930 608.490 2405.110 609.670 ;
        RECT 2403.930 430.090 2405.110 431.270 ;
        RECT 2403.930 428.490 2405.110 429.670 ;
        RECT 2403.930 250.090 2405.110 251.270 ;
        RECT 2403.930 248.490 2405.110 249.670 ;
        RECT 2403.930 70.090 2405.110 71.270 ;
        RECT 2403.930 68.490 2405.110 69.670 ;
        RECT 2403.930 -31.110 2405.110 -29.930 ;
        RECT 2403.930 -32.710 2405.110 -31.530 ;
        RECT 2583.930 3551.210 2585.110 3552.390 ;
        RECT 2583.930 3549.610 2585.110 3550.790 ;
        RECT 2583.930 3490.090 2585.110 3491.270 ;
        RECT 2583.930 3488.490 2585.110 3489.670 ;
        RECT 2583.930 3310.090 2585.110 3311.270 ;
        RECT 2583.930 3308.490 2585.110 3309.670 ;
        RECT 2583.930 3130.090 2585.110 3131.270 ;
        RECT 2583.930 3128.490 2585.110 3129.670 ;
        RECT 2583.930 2950.090 2585.110 2951.270 ;
        RECT 2583.930 2948.490 2585.110 2949.670 ;
        RECT 2583.930 2770.090 2585.110 2771.270 ;
        RECT 2583.930 2768.490 2585.110 2769.670 ;
        RECT 2583.930 2590.090 2585.110 2591.270 ;
        RECT 2583.930 2588.490 2585.110 2589.670 ;
        RECT 2583.930 2410.090 2585.110 2411.270 ;
        RECT 2583.930 2408.490 2585.110 2409.670 ;
        RECT 2583.930 2230.090 2585.110 2231.270 ;
        RECT 2583.930 2228.490 2585.110 2229.670 ;
        RECT 2583.930 2050.090 2585.110 2051.270 ;
        RECT 2583.930 2048.490 2585.110 2049.670 ;
        RECT 2583.930 1870.090 2585.110 1871.270 ;
        RECT 2583.930 1868.490 2585.110 1869.670 ;
        RECT 2583.930 1690.090 2585.110 1691.270 ;
        RECT 2583.930 1688.490 2585.110 1689.670 ;
        RECT 2583.930 1510.090 2585.110 1511.270 ;
        RECT 2583.930 1508.490 2585.110 1509.670 ;
        RECT 2583.930 1330.090 2585.110 1331.270 ;
        RECT 2583.930 1328.490 2585.110 1329.670 ;
        RECT 2583.930 1150.090 2585.110 1151.270 ;
        RECT 2583.930 1148.490 2585.110 1149.670 ;
        RECT 2583.930 970.090 2585.110 971.270 ;
        RECT 2583.930 968.490 2585.110 969.670 ;
        RECT 2583.930 790.090 2585.110 791.270 ;
        RECT 2583.930 788.490 2585.110 789.670 ;
        RECT 2583.930 610.090 2585.110 611.270 ;
        RECT 2583.930 608.490 2585.110 609.670 ;
        RECT 2583.930 430.090 2585.110 431.270 ;
        RECT 2583.930 428.490 2585.110 429.670 ;
        RECT 2583.930 250.090 2585.110 251.270 ;
        RECT 2583.930 248.490 2585.110 249.670 ;
        RECT 2583.930 70.090 2585.110 71.270 ;
        RECT 2583.930 68.490 2585.110 69.670 ;
        RECT 2583.930 -31.110 2585.110 -29.930 ;
        RECT 2583.930 -32.710 2585.110 -31.530 ;
        RECT 2763.930 3551.210 2765.110 3552.390 ;
        RECT 2763.930 3549.610 2765.110 3550.790 ;
        RECT 2763.930 3490.090 2765.110 3491.270 ;
        RECT 2763.930 3488.490 2765.110 3489.670 ;
        RECT 2763.930 3310.090 2765.110 3311.270 ;
        RECT 2763.930 3308.490 2765.110 3309.670 ;
        RECT 2763.930 3130.090 2765.110 3131.270 ;
        RECT 2763.930 3128.490 2765.110 3129.670 ;
        RECT 2763.930 2950.090 2765.110 2951.270 ;
        RECT 2763.930 2948.490 2765.110 2949.670 ;
        RECT 2763.930 2770.090 2765.110 2771.270 ;
        RECT 2763.930 2768.490 2765.110 2769.670 ;
        RECT 2763.930 2590.090 2765.110 2591.270 ;
        RECT 2763.930 2588.490 2765.110 2589.670 ;
        RECT 2763.930 2410.090 2765.110 2411.270 ;
        RECT 2763.930 2408.490 2765.110 2409.670 ;
        RECT 2763.930 2230.090 2765.110 2231.270 ;
        RECT 2763.930 2228.490 2765.110 2229.670 ;
        RECT 2763.930 2050.090 2765.110 2051.270 ;
        RECT 2763.930 2048.490 2765.110 2049.670 ;
        RECT 2763.930 1870.090 2765.110 1871.270 ;
        RECT 2763.930 1868.490 2765.110 1869.670 ;
        RECT 2763.930 1690.090 2765.110 1691.270 ;
        RECT 2763.930 1688.490 2765.110 1689.670 ;
        RECT 2763.930 1510.090 2765.110 1511.270 ;
        RECT 2763.930 1508.490 2765.110 1509.670 ;
        RECT 2763.930 1330.090 2765.110 1331.270 ;
        RECT 2763.930 1328.490 2765.110 1329.670 ;
        RECT 2763.930 1150.090 2765.110 1151.270 ;
        RECT 2763.930 1148.490 2765.110 1149.670 ;
        RECT 2763.930 970.090 2765.110 971.270 ;
        RECT 2763.930 968.490 2765.110 969.670 ;
        RECT 2763.930 790.090 2765.110 791.270 ;
        RECT 2763.930 788.490 2765.110 789.670 ;
        RECT 2763.930 610.090 2765.110 611.270 ;
        RECT 2763.930 608.490 2765.110 609.670 ;
        RECT 2763.930 430.090 2765.110 431.270 ;
        RECT 2763.930 428.490 2765.110 429.670 ;
        RECT 2763.930 250.090 2765.110 251.270 ;
        RECT 2763.930 248.490 2765.110 249.670 ;
        RECT 2763.930 70.090 2765.110 71.270 ;
        RECT 2763.930 68.490 2765.110 69.670 ;
        RECT 2763.930 -31.110 2765.110 -29.930 ;
        RECT 2763.930 -32.710 2765.110 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 3490.090 2956.890 3491.270 ;
        RECT 2955.710 3488.490 2956.890 3489.670 ;
        RECT 2955.710 3310.090 2956.890 3311.270 ;
        RECT 2955.710 3308.490 2956.890 3309.670 ;
        RECT 2955.710 3130.090 2956.890 3131.270 ;
        RECT 2955.710 3128.490 2956.890 3129.670 ;
        RECT 2955.710 2950.090 2956.890 2951.270 ;
        RECT 2955.710 2948.490 2956.890 2949.670 ;
        RECT 2955.710 2770.090 2956.890 2771.270 ;
        RECT 2955.710 2768.490 2956.890 2769.670 ;
        RECT 2955.710 2590.090 2956.890 2591.270 ;
        RECT 2955.710 2588.490 2956.890 2589.670 ;
        RECT 2955.710 2410.090 2956.890 2411.270 ;
        RECT 2955.710 2408.490 2956.890 2409.670 ;
        RECT 2955.710 2230.090 2956.890 2231.270 ;
        RECT 2955.710 2228.490 2956.890 2229.670 ;
        RECT 2955.710 2050.090 2956.890 2051.270 ;
        RECT 2955.710 2048.490 2956.890 2049.670 ;
        RECT 2955.710 1870.090 2956.890 1871.270 ;
        RECT 2955.710 1868.490 2956.890 1869.670 ;
        RECT 2955.710 1690.090 2956.890 1691.270 ;
        RECT 2955.710 1688.490 2956.890 1689.670 ;
        RECT 2955.710 1510.090 2956.890 1511.270 ;
        RECT 2955.710 1508.490 2956.890 1509.670 ;
        RECT 2955.710 1330.090 2956.890 1331.270 ;
        RECT 2955.710 1328.490 2956.890 1329.670 ;
        RECT 2955.710 1150.090 2956.890 1151.270 ;
        RECT 2955.710 1148.490 2956.890 1149.670 ;
        RECT 2955.710 970.090 2956.890 971.270 ;
        RECT 2955.710 968.490 2956.890 969.670 ;
        RECT 2955.710 790.090 2956.890 791.270 ;
        RECT 2955.710 788.490 2956.890 789.670 ;
        RECT 2955.710 610.090 2956.890 611.270 ;
        RECT 2955.710 608.490 2956.890 609.670 ;
        RECT 2955.710 430.090 2956.890 431.270 ;
        RECT 2955.710 428.490 2956.890 429.670 ;
        RECT 2955.710 250.090 2956.890 251.270 ;
        RECT 2955.710 248.490 2956.890 249.670 ;
        RECT 2955.710 70.090 2956.890 71.270 ;
        RECT 2955.710 68.490 2956.890 69.670 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 63.020 3552.500 66.020 3552.510 ;
        RECT 243.020 3552.500 246.020 3552.510 ;
        RECT 423.020 3552.500 426.020 3552.510 ;
        RECT 603.020 3552.500 606.020 3552.510 ;
        RECT 783.020 3552.500 786.020 3552.510 ;
        RECT 963.020 3552.500 966.020 3552.510 ;
        RECT 1143.020 3552.500 1146.020 3552.510 ;
        RECT 1323.020 3552.500 1326.020 3552.510 ;
        RECT 1503.020 3552.500 1506.020 3552.510 ;
        RECT 1683.020 3552.500 1686.020 3552.510 ;
        RECT 1863.020 3552.500 1866.020 3552.510 ;
        RECT 2043.020 3552.500 2046.020 3552.510 ;
        RECT 2223.020 3552.500 2226.020 3552.510 ;
        RECT 2403.020 3552.500 2406.020 3552.510 ;
        RECT 2583.020 3552.500 2586.020 3552.510 ;
        RECT 2763.020 3552.500 2766.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 63.020 3549.490 66.020 3549.500 ;
        RECT 243.020 3549.490 246.020 3549.500 ;
        RECT 423.020 3549.490 426.020 3549.500 ;
        RECT 603.020 3549.490 606.020 3549.500 ;
        RECT 783.020 3549.490 786.020 3549.500 ;
        RECT 963.020 3549.490 966.020 3549.500 ;
        RECT 1143.020 3549.490 1146.020 3549.500 ;
        RECT 1323.020 3549.490 1326.020 3549.500 ;
        RECT 1503.020 3549.490 1506.020 3549.500 ;
        RECT 1683.020 3549.490 1686.020 3549.500 ;
        RECT 1863.020 3549.490 1866.020 3549.500 ;
        RECT 2043.020 3549.490 2046.020 3549.500 ;
        RECT 2223.020 3549.490 2226.020 3549.500 ;
        RECT 2403.020 3549.490 2406.020 3549.500 ;
        RECT 2583.020 3549.490 2586.020 3549.500 ;
        RECT 2763.020 3549.490 2766.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3491.380 -35.180 3491.390 ;
        RECT 63.020 3491.380 66.020 3491.390 ;
        RECT 243.020 3491.380 246.020 3491.390 ;
        RECT 423.020 3491.380 426.020 3491.390 ;
        RECT 603.020 3491.380 606.020 3491.390 ;
        RECT 783.020 3491.380 786.020 3491.390 ;
        RECT 963.020 3491.380 966.020 3491.390 ;
        RECT 1143.020 3491.380 1146.020 3491.390 ;
        RECT 1323.020 3491.380 1326.020 3491.390 ;
        RECT 1503.020 3491.380 1506.020 3491.390 ;
        RECT 1683.020 3491.380 1686.020 3491.390 ;
        RECT 1863.020 3491.380 1866.020 3491.390 ;
        RECT 2043.020 3491.380 2046.020 3491.390 ;
        RECT 2223.020 3491.380 2226.020 3491.390 ;
        RECT 2403.020 3491.380 2406.020 3491.390 ;
        RECT 2583.020 3491.380 2586.020 3491.390 ;
        RECT 2763.020 3491.380 2766.020 3491.390 ;
        RECT 2954.800 3491.380 2957.800 3491.390 ;
        RECT -42.880 3488.380 2962.500 3491.380 ;
        RECT -38.180 3488.370 -35.180 3488.380 ;
        RECT 63.020 3488.370 66.020 3488.380 ;
        RECT 243.020 3488.370 246.020 3488.380 ;
        RECT 423.020 3488.370 426.020 3488.380 ;
        RECT 603.020 3488.370 606.020 3488.380 ;
        RECT 783.020 3488.370 786.020 3488.380 ;
        RECT 963.020 3488.370 966.020 3488.380 ;
        RECT 1143.020 3488.370 1146.020 3488.380 ;
        RECT 1323.020 3488.370 1326.020 3488.380 ;
        RECT 1503.020 3488.370 1506.020 3488.380 ;
        RECT 1683.020 3488.370 1686.020 3488.380 ;
        RECT 1863.020 3488.370 1866.020 3488.380 ;
        RECT 2043.020 3488.370 2046.020 3488.380 ;
        RECT 2223.020 3488.370 2226.020 3488.380 ;
        RECT 2403.020 3488.370 2406.020 3488.380 ;
        RECT 2583.020 3488.370 2586.020 3488.380 ;
        RECT 2763.020 3488.370 2766.020 3488.380 ;
        RECT 2954.800 3488.370 2957.800 3488.380 ;
        RECT -38.180 3311.380 -35.180 3311.390 ;
        RECT 63.020 3311.380 66.020 3311.390 ;
        RECT 243.020 3311.380 246.020 3311.390 ;
        RECT 423.020 3311.380 426.020 3311.390 ;
        RECT 603.020 3311.380 606.020 3311.390 ;
        RECT 783.020 3311.380 786.020 3311.390 ;
        RECT 963.020 3311.380 966.020 3311.390 ;
        RECT 1143.020 3311.380 1146.020 3311.390 ;
        RECT 1323.020 3311.380 1326.020 3311.390 ;
        RECT 1503.020 3311.380 1506.020 3311.390 ;
        RECT 1683.020 3311.380 1686.020 3311.390 ;
        RECT 1863.020 3311.380 1866.020 3311.390 ;
        RECT 2043.020 3311.380 2046.020 3311.390 ;
        RECT 2223.020 3311.380 2226.020 3311.390 ;
        RECT 2403.020 3311.380 2406.020 3311.390 ;
        RECT 2583.020 3311.380 2586.020 3311.390 ;
        RECT 2763.020 3311.380 2766.020 3311.390 ;
        RECT 2954.800 3311.380 2957.800 3311.390 ;
        RECT -42.880 3308.380 2962.500 3311.380 ;
        RECT -38.180 3308.370 -35.180 3308.380 ;
        RECT 63.020 3308.370 66.020 3308.380 ;
        RECT 243.020 3308.370 246.020 3308.380 ;
        RECT 423.020 3308.370 426.020 3308.380 ;
        RECT 603.020 3308.370 606.020 3308.380 ;
        RECT 783.020 3308.370 786.020 3308.380 ;
        RECT 963.020 3308.370 966.020 3308.380 ;
        RECT 1143.020 3308.370 1146.020 3308.380 ;
        RECT 1323.020 3308.370 1326.020 3308.380 ;
        RECT 1503.020 3308.370 1506.020 3308.380 ;
        RECT 1683.020 3308.370 1686.020 3308.380 ;
        RECT 1863.020 3308.370 1866.020 3308.380 ;
        RECT 2043.020 3308.370 2046.020 3308.380 ;
        RECT 2223.020 3308.370 2226.020 3308.380 ;
        RECT 2403.020 3308.370 2406.020 3308.380 ;
        RECT 2583.020 3308.370 2586.020 3308.380 ;
        RECT 2763.020 3308.370 2766.020 3308.380 ;
        RECT 2954.800 3308.370 2957.800 3308.380 ;
        RECT -38.180 3131.380 -35.180 3131.390 ;
        RECT 63.020 3131.380 66.020 3131.390 ;
        RECT 243.020 3131.380 246.020 3131.390 ;
        RECT 423.020 3131.380 426.020 3131.390 ;
        RECT 603.020 3131.380 606.020 3131.390 ;
        RECT 783.020 3131.380 786.020 3131.390 ;
        RECT 963.020 3131.380 966.020 3131.390 ;
        RECT 1143.020 3131.380 1146.020 3131.390 ;
        RECT 1323.020 3131.380 1326.020 3131.390 ;
        RECT 1503.020 3131.380 1506.020 3131.390 ;
        RECT 1683.020 3131.380 1686.020 3131.390 ;
        RECT 1863.020 3131.380 1866.020 3131.390 ;
        RECT 2043.020 3131.380 2046.020 3131.390 ;
        RECT 2223.020 3131.380 2226.020 3131.390 ;
        RECT 2403.020 3131.380 2406.020 3131.390 ;
        RECT 2583.020 3131.380 2586.020 3131.390 ;
        RECT 2763.020 3131.380 2766.020 3131.390 ;
        RECT 2954.800 3131.380 2957.800 3131.390 ;
        RECT -42.880 3128.380 2962.500 3131.380 ;
        RECT -38.180 3128.370 -35.180 3128.380 ;
        RECT 63.020 3128.370 66.020 3128.380 ;
        RECT 243.020 3128.370 246.020 3128.380 ;
        RECT 423.020 3128.370 426.020 3128.380 ;
        RECT 603.020 3128.370 606.020 3128.380 ;
        RECT 783.020 3128.370 786.020 3128.380 ;
        RECT 963.020 3128.370 966.020 3128.380 ;
        RECT 1143.020 3128.370 1146.020 3128.380 ;
        RECT 1323.020 3128.370 1326.020 3128.380 ;
        RECT 1503.020 3128.370 1506.020 3128.380 ;
        RECT 1683.020 3128.370 1686.020 3128.380 ;
        RECT 1863.020 3128.370 1866.020 3128.380 ;
        RECT 2043.020 3128.370 2046.020 3128.380 ;
        RECT 2223.020 3128.370 2226.020 3128.380 ;
        RECT 2403.020 3128.370 2406.020 3128.380 ;
        RECT 2583.020 3128.370 2586.020 3128.380 ;
        RECT 2763.020 3128.370 2766.020 3128.380 ;
        RECT 2954.800 3128.370 2957.800 3128.380 ;
        RECT -38.180 2951.380 -35.180 2951.390 ;
        RECT 63.020 2951.380 66.020 2951.390 ;
        RECT 243.020 2951.380 246.020 2951.390 ;
        RECT 423.020 2951.380 426.020 2951.390 ;
        RECT 603.020 2951.380 606.020 2951.390 ;
        RECT 783.020 2951.380 786.020 2951.390 ;
        RECT 963.020 2951.380 966.020 2951.390 ;
        RECT 1143.020 2951.380 1146.020 2951.390 ;
        RECT 1323.020 2951.380 1326.020 2951.390 ;
        RECT 1503.020 2951.380 1506.020 2951.390 ;
        RECT 1683.020 2951.380 1686.020 2951.390 ;
        RECT 1863.020 2951.380 1866.020 2951.390 ;
        RECT 2043.020 2951.380 2046.020 2951.390 ;
        RECT 2223.020 2951.380 2226.020 2951.390 ;
        RECT 2403.020 2951.380 2406.020 2951.390 ;
        RECT 2583.020 2951.380 2586.020 2951.390 ;
        RECT 2763.020 2951.380 2766.020 2951.390 ;
        RECT 2954.800 2951.380 2957.800 2951.390 ;
        RECT -42.880 2948.380 2962.500 2951.380 ;
        RECT -38.180 2948.370 -35.180 2948.380 ;
        RECT 63.020 2948.370 66.020 2948.380 ;
        RECT 243.020 2948.370 246.020 2948.380 ;
        RECT 423.020 2948.370 426.020 2948.380 ;
        RECT 603.020 2948.370 606.020 2948.380 ;
        RECT 783.020 2948.370 786.020 2948.380 ;
        RECT 963.020 2948.370 966.020 2948.380 ;
        RECT 1143.020 2948.370 1146.020 2948.380 ;
        RECT 1323.020 2948.370 1326.020 2948.380 ;
        RECT 1503.020 2948.370 1506.020 2948.380 ;
        RECT 1683.020 2948.370 1686.020 2948.380 ;
        RECT 1863.020 2948.370 1866.020 2948.380 ;
        RECT 2043.020 2948.370 2046.020 2948.380 ;
        RECT 2223.020 2948.370 2226.020 2948.380 ;
        RECT 2403.020 2948.370 2406.020 2948.380 ;
        RECT 2583.020 2948.370 2586.020 2948.380 ;
        RECT 2763.020 2948.370 2766.020 2948.380 ;
        RECT 2954.800 2948.370 2957.800 2948.380 ;
        RECT -38.180 2771.380 -35.180 2771.390 ;
        RECT 63.020 2771.380 66.020 2771.390 ;
        RECT 243.020 2771.380 246.020 2771.390 ;
        RECT 423.020 2771.380 426.020 2771.390 ;
        RECT 603.020 2771.380 606.020 2771.390 ;
        RECT 783.020 2771.380 786.020 2771.390 ;
        RECT 963.020 2771.380 966.020 2771.390 ;
        RECT 1143.020 2771.380 1146.020 2771.390 ;
        RECT 1323.020 2771.380 1326.020 2771.390 ;
        RECT 1503.020 2771.380 1506.020 2771.390 ;
        RECT 1683.020 2771.380 1686.020 2771.390 ;
        RECT 1863.020 2771.380 1866.020 2771.390 ;
        RECT 2043.020 2771.380 2046.020 2771.390 ;
        RECT 2223.020 2771.380 2226.020 2771.390 ;
        RECT 2403.020 2771.380 2406.020 2771.390 ;
        RECT 2583.020 2771.380 2586.020 2771.390 ;
        RECT 2763.020 2771.380 2766.020 2771.390 ;
        RECT 2954.800 2771.380 2957.800 2771.390 ;
        RECT -42.880 2768.380 2962.500 2771.380 ;
        RECT -38.180 2768.370 -35.180 2768.380 ;
        RECT 63.020 2768.370 66.020 2768.380 ;
        RECT 243.020 2768.370 246.020 2768.380 ;
        RECT 423.020 2768.370 426.020 2768.380 ;
        RECT 603.020 2768.370 606.020 2768.380 ;
        RECT 783.020 2768.370 786.020 2768.380 ;
        RECT 963.020 2768.370 966.020 2768.380 ;
        RECT 1143.020 2768.370 1146.020 2768.380 ;
        RECT 1323.020 2768.370 1326.020 2768.380 ;
        RECT 1503.020 2768.370 1506.020 2768.380 ;
        RECT 1683.020 2768.370 1686.020 2768.380 ;
        RECT 1863.020 2768.370 1866.020 2768.380 ;
        RECT 2043.020 2768.370 2046.020 2768.380 ;
        RECT 2223.020 2768.370 2226.020 2768.380 ;
        RECT 2403.020 2768.370 2406.020 2768.380 ;
        RECT 2583.020 2768.370 2586.020 2768.380 ;
        RECT 2763.020 2768.370 2766.020 2768.380 ;
        RECT 2954.800 2768.370 2957.800 2768.380 ;
        RECT -38.180 2591.380 -35.180 2591.390 ;
        RECT 63.020 2591.380 66.020 2591.390 ;
        RECT 243.020 2591.380 246.020 2591.390 ;
        RECT 423.020 2591.380 426.020 2591.390 ;
        RECT 603.020 2591.380 606.020 2591.390 ;
        RECT 783.020 2591.380 786.020 2591.390 ;
        RECT 963.020 2591.380 966.020 2591.390 ;
        RECT 1143.020 2591.380 1146.020 2591.390 ;
        RECT 1323.020 2591.380 1326.020 2591.390 ;
        RECT 1503.020 2591.380 1506.020 2591.390 ;
        RECT 1683.020 2591.380 1686.020 2591.390 ;
        RECT 1863.020 2591.380 1866.020 2591.390 ;
        RECT 2043.020 2591.380 2046.020 2591.390 ;
        RECT 2223.020 2591.380 2226.020 2591.390 ;
        RECT 2403.020 2591.380 2406.020 2591.390 ;
        RECT 2583.020 2591.380 2586.020 2591.390 ;
        RECT 2763.020 2591.380 2766.020 2591.390 ;
        RECT 2954.800 2591.380 2957.800 2591.390 ;
        RECT -42.880 2588.380 2962.500 2591.380 ;
        RECT -38.180 2588.370 -35.180 2588.380 ;
        RECT 63.020 2588.370 66.020 2588.380 ;
        RECT 243.020 2588.370 246.020 2588.380 ;
        RECT 423.020 2588.370 426.020 2588.380 ;
        RECT 603.020 2588.370 606.020 2588.380 ;
        RECT 783.020 2588.370 786.020 2588.380 ;
        RECT 963.020 2588.370 966.020 2588.380 ;
        RECT 1143.020 2588.370 1146.020 2588.380 ;
        RECT 1323.020 2588.370 1326.020 2588.380 ;
        RECT 1503.020 2588.370 1506.020 2588.380 ;
        RECT 1683.020 2588.370 1686.020 2588.380 ;
        RECT 1863.020 2588.370 1866.020 2588.380 ;
        RECT 2043.020 2588.370 2046.020 2588.380 ;
        RECT 2223.020 2588.370 2226.020 2588.380 ;
        RECT 2403.020 2588.370 2406.020 2588.380 ;
        RECT 2583.020 2588.370 2586.020 2588.380 ;
        RECT 2763.020 2588.370 2766.020 2588.380 ;
        RECT 2954.800 2588.370 2957.800 2588.380 ;
        RECT -38.180 2411.380 -35.180 2411.390 ;
        RECT 63.020 2411.380 66.020 2411.390 ;
        RECT 243.020 2411.380 246.020 2411.390 ;
        RECT 423.020 2411.380 426.020 2411.390 ;
        RECT 603.020 2411.380 606.020 2411.390 ;
        RECT 783.020 2411.380 786.020 2411.390 ;
        RECT 963.020 2411.380 966.020 2411.390 ;
        RECT 1143.020 2411.380 1146.020 2411.390 ;
        RECT 1323.020 2411.380 1326.020 2411.390 ;
        RECT 1503.020 2411.380 1506.020 2411.390 ;
        RECT 1683.020 2411.380 1686.020 2411.390 ;
        RECT 1863.020 2411.380 1866.020 2411.390 ;
        RECT 2043.020 2411.380 2046.020 2411.390 ;
        RECT 2223.020 2411.380 2226.020 2411.390 ;
        RECT 2403.020 2411.380 2406.020 2411.390 ;
        RECT 2583.020 2411.380 2586.020 2411.390 ;
        RECT 2763.020 2411.380 2766.020 2411.390 ;
        RECT 2954.800 2411.380 2957.800 2411.390 ;
        RECT -42.880 2408.380 2962.500 2411.380 ;
        RECT -38.180 2408.370 -35.180 2408.380 ;
        RECT 63.020 2408.370 66.020 2408.380 ;
        RECT 243.020 2408.370 246.020 2408.380 ;
        RECT 423.020 2408.370 426.020 2408.380 ;
        RECT 603.020 2408.370 606.020 2408.380 ;
        RECT 783.020 2408.370 786.020 2408.380 ;
        RECT 963.020 2408.370 966.020 2408.380 ;
        RECT 1143.020 2408.370 1146.020 2408.380 ;
        RECT 1323.020 2408.370 1326.020 2408.380 ;
        RECT 1503.020 2408.370 1506.020 2408.380 ;
        RECT 1683.020 2408.370 1686.020 2408.380 ;
        RECT 1863.020 2408.370 1866.020 2408.380 ;
        RECT 2043.020 2408.370 2046.020 2408.380 ;
        RECT 2223.020 2408.370 2226.020 2408.380 ;
        RECT 2403.020 2408.370 2406.020 2408.380 ;
        RECT 2583.020 2408.370 2586.020 2408.380 ;
        RECT 2763.020 2408.370 2766.020 2408.380 ;
        RECT 2954.800 2408.370 2957.800 2408.380 ;
        RECT -38.180 2231.380 -35.180 2231.390 ;
        RECT 63.020 2231.380 66.020 2231.390 ;
        RECT 243.020 2231.380 246.020 2231.390 ;
        RECT 423.020 2231.380 426.020 2231.390 ;
        RECT 603.020 2231.380 606.020 2231.390 ;
        RECT 783.020 2231.380 786.020 2231.390 ;
        RECT 963.020 2231.380 966.020 2231.390 ;
        RECT 1143.020 2231.380 1146.020 2231.390 ;
        RECT 1323.020 2231.380 1326.020 2231.390 ;
        RECT 1503.020 2231.380 1506.020 2231.390 ;
        RECT 1683.020 2231.380 1686.020 2231.390 ;
        RECT 1863.020 2231.380 1866.020 2231.390 ;
        RECT 2043.020 2231.380 2046.020 2231.390 ;
        RECT 2223.020 2231.380 2226.020 2231.390 ;
        RECT 2403.020 2231.380 2406.020 2231.390 ;
        RECT 2583.020 2231.380 2586.020 2231.390 ;
        RECT 2763.020 2231.380 2766.020 2231.390 ;
        RECT 2954.800 2231.380 2957.800 2231.390 ;
        RECT -42.880 2228.380 2962.500 2231.380 ;
        RECT -38.180 2228.370 -35.180 2228.380 ;
        RECT 63.020 2228.370 66.020 2228.380 ;
        RECT 243.020 2228.370 246.020 2228.380 ;
        RECT 423.020 2228.370 426.020 2228.380 ;
        RECT 603.020 2228.370 606.020 2228.380 ;
        RECT 783.020 2228.370 786.020 2228.380 ;
        RECT 963.020 2228.370 966.020 2228.380 ;
        RECT 1143.020 2228.370 1146.020 2228.380 ;
        RECT 1323.020 2228.370 1326.020 2228.380 ;
        RECT 1503.020 2228.370 1506.020 2228.380 ;
        RECT 1683.020 2228.370 1686.020 2228.380 ;
        RECT 1863.020 2228.370 1866.020 2228.380 ;
        RECT 2043.020 2228.370 2046.020 2228.380 ;
        RECT 2223.020 2228.370 2226.020 2228.380 ;
        RECT 2403.020 2228.370 2406.020 2228.380 ;
        RECT 2583.020 2228.370 2586.020 2228.380 ;
        RECT 2763.020 2228.370 2766.020 2228.380 ;
        RECT 2954.800 2228.370 2957.800 2228.380 ;
        RECT -38.180 2051.380 -35.180 2051.390 ;
        RECT 63.020 2051.380 66.020 2051.390 ;
        RECT 243.020 2051.380 246.020 2051.390 ;
        RECT 423.020 2051.380 426.020 2051.390 ;
        RECT 603.020 2051.380 606.020 2051.390 ;
        RECT 783.020 2051.380 786.020 2051.390 ;
        RECT 963.020 2051.380 966.020 2051.390 ;
        RECT 1143.020 2051.380 1146.020 2051.390 ;
        RECT 1323.020 2051.380 1326.020 2051.390 ;
        RECT 1503.020 2051.380 1506.020 2051.390 ;
        RECT 1683.020 2051.380 1686.020 2051.390 ;
        RECT 1863.020 2051.380 1866.020 2051.390 ;
        RECT 2043.020 2051.380 2046.020 2051.390 ;
        RECT 2223.020 2051.380 2226.020 2051.390 ;
        RECT 2403.020 2051.380 2406.020 2051.390 ;
        RECT 2583.020 2051.380 2586.020 2051.390 ;
        RECT 2763.020 2051.380 2766.020 2051.390 ;
        RECT 2954.800 2051.380 2957.800 2051.390 ;
        RECT -42.880 2048.380 2962.500 2051.380 ;
        RECT -38.180 2048.370 -35.180 2048.380 ;
        RECT 63.020 2048.370 66.020 2048.380 ;
        RECT 243.020 2048.370 246.020 2048.380 ;
        RECT 423.020 2048.370 426.020 2048.380 ;
        RECT 603.020 2048.370 606.020 2048.380 ;
        RECT 783.020 2048.370 786.020 2048.380 ;
        RECT 963.020 2048.370 966.020 2048.380 ;
        RECT 1143.020 2048.370 1146.020 2048.380 ;
        RECT 1323.020 2048.370 1326.020 2048.380 ;
        RECT 1503.020 2048.370 1506.020 2048.380 ;
        RECT 1683.020 2048.370 1686.020 2048.380 ;
        RECT 1863.020 2048.370 1866.020 2048.380 ;
        RECT 2043.020 2048.370 2046.020 2048.380 ;
        RECT 2223.020 2048.370 2226.020 2048.380 ;
        RECT 2403.020 2048.370 2406.020 2048.380 ;
        RECT 2583.020 2048.370 2586.020 2048.380 ;
        RECT 2763.020 2048.370 2766.020 2048.380 ;
        RECT 2954.800 2048.370 2957.800 2048.380 ;
        RECT -38.180 1871.380 -35.180 1871.390 ;
        RECT 63.020 1871.380 66.020 1871.390 ;
        RECT 243.020 1871.380 246.020 1871.390 ;
        RECT 423.020 1871.380 426.020 1871.390 ;
        RECT 603.020 1871.380 606.020 1871.390 ;
        RECT 783.020 1871.380 786.020 1871.390 ;
        RECT 963.020 1871.380 966.020 1871.390 ;
        RECT 1143.020 1871.380 1146.020 1871.390 ;
        RECT 1323.020 1871.380 1326.020 1871.390 ;
        RECT 1503.020 1871.380 1506.020 1871.390 ;
        RECT 1683.020 1871.380 1686.020 1871.390 ;
        RECT 1863.020 1871.380 1866.020 1871.390 ;
        RECT 2043.020 1871.380 2046.020 1871.390 ;
        RECT 2223.020 1871.380 2226.020 1871.390 ;
        RECT 2403.020 1871.380 2406.020 1871.390 ;
        RECT 2583.020 1871.380 2586.020 1871.390 ;
        RECT 2763.020 1871.380 2766.020 1871.390 ;
        RECT 2954.800 1871.380 2957.800 1871.390 ;
        RECT -42.880 1868.380 2962.500 1871.380 ;
        RECT -38.180 1868.370 -35.180 1868.380 ;
        RECT 63.020 1868.370 66.020 1868.380 ;
        RECT 243.020 1868.370 246.020 1868.380 ;
        RECT 423.020 1868.370 426.020 1868.380 ;
        RECT 603.020 1868.370 606.020 1868.380 ;
        RECT 783.020 1868.370 786.020 1868.380 ;
        RECT 963.020 1868.370 966.020 1868.380 ;
        RECT 1143.020 1868.370 1146.020 1868.380 ;
        RECT 1323.020 1868.370 1326.020 1868.380 ;
        RECT 1503.020 1868.370 1506.020 1868.380 ;
        RECT 1683.020 1868.370 1686.020 1868.380 ;
        RECT 1863.020 1868.370 1866.020 1868.380 ;
        RECT 2043.020 1868.370 2046.020 1868.380 ;
        RECT 2223.020 1868.370 2226.020 1868.380 ;
        RECT 2403.020 1868.370 2406.020 1868.380 ;
        RECT 2583.020 1868.370 2586.020 1868.380 ;
        RECT 2763.020 1868.370 2766.020 1868.380 ;
        RECT 2954.800 1868.370 2957.800 1868.380 ;
        RECT -38.180 1691.380 -35.180 1691.390 ;
        RECT 63.020 1691.380 66.020 1691.390 ;
        RECT 243.020 1691.380 246.020 1691.390 ;
        RECT 423.020 1691.380 426.020 1691.390 ;
        RECT 603.020 1691.380 606.020 1691.390 ;
        RECT 783.020 1691.380 786.020 1691.390 ;
        RECT 963.020 1691.380 966.020 1691.390 ;
        RECT 1143.020 1691.380 1146.020 1691.390 ;
        RECT 1323.020 1691.380 1326.020 1691.390 ;
        RECT 1503.020 1691.380 1506.020 1691.390 ;
        RECT 1683.020 1691.380 1686.020 1691.390 ;
        RECT 1863.020 1691.380 1866.020 1691.390 ;
        RECT 2043.020 1691.380 2046.020 1691.390 ;
        RECT 2223.020 1691.380 2226.020 1691.390 ;
        RECT 2403.020 1691.380 2406.020 1691.390 ;
        RECT 2583.020 1691.380 2586.020 1691.390 ;
        RECT 2763.020 1691.380 2766.020 1691.390 ;
        RECT 2954.800 1691.380 2957.800 1691.390 ;
        RECT -42.880 1688.380 2962.500 1691.380 ;
        RECT -38.180 1688.370 -35.180 1688.380 ;
        RECT 63.020 1688.370 66.020 1688.380 ;
        RECT 243.020 1688.370 246.020 1688.380 ;
        RECT 423.020 1688.370 426.020 1688.380 ;
        RECT 603.020 1688.370 606.020 1688.380 ;
        RECT 783.020 1688.370 786.020 1688.380 ;
        RECT 963.020 1688.370 966.020 1688.380 ;
        RECT 1143.020 1688.370 1146.020 1688.380 ;
        RECT 1323.020 1688.370 1326.020 1688.380 ;
        RECT 1503.020 1688.370 1506.020 1688.380 ;
        RECT 1683.020 1688.370 1686.020 1688.380 ;
        RECT 1863.020 1688.370 1866.020 1688.380 ;
        RECT 2043.020 1688.370 2046.020 1688.380 ;
        RECT 2223.020 1688.370 2226.020 1688.380 ;
        RECT 2403.020 1688.370 2406.020 1688.380 ;
        RECT 2583.020 1688.370 2586.020 1688.380 ;
        RECT 2763.020 1688.370 2766.020 1688.380 ;
        RECT 2954.800 1688.370 2957.800 1688.380 ;
        RECT -38.180 1511.380 -35.180 1511.390 ;
        RECT 63.020 1511.380 66.020 1511.390 ;
        RECT 243.020 1511.380 246.020 1511.390 ;
        RECT 423.020 1511.380 426.020 1511.390 ;
        RECT 603.020 1511.380 606.020 1511.390 ;
        RECT 783.020 1511.380 786.020 1511.390 ;
        RECT 963.020 1511.380 966.020 1511.390 ;
        RECT 1143.020 1511.380 1146.020 1511.390 ;
        RECT 1323.020 1511.380 1326.020 1511.390 ;
        RECT 1503.020 1511.380 1506.020 1511.390 ;
        RECT 1683.020 1511.380 1686.020 1511.390 ;
        RECT 1863.020 1511.380 1866.020 1511.390 ;
        RECT 2043.020 1511.380 2046.020 1511.390 ;
        RECT 2223.020 1511.380 2226.020 1511.390 ;
        RECT 2403.020 1511.380 2406.020 1511.390 ;
        RECT 2583.020 1511.380 2586.020 1511.390 ;
        RECT 2763.020 1511.380 2766.020 1511.390 ;
        RECT 2954.800 1511.380 2957.800 1511.390 ;
        RECT -42.880 1508.380 2962.500 1511.380 ;
        RECT -38.180 1508.370 -35.180 1508.380 ;
        RECT 63.020 1508.370 66.020 1508.380 ;
        RECT 243.020 1508.370 246.020 1508.380 ;
        RECT 423.020 1508.370 426.020 1508.380 ;
        RECT 603.020 1508.370 606.020 1508.380 ;
        RECT 783.020 1508.370 786.020 1508.380 ;
        RECT 963.020 1508.370 966.020 1508.380 ;
        RECT 1143.020 1508.370 1146.020 1508.380 ;
        RECT 1323.020 1508.370 1326.020 1508.380 ;
        RECT 1503.020 1508.370 1506.020 1508.380 ;
        RECT 1683.020 1508.370 1686.020 1508.380 ;
        RECT 1863.020 1508.370 1866.020 1508.380 ;
        RECT 2043.020 1508.370 2046.020 1508.380 ;
        RECT 2223.020 1508.370 2226.020 1508.380 ;
        RECT 2403.020 1508.370 2406.020 1508.380 ;
        RECT 2583.020 1508.370 2586.020 1508.380 ;
        RECT 2763.020 1508.370 2766.020 1508.380 ;
        RECT 2954.800 1508.370 2957.800 1508.380 ;
        RECT -38.180 1331.380 -35.180 1331.390 ;
        RECT 63.020 1331.380 66.020 1331.390 ;
        RECT 243.020 1331.380 246.020 1331.390 ;
        RECT 423.020 1331.380 426.020 1331.390 ;
        RECT 603.020 1331.380 606.020 1331.390 ;
        RECT 783.020 1331.380 786.020 1331.390 ;
        RECT 963.020 1331.380 966.020 1331.390 ;
        RECT 1143.020 1331.380 1146.020 1331.390 ;
        RECT 1323.020 1331.380 1326.020 1331.390 ;
        RECT 1503.020 1331.380 1506.020 1331.390 ;
        RECT 1683.020 1331.380 1686.020 1331.390 ;
        RECT 1863.020 1331.380 1866.020 1331.390 ;
        RECT 2043.020 1331.380 2046.020 1331.390 ;
        RECT 2223.020 1331.380 2226.020 1331.390 ;
        RECT 2403.020 1331.380 2406.020 1331.390 ;
        RECT 2583.020 1331.380 2586.020 1331.390 ;
        RECT 2763.020 1331.380 2766.020 1331.390 ;
        RECT 2954.800 1331.380 2957.800 1331.390 ;
        RECT -42.880 1328.380 2962.500 1331.380 ;
        RECT -38.180 1328.370 -35.180 1328.380 ;
        RECT 63.020 1328.370 66.020 1328.380 ;
        RECT 243.020 1328.370 246.020 1328.380 ;
        RECT 423.020 1328.370 426.020 1328.380 ;
        RECT 603.020 1328.370 606.020 1328.380 ;
        RECT 783.020 1328.370 786.020 1328.380 ;
        RECT 963.020 1328.370 966.020 1328.380 ;
        RECT 1143.020 1328.370 1146.020 1328.380 ;
        RECT 1323.020 1328.370 1326.020 1328.380 ;
        RECT 1503.020 1328.370 1506.020 1328.380 ;
        RECT 1683.020 1328.370 1686.020 1328.380 ;
        RECT 1863.020 1328.370 1866.020 1328.380 ;
        RECT 2043.020 1328.370 2046.020 1328.380 ;
        RECT 2223.020 1328.370 2226.020 1328.380 ;
        RECT 2403.020 1328.370 2406.020 1328.380 ;
        RECT 2583.020 1328.370 2586.020 1328.380 ;
        RECT 2763.020 1328.370 2766.020 1328.380 ;
        RECT 2954.800 1328.370 2957.800 1328.380 ;
        RECT -38.180 1151.380 -35.180 1151.390 ;
        RECT 63.020 1151.380 66.020 1151.390 ;
        RECT 243.020 1151.380 246.020 1151.390 ;
        RECT 423.020 1151.380 426.020 1151.390 ;
        RECT 603.020 1151.380 606.020 1151.390 ;
        RECT 783.020 1151.380 786.020 1151.390 ;
        RECT 963.020 1151.380 966.020 1151.390 ;
        RECT 1143.020 1151.380 1146.020 1151.390 ;
        RECT 1323.020 1151.380 1326.020 1151.390 ;
        RECT 1503.020 1151.380 1506.020 1151.390 ;
        RECT 1683.020 1151.380 1686.020 1151.390 ;
        RECT 1863.020 1151.380 1866.020 1151.390 ;
        RECT 2043.020 1151.380 2046.020 1151.390 ;
        RECT 2223.020 1151.380 2226.020 1151.390 ;
        RECT 2403.020 1151.380 2406.020 1151.390 ;
        RECT 2583.020 1151.380 2586.020 1151.390 ;
        RECT 2763.020 1151.380 2766.020 1151.390 ;
        RECT 2954.800 1151.380 2957.800 1151.390 ;
        RECT -42.880 1148.380 2962.500 1151.380 ;
        RECT -38.180 1148.370 -35.180 1148.380 ;
        RECT 63.020 1148.370 66.020 1148.380 ;
        RECT 243.020 1148.370 246.020 1148.380 ;
        RECT 423.020 1148.370 426.020 1148.380 ;
        RECT 603.020 1148.370 606.020 1148.380 ;
        RECT 783.020 1148.370 786.020 1148.380 ;
        RECT 963.020 1148.370 966.020 1148.380 ;
        RECT 1143.020 1148.370 1146.020 1148.380 ;
        RECT 1323.020 1148.370 1326.020 1148.380 ;
        RECT 1503.020 1148.370 1506.020 1148.380 ;
        RECT 1683.020 1148.370 1686.020 1148.380 ;
        RECT 1863.020 1148.370 1866.020 1148.380 ;
        RECT 2043.020 1148.370 2046.020 1148.380 ;
        RECT 2223.020 1148.370 2226.020 1148.380 ;
        RECT 2403.020 1148.370 2406.020 1148.380 ;
        RECT 2583.020 1148.370 2586.020 1148.380 ;
        RECT 2763.020 1148.370 2766.020 1148.380 ;
        RECT 2954.800 1148.370 2957.800 1148.380 ;
        RECT -38.180 971.380 -35.180 971.390 ;
        RECT 63.020 971.380 66.020 971.390 ;
        RECT 243.020 971.380 246.020 971.390 ;
        RECT 423.020 971.380 426.020 971.390 ;
        RECT 603.020 971.380 606.020 971.390 ;
        RECT 783.020 971.380 786.020 971.390 ;
        RECT 963.020 971.380 966.020 971.390 ;
        RECT 1143.020 971.380 1146.020 971.390 ;
        RECT 1323.020 971.380 1326.020 971.390 ;
        RECT 1503.020 971.380 1506.020 971.390 ;
        RECT 1683.020 971.380 1686.020 971.390 ;
        RECT 1863.020 971.380 1866.020 971.390 ;
        RECT 2043.020 971.380 2046.020 971.390 ;
        RECT 2223.020 971.380 2226.020 971.390 ;
        RECT 2403.020 971.380 2406.020 971.390 ;
        RECT 2583.020 971.380 2586.020 971.390 ;
        RECT 2763.020 971.380 2766.020 971.390 ;
        RECT 2954.800 971.380 2957.800 971.390 ;
        RECT -42.880 968.380 2962.500 971.380 ;
        RECT -38.180 968.370 -35.180 968.380 ;
        RECT 63.020 968.370 66.020 968.380 ;
        RECT 243.020 968.370 246.020 968.380 ;
        RECT 423.020 968.370 426.020 968.380 ;
        RECT 603.020 968.370 606.020 968.380 ;
        RECT 783.020 968.370 786.020 968.380 ;
        RECT 963.020 968.370 966.020 968.380 ;
        RECT 1143.020 968.370 1146.020 968.380 ;
        RECT 1323.020 968.370 1326.020 968.380 ;
        RECT 1503.020 968.370 1506.020 968.380 ;
        RECT 1683.020 968.370 1686.020 968.380 ;
        RECT 1863.020 968.370 1866.020 968.380 ;
        RECT 2043.020 968.370 2046.020 968.380 ;
        RECT 2223.020 968.370 2226.020 968.380 ;
        RECT 2403.020 968.370 2406.020 968.380 ;
        RECT 2583.020 968.370 2586.020 968.380 ;
        RECT 2763.020 968.370 2766.020 968.380 ;
        RECT 2954.800 968.370 2957.800 968.380 ;
        RECT -38.180 791.380 -35.180 791.390 ;
        RECT 63.020 791.380 66.020 791.390 ;
        RECT 243.020 791.380 246.020 791.390 ;
        RECT 423.020 791.380 426.020 791.390 ;
        RECT 603.020 791.380 606.020 791.390 ;
        RECT 783.020 791.380 786.020 791.390 ;
        RECT 963.020 791.380 966.020 791.390 ;
        RECT 1143.020 791.380 1146.020 791.390 ;
        RECT 1323.020 791.380 1326.020 791.390 ;
        RECT 1503.020 791.380 1506.020 791.390 ;
        RECT 1683.020 791.380 1686.020 791.390 ;
        RECT 1863.020 791.380 1866.020 791.390 ;
        RECT 2043.020 791.380 2046.020 791.390 ;
        RECT 2223.020 791.380 2226.020 791.390 ;
        RECT 2403.020 791.380 2406.020 791.390 ;
        RECT 2583.020 791.380 2586.020 791.390 ;
        RECT 2763.020 791.380 2766.020 791.390 ;
        RECT 2954.800 791.380 2957.800 791.390 ;
        RECT -42.880 788.380 2962.500 791.380 ;
        RECT -38.180 788.370 -35.180 788.380 ;
        RECT 63.020 788.370 66.020 788.380 ;
        RECT 243.020 788.370 246.020 788.380 ;
        RECT 423.020 788.370 426.020 788.380 ;
        RECT 603.020 788.370 606.020 788.380 ;
        RECT 783.020 788.370 786.020 788.380 ;
        RECT 963.020 788.370 966.020 788.380 ;
        RECT 1143.020 788.370 1146.020 788.380 ;
        RECT 1323.020 788.370 1326.020 788.380 ;
        RECT 1503.020 788.370 1506.020 788.380 ;
        RECT 1683.020 788.370 1686.020 788.380 ;
        RECT 1863.020 788.370 1866.020 788.380 ;
        RECT 2043.020 788.370 2046.020 788.380 ;
        RECT 2223.020 788.370 2226.020 788.380 ;
        RECT 2403.020 788.370 2406.020 788.380 ;
        RECT 2583.020 788.370 2586.020 788.380 ;
        RECT 2763.020 788.370 2766.020 788.380 ;
        RECT 2954.800 788.370 2957.800 788.380 ;
        RECT -38.180 611.380 -35.180 611.390 ;
        RECT 63.020 611.380 66.020 611.390 ;
        RECT 243.020 611.380 246.020 611.390 ;
        RECT 423.020 611.380 426.020 611.390 ;
        RECT 603.020 611.380 606.020 611.390 ;
        RECT 783.020 611.380 786.020 611.390 ;
        RECT 963.020 611.380 966.020 611.390 ;
        RECT 1143.020 611.380 1146.020 611.390 ;
        RECT 1323.020 611.380 1326.020 611.390 ;
        RECT 1503.020 611.380 1506.020 611.390 ;
        RECT 1683.020 611.380 1686.020 611.390 ;
        RECT 1863.020 611.380 1866.020 611.390 ;
        RECT 2043.020 611.380 2046.020 611.390 ;
        RECT 2223.020 611.380 2226.020 611.390 ;
        RECT 2403.020 611.380 2406.020 611.390 ;
        RECT 2583.020 611.380 2586.020 611.390 ;
        RECT 2763.020 611.380 2766.020 611.390 ;
        RECT 2954.800 611.380 2957.800 611.390 ;
        RECT -42.880 608.380 2962.500 611.380 ;
        RECT -38.180 608.370 -35.180 608.380 ;
        RECT 63.020 608.370 66.020 608.380 ;
        RECT 243.020 608.370 246.020 608.380 ;
        RECT 423.020 608.370 426.020 608.380 ;
        RECT 603.020 608.370 606.020 608.380 ;
        RECT 783.020 608.370 786.020 608.380 ;
        RECT 963.020 608.370 966.020 608.380 ;
        RECT 1143.020 608.370 1146.020 608.380 ;
        RECT 1323.020 608.370 1326.020 608.380 ;
        RECT 1503.020 608.370 1506.020 608.380 ;
        RECT 1683.020 608.370 1686.020 608.380 ;
        RECT 1863.020 608.370 1866.020 608.380 ;
        RECT 2043.020 608.370 2046.020 608.380 ;
        RECT 2223.020 608.370 2226.020 608.380 ;
        RECT 2403.020 608.370 2406.020 608.380 ;
        RECT 2583.020 608.370 2586.020 608.380 ;
        RECT 2763.020 608.370 2766.020 608.380 ;
        RECT 2954.800 608.370 2957.800 608.380 ;
        RECT -38.180 431.380 -35.180 431.390 ;
        RECT 63.020 431.380 66.020 431.390 ;
        RECT 243.020 431.380 246.020 431.390 ;
        RECT 423.020 431.380 426.020 431.390 ;
        RECT 603.020 431.380 606.020 431.390 ;
        RECT 783.020 431.380 786.020 431.390 ;
        RECT 963.020 431.380 966.020 431.390 ;
        RECT 1143.020 431.380 1146.020 431.390 ;
        RECT 1323.020 431.380 1326.020 431.390 ;
        RECT 1503.020 431.380 1506.020 431.390 ;
        RECT 1683.020 431.380 1686.020 431.390 ;
        RECT 1863.020 431.380 1866.020 431.390 ;
        RECT 2043.020 431.380 2046.020 431.390 ;
        RECT 2223.020 431.380 2226.020 431.390 ;
        RECT 2403.020 431.380 2406.020 431.390 ;
        RECT 2583.020 431.380 2586.020 431.390 ;
        RECT 2763.020 431.380 2766.020 431.390 ;
        RECT 2954.800 431.380 2957.800 431.390 ;
        RECT -42.880 428.380 2962.500 431.380 ;
        RECT -38.180 428.370 -35.180 428.380 ;
        RECT 63.020 428.370 66.020 428.380 ;
        RECT 243.020 428.370 246.020 428.380 ;
        RECT 423.020 428.370 426.020 428.380 ;
        RECT 603.020 428.370 606.020 428.380 ;
        RECT 783.020 428.370 786.020 428.380 ;
        RECT 963.020 428.370 966.020 428.380 ;
        RECT 1143.020 428.370 1146.020 428.380 ;
        RECT 1323.020 428.370 1326.020 428.380 ;
        RECT 1503.020 428.370 1506.020 428.380 ;
        RECT 1683.020 428.370 1686.020 428.380 ;
        RECT 1863.020 428.370 1866.020 428.380 ;
        RECT 2043.020 428.370 2046.020 428.380 ;
        RECT 2223.020 428.370 2226.020 428.380 ;
        RECT 2403.020 428.370 2406.020 428.380 ;
        RECT 2583.020 428.370 2586.020 428.380 ;
        RECT 2763.020 428.370 2766.020 428.380 ;
        RECT 2954.800 428.370 2957.800 428.380 ;
        RECT -38.180 251.380 -35.180 251.390 ;
        RECT 63.020 251.380 66.020 251.390 ;
        RECT 243.020 251.380 246.020 251.390 ;
        RECT 423.020 251.380 426.020 251.390 ;
        RECT 603.020 251.380 606.020 251.390 ;
        RECT 783.020 251.380 786.020 251.390 ;
        RECT 963.020 251.380 966.020 251.390 ;
        RECT 1143.020 251.380 1146.020 251.390 ;
        RECT 1323.020 251.380 1326.020 251.390 ;
        RECT 1503.020 251.380 1506.020 251.390 ;
        RECT 1683.020 251.380 1686.020 251.390 ;
        RECT 1863.020 251.380 1866.020 251.390 ;
        RECT 2043.020 251.380 2046.020 251.390 ;
        RECT 2223.020 251.380 2226.020 251.390 ;
        RECT 2403.020 251.380 2406.020 251.390 ;
        RECT 2583.020 251.380 2586.020 251.390 ;
        RECT 2763.020 251.380 2766.020 251.390 ;
        RECT 2954.800 251.380 2957.800 251.390 ;
        RECT -42.880 248.380 2962.500 251.380 ;
        RECT -38.180 248.370 -35.180 248.380 ;
        RECT 63.020 248.370 66.020 248.380 ;
        RECT 243.020 248.370 246.020 248.380 ;
        RECT 423.020 248.370 426.020 248.380 ;
        RECT 603.020 248.370 606.020 248.380 ;
        RECT 783.020 248.370 786.020 248.380 ;
        RECT 963.020 248.370 966.020 248.380 ;
        RECT 1143.020 248.370 1146.020 248.380 ;
        RECT 1323.020 248.370 1326.020 248.380 ;
        RECT 1503.020 248.370 1506.020 248.380 ;
        RECT 1683.020 248.370 1686.020 248.380 ;
        RECT 1863.020 248.370 1866.020 248.380 ;
        RECT 2043.020 248.370 2046.020 248.380 ;
        RECT 2223.020 248.370 2226.020 248.380 ;
        RECT 2403.020 248.370 2406.020 248.380 ;
        RECT 2583.020 248.370 2586.020 248.380 ;
        RECT 2763.020 248.370 2766.020 248.380 ;
        RECT 2954.800 248.370 2957.800 248.380 ;
        RECT -38.180 71.380 -35.180 71.390 ;
        RECT 63.020 71.380 66.020 71.390 ;
        RECT 243.020 71.380 246.020 71.390 ;
        RECT 423.020 71.380 426.020 71.390 ;
        RECT 603.020 71.380 606.020 71.390 ;
        RECT 783.020 71.380 786.020 71.390 ;
        RECT 963.020 71.380 966.020 71.390 ;
        RECT 1143.020 71.380 1146.020 71.390 ;
        RECT 1323.020 71.380 1326.020 71.390 ;
        RECT 1503.020 71.380 1506.020 71.390 ;
        RECT 1683.020 71.380 1686.020 71.390 ;
        RECT 1863.020 71.380 1866.020 71.390 ;
        RECT 2043.020 71.380 2046.020 71.390 ;
        RECT 2223.020 71.380 2226.020 71.390 ;
        RECT 2403.020 71.380 2406.020 71.390 ;
        RECT 2583.020 71.380 2586.020 71.390 ;
        RECT 2763.020 71.380 2766.020 71.390 ;
        RECT 2954.800 71.380 2957.800 71.390 ;
        RECT -42.880 68.380 2962.500 71.380 ;
        RECT -38.180 68.370 -35.180 68.380 ;
        RECT 63.020 68.370 66.020 68.380 ;
        RECT 243.020 68.370 246.020 68.380 ;
        RECT 423.020 68.370 426.020 68.380 ;
        RECT 603.020 68.370 606.020 68.380 ;
        RECT 783.020 68.370 786.020 68.380 ;
        RECT 963.020 68.370 966.020 68.380 ;
        RECT 1143.020 68.370 1146.020 68.380 ;
        RECT 1323.020 68.370 1326.020 68.380 ;
        RECT 1503.020 68.370 1506.020 68.380 ;
        RECT 1683.020 68.370 1686.020 68.380 ;
        RECT 1863.020 68.370 1866.020 68.380 ;
        RECT 2043.020 68.370 2046.020 68.380 ;
        RECT 2223.020 68.370 2226.020 68.380 ;
        RECT 2403.020 68.370 2406.020 68.380 ;
        RECT 2583.020 68.370 2586.020 68.380 ;
        RECT 2763.020 68.370 2766.020 68.380 ;
        RECT 2954.800 68.370 2957.800 68.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 63.020 -29.820 66.020 -29.810 ;
        RECT 243.020 -29.820 246.020 -29.810 ;
        RECT 423.020 -29.820 426.020 -29.810 ;
        RECT 603.020 -29.820 606.020 -29.810 ;
        RECT 783.020 -29.820 786.020 -29.810 ;
        RECT 963.020 -29.820 966.020 -29.810 ;
        RECT 1143.020 -29.820 1146.020 -29.810 ;
        RECT 1323.020 -29.820 1326.020 -29.810 ;
        RECT 1503.020 -29.820 1506.020 -29.810 ;
        RECT 1683.020 -29.820 1686.020 -29.810 ;
        RECT 1863.020 -29.820 1866.020 -29.810 ;
        RECT 2043.020 -29.820 2046.020 -29.810 ;
        RECT 2223.020 -29.820 2226.020 -29.810 ;
        RECT 2403.020 -29.820 2406.020 -29.810 ;
        RECT 2583.020 -29.820 2586.020 -29.810 ;
        RECT 2763.020 -29.820 2766.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 63.020 -32.830 66.020 -32.820 ;
        RECT 243.020 -32.830 246.020 -32.820 ;
        RECT 423.020 -32.830 426.020 -32.820 ;
        RECT 603.020 -32.830 606.020 -32.820 ;
        RECT 783.020 -32.830 786.020 -32.820 ;
        RECT 963.020 -32.830 966.020 -32.820 ;
        RECT 1143.020 -32.830 1146.020 -32.820 ;
        RECT 1323.020 -32.830 1326.020 -32.820 ;
        RECT 1503.020 -32.830 1506.020 -32.820 ;
        RECT 1683.020 -32.830 1686.020 -32.820 ;
        RECT 1863.020 -32.830 1866.020 -32.820 ;
        RECT 2043.020 -32.830 2046.020 -32.820 ;
        RECT 2223.020 -32.830 2226.020 -32.820 ;
        RECT 2403.020 -32.830 2406.020 -32.820 ;
        RECT 2583.020 -32.830 2586.020 -32.820 ;
        RECT 2763.020 -32.830 2766.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 153.020 -37.520 156.020 3557.200 ;
        RECT 333.020 -37.520 336.020 3557.200 ;
        RECT 513.020 -37.520 516.020 3557.200 ;
        RECT 693.020 -37.520 696.020 3557.200 ;
        RECT 873.020 -37.520 876.020 3557.200 ;
        RECT 1053.020 -37.520 1056.020 3557.200 ;
        RECT 1233.020 -37.520 1236.020 3557.200 ;
        RECT 1413.020 -37.520 1416.020 3557.200 ;
        RECT 1593.020 -37.520 1596.020 3557.200 ;
        RECT 1773.020 -37.520 1776.020 3557.200 ;
        RECT 1953.020 -37.520 1956.020 3557.200 ;
        RECT 2133.020 -37.520 2136.020 3557.200 ;
        RECT 2313.020 -37.520 2316.020 3557.200 ;
        RECT 2493.020 -37.520 2496.020 3557.200 ;
        RECT 2673.020 -37.520 2676.020 3557.200 ;
        RECT 2853.020 -37.520 2856.020 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 3400.090 -40.790 3401.270 ;
        RECT -41.970 3398.490 -40.790 3399.670 ;
        RECT -41.970 3220.090 -40.790 3221.270 ;
        RECT -41.970 3218.490 -40.790 3219.670 ;
        RECT -41.970 3040.090 -40.790 3041.270 ;
        RECT -41.970 3038.490 -40.790 3039.670 ;
        RECT -41.970 2860.090 -40.790 2861.270 ;
        RECT -41.970 2858.490 -40.790 2859.670 ;
        RECT -41.970 2680.090 -40.790 2681.270 ;
        RECT -41.970 2678.490 -40.790 2679.670 ;
        RECT -41.970 2500.090 -40.790 2501.270 ;
        RECT -41.970 2498.490 -40.790 2499.670 ;
        RECT -41.970 2320.090 -40.790 2321.270 ;
        RECT -41.970 2318.490 -40.790 2319.670 ;
        RECT -41.970 2140.090 -40.790 2141.270 ;
        RECT -41.970 2138.490 -40.790 2139.670 ;
        RECT -41.970 1960.090 -40.790 1961.270 ;
        RECT -41.970 1958.490 -40.790 1959.670 ;
        RECT -41.970 1780.090 -40.790 1781.270 ;
        RECT -41.970 1778.490 -40.790 1779.670 ;
        RECT -41.970 1600.090 -40.790 1601.270 ;
        RECT -41.970 1598.490 -40.790 1599.670 ;
        RECT -41.970 1420.090 -40.790 1421.270 ;
        RECT -41.970 1418.490 -40.790 1419.670 ;
        RECT -41.970 1240.090 -40.790 1241.270 ;
        RECT -41.970 1238.490 -40.790 1239.670 ;
        RECT -41.970 1060.090 -40.790 1061.270 ;
        RECT -41.970 1058.490 -40.790 1059.670 ;
        RECT -41.970 880.090 -40.790 881.270 ;
        RECT -41.970 878.490 -40.790 879.670 ;
        RECT -41.970 700.090 -40.790 701.270 ;
        RECT -41.970 698.490 -40.790 699.670 ;
        RECT -41.970 520.090 -40.790 521.270 ;
        RECT -41.970 518.490 -40.790 519.670 ;
        RECT -41.970 340.090 -40.790 341.270 ;
        RECT -41.970 338.490 -40.790 339.670 ;
        RECT -41.970 160.090 -40.790 161.270 ;
        RECT -41.970 158.490 -40.790 159.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 153.930 3555.910 155.110 3557.090 ;
        RECT 153.930 3554.310 155.110 3555.490 ;
        RECT 153.930 3400.090 155.110 3401.270 ;
        RECT 153.930 3398.490 155.110 3399.670 ;
        RECT 153.930 3220.090 155.110 3221.270 ;
        RECT 153.930 3218.490 155.110 3219.670 ;
        RECT 153.930 3040.090 155.110 3041.270 ;
        RECT 153.930 3038.490 155.110 3039.670 ;
        RECT 153.930 2860.090 155.110 2861.270 ;
        RECT 153.930 2858.490 155.110 2859.670 ;
        RECT 153.930 2680.090 155.110 2681.270 ;
        RECT 153.930 2678.490 155.110 2679.670 ;
        RECT 153.930 2500.090 155.110 2501.270 ;
        RECT 153.930 2498.490 155.110 2499.670 ;
        RECT 153.930 2320.090 155.110 2321.270 ;
        RECT 153.930 2318.490 155.110 2319.670 ;
        RECT 153.930 2140.090 155.110 2141.270 ;
        RECT 153.930 2138.490 155.110 2139.670 ;
        RECT 153.930 1960.090 155.110 1961.270 ;
        RECT 153.930 1958.490 155.110 1959.670 ;
        RECT 153.930 1780.090 155.110 1781.270 ;
        RECT 153.930 1778.490 155.110 1779.670 ;
        RECT 153.930 1600.090 155.110 1601.270 ;
        RECT 153.930 1598.490 155.110 1599.670 ;
        RECT 153.930 1420.090 155.110 1421.270 ;
        RECT 153.930 1418.490 155.110 1419.670 ;
        RECT 153.930 1240.090 155.110 1241.270 ;
        RECT 153.930 1238.490 155.110 1239.670 ;
        RECT 153.930 1060.090 155.110 1061.270 ;
        RECT 153.930 1058.490 155.110 1059.670 ;
        RECT 153.930 880.090 155.110 881.270 ;
        RECT 153.930 878.490 155.110 879.670 ;
        RECT 153.930 700.090 155.110 701.270 ;
        RECT 153.930 698.490 155.110 699.670 ;
        RECT 153.930 520.090 155.110 521.270 ;
        RECT 153.930 518.490 155.110 519.670 ;
        RECT 153.930 340.090 155.110 341.270 ;
        RECT 153.930 338.490 155.110 339.670 ;
        RECT 153.930 160.090 155.110 161.270 ;
        RECT 153.930 158.490 155.110 159.670 ;
        RECT 153.930 -35.810 155.110 -34.630 ;
        RECT 153.930 -37.410 155.110 -36.230 ;
        RECT 333.930 3555.910 335.110 3557.090 ;
        RECT 333.930 3554.310 335.110 3555.490 ;
        RECT 333.930 3400.090 335.110 3401.270 ;
        RECT 333.930 3398.490 335.110 3399.670 ;
        RECT 333.930 3220.090 335.110 3221.270 ;
        RECT 333.930 3218.490 335.110 3219.670 ;
        RECT 333.930 3040.090 335.110 3041.270 ;
        RECT 333.930 3038.490 335.110 3039.670 ;
        RECT 333.930 2860.090 335.110 2861.270 ;
        RECT 333.930 2858.490 335.110 2859.670 ;
        RECT 333.930 2680.090 335.110 2681.270 ;
        RECT 333.930 2678.490 335.110 2679.670 ;
        RECT 333.930 2500.090 335.110 2501.270 ;
        RECT 333.930 2498.490 335.110 2499.670 ;
        RECT 333.930 2320.090 335.110 2321.270 ;
        RECT 333.930 2318.490 335.110 2319.670 ;
        RECT 333.930 2140.090 335.110 2141.270 ;
        RECT 333.930 2138.490 335.110 2139.670 ;
        RECT 333.930 1960.090 335.110 1961.270 ;
        RECT 333.930 1958.490 335.110 1959.670 ;
        RECT 333.930 1780.090 335.110 1781.270 ;
        RECT 333.930 1778.490 335.110 1779.670 ;
        RECT 333.930 1600.090 335.110 1601.270 ;
        RECT 333.930 1598.490 335.110 1599.670 ;
        RECT 333.930 1420.090 335.110 1421.270 ;
        RECT 333.930 1418.490 335.110 1419.670 ;
        RECT 333.930 1240.090 335.110 1241.270 ;
        RECT 333.930 1238.490 335.110 1239.670 ;
        RECT 333.930 1060.090 335.110 1061.270 ;
        RECT 333.930 1058.490 335.110 1059.670 ;
        RECT 333.930 880.090 335.110 881.270 ;
        RECT 333.930 878.490 335.110 879.670 ;
        RECT 333.930 700.090 335.110 701.270 ;
        RECT 333.930 698.490 335.110 699.670 ;
        RECT 333.930 520.090 335.110 521.270 ;
        RECT 333.930 518.490 335.110 519.670 ;
        RECT 333.930 340.090 335.110 341.270 ;
        RECT 333.930 338.490 335.110 339.670 ;
        RECT 333.930 160.090 335.110 161.270 ;
        RECT 333.930 158.490 335.110 159.670 ;
        RECT 333.930 -35.810 335.110 -34.630 ;
        RECT 333.930 -37.410 335.110 -36.230 ;
        RECT 513.930 3555.910 515.110 3557.090 ;
        RECT 513.930 3554.310 515.110 3555.490 ;
        RECT 513.930 3400.090 515.110 3401.270 ;
        RECT 513.930 3398.490 515.110 3399.670 ;
        RECT 513.930 3220.090 515.110 3221.270 ;
        RECT 513.930 3218.490 515.110 3219.670 ;
        RECT 513.930 3040.090 515.110 3041.270 ;
        RECT 513.930 3038.490 515.110 3039.670 ;
        RECT 513.930 2860.090 515.110 2861.270 ;
        RECT 513.930 2858.490 515.110 2859.670 ;
        RECT 513.930 2680.090 515.110 2681.270 ;
        RECT 513.930 2678.490 515.110 2679.670 ;
        RECT 513.930 2500.090 515.110 2501.270 ;
        RECT 513.930 2498.490 515.110 2499.670 ;
        RECT 513.930 2320.090 515.110 2321.270 ;
        RECT 513.930 2318.490 515.110 2319.670 ;
        RECT 513.930 2140.090 515.110 2141.270 ;
        RECT 513.930 2138.490 515.110 2139.670 ;
        RECT 513.930 1960.090 515.110 1961.270 ;
        RECT 513.930 1958.490 515.110 1959.670 ;
        RECT 513.930 1780.090 515.110 1781.270 ;
        RECT 513.930 1778.490 515.110 1779.670 ;
        RECT 513.930 1600.090 515.110 1601.270 ;
        RECT 513.930 1598.490 515.110 1599.670 ;
        RECT 513.930 1420.090 515.110 1421.270 ;
        RECT 513.930 1418.490 515.110 1419.670 ;
        RECT 513.930 1240.090 515.110 1241.270 ;
        RECT 513.930 1238.490 515.110 1239.670 ;
        RECT 513.930 1060.090 515.110 1061.270 ;
        RECT 513.930 1058.490 515.110 1059.670 ;
        RECT 513.930 880.090 515.110 881.270 ;
        RECT 513.930 878.490 515.110 879.670 ;
        RECT 513.930 700.090 515.110 701.270 ;
        RECT 513.930 698.490 515.110 699.670 ;
        RECT 513.930 520.090 515.110 521.270 ;
        RECT 513.930 518.490 515.110 519.670 ;
        RECT 513.930 340.090 515.110 341.270 ;
        RECT 513.930 338.490 515.110 339.670 ;
        RECT 513.930 160.090 515.110 161.270 ;
        RECT 513.930 158.490 515.110 159.670 ;
        RECT 513.930 -35.810 515.110 -34.630 ;
        RECT 513.930 -37.410 515.110 -36.230 ;
        RECT 693.930 3555.910 695.110 3557.090 ;
        RECT 693.930 3554.310 695.110 3555.490 ;
        RECT 693.930 3400.090 695.110 3401.270 ;
        RECT 693.930 3398.490 695.110 3399.670 ;
        RECT 693.930 3220.090 695.110 3221.270 ;
        RECT 693.930 3218.490 695.110 3219.670 ;
        RECT 693.930 3040.090 695.110 3041.270 ;
        RECT 693.930 3038.490 695.110 3039.670 ;
        RECT 693.930 2860.090 695.110 2861.270 ;
        RECT 693.930 2858.490 695.110 2859.670 ;
        RECT 693.930 2680.090 695.110 2681.270 ;
        RECT 693.930 2678.490 695.110 2679.670 ;
        RECT 693.930 2500.090 695.110 2501.270 ;
        RECT 693.930 2498.490 695.110 2499.670 ;
        RECT 693.930 2320.090 695.110 2321.270 ;
        RECT 693.930 2318.490 695.110 2319.670 ;
        RECT 693.930 2140.090 695.110 2141.270 ;
        RECT 693.930 2138.490 695.110 2139.670 ;
        RECT 693.930 1960.090 695.110 1961.270 ;
        RECT 693.930 1958.490 695.110 1959.670 ;
        RECT 693.930 1780.090 695.110 1781.270 ;
        RECT 693.930 1778.490 695.110 1779.670 ;
        RECT 693.930 1600.090 695.110 1601.270 ;
        RECT 693.930 1598.490 695.110 1599.670 ;
        RECT 693.930 1420.090 695.110 1421.270 ;
        RECT 693.930 1418.490 695.110 1419.670 ;
        RECT 693.930 1240.090 695.110 1241.270 ;
        RECT 693.930 1238.490 695.110 1239.670 ;
        RECT 693.930 1060.090 695.110 1061.270 ;
        RECT 693.930 1058.490 695.110 1059.670 ;
        RECT 693.930 880.090 695.110 881.270 ;
        RECT 693.930 878.490 695.110 879.670 ;
        RECT 693.930 700.090 695.110 701.270 ;
        RECT 693.930 698.490 695.110 699.670 ;
        RECT 693.930 520.090 695.110 521.270 ;
        RECT 693.930 518.490 695.110 519.670 ;
        RECT 693.930 340.090 695.110 341.270 ;
        RECT 693.930 338.490 695.110 339.670 ;
        RECT 693.930 160.090 695.110 161.270 ;
        RECT 693.930 158.490 695.110 159.670 ;
        RECT 693.930 -35.810 695.110 -34.630 ;
        RECT 693.930 -37.410 695.110 -36.230 ;
        RECT 873.930 3555.910 875.110 3557.090 ;
        RECT 873.930 3554.310 875.110 3555.490 ;
        RECT 873.930 3400.090 875.110 3401.270 ;
        RECT 873.930 3398.490 875.110 3399.670 ;
        RECT 873.930 3220.090 875.110 3221.270 ;
        RECT 873.930 3218.490 875.110 3219.670 ;
        RECT 873.930 3040.090 875.110 3041.270 ;
        RECT 873.930 3038.490 875.110 3039.670 ;
        RECT 873.930 2860.090 875.110 2861.270 ;
        RECT 873.930 2858.490 875.110 2859.670 ;
        RECT 873.930 2680.090 875.110 2681.270 ;
        RECT 873.930 2678.490 875.110 2679.670 ;
        RECT 873.930 2500.090 875.110 2501.270 ;
        RECT 873.930 2498.490 875.110 2499.670 ;
        RECT 873.930 2320.090 875.110 2321.270 ;
        RECT 873.930 2318.490 875.110 2319.670 ;
        RECT 873.930 2140.090 875.110 2141.270 ;
        RECT 873.930 2138.490 875.110 2139.670 ;
        RECT 873.930 1960.090 875.110 1961.270 ;
        RECT 873.930 1958.490 875.110 1959.670 ;
        RECT 873.930 1780.090 875.110 1781.270 ;
        RECT 873.930 1778.490 875.110 1779.670 ;
        RECT 873.930 1600.090 875.110 1601.270 ;
        RECT 873.930 1598.490 875.110 1599.670 ;
        RECT 873.930 1420.090 875.110 1421.270 ;
        RECT 873.930 1418.490 875.110 1419.670 ;
        RECT 873.930 1240.090 875.110 1241.270 ;
        RECT 873.930 1238.490 875.110 1239.670 ;
        RECT 873.930 1060.090 875.110 1061.270 ;
        RECT 873.930 1058.490 875.110 1059.670 ;
        RECT 873.930 880.090 875.110 881.270 ;
        RECT 873.930 878.490 875.110 879.670 ;
        RECT 873.930 700.090 875.110 701.270 ;
        RECT 873.930 698.490 875.110 699.670 ;
        RECT 873.930 520.090 875.110 521.270 ;
        RECT 873.930 518.490 875.110 519.670 ;
        RECT 873.930 340.090 875.110 341.270 ;
        RECT 873.930 338.490 875.110 339.670 ;
        RECT 873.930 160.090 875.110 161.270 ;
        RECT 873.930 158.490 875.110 159.670 ;
        RECT 873.930 -35.810 875.110 -34.630 ;
        RECT 873.930 -37.410 875.110 -36.230 ;
        RECT 1053.930 3555.910 1055.110 3557.090 ;
        RECT 1053.930 3554.310 1055.110 3555.490 ;
        RECT 1053.930 3400.090 1055.110 3401.270 ;
        RECT 1053.930 3398.490 1055.110 3399.670 ;
        RECT 1053.930 3220.090 1055.110 3221.270 ;
        RECT 1053.930 3218.490 1055.110 3219.670 ;
        RECT 1053.930 3040.090 1055.110 3041.270 ;
        RECT 1053.930 3038.490 1055.110 3039.670 ;
        RECT 1053.930 2860.090 1055.110 2861.270 ;
        RECT 1053.930 2858.490 1055.110 2859.670 ;
        RECT 1053.930 2680.090 1055.110 2681.270 ;
        RECT 1053.930 2678.490 1055.110 2679.670 ;
        RECT 1053.930 2500.090 1055.110 2501.270 ;
        RECT 1053.930 2498.490 1055.110 2499.670 ;
        RECT 1053.930 2320.090 1055.110 2321.270 ;
        RECT 1053.930 2318.490 1055.110 2319.670 ;
        RECT 1053.930 2140.090 1055.110 2141.270 ;
        RECT 1053.930 2138.490 1055.110 2139.670 ;
        RECT 1053.930 1960.090 1055.110 1961.270 ;
        RECT 1053.930 1958.490 1055.110 1959.670 ;
        RECT 1053.930 1780.090 1055.110 1781.270 ;
        RECT 1053.930 1778.490 1055.110 1779.670 ;
        RECT 1053.930 1600.090 1055.110 1601.270 ;
        RECT 1053.930 1598.490 1055.110 1599.670 ;
        RECT 1053.930 1420.090 1055.110 1421.270 ;
        RECT 1053.930 1418.490 1055.110 1419.670 ;
        RECT 1053.930 1240.090 1055.110 1241.270 ;
        RECT 1053.930 1238.490 1055.110 1239.670 ;
        RECT 1053.930 1060.090 1055.110 1061.270 ;
        RECT 1053.930 1058.490 1055.110 1059.670 ;
        RECT 1053.930 880.090 1055.110 881.270 ;
        RECT 1053.930 878.490 1055.110 879.670 ;
        RECT 1053.930 700.090 1055.110 701.270 ;
        RECT 1053.930 698.490 1055.110 699.670 ;
        RECT 1053.930 520.090 1055.110 521.270 ;
        RECT 1053.930 518.490 1055.110 519.670 ;
        RECT 1053.930 340.090 1055.110 341.270 ;
        RECT 1053.930 338.490 1055.110 339.670 ;
        RECT 1053.930 160.090 1055.110 161.270 ;
        RECT 1053.930 158.490 1055.110 159.670 ;
        RECT 1053.930 -35.810 1055.110 -34.630 ;
        RECT 1053.930 -37.410 1055.110 -36.230 ;
        RECT 1233.930 3555.910 1235.110 3557.090 ;
        RECT 1233.930 3554.310 1235.110 3555.490 ;
        RECT 1233.930 3400.090 1235.110 3401.270 ;
        RECT 1233.930 3398.490 1235.110 3399.670 ;
        RECT 1233.930 3220.090 1235.110 3221.270 ;
        RECT 1233.930 3218.490 1235.110 3219.670 ;
        RECT 1233.930 3040.090 1235.110 3041.270 ;
        RECT 1233.930 3038.490 1235.110 3039.670 ;
        RECT 1233.930 2860.090 1235.110 2861.270 ;
        RECT 1233.930 2858.490 1235.110 2859.670 ;
        RECT 1233.930 2680.090 1235.110 2681.270 ;
        RECT 1233.930 2678.490 1235.110 2679.670 ;
        RECT 1233.930 2500.090 1235.110 2501.270 ;
        RECT 1233.930 2498.490 1235.110 2499.670 ;
        RECT 1233.930 2320.090 1235.110 2321.270 ;
        RECT 1233.930 2318.490 1235.110 2319.670 ;
        RECT 1233.930 2140.090 1235.110 2141.270 ;
        RECT 1233.930 2138.490 1235.110 2139.670 ;
        RECT 1233.930 1960.090 1235.110 1961.270 ;
        RECT 1233.930 1958.490 1235.110 1959.670 ;
        RECT 1233.930 1780.090 1235.110 1781.270 ;
        RECT 1233.930 1778.490 1235.110 1779.670 ;
        RECT 1233.930 1600.090 1235.110 1601.270 ;
        RECT 1233.930 1598.490 1235.110 1599.670 ;
        RECT 1233.930 1420.090 1235.110 1421.270 ;
        RECT 1233.930 1418.490 1235.110 1419.670 ;
        RECT 1233.930 1240.090 1235.110 1241.270 ;
        RECT 1233.930 1238.490 1235.110 1239.670 ;
        RECT 1233.930 1060.090 1235.110 1061.270 ;
        RECT 1233.930 1058.490 1235.110 1059.670 ;
        RECT 1233.930 880.090 1235.110 881.270 ;
        RECT 1233.930 878.490 1235.110 879.670 ;
        RECT 1233.930 700.090 1235.110 701.270 ;
        RECT 1233.930 698.490 1235.110 699.670 ;
        RECT 1233.930 520.090 1235.110 521.270 ;
        RECT 1233.930 518.490 1235.110 519.670 ;
        RECT 1233.930 340.090 1235.110 341.270 ;
        RECT 1233.930 338.490 1235.110 339.670 ;
        RECT 1233.930 160.090 1235.110 161.270 ;
        RECT 1233.930 158.490 1235.110 159.670 ;
        RECT 1233.930 -35.810 1235.110 -34.630 ;
        RECT 1233.930 -37.410 1235.110 -36.230 ;
        RECT 1413.930 3555.910 1415.110 3557.090 ;
        RECT 1413.930 3554.310 1415.110 3555.490 ;
        RECT 1413.930 3400.090 1415.110 3401.270 ;
        RECT 1413.930 3398.490 1415.110 3399.670 ;
        RECT 1413.930 3220.090 1415.110 3221.270 ;
        RECT 1413.930 3218.490 1415.110 3219.670 ;
        RECT 1413.930 3040.090 1415.110 3041.270 ;
        RECT 1413.930 3038.490 1415.110 3039.670 ;
        RECT 1413.930 2860.090 1415.110 2861.270 ;
        RECT 1413.930 2858.490 1415.110 2859.670 ;
        RECT 1413.930 2680.090 1415.110 2681.270 ;
        RECT 1413.930 2678.490 1415.110 2679.670 ;
        RECT 1413.930 2500.090 1415.110 2501.270 ;
        RECT 1413.930 2498.490 1415.110 2499.670 ;
        RECT 1413.930 2320.090 1415.110 2321.270 ;
        RECT 1413.930 2318.490 1415.110 2319.670 ;
        RECT 1413.930 2140.090 1415.110 2141.270 ;
        RECT 1413.930 2138.490 1415.110 2139.670 ;
        RECT 1413.930 1960.090 1415.110 1961.270 ;
        RECT 1413.930 1958.490 1415.110 1959.670 ;
        RECT 1413.930 1780.090 1415.110 1781.270 ;
        RECT 1413.930 1778.490 1415.110 1779.670 ;
        RECT 1413.930 1600.090 1415.110 1601.270 ;
        RECT 1413.930 1598.490 1415.110 1599.670 ;
        RECT 1413.930 1420.090 1415.110 1421.270 ;
        RECT 1413.930 1418.490 1415.110 1419.670 ;
        RECT 1413.930 1240.090 1415.110 1241.270 ;
        RECT 1413.930 1238.490 1415.110 1239.670 ;
        RECT 1413.930 1060.090 1415.110 1061.270 ;
        RECT 1413.930 1058.490 1415.110 1059.670 ;
        RECT 1413.930 880.090 1415.110 881.270 ;
        RECT 1413.930 878.490 1415.110 879.670 ;
        RECT 1413.930 700.090 1415.110 701.270 ;
        RECT 1413.930 698.490 1415.110 699.670 ;
        RECT 1413.930 520.090 1415.110 521.270 ;
        RECT 1413.930 518.490 1415.110 519.670 ;
        RECT 1413.930 340.090 1415.110 341.270 ;
        RECT 1413.930 338.490 1415.110 339.670 ;
        RECT 1413.930 160.090 1415.110 161.270 ;
        RECT 1413.930 158.490 1415.110 159.670 ;
        RECT 1413.930 -35.810 1415.110 -34.630 ;
        RECT 1413.930 -37.410 1415.110 -36.230 ;
        RECT 1593.930 3555.910 1595.110 3557.090 ;
        RECT 1593.930 3554.310 1595.110 3555.490 ;
        RECT 1593.930 3400.090 1595.110 3401.270 ;
        RECT 1593.930 3398.490 1595.110 3399.670 ;
        RECT 1593.930 3220.090 1595.110 3221.270 ;
        RECT 1593.930 3218.490 1595.110 3219.670 ;
        RECT 1593.930 3040.090 1595.110 3041.270 ;
        RECT 1593.930 3038.490 1595.110 3039.670 ;
        RECT 1593.930 2860.090 1595.110 2861.270 ;
        RECT 1593.930 2858.490 1595.110 2859.670 ;
        RECT 1593.930 2680.090 1595.110 2681.270 ;
        RECT 1593.930 2678.490 1595.110 2679.670 ;
        RECT 1593.930 2500.090 1595.110 2501.270 ;
        RECT 1593.930 2498.490 1595.110 2499.670 ;
        RECT 1593.930 2320.090 1595.110 2321.270 ;
        RECT 1593.930 2318.490 1595.110 2319.670 ;
        RECT 1593.930 2140.090 1595.110 2141.270 ;
        RECT 1593.930 2138.490 1595.110 2139.670 ;
        RECT 1593.930 1960.090 1595.110 1961.270 ;
        RECT 1593.930 1958.490 1595.110 1959.670 ;
        RECT 1593.930 1780.090 1595.110 1781.270 ;
        RECT 1593.930 1778.490 1595.110 1779.670 ;
        RECT 1593.930 1600.090 1595.110 1601.270 ;
        RECT 1593.930 1598.490 1595.110 1599.670 ;
        RECT 1593.930 1420.090 1595.110 1421.270 ;
        RECT 1593.930 1418.490 1595.110 1419.670 ;
        RECT 1593.930 1240.090 1595.110 1241.270 ;
        RECT 1593.930 1238.490 1595.110 1239.670 ;
        RECT 1593.930 1060.090 1595.110 1061.270 ;
        RECT 1593.930 1058.490 1595.110 1059.670 ;
        RECT 1593.930 880.090 1595.110 881.270 ;
        RECT 1593.930 878.490 1595.110 879.670 ;
        RECT 1593.930 700.090 1595.110 701.270 ;
        RECT 1593.930 698.490 1595.110 699.670 ;
        RECT 1593.930 520.090 1595.110 521.270 ;
        RECT 1593.930 518.490 1595.110 519.670 ;
        RECT 1593.930 340.090 1595.110 341.270 ;
        RECT 1593.930 338.490 1595.110 339.670 ;
        RECT 1593.930 160.090 1595.110 161.270 ;
        RECT 1593.930 158.490 1595.110 159.670 ;
        RECT 1593.930 -35.810 1595.110 -34.630 ;
        RECT 1593.930 -37.410 1595.110 -36.230 ;
        RECT 1773.930 3555.910 1775.110 3557.090 ;
        RECT 1773.930 3554.310 1775.110 3555.490 ;
        RECT 1773.930 3400.090 1775.110 3401.270 ;
        RECT 1773.930 3398.490 1775.110 3399.670 ;
        RECT 1773.930 3220.090 1775.110 3221.270 ;
        RECT 1773.930 3218.490 1775.110 3219.670 ;
        RECT 1773.930 3040.090 1775.110 3041.270 ;
        RECT 1773.930 3038.490 1775.110 3039.670 ;
        RECT 1773.930 2860.090 1775.110 2861.270 ;
        RECT 1773.930 2858.490 1775.110 2859.670 ;
        RECT 1773.930 2680.090 1775.110 2681.270 ;
        RECT 1773.930 2678.490 1775.110 2679.670 ;
        RECT 1773.930 2500.090 1775.110 2501.270 ;
        RECT 1773.930 2498.490 1775.110 2499.670 ;
        RECT 1773.930 2320.090 1775.110 2321.270 ;
        RECT 1773.930 2318.490 1775.110 2319.670 ;
        RECT 1773.930 2140.090 1775.110 2141.270 ;
        RECT 1773.930 2138.490 1775.110 2139.670 ;
        RECT 1773.930 1960.090 1775.110 1961.270 ;
        RECT 1773.930 1958.490 1775.110 1959.670 ;
        RECT 1773.930 1780.090 1775.110 1781.270 ;
        RECT 1773.930 1778.490 1775.110 1779.670 ;
        RECT 1773.930 1600.090 1775.110 1601.270 ;
        RECT 1773.930 1598.490 1775.110 1599.670 ;
        RECT 1773.930 1420.090 1775.110 1421.270 ;
        RECT 1773.930 1418.490 1775.110 1419.670 ;
        RECT 1773.930 1240.090 1775.110 1241.270 ;
        RECT 1773.930 1238.490 1775.110 1239.670 ;
        RECT 1773.930 1060.090 1775.110 1061.270 ;
        RECT 1773.930 1058.490 1775.110 1059.670 ;
        RECT 1773.930 880.090 1775.110 881.270 ;
        RECT 1773.930 878.490 1775.110 879.670 ;
        RECT 1773.930 700.090 1775.110 701.270 ;
        RECT 1773.930 698.490 1775.110 699.670 ;
        RECT 1773.930 520.090 1775.110 521.270 ;
        RECT 1773.930 518.490 1775.110 519.670 ;
        RECT 1773.930 340.090 1775.110 341.270 ;
        RECT 1773.930 338.490 1775.110 339.670 ;
        RECT 1773.930 160.090 1775.110 161.270 ;
        RECT 1773.930 158.490 1775.110 159.670 ;
        RECT 1773.930 -35.810 1775.110 -34.630 ;
        RECT 1773.930 -37.410 1775.110 -36.230 ;
        RECT 1953.930 3555.910 1955.110 3557.090 ;
        RECT 1953.930 3554.310 1955.110 3555.490 ;
        RECT 1953.930 3400.090 1955.110 3401.270 ;
        RECT 1953.930 3398.490 1955.110 3399.670 ;
        RECT 1953.930 3220.090 1955.110 3221.270 ;
        RECT 1953.930 3218.490 1955.110 3219.670 ;
        RECT 1953.930 3040.090 1955.110 3041.270 ;
        RECT 1953.930 3038.490 1955.110 3039.670 ;
        RECT 1953.930 2860.090 1955.110 2861.270 ;
        RECT 1953.930 2858.490 1955.110 2859.670 ;
        RECT 1953.930 2680.090 1955.110 2681.270 ;
        RECT 1953.930 2678.490 1955.110 2679.670 ;
        RECT 1953.930 2500.090 1955.110 2501.270 ;
        RECT 1953.930 2498.490 1955.110 2499.670 ;
        RECT 1953.930 2320.090 1955.110 2321.270 ;
        RECT 1953.930 2318.490 1955.110 2319.670 ;
        RECT 1953.930 2140.090 1955.110 2141.270 ;
        RECT 1953.930 2138.490 1955.110 2139.670 ;
        RECT 1953.930 1960.090 1955.110 1961.270 ;
        RECT 1953.930 1958.490 1955.110 1959.670 ;
        RECT 1953.930 1780.090 1955.110 1781.270 ;
        RECT 1953.930 1778.490 1955.110 1779.670 ;
        RECT 1953.930 1600.090 1955.110 1601.270 ;
        RECT 1953.930 1598.490 1955.110 1599.670 ;
        RECT 1953.930 1420.090 1955.110 1421.270 ;
        RECT 1953.930 1418.490 1955.110 1419.670 ;
        RECT 1953.930 1240.090 1955.110 1241.270 ;
        RECT 1953.930 1238.490 1955.110 1239.670 ;
        RECT 1953.930 1060.090 1955.110 1061.270 ;
        RECT 1953.930 1058.490 1955.110 1059.670 ;
        RECT 1953.930 880.090 1955.110 881.270 ;
        RECT 1953.930 878.490 1955.110 879.670 ;
        RECT 1953.930 700.090 1955.110 701.270 ;
        RECT 1953.930 698.490 1955.110 699.670 ;
        RECT 1953.930 520.090 1955.110 521.270 ;
        RECT 1953.930 518.490 1955.110 519.670 ;
        RECT 1953.930 340.090 1955.110 341.270 ;
        RECT 1953.930 338.490 1955.110 339.670 ;
        RECT 1953.930 160.090 1955.110 161.270 ;
        RECT 1953.930 158.490 1955.110 159.670 ;
        RECT 1953.930 -35.810 1955.110 -34.630 ;
        RECT 1953.930 -37.410 1955.110 -36.230 ;
        RECT 2133.930 3555.910 2135.110 3557.090 ;
        RECT 2133.930 3554.310 2135.110 3555.490 ;
        RECT 2133.930 3400.090 2135.110 3401.270 ;
        RECT 2133.930 3398.490 2135.110 3399.670 ;
        RECT 2133.930 3220.090 2135.110 3221.270 ;
        RECT 2133.930 3218.490 2135.110 3219.670 ;
        RECT 2133.930 3040.090 2135.110 3041.270 ;
        RECT 2133.930 3038.490 2135.110 3039.670 ;
        RECT 2133.930 2860.090 2135.110 2861.270 ;
        RECT 2133.930 2858.490 2135.110 2859.670 ;
        RECT 2133.930 2680.090 2135.110 2681.270 ;
        RECT 2133.930 2678.490 2135.110 2679.670 ;
        RECT 2133.930 2500.090 2135.110 2501.270 ;
        RECT 2133.930 2498.490 2135.110 2499.670 ;
        RECT 2133.930 2320.090 2135.110 2321.270 ;
        RECT 2133.930 2318.490 2135.110 2319.670 ;
        RECT 2133.930 2140.090 2135.110 2141.270 ;
        RECT 2133.930 2138.490 2135.110 2139.670 ;
        RECT 2133.930 1960.090 2135.110 1961.270 ;
        RECT 2133.930 1958.490 2135.110 1959.670 ;
        RECT 2133.930 1780.090 2135.110 1781.270 ;
        RECT 2133.930 1778.490 2135.110 1779.670 ;
        RECT 2133.930 1600.090 2135.110 1601.270 ;
        RECT 2133.930 1598.490 2135.110 1599.670 ;
        RECT 2133.930 1420.090 2135.110 1421.270 ;
        RECT 2133.930 1418.490 2135.110 1419.670 ;
        RECT 2133.930 1240.090 2135.110 1241.270 ;
        RECT 2133.930 1238.490 2135.110 1239.670 ;
        RECT 2133.930 1060.090 2135.110 1061.270 ;
        RECT 2133.930 1058.490 2135.110 1059.670 ;
        RECT 2133.930 880.090 2135.110 881.270 ;
        RECT 2133.930 878.490 2135.110 879.670 ;
        RECT 2133.930 700.090 2135.110 701.270 ;
        RECT 2133.930 698.490 2135.110 699.670 ;
        RECT 2133.930 520.090 2135.110 521.270 ;
        RECT 2133.930 518.490 2135.110 519.670 ;
        RECT 2133.930 340.090 2135.110 341.270 ;
        RECT 2133.930 338.490 2135.110 339.670 ;
        RECT 2133.930 160.090 2135.110 161.270 ;
        RECT 2133.930 158.490 2135.110 159.670 ;
        RECT 2133.930 -35.810 2135.110 -34.630 ;
        RECT 2133.930 -37.410 2135.110 -36.230 ;
        RECT 2313.930 3555.910 2315.110 3557.090 ;
        RECT 2313.930 3554.310 2315.110 3555.490 ;
        RECT 2313.930 3400.090 2315.110 3401.270 ;
        RECT 2313.930 3398.490 2315.110 3399.670 ;
        RECT 2313.930 3220.090 2315.110 3221.270 ;
        RECT 2313.930 3218.490 2315.110 3219.670 ;
        RECT 2313.930 3040.090 2315.110 3041.270 ;
        RECT 2313.930 3038.490 2315.110 3039.670 ;
        RECT 2313.930 2860.090 2315.110 2861.270 ;
        RECT 2313.930 2858.490 2315.110 2859.670 ;
        RECT 2313.930 2680.090 2315.110 2681.270 ;
        RECT 2313.930 2678.490 2315.110 2679.670 ;
        RECT 2313.930 2500.090 2315.110 2501.270 ;
        RECT 2313.930 2498.490 2315.110 2499.670 ;
        RECT 2313.930 2320.090 2315.110 2321.270 ;
        RECT 2313.930 2318.490 2315.110 2319.670 ;
        RECT 2313.930 2140.090 2315.110 2141.270 ;
        RECT 2313.930 2138.490 2315.110 2139.670 ;
        RECT 2313.930 1960.090 2315.110 1961.270 ;
        RECT 2313.930 1958.490 2315.110 1959.670 ;
        RECT 2313.930 1780.090 2315.110 1781.270 ;
        RECT 2313.930 1778.490 2315.110 1779.670 ;
        RECT 2313.930 1600.090 2315.110 1601.270 ;
        RECT 2313.930 1598.490 2315.110 1599.670 ;
        RECT 2313.930 1420.090 2315.110 1421.270 ;
        RECT 2313.930 1418.490 2315.110 1419.670 ;
        RECT 2313.930 1240.090 2315.110 1241.270 ;
        RECT 2313.930 1238.490 2315.110 1239.670 ;
        RECT 2313.930 1060.090 2315.110 1061.270 ;
        RECT 2313.930 1058.490 2315.110 1059.670 ;
        RECT 2313.930 880.090 2315.110 881.270 ;
        RECT 2313.930 878.490 2315.110 879.670 ;
        RECT 2313.930 700.090 2315.110 701.270 ;
        RECT 2313.930 698.490 2315.110 699.670 ;
        RECT 2313.930 520.090 2315.110 521.270 ;
        RECT 2313.930 518.490 2315.110 519.670 ;
        RECT 2313.930 340.090 2315.110 341.270 ;
        RECT 2313.930 338.490 2315.110 339.670 ;
        RECT 2313.930 160.090 2315.110 161.270 ;
        RECT 2313.930 158.490 2315.110 159.670 ;
        RECT 2313.930 -35.810 2315.110 -34.630 ;
        RECT 2313.930 -37.410 2315.110 -36.230 ;
        RECT 2493.930 3555.910 2495.110 3557.090 ;
        RECT 2493.930 3554.310 2495.110 3555.490 ;
        RECT 2493.930 3400.090 2495.110 3401.270 ;
        RECT 2493.930 3398.490 2495.110 3399.670 ;
        RECT 2493.930 3220.090 2495.110 3221.270 ;
        RECT 2493.930 3218.490 2495.110 3219.670 ;
        RECT 2493.930 3040.090 2495.110 3041.270 ;
        RECT 2493.930 3038.490 2495.110 3039.670 ;
        RECT 2493.930 2860.090 2495.110 2861.270 ;
        RECT 2493.930 2858.490 2495.110 2859.670 ;
        RECT 2493.930 2680.090 2495.110 2681.270 ;
        RECT 2493.930 2678.490 2495.110 2679.670 ;
        RECT 2493.930 2500.090 2495.110 2501.270 ;
        RECT 2493.930 2498.490 2495.110 2499.670 ;
        RECT 2493.930 2320.090 2495.110 2321.270 ;
        RECT 2493.930 2318.490 2495.110 2319.670 ;
        RECT 2493.930 2140.090 2495.110 2141.270 ;
        RECT 2493.930 2138.490 2495.110 2139.670 ;
        RECT 2493.930 1960.090 2495.110 1961.270 ;
        RECT 2493.930 1958.490 2495.110 1959.670 ;
        RECT 2493.930 1780.090 2495.110 1781.270 ;
        RECT 2493.930 1778.490 2495.110 1779.670 ;
        RECT 2493.930 1600.090 2495.110 1601.270 ;
        RECT 2493.930 1598.490 2495.110 1599.670 ;
        RECT 2493.930 1420.090 2495.110 1421.270 ;
        RECT 2493.930 1418.490 2495.110 1419.670 ;
        RECT 2493.930 1240.090 2495.110 1241.270 ;
        RECT 2493.930 1238.490 2495.110 1239.670 ;
        RECT 2493.930 1060.090 2495.110 1061.270 ;
        RECT 2493.930 1058.490 2495.110 1059.670 ;
        RECT 2493.930 880.090 2495.110 881.270 ;
        RECT 2493.930 878.490 2495.110 879.670 ;
        RECT 2493.930 700.090 2495.110 701.270 ;
        RECT 2493.930 698.490 2495.110 699.670 ;
        RECT 2493.930 520.090 2495.110 521.270 ;
        RECT 2493.930 518.490 2495.110 519.670 ;
        RECT 2493.930 340.090 2495.110 341.270 ;
        RECT 2493.930 338.490 2495.110 339.670 ;
        RECT 2493.930 160.090 2495.110 161.270 ;
        RECT 2493.930 158.490 2495.110 159.670 ;
        RECT 2493.930 -35.810 2495.110 -34.630 ;
        RECT 2493.930 -37.410 2495.110 -36.230 ;
        RECT 2673.930 3555.910 2675.110 3557.090 ;
        RECT 2673.930 3554.310 2675.110 3555.490 ;
        RECT 2673.930 3400.090 2675.110 3401.270 ;
        RECT 2673.930 3398.490 2675.110 3399.670 ;
        RECT 2673.930 3220.090 2675.110 3221.270 ;
        RECT 2673.930 3218.490 2675.110 3219.670 ;
        RECT 2673.930 3040.090 2675.110 3041.270 ;
        RECT 2673.930 3038.490 2675.110 3039.670 ;
        RECT 2673.930 2860.090 2675.110 2861.270 ;
        RECT 2673.930 2858.490 2675.110 2859.670 ;
        RECT 2673.930 2680.090 2675.110 2681.270 ;
        RECT 2673.930 2678.490 2675.110 2679.670 ;
        RECT 2673.930 2500.090 2675.110 2501.270 ;
        RECT 2673.930 2498.490 2675.110 2499.670 ;
        RECT 2673.930 2320.090 2675.110 2321.270 ;
        RECT 2673.930 2318.490 2675.110 2319.670 ;
        RECT 2673.930 2140.090 2675.110 2141.270 ;
        RECT 2673.930 2138.490 2675.110 2139.670 ;
        RECT 2673.930 1960.090 2675.110 1961.270 ;
        RECT 2673.930 1958.490 2675.110 1959.670 ;
        RECT 2673.930 1780.090 2675.110 1781.270 ;
        RECT 2673.930 1778.490 2675.110 1779.670 ;
        RECT 2673.930 1600.090 2675.110 1601.270 ;
        RECT 2673.930 1598.490 2675.110 1599.670 ;
        RECT 2673.930 1420.090 2675.110 1421.270 ;
        RECT 2673.930 1418.490 2675.110 1419.670 ;
        RECT 2673.930 1240.090 2675.110 1241.270 ;
        RECT 2673.930 1238.490 2675.110 1239.670 ;
        RECT 2673.930 1060.090 2675.110 1061.270 ;
        RECT 2673.930 1058.490 2675.110 1059.670 ;
        RECT 2673.930 880.090 2675.110 881.270 ;
        RECT 2673.930 878.490 2675.110 879.670 ;
        RECT 2673.930 700.090 2675.110 701.270 ;
        RECT 2673.930 698.490 2675.110 699.670 ;
        RECT 2673.930 520.090 2675.110 521.270 ;
        RECT 2673.930 518.490 2675.110 519.670 ;
        RECT 2673.930 340.090 2675.110 341.270 ;
        RECT 2673.930 338.490 2675.110 339.670 ;
        RECT 2673.930 160.090 2675.110 161.270 ;
        RECT 2673.930 158.490 2675.110 159.670 ;
        RECT 2673.930 -35.810 2675.110 -34.630 ;
        RECT 2673.930 -37.410 2675.110 -36.230 ;
        RECT 2853.930 3555.910 2855.110 3557.090 ;
        RECT 2853.930 3554.310 2855.110 3555.490 ;
        RECT 2853.930 3400.090 2855.110 3401.270 ;
        RECT 2853.930 3398.490 2855.110 3399.670 ;
        RECT 2853.930 3220.090 2855.110 3221.270 ;
        RECT 2853.930 3218.490 2855.110 3219.670 ;
        RECT 2853.930 3040.090 2855.110 3041.270 ;
        RECT 2853.930 3038.490 2855.110 3039.670 ;
        RECT 2853.930 2860.090 2855.110 2861.270 ;
        RECT 2853.930 2858.490 2855.110 2859.670 ;
        RECT 2853.930 2680.090 2855.110 2681.270 ;
        RECT 2853.930 2678.490 2855.110 2679.670 ;
        RECT 2853.930 2500.090 2855.110 2501.270 ;
        RECT 2853.930 2498.490 2855.110 2499.670 ;
        RECT 2853.930 2320.090 2855.110 2321.270 ;
        RECT 2853.930 2318.490 2855.110 2319.670 ;
        RECT 2853.930 2140.090 2855.110 2141.270 ;
        RECT 2853.930 2138.490 2855.110 2139.670 ;
        RECT 2853.930 1960.090 2855.110 1961.270 ;
        RECT 2853.930 1958.490 2855.110 1959.670 ;
        RECT 2853.930 1780.090 2855.110 1781.270 ;
        RECT 2853.930 1778.490 2855.110 1779.670 ;
        RECT 2853.930 1600.090 2855.110 1601.270 ;
        RECT 2853.930 1598.490 2855.110 1599.670 ;
        RECT 2853.930 1420.090 2855.110 1421.270 ;
        RECT 2853.930 1418.490 2855.110 1419.670 ;
        RECT 2853.930 1240.090 2855.110 1241.270 ;
        RECT 2853.930 1238.490 2855.110 1239.670 ;
        RECT 2853.930 1060.090 2855.110 1061.270 ;
        RECT 2853.930 1058.490 2855.110 1059.670 ;
        RECT 2853.930 880.090 2855.110 881.270 ;
        RECT 2853.930 878.490 2855.110 879.670 ;
        RECT 2853.930 700.090 2855.110 701.270 ;
        RECT 2853.930 698.490 2855.110 699.670 ;
        RECT 2853.930 520.090 2855.110 521.270 ;
        RECT 2853.930 518.490 2855.110 519.670 ;
        RECT 2853.930 340.090 2855.110 341.270 ;
        RECT 2853.930 338.490 2855.110 339.670 ;
        RECT 2853.930 160.090 2855.110 161.270 ;
        RECT 2853.930 158.490 2855.110 159.670 ;
        RECT 2853.930 -35.810 2855.110 -34.630 ;
        RECT 2853.930 -37.410 2855.110 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 3400.090 2961.590 3401.270 ;
        RECT 2960.410 3398.490 2961.590 3399.670 ;
        RECT 2960.410 3220.090 2961.590 3221.270 ;
        RECT 2960.410 3218.490 2961.590 3219.670 ;
        RECT 2960.410 3040.090 2961.590 3041.270 ;
        RECT 2960.410 3038.490 2961.590 3039.670 ;
        RECT 2960.410 2860.090 2961.590 2861.270 ;
        RECT 2960.410 2858.490 2961.590 2859.670 ;
        RECT 2960.410 2680.090 2961.590 2681.270 ;
        RECT 2960.410 2678.490 2961.590 2679.670 ;
        RECT 2960.410 2500.090 2961.590 2501.270 ;
        RECT 2960.410 2498.490 2961.590 2499.670 ;
        RECT 2960.410 2320.090 2961.590 2321.270 ;
        RECT 2960.410 2318.490 2961.590 2319.670 ;
        RECT 2960.410 2140.090 2961.590 2141.270 ;
        RECT 2960.410 2138.490 2961.590 2139.670 ;
        RECT 2960.410 1960.090 2961.590 1961.270 ;
        RECT 2960.410 1958.490 2961.590 1959.670 ;
        RECT 2960.410 1780.090 2961.590 1781.270 ;
        RECT 2960.410 1778.490 2961.590 1779.670 ;
        RECT 2960.410 1600.090 2961.590 1601.270 ;
        RECT 2960.410 1598.490 2961.590 1599.670 ;
        RECT 2960.410 1420.090 2961.590 1421.270 ;
        RECT 2960.410 1418.490 2961.590 1419.670 ;
        RECT 2960.410 1240.090 2961.590 1241.270 ;
        RECT 2960.410 1238.490 2961.590 1239.670 ;
        RECT 2960.410 1060.090 2961.590 1061.270 ;
        RECT 2960.410 1058.490 2961.590 1059.670 ;
        RECT 2960.410 880.090 2961.590 881.270 ;
        RECT 2960.410 878.490 2961.590 879.670 ;
        RECT 2960.410 700.090 2961.590 701.270 ;
        RECT 2960.410 698.490 2961.590 699.670 ;
        RECT 2960.410 520.090 2961.590 521.270 ;
        RECT 2960.410 518.490 2961.590 519.670 ;
        RECT 2960.410 340.090 2961.590 341.270 ;
        RECT 2960.410 338.490 2961.590 339.670 ;
        RECT 2960.410 160.090 2961.590 161.270 ;
        RECT 2960.410 158.490 2961.590 159.670 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 153.020 3557.200 156.020 3557.210 ;
        RECT 333.020 3557.200 336.020 3557.210 ;
        RECT 513.020 3557.200 516.020 3557.210 ;
        RECT 693.020 3557.200 696.020 3557.210 ;
        RECT 873.020 3557.200 876.020 3557.210 ;
        RECT 1053.020 3557.200 1056.020 3557.210 ;
        RECT 1233.020 3557.200 1236.020 3557.210 ;
        RECT 1413.020 3557.200 1416.020 3557.210 ;
        RECT 1593.020 3557.200 1596.020 3557.210 ;
        RECT 1773.020 3557.200 1776.020 3557.210 ;
        RECT 1953.020 3557.200 1956.020 3557.210 ;
        RECT 2133.020 3557.200 2136.020 3557.210 ;
        RECT 2313.020 3557.200 2316.020 3557.210 ;
        RECT 2493.020 3557.200 2496.020 3557.210 ;
        RECT 2673.020 3557.200 2676.020 3557.210 ;
        RECT 2853.020 3557.200 2856.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 153.020 3554.190 156.020 3554.200 ;
        RECT 333.020 3554.190 336.020 3554.200 ;
        RECT 513.020 3554.190 516.020 3554.200 ;
        RECT 693.020 3554.190 696.020 3554.200 ;
        RECT 873.020 3554.190 876.020 3554.200 ;
        RECT 1053.020 3554.190 1056.020 3554.200 ;
        RECT 1233.020 3554.190 1236.020 3554.200 ;
        RECT 1413.020 3554.190 1416.020 3554.200 ;
        RECT 1593.020 3554.190 1596.020 3554.200 ;
        RECT 1773.020 3554.190 1776.020 3554.200 ;
        RECT 1953.020 3554.190 1956.020 3554.200 ;
        RECT 2133.020 3554.190 2136.020 3554.200 ;
        RECT 2313.020 3554.190 2316.020 3554.200 ;
        RECT 2493.020 3554.190 2496.020 3554.200 ;
        RECT 2673.020 3554.190 2676.020 3554.200 ;
        RECT 2853.020 3554.190 2856.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3401.380 -39.880 3401.390 ;
        RECT 153.020 3401.380 156.020 3401.390 ;
        RECT 333.020 3401.380 336.020 3401.390 ;
        RECT 513.020 3401.380 516.020 3401.390 ;
        RECT 693.020 3401.380 696.020 3401.390 ;
        RECT 873.020 3401.380 876.020 3401.390 ;
        RECT 1053.020 3401.380 1056.020 3401.390 ;
        RECT 1233.020 3401.380 1236.020 3401.390 ;
        RECT 1413.020 3401.380 1416.020 3401.390 ;
        RECT 1593.020 3401.380 1596.020 3401.390 ;
        RECT 1773.020 3401.380 1776.020 3401.390 ;
        RECT 1953.020 3401.380 1956.020 3401.390 ;
        RECT 2133.020 3401.380 2136.020 3401.390 ;
        RECT 2313.020 3401.380 2316.020 3401.390 ;
        RECT 2493.020 3401.380 2496.020 3401.390 ;
        RECT 2673.020 3401.380 2676.020 3401.390 ;
        RECT 2853.020 3401.380 2856.020 3401.390 ;
        RECT 2959.500 3401.380 2962.500 3401.390 ;
        RECT -42.880 3398.380 2962.500 3401.380 ;
        RECT -42.880 3398.370 -39.880 3398.380 ;
        RECT 153.020 3398.370 156.020 3398.380 ;
        RECT 333.020 3398.370 336.020 3398.380 ;
        RECT 513.020 3398.370 516.020 3398.380 ;
        RECT 693.020 3398.370 696.020 3398.380 ;
        RECT 873.020 3398.370 876.020 3398.380 ;
        RECT 1053.020 3398.370 1056.020 3398.380 ;
        RECT 1233.020 3398.370 1236.020 3398.380 ;
        RECT 1413.020 3398.370 1416.020 3398.380 ;
        RECT 1593.020 3398.370 1596.020 3398.380 ;
        RECT 1773.020 3398.370 1776.020 3398.380 ;
        RECT 1953.020 3398.370 1956.020 3398.380 ;
        RECT 2133.020 3398.370 2136.020 3398.380 ;
        RECT 2313.020 3398.370 2316.020 3398.380 ;
        RECT 2493.020 3398.370 2496.020 3398.380 ;
        RECT 2673.020 3398.370 2676.020 3398.380 ;
        RECT 2853.020 3398.370 2856.020 3398.380 ;
        RECT 2959.500 3398.370 2962.500 3398.380 ;
        RECT -42.880 3221.380 -39.880 3221.390 ;
        RECT 153.020 3221.380 156.020 3221.390 ;
        RECT 333.020 3221.380 336.020 3221.390 ;
        RECT 513.020 3221.380 516.020 3221.390 ;
        RECT 693.020 3221.380 696.020 3221.390 ;
        RECT 873.020 3221.380 876.020 3221.390 ;
        RECT 1053.020 3221.380 1056.020 3221.390 ;
        RECT 1233.020 3221.380 1236.020 3221.390 ;
        RECT 1413.020 3221.380 1416.020 3221.390 ;
        RECT 1593.020 3221.380 1596.020 3221.390 ;
        RECT 1773.020 3221.380 1776.020 3221.390 ;
        RECT 1953.020 3221.380 1956.020 3221.390 ;
        RECT 2133.020 3221.380 2136.020 3221.390 ;
        RECT 2313.020 3221.380 2316.020 3221.390 ;
        RECT 2493.020 3221.380 2496.020 3221.390 ;
        RECT 2673.020 3221.380 2676.020 3221.390 ;
        RECT 2853.020 3221.380 2856.020 3221.390 ;
        RECT 2959.500 3221.380 2962.500 3221.390 ;
        RECT -42.880 3218.380 2962.500 3221.380 ;
        RECT -42.880 3218.370 -39.880 3218.380 ;
        RECT 153.020 3218.370 156.020 3218.380 ;
        RECT 333.020 3218.370 336.020 3218.380 ;
        RECT 513.020 3218.370 516.020 3218.380 ;
        RECT 693.020 3218.370 696.020 3218.380 ;
        RECT 873.020 3218.370 876.020 3218.380 ;
        RECT 1053.020 3218.370 1056.020 3218.380 ;
        RECT 1233.020 3218.370 1236.020 3218.380 ;
        RECT 1413.020 3218.370 1416.020 3218.380 ;
        RECT 1593.020 3218.370 1596.020 3218.380 ;
        RECT 1773.020 3218.370 1776.020 3218.380 ;
        RECT 1953.020 3218.370 1956.020 3218.380 ;
        RECT 2133.020 3218.370 2136.020 3218.380 ;
        RECT 2313.020 3218.370 2316.020 3218.380 ;
        RECT 2493.020 3218.370 2496.020 3218.380 ;
        RECT 2673.020 3218.370 2676.020 3218.380 ;
        RECT 2853.020 3218.370 2856.020 3218.380 ;
        RECT 2959.500 3218.370 2962.500 3218.380 ;
        RECT -42.880 3041.380 -39.880 3041.390 ;
        RECT 153.020 3041.380 156.020 3041.390 ;
        RECT 333.020 3041.380 336.020 3041.390 ;
        RECT 513.020 3041.380 516.020 3041.390 ;
        RECT 693.020 3041.380 696.020 3041.390 ;
        RECT 873.020 3041.380 876.020 3041.390 ;
        RECT 1053.020 3041.380 1056.020 3041.390 ;
        RECT 1233.020 3041.380 1236.020 3041.390 ;
        RECT 1413.020 3041.380 1416.020 3041.390 ;
        RECT 1593.020 3041.380 1596.020 3041.390 ;
        RECT 1773.020 3041.380 1776.020 3041.390 ;
        RECT 1953.020 3041.380 1956.020 3041.390 ;
        RECT 2133.020 3041.380 2136.020 3041.390 ;
        RECT 2313.020 3041.380 2316.020 3041.390 ;
        RECT 2493.020 3041.380 2496.020 3041.390 ;
        RECT 2673.020 3041.380 2676.020 3041.390 ;
        RECT 2853.020 3041.380 2856.020 3041.390 ;
        RECT 2959.500 3041.380 2962.500 3041.390 ;
        RECT -42.880 3038.380 2962.500 3041.380 ;
        RECT -42.880 3038.370 -39.880 3038.380 ;
        RECT 153.020 3038.370 156.020 3038.380 ;
        RECT 333.020 3038.370 336.020 3038.380 ;
        RECT 513.020 3038.370 516.020 3038.380 ;
        RECT 693.020 3038.370 696.020 3038.380 ;
        RECT 873.020 3038.370 876.020 3038.380 ;
        RECT 1053.020 3038.370 1056.020 3038.380 ;
        RECT 1233.020 3038.370 1236.020 3038.380 ;
        RECT 1413.020 3038.370 1416.020 3038.380 ;
        RECT 1593.020 3038.370 1596.020 3038.380 ;
        RECT 1773.020 3038.370 1776.020 3038.380 ;
        RECT 1953.020 3038.370 1956.020 3038.380 ;
        RECT 2133.020 3038.370 2136.020 3038.380 ;
        RECT 2313.020 3038.370 2316.020 3038.380 ;
        RECT 2493.020 3038.370 2496.020 3038.380 ;
        RECT 2673.020 3038.370 2676.020 3038.380 ;
        RECT 2853.020 3038.370 2856.020 3038.380 ;
        RECT 2959.500 3038.370 2962.500 3038.380 ;
        RECT -42.880 2861.380 -39.880 2861.390 ;
        RECT 153.020 2861.380 156.020 2861.390 ;
        RECT 333.020 2861.380 336.020 2861.390 ;
        RECT 513.020 2861.380 516.020 2861.390 ;
        RECT 693.020 2861.380 696.020 2861.390 ;
        RECT 873.020 2861.380 876.020 2861.390 ;
        RECT 1053.020 2861.380 1056.020 2861.390 ;
        RECT 1233.020 2861.380 1236.020 2861.390 ;
        RECT 1413.020 2861.380 1416.020 2861.390 ;
        RECT 1593.020 2861.380 1596.020 2861.390 ;
        RECT 1773.020 2861.380 1776.020 2861.390 ;
        RECT 1953.020 2861.380 1956.020 2861.390 ;
        RECT 2133.020 2861.380 2136.020 2861.390 ;
        RECT 2313.020 2861.380 2316.020 2861.390 ;
        RECT 2493.020 2861.380 2496.020 2861.390 ;
        RECT 2673.020 2861.380 2676.020 2861.390 ;
        RECT 2853.020 2861.380 2856.020 2861.390 ;
        RECT 2959.500 2861.380 2962.500 2861.390 ;
        RECT -42.880 2858.380 2962.500 2861.380 ;
        RECT -42.880 2858.370 -39.880 2858.380 ;
        RECT 153.020 2858.370 156.020 2858.380 ;
        RECT 333.020 2858.370 336.020 2858.380 ;
        RECT 513.020 2858.370 516.020 2858.380 ;
        RECT 693.020 2858.370 696.020 2858.380 ;
        RECT 873.020 2858.370 876.020 2858.380 ;
        RECT 1053.020 2858.370 1056.020 2858.380 ;
        RECT 1233.020 2858.370 1236.020 2858.380 ;
        RECT 1413.020 2858.370 1416.020 2858.380 ;
        RECT 1593.020 2858.370 1596.020 2858.380 ;
        RECT 1773.020 2858.370 1776.020 2858.380 ;
        RECT 1953.020 2858.370 1956.020 2858.380 ;
        RECT 2133.020 2858.370 2136.020 2858.380 ;
        RECT 2313.020 2858.370 2316.020 2858.380 ;
        RECT 2493.020 2858.370 2496.020 2858.380 ;
        RECT 2673.020 2858.370 2676.020 2858.380 ;
        RECT 2853.020 2858.370 2856.020 2858.380 ;
        RECT 2959.500 2858.370 2962.500 2858.380 ;
        RECT -42.880 2681.380 -39.880 2681.390 ;
        RECT 153.020 2681.380 156.020 2681.390 ;
        RECT 333.020 2681.380 336.020 2681.390 ;
        RECT 513.020 2681.380 516.020 2681.390 ;
        RECT 693.020 2681.380 696.020 2681.390 ;
        RECT 873.020 2681.380 876.020 2681.390 ;
        RECT 1053.020 2681.380 1056.020 2681.390 ;
        RECT 1233.020 2681.380 1236.020 2681.390 ;
        RECT 1413.020 2681.380 1416.020 2681.390 ;
        RECT 1593.020 2681.380 1596.020 2681.390 ;
        RECT 1773.020 2681.380 1776.020 2681.390 ;
        RECT 1953.020 2681.380 1956.020 2681.390 ;
        RECT 2133.020 2681.380 2136.020 2681.390 ;
        RECT 2313.020 2681.380 2316.020 2681.390 ;
        RECT 2493.020 2681.380 2496.020 2681.390 ;
        RECT 2673.020 2681.380 2676.020 2681.390 ;
        RECT 2853.020 2681.380 2856.020 2681.390 ;
        RECT 2959.500 2681.380 2962.500 2681.390 ;
        RECT -42.880 2678.380 2962.500 2681.380 ;
        RECT -42.880 2678.370 -39.880 2678.380 ;
        RECT 153.020 2678.370 156.020 2678.380 ;
        RECT 333.020 2678.370 336.020 2678.380 ;
        RECT 513.020 2678.370 516.020 2678.380 ;
        RECT 693.020 2678.370 696.020 2678.380 ;
        RECT 873.020 2678.370 876.020 2678.380 ;
        RECT 1053.020 2678.370 1056.020 2678.380 ;
        RECT 1233.020 2678.370 1236.020 2678.380 ;
        RECT 1413.020 2678.370 1416.020 2678.380 ;
        RECT 1593.020 2678.370 1596.020 2678.380 ;
        RECT 1773.020 2678.370 1776.020 2678.380 ;
        RECT 1953.020 2678.370 1956.020 2678.380 ;
        RECT 2133.020 2678.370 2136.020 2678.380 ;
        RECT 2313.020 2678.370 2316.020 2678.380 ;
        RECT 2493.020 2678.370 2496.020 2678.380 ;
        RECT 2673.020 2678.370 2676.020 2678.380 ;
        RECT 2853.020 2678.370 2856.020 2678.380 ;
        RECT 2959.500 2678.370 2962.500 2678.380 ;
        RECT -42.880 2501.380 -39.880 2501.390 ;
        RECT 153.020 2501.380 156.020 2501.390 ;
        RECT 333.020 2501.380 336.020 2501.390 ;
        RECT 513.020 2501.380 516.020 2501.390 ;
        RECT 693.020 2501.380 696.020 2501.390 ;
        RECT 873.020 2501.380 876.020 2501.390 ;
        RECT 1053.020 2501.380 1056.020 2501.390 ;
        RECT 1233.020 2501.380 1236.020 2501.390 ;
        RECT 1413.020 2501.380 1416.020 2501.390 ;
        RECT 1593.020 2501.380 1596.020 2501.390 ;
        RECT 1773.020 2501.380 1776.020 2501.390 ;
        RECT 1953.020 2501.380 1956.020 2501.390 ;
        RECT 2133.020 2501.380 2136.020 2501.390 ;
        RECT 2313.020 2501.380 2316.020 2501.390 ;
        RECT 2493.020 2501.380 2496.020 2501.390 ;
        RECT 2673.020 2501.380 2676.020 2501.390 ;
        RECT 2853.020 2501.380 2856.020 2501.390 ;
        RECT 2959.500 2501.380 2962.500 2501.390 ;
        RECT -42.880 2498.380 2962.500 2501.380 ;
        RECT -42.880 2498.370 -39.880 2498.380 ;
        RECT 153.020 2498.370 156.020 2498.380 ;
        RECT 333.020 2498.370 336.020 2498.380 ;
        RECT 513.020 2498.370 516.020 2498.380 ;
        RECT 693.020 2498.370 696.020 2498.380 ;
        RECT 873.020 2498.370 876.020 2498.380 ;
        RECT 1053.020 2498.370 1056.020 2498.380 ;
        RECT 1233.020 2498.370 1236.020 2498.380 ;
        RECT 1413.020 2498.370 1416.020 2498.380 ;
        RECT 1593.020 2498.370 1596.020 2498.380 ;
        RECT 1773.020 2498.370 1776.020 2498.380 ;
        RECT 1953.020 2498.370 1956.020 2498.380 ;
        RECT 2133.020 2498.370 2136.020 2498.380 ;
        RECT 2313.020 2498.370 2316.020 2498.380 ;
        RECT 2493.020 2498.370 2496.020 2498.380 ;
        RECT 2673.020 2498.370 2676.020 2498.380 ;
        RECT 2853.020 2498.370 2856.020 2498.380 ;
        RECT 2959.500 2498.370 2962.500 2498.380 ;
        RECT -42.880 2321.380 -39.880 2321.390 ;
        RECT 153.020 2321.380 156.020 2321.390 ;
        RECT 333.020 2321.380 336.020 2321.390 ;
        RECT 513.020 2321.380 516.020 2321.390 ;
        RECT 693.020 2321.380 696.020 2321.390 ;
        RECT 873.020 2321.380 876.020 2321.390 ;
        RECT 1053.020 2321.380 1056.020 2321.390 ;
        RECT 1233.020 2321.380 1236.020 2321.390 ;
        RECT 1413.020 2321.380 1416.020 2321.390 ;
        RECT 1593.020 2321.380 1596.020 2321.390 ;
        RECT 1773.020 2321.380 1776.020 2321.390 ;
        RECT 1953.020 2321.380 1956.020 2321.390 ;
        RECT 2133.020 2321.380 2136.020 2321.390 ;
        RECT 2313.020 2321.380 2316.020 2321.390 ;
        RECT 2493.020 2321.380 2496.020 2321.390 ;
        RECT 2673.020 2321.380 2676.020 2321.390 ;
        RECT 2853.020 2321.380 2856.020 2321.390 ;
        RECT 2959.500 2321.380 2962.500 2321.390 ;
        RECT -42.880 2318.380 2962.500 2321.380 ;
        RECT -42.880 2318.370 -39.880 2318.380 ;
        RECT 153.020 2318.370 156.020 2318.380 ;
        RECT 333.020 2318.370 336.020 2318.380 ;
        RECT 513.020 2318.370 516.020 2318.380 ;
        RECT 693.020 2318.370 696.020 2318.380 ;
        RECT 873.020 2318.370 876.020 2318.380 ;
        RECT 1053.020 2318.370 1056.020 2318.380 ;
        RECT 1233.020 2318.370 1236.020 2318.380 ;
        RECT 1413.020 2318.370 1416.020 2318.380 ;
        RECT 1593.020 2318.370 1596.020 2318.380 ;
        RECT 1773.020 2318.370 1776.020 2318.380 ;
        RECT 1953.020 2318.370 1956.020 2318.380 ;
        RECT 2133.020 2318.370 2136.020 2318.380 ;
        RECT 2313.020 2318.370 2316.020 2318.380 ;
        RECT 2493.020 2318.370 2496.020 2318.380 ;
        RECT 2673.020 2318.370 2676.020 2318.380 ;
        RECT 2853.020 2318.370 2856.020 2318.380 ;
        RECT 2959.500 2318.370 2962.500 2318.380 ;
        RECT -42.880 2141.380 -39.880 2141.390 ;
        RECT 153.020 2141.380 156.020 2141.390 ;
        RECT 333.020 2141.380 336.020 2141.390 ;
        RECT 513.020 2141.380 516.020 2141.390 ;
        RECT 693.020 2141.380 696.020 2141.390 ;
        RECT 873.020 2141.380 876.020 2141.390 ;
        RECT 1053.020 2141.380 1056.020 2141.390 ;
        RECT 1233.020 2141.380 1236.020 2141.390 ;
        RECT 1413.020 2141.380 1416.020 2141.390 ;
        RECT 1593.020 2141.380 1596.020 2141.390 ;
        RECT 1773.020 2141.380 1776.020 2141.390 ;
        RECT 1953.020 2141.380 1956.020 2141.390 ;
        RECT 2133.020 2141.380 2136.020 2141.390 ;
        RECT 2313.020 2141.380 2316.020 2141.390 ;
        RECT 2493.020 2141.380 2496.020 2141.390 ;
        RECT 2673.020 2141.380 2676.020 2141.390 ;
        RECT 2853.020 2141.380 2856.020 2141.390 ;
        RECT 2959.500 2141.380 2962.500 2141.390 ;
        RECT -42.880 2138.380 2962.500 2141.380 ;
        RECT -42.880 2138.370 -39.880 2138.380 ;
        RECT 153.020 2138.370 156.020 2138.380 ;
        RECT 333.020 2138.370 336.020 2138.380 ;
        RECT 513.020 2138.370 516.020 2138.380 ;
        RECT 693.020 2138.370 696.020 2138.380 ;
        RECT 873.020 2138.370 876.020 2138.380 ;
        RECT 1053.020 2138.370 1056.020 2138.380 ;
        RECT 1233.020 2138.370 1236.020 2138.380 ;
        RECT 1413.020 2138.370 1416.020 2138.380 ;
        RECT 1593.020 2138.370 1596.020 2138.380 ;
        RECT 1773.020 2138.370 1776.020 2138.380 ;
        RECT 1953.020 2138.370 1956.020 2138.380 ;
        RECT 2133.020 2138.370 2136.020 2138.380 ;
        RECT 2313.020 2138.370 2316.020 2138.380 ;
        RECT 2493.020 2138.370 2496.020 2138.380 ;
        RECT 2673.020 2138.370 2676.020 2138.380 ;
        RECT 2853.020 2138.370 2856.020 2138.380 ;
        RECT 2959.500 2138.370 2962.500 2138.380 ;
        RECT -42.880 1961.380 -39.880 1961.390 ;
        RECT 153.020 1961.380 156.020 1961.390 ;
        RECT 333.020 1961.380 336.020 1961.390 ;
        RECT 513.020 1961.380 516.020 1961.390 ;
        RECT 693.020 1961.380 696.020 1961.390 ;
        RECT 873.020 1961.380 876.020 1961.390 ;
        RECT 1053.020 1961.380 1056.020 1961.390 ;
        RECT 1233.020 1961.380 1236.020 1961.390 ;
        RECT 1413.020 1961.380 1416.020 1961.390 ;
        RECT 1593.020 1961.380 1596.020 1961.390 ;
        RECT 1773.020 1961.380 1776.020 1961.390 ;
        RECT 1953.020 1961.380 1956.020 1961.390 ;
        RECT 2133.020 1961.380 2136.020 1961.390 ;
        RECT 2313.020 1961.380 2316.020 1961.390 ;
        RECT 2493.020 1961.380 2496.020 1961.390 ;
        RECT 2673.020 1961.380 2676.020 1961.390 ;
        RECT 2853.020 1961.380 2856.020 1961.390 ;
        RECT 2959.500 1961.380 2962.500 1961.390 ;
        RECT -42.880 1958.380 2962.500 1961.380 ;
        RECT -42.880 1958.370 -39.880 1958.380 ;
        RECT 153.020 1958.370 156.020 1958.380 ;
        RECT 333.020 1958.370 336.020 1958.380 ;
        RECT 513.020 1958.370 516.020 1958.380 ;
        RECT 693.020 1958.370 696.020 1958.380 ;
        RECT 873.020 1958.370 876.020 1958.380 ;
        RECT 1053.020 1958.370 1056.020 1958.380 ;
        RECT 1233.020 1958.370 1236.020 1958.380 ;
        RECT 1413.020 1958.370 1416.020 1958.380 ;
        RECT 1593.020 1958.370 1596.020 1958.380 ;
        RECT 1773.020 1958.370 1776.020 1958.380 ;
        RECT 1953.020 1958.370 1956.020 1958.380 ;
        RECT 2133.020 1958.370 2136.020 1958.380 ;
        RECT 2313.020 1958.370 2316.020 1958.380 ;
        RECT 2493.020 1958.370 2496.020 1958.380 ;
        RECT 2673.020 1958.370 2676.020 1958.380 ;
        RECT 2853.020 1958.370 2856.020 1958.380 ;
        RECT 2959.500 1958.370 2962.500 1958.380 ;
        RECT -42.880 1781.380 -39.880 1781.390 ;
        RECT 153.020 1781.380 156.020 1781.390 ;
        RECT 333.020 1781.380 336.020 1781.390 ;
        RECT 513.020 1781.380 516.020 1781.390 ;
        RECT 693.020 1781.380 696.020 1781.390 ;
        RECT 873.020 1781.380 876.020 1781.390 ;
        RECT 1053.020 1781.380 1056.020 1781.390 ;
        RECT 1233.020 1781.380 1236.020 1781.390 ;
        RECT 1413.020 1781.380 1416.020 1781.390 ;
        RECT 1593.020 1781.380 1596.020 1781.390 ;
        RECT 1773.020 1781.380 1776.020 1781.390 ;
        RECT 1953.020 1781.380 1956.020 1781.390 ;
        RECT 2133.020 1781.380 2136.020 1781.390 ;
        RECT 2313.020 1781.380 2316.020 1781.390 ;
        RECT 2493.020 1781.380 2496.020 1781.390 ;
        RECT 2673.020 1781.380 2676.020 1781.390 ;
        RECT 2853.020 1781.380 2856.020 1781.390 ;
        RECT 2959.500 1781.380 2962.500 1781.390 ;
        RECT -42.880 1778.380 2962.500 1781.380 ;
        RECT -42.880 1778.370 -39.880 1778.380 ;
        RECT 153.020 1778.370 156.020 1778.380 ;
        RECT 333.020 1778.370 336.020 1778.380 ;
        RECT 513.020 1778.370 516.020 1778.380 ;
        RECT 693.020 1778.370 696.020 1778.380 ;
        RECT 873.020 1778.370 876.020 1778.380 ;
        RECT 1053.020 1778.370 1056.020 1778.380 ;
        RECT 1233.020 1778.370 1236.020 1778.380 ;
        RECT 1413.020 1778.370 1416.020 1778.380 ;
        RECT 1593.020 1778.370 1596.020 1778.380 ;
        RECT 1773.020 1778.370 1776.020 1778.380 ;
        RECT 1953.020 1778.370 1956.020 1778.380 ;
        RECT 2133.020 1778.370 2136.020 1778.380 ;
        RECT 2313.020 1778.370 2316.020 1778.380 ;
        RECT 2493.020 1778.370 2496.020 1778.380 ;
        RECT 2673.020 1778.370 2676.020 1778.380 ;
        RECT 2853.020 1778.370 2856.020 1778.380 ;
        RECT 2959.500 1778.370 2962.500 1778.380 ;
        RECT -42.880 1601.380 -39.880 1601.390 ;
        RECT 153.020 1601.380 156.020 1601.390 ;
        RECT 333.020 1601.380 336.020 1601.390 ;
        RECT 513.020 1601.380 516.020 1601.390 ;
        RECT 693.020 1601.380 696.020 1601.390 ;
        RECT 873.020 1601.380 876.020 1601.390 ;
        RECT 1053.020 1601.380 1056.020 1601.390 ;
        RECT 1233.020 1601.380 1236.020 1601.390 ;
        RECT 1413.020 1601.380 1416.020 1601.390 ;
        RECT 1593.020 1601.380 1596.020 1601.390 ;
        RECT 1773.020 1601.380 1776.020 1601.390 ;
        RECT 1953.020 1601.380 1956.020 1601.390 ;
        RECT 2133.020 1601.380 2136.020 1601.390 ;
        RECT 2313.020 1601.380 2316.020 1601.390 ;
        RECT 2493.020 1601.380 2496.020 1601.390 ;
        RECT 2673.020 1601.380 2676.020 1601.390 ;
        RECT 2853.020 1601.380 2856.020 1601.390 ;
        RECT 2959.500 1601.380 2962.500 1601.390 ;
        RECT -42.880 1598.380 2962.500 1601.380 ;
        RECT -42.880 1598.370 -39.880 1598.380 ;
        RECT 153.020 1598.370 156.020 1598.380 ;
        RECT 333.020 1598.370 336.020 1598.380 ;
        RECT 513.020 1598.370 516.020 1598.380 ;
        RECT 693.020 1598.370 696.020 1598.380 ;
        RECT 873.020 1598.370 876.020 1598.380 ;
        RECT 1053.020 1598.370 1056.020 1598.380 ;
        RECT 1233.020 1598.370 1236.020 1598.380 ;
        RECT 1413.020 1598.370 1416.020 1598.380 ;
        RECT 1593.020 1598.370 1596.020 1598.380 ;
        RECT 1773.020 1598.370 1776.020 1598.380 ;
        RECT 1953.020 1598.370 1956.020 1598.380 ;
        RECT 2133.020 1598.370 2136.020 1598.380 ;
        RECT 2313.020 1598.370 2316.020 1598.380 ;
        RECT 2493.020 1598.370 2496.020 1598.380 ;
        RECT 2673.020 1598.370 2676.020 1598.380 ;
        RECT 2853.020 1598.370 2856.020 1598.380 ;
        RECT 2959.500 1598.370 2962.500 1598.380 ;
        RECT -42.880 1421.380 -39.880 1421.390 ;
        RECT 153.020 1421.380 156.020 1421.390 ;
        RECT 333.020 1421.380 336.020 1421.390 ;
        RECT 513.020 1421.380 516.020 1421.390 ;
        RECT 693.020 1421.380 696.020 1421.390 ;
        RECT 873.020 1421.380 876.020 1421.390 ;
        RECT 1053.020 1421.380 1056.020 1421.390 ;
        RECT 1233.020 1421.380 1236.020 1421.390 ;
        RECT 1413.020 1421.380 1416.020 1421.390 ;
        RECT 1593.020 1421.380 1596.020 1421.390 ;
        RECT 1773.020 1421.380 1776.020 1421.390 ;
        RECT 1953.020 1421.380 1956.020 1421.390 ;
        RECT 2133.020 1421.380 2136.020 1421.390 ;
        RECT 2313.020 1421.380 2316.020 1421.390 ;
        RECT 2493.020 1421.380 2496.020 1421.390 ;
        RECT 2673.020 1421.380 2676.020 1421.390 ;
        RECT 2853.020 1421.380 2856.020 1421.390 ;
        RECT 2959.500 1421.380 2962.500 1421.390 ;
        RECT -42.880 1418.380 2962.500 1421.380 ;
        RECT -42.880 1418.370 -39.880 1418.380 ;
        RECT 153.020 1418.370 156.020 1418.380 ;
        RECT 333.020 1418.370 336.020 1418.380 ;
        RECT 513.020 1418.370 516.020 1418.380 ;
        RECT 693.020 1418.370 696.020 1418.380 ;
        RECT 873.020 1418.370 876.020 1418.380 ;
        RECT 1053.020 1418.370 1056.020 1418.380 ;
        RECT 1233.020 1418.370 1236.020 1418.380 ;
        RECT 1413.020 1418.370 1416.020 1418.380 ;
        RECT 1593.020 1418.370 1596.020 1418.380 ;
        RECT 1773.020 1418.370 1776.020 1418.380 ;
        RECT 1953.020 1418.370 1956.020 1418.380 ;
        RECT 2133.020 1418.370 2136.020 1418.380 ;
        RECT 2313.020 1418.370 2316.020 1418.380 ;
        RECT 2493.020 1418.370 2496.020 1418.380 ;
        RECT 2673.020 1418.370 2676.020 1418.380 ;
        RECT 2853.020 1418.370 2856.020 1418.380 ;
        RECT 2959.500 1418.370 2962.500 1418.380 ;
        RECT -42.880 1241.380 -39.880 1241.390 ;
        RECT 153.020 1241.380 156.020 1241.390 ;
        RECT 333.020 1241.380 336.020 1241.390 ;
        RECT 513.020 1241.380 516.020 1241.390 ;
        RECT 693.020 1241.380 696.020 1241.390 ;
        RECT 873.020 1241.380 876.020 1241.390 ;
        RECT 1053.020 1241.380 1056.020 1241.390 ;
        RECT 1233.020 1241.380 1236.020 1241.390 ;
        RECT 1413.020 1241.380 1416.020 1241.390 ;
        RECT 1593.020 1241.380 1596.020 1241.390 ;
        RECT 1773.020 1241.380 1776.020 1241.390 ;
        RECT 1953.020 1241.380 1956.020 1241.390 ;
        RECT 2133.020 1241.380 2136.020 1241.390 ;
        RECT 2313.020 1241.380 2316.020 1241.390 ;
        RECT 2493.020 1241.380 2496.020 1241.390 ;
        RECT 2673.020 1241.380 2676.020 1241.390 ;
        RECT 2853.020 1241.380 2856.020 1241.390 ;
        RECT 2959.500 1241.380 2962.500 1241.390 ;
        RECT -42.880 1238.380 2962.500 1241.380 ;
        RECT -42.880 1238.370 -39.880 1238.380 ;
        RECT 153.020 1238.370 156.020 1238.380 ;
        RECT 333.020 1238.370 336.020 1238.380 ;
        RECT 513.020 1238.370 516.020 1238.380 ;
        RECT 693.020 1238.370 696.020 1238.380 ;
        RECT 873.020 1238.370 876.020 1238.380 ;
        RECT 1053.020 1238.370 1056.020 1238.380 ;
        RECT 1233.020 1238.370 1236.020 1238.380 ;
        RECT 1413.020 1238.370 1416.020 1238.380 ;
        RECT 1593.020 1238.370 1596.020 1238.380 ;
        RECT 1773.020 1238.370 1776.020 1238.380 ;
        RECT 1953.020 1238.370 1956.020 1238.380 ;
        RECT 2133.020 1238.370 2136.020 1238.380 ;
        RECT 2313.020 1238.370 2316.020 1238.380 ;
        RECT 2493.020 1238.370 2496.020 1238.380 ;
        RECT 2673.020 1238.370 2676.020 1238.380 ;
        RECT 2853.020 1238.370 2856.020 1238.380 ;
        RECT 2959.500 1238.370 2962.500 1238.380 ;
        RECT -42.880 1061.380 -39.880 1061.390 ;
        RECT 153.020 1061.380 156.020 1061.390 ;
        RECT 333.020 1061.380 336.020 1061.390 ;
        RECT 513.020 1061.380 516.020 1061.390 ;
        RECT 693.020 1061.380 696.020 1061.390 ;
        RECT 873.020 1061.380 876.020 1061.390 ;
        RECT 1053.020 1061.380 1056.020 1061.390 ;
        RECT 1233.020 1061.380 1236.020 1061.390 ;
        RECT 1413.020 1061.380 1416.020 1061.390 ;
        RECT 1593.020 1061.380 1596.020 1061.390 ;
        RECT 1773.020 1061.380 1776.020 1061.390 ;
        RECT 1953.020 1061.380 1956.020 1061.390 ;
        RECT 2133.020 1061.380 2136.020 1061.390 ;
        RECT 2313.020 1061.380 2316.020 1061.390 ;
        RECT 2493.020 1061.380 2496.020 1061.390 ;
        RECT 2673.020 1061.380 2676.020 1061.390 ;
        RECT 2853.020 1061.380 2856.020 1061.390 ;
        RECT 2959.500 1061.380 2962.500 1061.390 ;
        RECT -42.880 1058.380 2962.500 1061.380 ;
        RECT -42.880 1058.370 -39.880 1058.380 ;
        RECT 153.020 1058.370 156.020 1058.380 ;
        RECT 333.020 1058.370 336.020 1058.380 ;
        RECT 513.020 1058.370 516.020 1058.380 ;
        RECT 693.020 1058.370 696.020 1058.380 ;
        RECT 873.020 1058.370 876.020 1058.380 ;
        RECT 1053.020 1058.370 1056.020 1058.380 ;
        RECT 1233.020 1058.370 1236.020 1058.380 ;
        RECT 1413.020 1058.370 1416.020 1058.380 ;
        RECT 1593.020 1058.370 1596.020 1058.380 ;
        RECT 1773.020 1058.370 1776.020 1058.380 ;
        RECT 1953.020 1058.370 1956.020 1058.380 ;
        RECT 2133.020 1058.370 2136.020 1058.380 ;
        RECT 2313.020 1058.370 2316.020 1058.380 ;
        RECT 2493.020 1058.370 2496.020 1058.380 ;
        RECT 2673.020 1058.370 2676.020 1058.380 ;
        RECT 2853.020 1058.370 2856.020 1058.380 ;
        RECT 2959.500 1058.370 2962.500 1058.380 ;
        RECT -42.880 881.380 -39.880 881.390 ;
        RECT 153.020 881.380 156.020 881.390 ;
        RECT 333.020 881.380 336.020 881.390 ;
        RECT 513.020 881.380 516.020 881.390 ;
        RECT 693.020 881.380 696.020 881.390 ;
        RECT 873.020 881.380 876.020 881.390 ;
        RECT 1053.020 881.380 1056.020 881.390 ;
        RECT 1233.020 881.380 1236.020 881.390 ;
        RECT 1413.020 881.380 1416.020 881.390 ;
        RECT 1593.020 881.380 1596.020 881.390 ;
        RECT 1773.020 881.380 1776.020 881.390 ;
        RECT 1953.020 881.380 1956.020 881.390 ;
        RECT 2133.020 881.380 2136.020 881.390 ;
        RECT 2313.020 881.380 2316.020 881.390 ;
        RECT 2493.020 881.380 2496.020 881.390 ;
        RECT 2673.020 881.380 2676.020 881.390 ;
        RECT 2853.020 881.380 2856.020 881.390 ;
        RECT 2959.500 881.380 2962.500 881.390 ;
        RECT -42.880 878.380 2962.500 881.380 ;
        RECT -42.880 878.370 -39.880 878.380 ;
        RECT 153.020 878.370 156.020 878.380 ;
        RECT 333.020 878.370 336.020 878.380 ;
        RECT 513.020 878.370 516.020 878.380 ;
        RECT 693.020 878.370 696.020 878.380 ;
        RECT 873.020 878.370 876.020 878.380 ;
        RECT 1053.020 878.370 1056.020 878.380 ;
        RECT 1233.020 878.370 1236.020 878.380 ;
        RECT 1413.020 878.370 1416.020 878.380 ;
        RECT 1593.020 878.370 1596.020 878.380 ;
        RECT 1773.020 878.370 1776.020 878.380 ;
        RECT 1953.020 878.370 1956.020 878.380 ;
        RECT 2133.020 878.370 2136.020 878.380 ;
        RECT 2313.020 878.370 2316.020 878.380 ;
        RECT 2493.020 878.370 2496.020 878.380 ;
        RECT 2673.020 878.370 2676.020 878.380 ;
        RECT 2853.020 878.370 2856.020 878.380 ;
        RECT 2959.500 878.370 2962.500 878.380 ;
        RECT -42.880 701.380 -39.880 701.390 ;
        RECT 153.020 701.380 156.020 701.390 ;
        RECT 333.020 701.380 336.020 701.390 ;
        RECT 513.020 701.380 516.020 701.390 ;
        RECT 693.020 701.380 696.020 701.390 ;
        RECT 873.020 701.380 876.020 701.390 ;
        RECT 1053.020 701.380 1056.020 701.390 ;
        RECT 1233.020 701.380 1236.020 701.390 ;
        RECT 1413.020 701.380 1416.020 701.390 ;
        RECT 1593.020 701.380 1596.020 701.390 ;
        RECT 1773.020 701.380 1776.020 701.390 ;
        RECT 1953.020 701.380 1956.020 701.390 ;
        RECT 2133.020 701.380 2136.020 701.390 ;
        RECT 2313.020 701.380 2316.020 701.390 ;
        RECT 2493.020 701.380 2496.020 701.390 ;
        RECT 2673.020 701.380 2676.020 701.390 ;
        RECT 2853.020 701.380 2856.020 701.390 ;
        RECT 2959.500 701.380 2962.500 701.390 ;
        RECT -42.880 698.380 2962.500 701.380 ;
        RECT -42.880 698.370 -39.880 698.380 ;
        RECT 153.020 698.370 156.020 698.380 ;
        RECT 333.020 698.370 336.020 698.380 ;
        RECT 513.020 698.370 516.020 698.380 ;
        RECT 693.020 698.370 696.020 698.380 ;
        RECT 873.020 698.370 876.020 698.380 ;
        RECT 1053.020 698.370 1056.020 698.380 ;
        RECT 1233.020 698.370 1236.020 698.380 ;
        RECT 1413.020 698.370 1416.020 698.380 ;
        RECT 1593.020 698.370 1596.020 698.380 ;
        RECT 1773.020 698.370 1776.020 698.380 ;
        RECT 1953.020 698.370 1956.020 698.380 ;
        RECT 2133.020 698.370 2136.020 698.380 ;
        RECT 2313.020 698.370 2316.020 698.380 ;
        RECT 2493.020 698.370 2496.020 698.380 ;
        RECT 2673.020 698.370 2676.020 698.380 ;
        RECT 2853.020 698.370 2856.020 698.380 ;
        RECT 2959.500 698.370 2962.500 698.380 ;
        RECT -42.880 521.380 -39.880 521.390 ;
        RECT 153.020 521.380 156.020 521.390 ;
        RECT 333.020 521.380 336.020 521.390 ;
        RECT 513.020 521.380 516.020 521.390 ;
        RECT 693.020 521.380 696.020 521.390 ;
        RECT 873.020 521.380 876.020 521.390 ;
        RECT 1053.020 521.380 1056.020 521.390 ;
        RECT 1233.020 521.380 1236.020 521.390 ;
        RECT 1413.020 521.380 1416.020 521.390 ;
        RECT 1593.020 521.380 1596.020 521.390 ;
        RECT 1773.020 521.380 1776.020 521.390 ;
        RECT 1953.020 521.380 1956.020 521.390 ;
        RECT 2133.020 521.380 2136.020 521.390 ;
        RECT 2313.020 521.380 2316.020 521.390 ;
        RECT 2493.020 521.380 2496.020 521.390 ;
        RECT 2673.020 521.380 2676.020 521.390 ;
        RECT 2853.020 521.380 2856.020 521.390 ;
        RECT 2959.500 521.380 2962.500 521.390 ;
        RECT -42.880 518.380 2962.500 521.380 ;
        RECT -42.880 518.370 -39.880 518.380 ;
        RECT 153.020 518.370 156.020 518.380 ;
        RECT 333.020 518.370 336.020 518.380 ;
        RECT 513.020 518.370 516.020 518.380 ;
        RECT 693.020 518.370 696.020 518.380 ;
        RECT 873.020 518.370 876.020 518.380 ;
        RECT 1053.020 518.370 1056.020 518.380 ;
        RECT 1233.020 518.370 1236.020 518.380 ;
        RECT 1413.020 518.370 1416.020 518.380 ;
        RECT 1593.020 518.370 1596.020 518.380 ;
        RECT 1773.020 518.370 1776.020 518.380 ;
        RECT 1953.020 518.370 1956.020 518.380 ;
        RECT 2133.020 518.370 2136.020 518.380 ;
        RECT 2313.020 518.370 2316.020 518.380 ;
        RECT 2493.020 518.370 2496.020 518.380 ;
        RECT 2673.020 518.370 2676.020 518.380 ;
        RECT 2853.020 518.370 2856.020 518.380 ;
        RECT 2959.500 518.370 2962.500 518.380 ;
        RECT -42.880 341.380 -39.880 341.390 ;
        RECT 153.020 341.380 156.020 341.390 ;
        RECT 333.020 341.380 336.020 341.390 ;
        RECT 513.020 341.380 516.020 341.390 ;
        RECT 693.020 341.380 696.020 341.390 ;
        RECT 873.020 341.380 876.020 341.390 ;
        RECT 1053.020 341.380 1056.020 341.390 ;
        RECT 1233.020 341.380 1236.020 341.390 ;
        RECT 1413.020 341.380 1416.020 341.390 ;
        RECT 1593.020 341.380 1596.020 341.390 ;
        RECT 1773.020 341.380 1776.020 341.390 ;
        RECT 1953.020 341.380 1956.020 341.390 ;
        RECT 2133.020 341.380 2136.020 341.390 ;
        RECT 2313.020 341.380 2316.020 341.390 ;
        RECT 2493.020 341.380 2496.020 341.390 ;
        RECT 2673.020 341.380 2676.020 341.390 ;
        RECT 2853.020 341.380 2856.020 341.390 ;
        RECT 2959.500 341.380 2962.500 341.390 ;
        RECT -42.880 338.380 2962.500 341.380 ;
        RECT -42.880 338.370 -39.880 338.380 ;
        RECT 153.020 338.370 156.020 338.380 ;
        RECT 333.020 338.370 336.020 338.380 ;
        RECT 513.020 338.370 516.020 338.380 ;
        RECT 693.020 338.370 696.020 338.380 ;
        RECT 873.020 338.370 876.020 338.380 ;
        RECT 1053.020 338.370 1056.020 338.380 ;
        RECT 1233.020 338.370 1236.020 338.380 ;
        RECT 1413.020 338.370 1416.020 338.380 ;
        RECT 1593.020 338.370 1596.020 338.380 ;
        RECT 1773.020 338.370 1776.020 338.380 ;
        RECT 1953.020 338.370 1956.020 338.380 ;
        RECT 2133.020 338.370 2136.020 338.380 ;
        RECT 2313.020 338.370 2316.020 338.380 ;
        RECT 2493.020 338.370 2496.020 338.380 ;
        RECT 2673.020 338.370 2676.020 338.380 ;
        RECT 2853.020 338.370 2856.020 338.380 ;
        RECT 2959.500 338.370 2962.500 338.380 ;
        RECT -42.880 161.380 -39.880 161.390 ;
        RECT 153.020 161.380 156.020 161.390 ;
        RECT 333.020 161.380 336.020 161.390 ;
        RECT 513.020 161.380 516.020 161.390 ;
        RECT 693.020 161.380 696.020 161.390 ;
        RECT 873.020 161.380 876.020 161.390 ;
        RECT 1053.020 161.380 1056.020 161.390 ;
        RECT 1233.020 161.380 1236.020 161.390 ;
        RECT 1413.020 161.380 1416.020 161.390 ;
        RECT 1593.020 161.380 1596.020 161.390 ;
        RECT 1773.020 161.380 1776.020 161.390 ;
        RECT 1953.020 161.380 1956.020 161.390 ;
        RECT 2133.020 161.380 2136.020 161.390 ;
        RECT 2313.020 161.380 2316.020 161.390 ;
        RECT 2493.020 161.380 2496.020 161.390 ;
        RECT 2673.020 161.380 2676.020 161.390 ;
        RECT 2853.020 161.380 2856.020 161.390 ;
        RECT 2959.500 161.380 2962.500 161.390 ;
        RECT -42.880 158.380 2962.500 161.380 ;
        RECT -42.880 158.370 -39.880 158.380 ;
        RECT 153.020 158.370 156.020 158.380 ;
        RECT 333.020 158.370 336.020 158.380 ;
        RECT 513.020 158.370 516.020 158.380 ;
        RECT 693.020 158.370 696.020 158.380 ;
        RECT 873.020 158.370 876.020 158.380 ;
        RECT 1053.020 158.370 1056.020 158.380 ;
        RECT 1233.020 158.370 1236.020 158.380 ;
        RECT 1413.020 158.370 1416.020 158.380 ;
        RECT 1593.020 158.370 1596.020 158.380 ;
        RECT 1773.020 158.370 1776.020 158.380 ;
        RECT 1953.020 158.370 1956.020 158.380 ;
        RECT 2133.020 158.370 2136.020 158.380 ;
        RECT 2313.020 158.370 2316.020 158.380 ;
        RECT 2493.020 158.370 2496.020 158.380 ;
        RECT 2673.020 158.370 2676.020 158.380 ;
        RECT 2853.020 158.370 2856.020 158.380 ;
        RECT 2959.500 158.370 2962.500 158.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 153.020 -34.520 156.020 -34.510 ;
        RECT 333.020 -34.520 336.020 -34.510 ;
        RECT 513.020 -34.520 516.020 -34.510 ;
        RECT 693.020 -34.520 696.020 -34.510 ;
        RECT 873.020 -34.520 876.020 -34.510 ;
        RECT 1053.020 -34.520 1056.020 -34.510 ;
        RECT 1233.020 -34.520 1236.020 -34.510 ;
        RECT 1413.020 -34.520 1416.020 -34.510 ;
        RECT 1593.020 -34.520 1596.020 -34.510 ;
        RECT 1773.020 -34.520 1776.020 -34.510 ;
        RECT 1953.020 -34.520 1956.020 -34.510 ;
        RECT 2133.020 -34.520 2136.020 -34.510 ;
        RECT 2313.020 -34.520 2316.020 -34.510 ;
        RECT 2493.020 -34.520 2496.020 -34.510 ;
        RECT 2673.020 -34.520 2676.020 -34.510 ;
        RECT 2853.020 -34.520 2856.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 153.020 -37.530 156.020 -37.520 ;
        RECT 333.020 -37.530 336.020 -37.520 ;
        RECT 513.020 -37.530 516.020 -37.520 ;
        RECT 693.020 -37.530 696.020 -37.520 ;
        RECT 873.020 -37.530 876.020 -37.520 ;
        RECT 1053.020 -37.530 1056.020 -37.520 ;
        RECT 1233.020 -37.530 1236.020 -37.520 ;
        RECT 1413.020 -37.530 1416.020 -37.520 ;
        RECT 1593.020 -37.530 1596.020 -37.520 ;
        RECT 1773.020 -37.530 1776.020 -37.520 ;
        RECT 1953.020 -37.530 1956.020 -37.520 ;
        RECT 2133.020 -37.530 2136.020 -37.520 ;
        RECT 2313.020 -37.530 2316.020 -37.520 ;
        RECT 2493.020 -37.530 2496.020 -37.520 ;
        RECT 2673.020 -37.530 2676.020 -37.520 ;
        RECT 2853.020 -37.530 2856.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
END user_project_wrapper
END LIBRARY

