magic
tech sky130A
magscale 1 2
timestamp 1606424343
<< pwell >>
rect -3867 -1778 3867 1778
<< nmos >>
rect -3671 668 -3581 1568
rect -3523 668 -3433 1568
rect -3375 668 -3285 1568
rect -3227 668 -3137 1568
rect -3079 668 -2989 1568
rect -2931 668 -2841 1568
rect -2783 668 -2693 1568
rect -2635 668 -2545 1568
rect -2487 668 -2397 1568
rect -2339 668 -2249 1568
rect -2191 668 -2101 1568
rect -2043 668 -1953 1568
rect -1895 668 -1805 1568
rect -1747 668 -1657 1568
rect -1599 668 -1509 1568
rect -1451 668 -1361 1568
rect -1303 668 -1213 1568
rect -1155 668 -1065 1568
rect -1007 668 -917 1568
rect -859 668 -769 1568
rect -711 668 -621 1568
rect -563 668 -473 1568
rect -415 668 -325 1568
rect -267 668 -177 1568
rect -119 668 -29 1568
rect 29 668 119 1568
rect 177 668 267 1568
rect 325 668 415 1568
rect 473 668 563 1568
rect 621 668 711 1568
rect 769 668 859 1568
rect 917 668 1007 1568
rect 1065 668 1155 1568
rect 1213 668 1303 1568
rect 1361 668 1451 1568
rect 1509 668 1599 1568
rect 1657 668 1747 1568
rect 1805 668 1895 1568
rect 1953 668 2043 1568
rect 2101 668 2191 1568
rect 2249 668 2339 1568
rect 2397 668 2487 1568
rect 2545 668 2635 1568
rect 2693 668 2783 1568
rect 2841 668 2931 1568
rect 2989 668 3079 1568
rect 3137 668 3227 1568
rect 3285 668 3375 1568
rect 3433 668 3523 1568
rect 3581 668 3671 1568
rect -3671 -450 -3581 450
rect -3523 -450 -3433 450
rect -3375 -450 -3285 450
rect -3227 -450 -3137 450
rect -3079 -450 -2989 450
rect -2931 -450 -2841 450
rect -2783 -450 -2693 450
rect -2635 -450 -2545 450
rect -2487 -450 -2397 450
rect -2339 -450 -2249 450
rect -2191 -450 -2101 450
rect -2043 -450 -1953 450
rect -1895 -450 -1805 450
rect -1747 -450 -1657 450
rect -1599 -450 -1509 450
rect -1451 -450 -1361 450
rect -1303 -450 -1213 450
rect -1155 -450 -1065 450
rect -1007 -450 -917 450
rect -859 -450 -769 450
rect -711 -450 -621 450
rect -563 -450 -473 450
rect -415 -450 -325 450
rect -267 -450 -177 450
rect -119 -450 -29 450
rect 29 -450 119 450
rect 177 -450 267 450
rect 325 -450 415 450
rect 473 -450 563 450
rect 621 -450 711 450
rect 769 -450 859 450
rect 917 -450 1007 450
rect 1065 -450 1155 450
rect 1213 -450 1303 450
rect 1361 -450 1451 450
rect 1509 -450 1599 450
rect 1657 -450 1747 450
rect 1805 -450 1895 450
rect 1953 -450 2043 450
rect 2101 -450 2191 450
rect 2249 -450 2339 450
rect 2397 -450 2487 450
rect 2545 -450 2635 450
rect 2693 -450 2783 450
rect 2841 -450 2931 450
rect 2989 -450 3079 450
rect 3137 -450 3227 450
rect 3285 -450 3375 450
rect 3433 -450 3523 450
rect 3581 -450 3671 450
rect -3671 -1568 -3581 -668
rect -3523 -1568 -3433 -668
rect -3375 -1568 -3285 -668
rect -3227 -1568 -3137 -668
rect -3079 -1568 -2989 -668
rect -2931 -1568 -2841 -668
rect -2783 -1568 -2693 -668
rect -2635 -1568 -2545 -668
rect -2487 -1568 -2397 -668
rect -2339 -1568 -2249 -668
rect -2191 -1568 -2101 -668
rect -2043 -1568 -1953 -668
rect -1895 -1568 -1805 -668
rect -1747 -1568 -1657 -668
rect -1599 -1568 -1509 -668
rect -1451 -1568 -1361 -668
rect -1303 -1568 -1213 -668
rect -1155 -1568 -1065 -668
rect -1007 -1568 -917 -668
rect -859 -1568 -769 -668
rect -711 -1568 -621 -668
rect -563 -1568 -473 -668
rect -415 -1568 -325 -668
rect -267 -1568 -177 -668
rect -119 -1568 -29 -668
rect 29 -1568 119 -668
rect 177 -1568 267 -668
rect 325 -1568 415 -668
rect 473 -1568 563 -668
rect 621 -1568 711 -668
rect 769 -1568 859 -668
rect 917 -1568 1007 -668
rect 1065 -1568 1155 -668
rect 1213 -1568 1303 -668
rect 1361 -1568 1451 -668
rect 1509 -1568 1599 -668
rect 1657 -1568 1747 -668
rect 1805 -1568 1895 -668
rect 1953 -1568 2043 -668
rect 2101 -1568 2191 -668
rect 2249 -1568 2339 -668
rect 2397 -1568 2487 -668
rect 2545 -1568 2635 -668
rect 2693 -1568 2783 -668
rect 2841 -1568 2931 -668
rect 2989 -1568 3079 -668
rect 3137 -1568 3227 -668
rect 3285 -1568 3375 -668
rect 3433 -1568 3523 -668
rect 3581 -1568 3671 -668
<< ndiff >>
rect -3729 1556 -3671 1568
rect -3729 680 -3717 1556
rect -3683 680 -3671 1556
rect -3729 668 -3671 680
rect -3581 1556 -3523 1568
rect -3581 680 -3569 1556
rect -3535 680 -3523 1556
rect -3581 668 -3523 680
rect -3433 1556 -3375 1568
rect -3433 680 -3421 1556
rect -3387 680 -3375 1556
rect -3433 668 -3375 680
rect -3285 1556 -3227 1568
rect -3285 680 -3273 1556
rect -3239 680 -3227 1556
rect -3285 668 -3227 680
rect -3137 1556 -3079 1568
rect -3137 680 -3125 1556
rect -3091 680 -3079 1556
rect -3137 668 -3079 680
rect -2989 1556 -2931 1568
rect -2989 680 -2977 1556
rect -2943 680 -2931 1556
rect -2989 668 -2931 680
rect -2841 1556 -2783 1568
rect -2841 680 -2829 1556
rect -2795 680 -2783 1556
rect -2841 668 -2783 680
rect -2693 1556 -2635 1568
rect -2693 680 -2681 1556
rect -2647 680 -2635 1556
rect -2693 668 -2635 680
rect -2545 1556 -2487 1568
rect -2545 680 -2533 1556
rect -2499 680 -2487 1556
rect -2545 668 -2487 680
rect -2397 1556 -2339 1568
rect -2397 680 -2385 1556
rect -2351 680 -2339 1556
rect -2397 668 -2339 680
rect -2249 1556 -2191 1568
rect -2249 680 -2237 1556
rect -2203 680 -2191 1556
rect -2249 668 -2191 680
rect -2101 1556 -2043 1568
rect -2101 680 -2089 1556
rect -2055 680 -2043 1556
rect -2101 668 -2043 680
rect -1953 1556 -1895 1568
rect -1953 680 -1941 1556
rect -1907 680 -1895 1556
rect -1953 668 -1895 680
rect -1805 1556 -1747 1568
rect -1805 680 -1793 1556
rect -1759 680 -1747 1556
rect -1805 668 -1747 680
rect -1657 1556 -1599 1568
rect -1657 680 -1645 1556
rect -1611 680 -1599 1556
rect -1657 668 -1599 680
rect -1509 1556 -1451 1568
rect -1509 680 -1497 1556
rect -1463 680 -1451 1556
rect -1509 668 -1451 680
rect -1361 1556 -1303 1568
rect -1361 680 -1349 1556
rect -1315 680 -1303 1556
rect -1361 668 -1303 680
rect -1213 1556 -1155 1568
rect -1213 680 -1201 1556
rect -1167 680 -1155 1556
rect -1213 668 -1155 680
rect -1065 1556 -1007 1568
rect -1065 680 -1053 1556
rect -1019 680 -1007 1556
rect -1065 668 -1007 680
rect -917 1556 -859 1568
rect -917 680 -905 1556
rect -871 680 -859 1556
rect -917 668 -859 680
rect -769 1556 -711 1568
rect -769 680 -757 1556
rect -723 680 -711 1556
rect -769 668 -711 680
rect -621 1556 -563 1568
rect -621 680 -609 1556
rect -575 680 -563 1556
rect -621 668 -563 680
rect -473 1556 -415 1568
rect -473 680 -461 1556
rect -427 680 -415 1556
rect -473 668 -415 680
rect -325 1556 -267 1568
rect -325 680 -313 1556
rect -279 680 -267 1556
rect -325 668 -267 680
rect -177 1556 -119 1568
rect -177 680 -165 1556
rect -131 680 -119 1556
rect -177 668 -119 680
rect -29 1556 29 1568
rect -29 680 -17 1556
rect 17 680 29 1556
rect -29 668 29 680
rect 119 1556 177 1568
rect 119 680 131 1556
rect 165 680 177 1556
rect 119 668 177 680
rect 267 1556 325 1568
rect 267 680 279 1556
rect 313 680 325 1556
rect 267 668 325 680
rect 415 1556 473 1568
rect 415 680 427 1556
rect 461 680 473 1556
rect 415 668 473 680
rect 563 1556 621 1568
rect 563 680 575 1556
rect 609 680 621 1556
rect 563 668 621 680
rect 711 1556 769 1568
rect 711 680 723 1556
rect 757 680 769 1556
rect 711 668 769 680
rect 859 1556 917 1568
rect 859 680 871 1556
rect 905 680 917 1556
rect 859 668 917 680
rect 1007 1556 1065 1568
rect 1007 680 1019 1556
rect 1053 680 1065 1556
rect 1007 668 1065 680
rect 1155 1556 1213 1568
rect 1155 680 1167 1556
rect 1201 680 1213 1556
rect 1155 668 1213 680
rect 1303 1556 1361 1568
rect 1303 680 1315 1556
rect 1349 680 1361 1556
rect 1303 668 1361 680
rect 1451 1556 1509 1568
rect 1451 680 1463 1556
rect 1497 680 1509 1556
rect 1451 668 1509 680
rect 1599 1556 1657 1568
rect 1599 680 1611 1556
rect 1645 680 1657 1556
rect 1599 668 1657 680
rect 1747 1556 1805 1568
rect 1747 680 1759 1556
rect 1793 680 1805 1556
rect 1747 668 1805 680
rect 1895 1556 1953 1568
rect 1895 680 1907 1556
rect 1941 680 1953 1556
rect 1895 668 1953 680
rect 2043 1556 2101 1568
rect 2043 680 2055 1556
rect 2089 680 2101 1556
rect 2043 668 2101 680
rect 2191 1556 2249 1568
rect 2191 680 2203 1556
rect 2237 680 2249 1556
rect 2191 668 2249 680
rect 2339 1556 2397 1568
rect 2339 680 2351 1556
rect 2385 680 2397 1556
rect 2339 668 2397 680
rect 2487 1556 2545 1568
rect 2487 680 2499 1556
rect 2533 680 2545 1556
rect 2487 668 2545 680
rect 2635 1556 2693 1568
rect 2635 680 2647 1556
rect 2681 680 2693 1556
rect 2635 668 2693 680
rect 2783 1556 2841 1568
rect 2783 680 2795 1556
rect 2829 680 2841 1556
rect 2783 668 2841 680
rect 2931 1556 2989 1568
rect 2931 680 2943 1556
rect 2977 680 2989 1556
rect 2931 668 2989 680
rect 3079 1556 3137 1568
rect 3079 680 3091 1556
rect 3125 680 3137 1556
rect 3079 668 3137 680
rect 3227 1556 3285 1568
rect 3227 680 3239 1556
rect 3273 680 3285 1556
rect 3227 668 3285 680
rect 3375 1556 3433 1568
rect 3375 680 3387 1556
rect 3421 680 3433 1556
rect 3375 668 3433 680
rect 3523 1556 3581 1568
rect 3523 680 3535 1556
rect 3569 680 3581 1556
rect 3523 668 3581 680
rect 3671 1556 3729 1568
rect 3671 680 3683 1556
rect 3717 680 3729 1556
rect 3671 668 3729 680
rect -3729 438 -3671 450
rect -3729 -438 -3717 438
rect -3683 -438 -3671 438
rect -3729 -450 -3671 -438
rect -3581 438 -3523 450
rect -3581 -438 -3569 438
rect -3535 -438 -3523 438
rect -3581 -450 -3523 -438
rect -3433 438 -3375 450
rect -3433 -438 -3421 438
rect -3387 -438 -3375 438
rect -3433 -450 -3375 -438
rect -3285 438 -3227 450
rect -3285 -438 -3273 438
rect -3239 -438 -3227 438
rect -3285 -450 -3227 -438
rect -3137 438 -3079 450
rect -3137 -438 -3125 438
rect -3091 -438 -3079 438
rect -3137 -450 -3079 -438
rect -2989 438 -2931 450
rect -2989 -438 -2977 438
rect -2943 -438 -2931 438
rect -2989 -450 -2931 -438
rect -2841 438 -2783 450
rect -2841 -438 -2829 438
rect -2795 -438 -2783 438
rect -2841 -450 -2783 -438
rect -2693 438 -2635 450
rect -2693 -438 -2681 438
rect -2647 -438 -2635 438
rect -2693 -450 -2635 -438
rect -2545 438 -2487 450
rect -2545 -438 -2533 438
rect -2499 -438 -2487 438
rect -2545 -450 -2487 -438
rect -2397 438 -2339 450
rect -2397 -438 -2385 438
rect -2351 -438 -2339 438
rect -2397 -450 -2339 -438
rect -2249 438 -2191 450
rect -2249 -438 -2237 438
rect -2203 -438 -2191 438
rect -2249 -450 -2191 -438
rect -2101 438 -2043 450
rect -2101 -438 -2089 438
rect -2055 -438 -2043 438
rect -2101 -450 -2043 -438
rect -1953 438 -1895 450
rect -1953 -438 -1941 438
rect -1907 -438 -1895 438
rect -1953 -450 -1895 -438
rect -1805 438 -1747 450
rect -1805 -438 -1793 438
rect -1759 -438 -1747 438
rect -1805 -450 -1747 -438
rect -1657 438 -1599 450
rect -1657 -438 -1645 438
rect -1611 -438 -1599 438
rect -1657 -450 -1599 -438
rect -1509 438 -1451 450
rect -1509 -438 -1497 438
rect -1463 -438 -1451 438
rect -1509 -450 -1451 -438
rect -1361 438 -1303 450
rect -1361 -438 -1349 438
rect -1315 -438 -1303 438
rect -1361 -450 -1303 -438
rect -1213 438 -1155 450
rect -1213 -438 -1201 438
rect -1167 -438 -1155 438
rect -1213 -450 -1155 -438
rect -1065 438 -1007 450
rect -1065 -438 -1053 438
rect -1019 -438 -1007 438
rect -1065 -450 -1007 -438
rect -917 438 -859 450
rect -917 -438 -905 438
rect -871 -438 -859 438
rect -917 -450 -859 -438
rect -769 438 -711 450
rect -769 -438 -757 438
rect -723 -438 -711 438
rect -769 -450 -711 -438
rect -621 438 -563 450
rect -621 -438 -609 438
rect -575 -438 -563 438
rect -621 -450 -563 -438
rect -473 438 -415 450
rect -473 -438 -461 438
rect -427 -438 -415 438
rect -473 -450 -415 -438
rect -325 438 -267 450
rect -325 -438 -313 438
rect -279 -438 -267 438
rect -325 -450 -267 -438
rect -177 438 -119 450
rect -177 -438 -165 438
rect -131 -438 -119 438
rect -177 -450 -119 -438
rect -29 438 29 450
rect -29 -438 -17 438
rect 17 -438 29 438
rect -29 -450 29 -438
rect 119 438 177 450
rect 119 -438 131 438
rect 165 -438 177 438
rect 119 -450 177 -438
rect 267 438 325 450
rect 267 -438 279 438
rect 313 -438 325 438
rect 267 -450 325 -438
rect 415 438 473 450
rect 415 -438 427 438
rect 461 -438 473 438
rect 415 -450 473 -438
rect 563 438 621 450
rect 563 -438 575 438
rect 609 -438 621 438
rect 563 -450 621 -438
rect 711 438 769 450
rect 711 -438 723 438
rect 757 -438 769 438
rect 711 -450 769 -438
rect 859 438 917 450
rect 859 -438 871 438
rect 905 -438 917 438
rect 859 -450 917 -438
rect 1007 438 1065 450
rect 1007 -438 1019 438
rect 1053 -438 1065 438
rect 1007 -450 1065 -438
rect 1155 438 1213 450
rect 1155 -438 1167 438
rect 1201 -438 1213 438
rect 1155 -450 1213 -438
rect 1303 438 1361 450
rect 1303 -438 1315 438
rect 1349 -438 1361 438
rect 1303 -450 1361 -438
rect 1451 438 1509 450
rect 1451 -438 1463 438
rect 1497 -438 1509 438
rect 1451 -450 1509 -438
rect 1599 438 1657 450
rect 1599 -438 1611 438
rect 1645 -438 1657 438
rect 1599 -450 1657 -438
rect 1747 438 1805 450
rect 1747 -438 1759 438
rect 1793 -438 1805 438
rect 1747 -450 1805 -438
rect 1895 438 1953 450
rect 1895 -438 1907 438
rect 1941 -438 1953 438
rect 1895 -450 1953 -438
rect 2043 438 2101 450
rect 2043 -438 2055 438
rect 2089 -438 2101 438
rect 2043 -450 2101 -438
rect 2191 438 2249 450
rect 2191 -438 2203 438
rect 2237 -438 2249 438
rect 2191 -450 2249 -438
rect 2339 438 2397 450
rect 2339 -438 2351 438
rect 2385 -438 2397 438
rect 2339 -450 2397 -438
rect 2487 438 2545 450
rect 2487 -438 2499 438
rect 2533 -438 2545 438
rect 2487 -450 2545 -438
rect 2635 438 2693 450
rect 2635 -438 2647 438
rect 2681 -438 2693 438
rect 2635 -450 2693 -438
rect 2783 438 2841 450
rect 2783 -438 2795 438
rect 2829 -438 2841 438
rect 2783 -450 2841 -438
rect 2931 438 2989 450
rect 2931 -438 2943 438
rect 2977 -438 2989 438
rect 2931 -450 2989 -438
rect 3079 438 3137 450
rect 3079 -438 3091 438
rect 3125 -438 3137 438
rect 3079 -450 3137 -438
rect 3227 438 3285 450
rect 3227 -438 3239 438
rect 3273 -438 3285 438
rect 3227 -450 3285 -438
rect 3375 438 3433 450
rect 3375 -438 3387 438
rect 3421 -438 3433 438
rect 3375 -450 3433 -438
rect 3523 438 3581 450
rect 3523 -438 3535 438
rect 3569 -438 3581 438
rect 3523 -450 3581 -438
rect 3671 438 3729 450
rect 3671 -438 3683 438
rect 3717 -438 3729 438
rect 3671 -450 3729 -438
rect -3729 -680 -3671 -668
rect -3729 -1556 -3717 -680
rect -3683 -1556 -3671 -680
rect -3729 -1568 -3671 -1556
rect -3581 -680 -3523 -668
rect -3581 -1556 -3569 -680
rect -3535 -1556 -3523 -680
rect -3581 -1568 -3523 -1556
rect -3433 -680 -3375 -668
rect -3433 -1556 -3421 -680
rect -3387 -1556 -3375 -680
rect -3433 -1568 -3375 -1556
rect -3285 -680 -3227 -668
rect -3285 -1556 -3273 -680
rect -3239 -1556 -3227 -680
rect -3285 -1568 -3227 -1556
rect -3137 -680 -3079 -668
rect -3137 -1556 -3125 -680
rect -3091 -1556 -3079 -680
rect -3137 -1568 -3079 -1556
rect -2989 -680 -2931 -668
rect -2989 -1556 -2977 -680
rect -2943 -1556 -2931 -680
rect -2989 -1568 -2931 -1556
rect -2841 -680 -2783 -668
rect -2841 -1556 -2829 -680
rect -2795 -1556 -2783 -680
rect -2841 -1568 -2783 -1556
rect -2693 -680 -2635 -668
rect -2693 -1556 -2681 -680
rect -2647 -1556 -2635 -680
rect -2693 -1568 -2635 -1556
rect -2545 -680 -2487 -668
rect -2545 -1556 -2533 -680
rect -2499 -1556 -2487 -680
rect -2545 -1568 -2487 -1556
rect -2397 -680 -2339 -668
rect -2397 -1556 -2385 -680
rect -2351 -1556 -2339 -680
rect -2397 -1568 -2339 -1556
rect -2249 -680 -2191 -668
rect -2249 -1556 -2237 -680
rect -2203 -1556 -2191 -680
rect -2249 -1568 -2191 -1556
rect -2101 -680 -2043 -668
rect -2101 -1556 -2089 -680
rect -2055 -1556 -2043 -680
rect -2101 -1568 -2043 -1556
rect -1953 -680 -1895 -668
rect -1953 -1556 -1941 -680
rect -1907 -1556 -1895 -680
rect -1953 -1568 -1895 -1556
rect -1805 -680 -1747 -668
rect -1805 -1556 -1793 -680
rect -1759 -1556 -1747 -680
rect -1805 -1568 -1747 -1556
rect -1657 -680 -1599 -668
rect -1657 -1556 -1645 -680
rect -1611 -1556 -1599 -680
rect -1657 -1568 -1599 -1556
rect -1509 -680 -1451 -668
rect -1509 -1556 -1497 -680
rect -1463 -1556 -1451 -680
rect -1509 -1568 -1451 -1556
rect -1361 -680 -1303 -668
rect -1361 -1556 -1349 -680
rect -1315 -1556 -1303 -680
rect -1361 -1568 -1303 -1556
rect -1213 -680 -1155 -668
rect -1213 -1556 -1201 -680
rect -1167 -1556 -1155 -680
rect -1213 -1568 -1155 -1556
rect -1065 -680 -1007 -668
rect -1065 -1556 -1053 -680
rect -1019 -1556 -1007 -680
rect -1065 -1568 -1007 -1556
rect -917 -680 -859 -668
rect -917 -1556 -905 -680
rect -871 -1556 -859 -680
rect -917 -1568 -859 -1556
rect -769 -680 -711 -668
rect -769 -1556 -757 -680
rect -723 -1556 -711 -680
rect -769 -1568 -711 -1556
rect -621 -680 -563 -668
rect -621 -1556 -609 -680
rect -575 -1556 -563 -680
rect -621 -1568 -563 -1556
rect -473 -680 -415 -668
rect -473 -1556 -461 -680
rect -427 -1556 -415 -680
rect -473 -1568 -415 -1556
rect -325 -680 -267 -668
rect -325 -1556 -313 -680
rect -279 -1556 -267 -680
rect -325 -1568 -267 -1556
rect -177 -680 -119 -668
rect -177 -1556 -165 -680
rect -131 -1556 -119 -680
rect -177 -1568 -119 -1556
rect -29 -680 29 -668
rect -29 -1556 -17 -680
rect 17 -1556 29 -680
rect -29 -1568 29 -1556
rect 119 -680 177 -668
rect 119 -1556 131 -680
rect 165 -1556 177 -680
rect 119 -1568 177 -1556
rect 267 -680 325 -668
rect 267 -1556 279 -680
rect 313 -1556 325 -680
rect 267 -1568 325 -1556
rect 415 -680 473 -668
rect 415 -1556 427 -680
rect 461 -1556 473 -680
rect 415 -1568 473 -1556
rect 563 -680 621 -668
rect 563 -1556 575 -680
rect 609 -1556 621 -680
rect 563 -1568 621 -1556
rect 711 -680 769 -668
rect 711 -1556 723 -680
rect 757 -1556 769 -680
rect 711 -1568 769 -1556
rect 859 -680 917 -668
rect 859 -1556 871 -680
rect 905 -1556 917 -680
rect 859 -1568 917 -1556
rect 1007 -680 1065 -668
rect 1007 -1556 1019 -680
rect 1053 -1556 1065 -680
rect 1007 -1568 1065 -1556
rect 1155 -680 1213 -668
rect 1155 -1556 1167 -680
rect 1201 -1556 1213 -680
rect 1155 -1568 1213 -1556
rect 1303 -680 1361 -668
rect 1303 -1556 1315 -680
rect 1349 -1556 1361 -680
rect 1303 -1568 1361 -1556
rect 1451 -680 1509 -668
rect 1451 -1556 1463 -680
rect 1497 -1556 1509 -680
rect 1451 -1568 1509 -1556
rect 1599 -680 1657 -668
rect 1599 -1556 1611 -680
rect 1645 -1556 1657 -680
rect 1599 -1568 1657 -1556
rect 1747 -680 1805 -668
rect 1747 -1556 1759 -680
rect 1793 -1556 1805 -680
rect 1747 -1568 1805 -1556
rect 1895 -680 1953 -668
rect 1895 -1556 1907 -680
rect 1941 -1556 1953 -680
rect 1895 -1568 1953 -1556
rect 2043 -680 2101 -668
rect 2043 -1556 2055 -680
rect 2089 -1556 2101 -680
rect 2043 -1568 2101 -1556
rect 2191 -680 2249 -668
rect 2191 -1556 2203 -680
rect 2237 -1556 2249 -680
rect 2191 -1568 2249 -1556
rect 2339 -680 2397 -668
rect 2339 -1556 2351 -680
rect 2385 -1556 2397 -680
rect 2339 -1568 2397 -1556
rect 2487 -680 2545 -668
rect 2487 -1556 2499 -680
rect 2533 -1556 2545 -680
rect 2487 -1568 2545 -1556
rect 2635 -680 2693 -668
rect 2635 -1556 2647 -680
rect 2681 -1556 2693 -680
rect 2635 -1568 2693 -1556
rect 2783 -680 2841 -668
rect 2783 -1556 2795 -680
rect 2829 -1556 2841 -680
rect 2783 -1568 2841 -1556
rect 2931 -680 2989 -668
rect 2931 -1556 2943 -680
rect 2977 -1556 2989 -680
rect 2931 -1568 2989 -1556
rect 3079 -680 3137 -668
rect 3079 -1556 3091 -680
rect 3125 -1556 3137 -680
rect 3079 -1568 3137 -1556
rect 3227 -680 3285 -668
rect 3227 -1556 3239 -680
rect 3273 -1556 3285 -680
rect 3227 -1568 3285 -1556
rect 3375 -680 3433 -668
rect 3375 -1556 3387 -680
rect 3421 -1556 3433 -680
rect 3375 -1568 3433 -1556
rect 3523 -680 3581 -668
rect 3523 -1556 3535 -680
rect 3569 -1556 3581 -680
rect 3523 -1568 3581 -1556
rect 3671 -680 3729 -668
rect 3671 -1556 3683 -680
rect 3717 -1556 3729 -680
rect 3671 -1568 3729 -1556
<< ndiffc >>
rect -3717 680 -3683 1556
rect -3569 680 -3535 1556
rect -3421 680 -3387 1556
rect -3273 680 -3239 1556
rect -3125 680 -3091 1556
rect -2977 680 -2943 1556
rect -2829 680 -2795 1556
rect -2681 680 -2647 1556
rect -2533 680 -2499 1556
rect -2385 680 -2351 1556
rect -2237 680 -2203 1556
rect -2089 680 -2055 1556
rect -1941 680 -1907 1556
rect -1793 680 -1759 1556
rect -1645 680 -1611 1556
rect -1497 680 -1463 1556
rect -1349 680 -1315 1556
rect -1201 680 -1167 1556
rect -1053 680 -1019 1556
rect -905 680 -871 1556
rect -757 680 -723 1556
rect -609 680 -575 1556
rect -461 680 -427 1556
rect -313 680 -279 1556
rect -165 680 -131 1556
rect -17 680 17 1556
rect 131 680 165 1556
rect 279 680 313 1556
rect 427 680 461 1556
rect 575 680 609 1556
rect 723 680 757 1556
rect 871 680 905 1556
rect 1019 680 1053 1556
rect 1167 680 1201 1556
rect 1315 680 1349 1556
rect 1463 680 1497 1556
rect 1611 680 1645 1556
rect 1759 680 1793 1556
rect 1907 680 1941 1556
rect 2055 680 2089 1556
rect 2203 680 2237 1556
rect 2351 680 2385 1556
rect 2499 680 2533 1556
rect 2647 680 2681 1556
rect 2795 680 2829 1556
rect 2943 680 2977 1556
rect 3091 680 3125 1556
rect 3239 680 3273 1556
rect 3387 680 3421 1556
rect 3535 680 3569 1556
rect 3683 680 3717 1556
rect -3717 -438 -3683 438
rect -3569 -438 -3535 438
rect -3421 -438 -3387 438
rect -3273 -438 -3239 438
rect -3125 -438 -3091 438
rect -2977 -438 -2943 438
rect -2829 -438 -2795 438
rect -2681 -438 -2647 438
rect -2533 -438 -2499 438
rect -2385 -438 -2351 438
rect -2237 -438 -2203 438
rect -2089 -438 -2055 438
rect -1941 -438 -1907 438
rect -1793 -438 -1759 438
rect -1645 -438 -1611 438
rect -1497 -438 -1463 438
rect -1349 -438 -1315 438
rect -1201 -438 -1167 438
rect -1053 -438 -1019 438
rect -905 -438 -871 438
rect -757 -438 -723 438
rect -609 -438 -575 438
rect -461 -438 -427 438
rect -313 -438 -279 438
rect -165 -438 -131 438
rect -17 -438 17 438
rect 131 -438 165 438
rect 279 -438 313 438
rect 427 -438 461 438
rect 575 -438 609 438
rect 723 -438 757 438
rect 871 -438 905 438
rect 1019 -438 1053 438
rect 1167 -438 1201 438
rect 1315 -438 1349 438
rect 1463 -438 1497 438
rect 1611 -438 1645 438
rect 1759 -438 1793 438
rect 1907 -438 1941 438
rect 2055 -438 2089 438
rect 2203 -438 2237 438
rect 2351 -438 2385 438
rect 2499 -438 2533 438
rect 2647 -438 2681 438
rect 2795 -438 2829 438
rect 2943 -438 2977 438
rect 3091 -438 3125 438
rect 3239 -438 3273 438
rect 3387 -438 3421 438
rect 3535 -438 3569 438
rect 3683 -438 3717 438
rect -3717 -1556 -3683 -680
rect -3569 -1556 -3535 -680
rect -3421 -1556 -3387 -680
rect -3273 -1556 -3239 -680
rect -3125 -1556 -3091 -680
rect -2977 -1556 -2943 -680
rect -2829 -1556 -2795 -680
rect -2681 -1556 -2647 -680
rect -2533 -1556 -2499 -680
rect -2385 -1556 -2351 -680
rect -2237 -1556 -2203 -680
rect -2089 -1556 -2055 -680
rect -1941 -1556 -1907 -680
rect -1793 -1556 -1759 -680
rect -1645 -1556 -1611 -680
rect -1497 -1556 -1463 -680
rect -1349 -1556 -1315 -680
rect -1201 -1556 -1167 -680
rect -1053 -1556 -1019 -680
rect -905 -1556 -871 -680
rect -757 -1556 -723 -680
rect -609 -1556 -575 -680
rect -461 -1556 -427 -680
rect -313 -1556 -279 -680
rect -165 -1556 -131 -680
rect -17 -1556 17 -680
rect 131 -1556 165 -680
rect 279 -1556 313 -680
rect 427 -1556 461 -680
rect 575 -1556 609 -680
rect 723 -1556 757 -680
rect 871 -1556 905 -680
rect 1019 -1556 1053 -680
rect 1167 -1556 1201 -680
rect 1315 -1556 1349 -680
rect 1463 -1556 1497 -680
rect 1611 -1556 1645 -680
rect 1759 -1556 1793 -680
rect 1907 -1556 1941 -680
rect 2055 -1556 2089 -680
rect 2203 -1556 2237 -680
rect 2351 -1556 2385 -680
rect 2499 -1556 2533 -680
rect 2647 -1556 2681 -680
rect 2795 -1556 2829 -680
rect 2943 -1556 2977 -680
rect 3091 -1556 3125 -680
rect 3239 -1556 3273 -680
rect 3387 -1556 3421 -680
rect 3535 -1556 3569 -680
rect 3683 -1556 3717 -680
<< psubdiff >>
rect -3831 1708 -3735 1742
rect 3735 1708 3831 1742
rect -3831 1646 -3797 1708
rect 3797 1646 3831 1708
rect -3831 -1708 -3797 -1646
rect 3797 -1708 3831 -1646
rect -3831 -1742 -3735 -1708
rect 3735 -1742 3831 -1708
<< psubdiffcont >>
rect -3735 1708 3735 1742
rect -3831 -1646 -3797 1646
rect 3797 -1646 3831 1646
rect -3735 -1742 3735 -1708
<< poly >>
rect -3671 1640 -3581 1656
rect -3671 1606 -3655 1640
rect -3597 1606 -3581 1640
rect -3671 1568 -3581 1606
rect -3523 1640 -3433 1656
rect -3523 1606 -3507 1640
rect -3449 1606 -3433 1640
rect -3523 1568 -3433 1606
rect -3375 1640 -3285 1656
rect -3375 1606 -3359 1640
rect -3301 1606 -3285 1640
rect -3375 1568 -3285 1606
rect -3227 1640 -3137 1656
rect -3227 1606 -3211 1640
rect -3153 1606 -3137 1640
rect -3227 1568 -3137 1606
rect -3079 1640 -2989 1656
rect -3079 1606 -3063 1640
rect -3005 1606 -2989 1640
rect -3079 1568 -2989 1606
rect -2931 1640 -2841 1656
rect -2931 1606 -2915 1640
rect -2857 1606 -2841 1640
rect -2931 1568 -2841 1606
rect -2783 1640 -2693 1656
rect -2783 1606 -2767 1640
rect -2709 1606 -2693 1640
rect -2783 1568 -2693 1606
rect -2635 1640 -2545 1656
rect -2635 1606 -2619 1640
rect -2561 1606 -2545 1640
rect -2635 1568 -2545 1606
rect -2487 1640 -2397 1656
rect -2487 1606 -2471 1640
rect -2413 1606 -2397 1640
rect -2487 1568 -2397 1606
rect -2339 1640 -2249 1656
rect -2339 1606 -2323 1640
rect -2265 1606 -2249 1640
rect -2339 1568 -2249 1606
rect -2191 1640 -2101 1656
rect -2191 1606 -2175 1640
rect -2117 1606 -2101 1640
rect -2191 1568 -2101 1606
rect -2043 1640 -1953 1656
rect -2043 1606 -2027 1640
rect -1969 1606 -1953 1640
rect -2043 1568 -1953 1606
rect -1895 1640 -1805 1656
rect -1895 1606 -1879 1640
rect -1821 1606 -1805 1640
rect -1895 1568 -1805 1606
rect -1747 1640 -1657 1656
rect -1747 1606 -1731 1640
rect -1673 1606 -1657 1640
rect -1747 1568 -1657 1606
rect -1599 1640 -1509 1656
rect -1599 1606 -1583 1640
rect -1525 1606 -1509 1640
rect -1599 1568 -1509 1606
rect -1451 1640 -1361 1656
rect -1451 1606 -1435 1640
rect -1377 1606 -1361 1640
rect -1451 1568 -1361 1606
rect -1303 1640 -1213 1656
rect -1303 1606 -1287 1640
rect -1229 1606 -1213 1640
rect -1303 1568 -1213 1606
rect -1155 1640 -1065 1656
rect -1155 1606 -1139 1640
rect -1081 1606 -1065 1640
rect -1155 1568 -1065 1606
rect -1007 1640 -917 1656
rect -1007 1606 -991 1640
rect -933 1606 -917 1640
rect -1007 1568 -917 1606
rect -859 1640 -769 1656
rect -859 1606 -843 1640
rect -785 1606 -769 1640
rect -859 1568 -769 1606
rect -711 1640 -621 1656
rect -711 1606 -695 1640
rect -637 1606 -621 1640
rect -711 1568 -621 1606
rect -563 1640 -473 1656
rect -563 1606 -547 1640
rect -489 1606 -473 1640
rect -563 1568 -473 1606
rect -415 1640 -325 1656
rect -415 1606 -399 1640
rect -341 1606 -325 1640
rect -415 1568 -325 1606
rect -267 1640 -177 1656
rect -267 1606 -251 1640
rect -193 1606 -177 1640
rect -267 1568 -177 1606
rect -119 1640 -29 1656
rect -119 1606 -103 1640
rect -45 1606 -29 1640
rect -119 1568 -29 1606
rect 29 1640 119 1656
rect 29 1606 45 1640
rect 103 1606 119 1640
rect 29 1568 119 1606
rect 177 1640 267 1656
rect 177 1606 193 1640
rect 251 1606 267 1640
rect 177 1568 267 1606
rect 325 1640 415 1656
rect 325 1606 341 1640
rect 399 1606 415 1640
rect 325 1568 415 1606
rect 473 1640 563 1656
rect 473 1606 489 1640
rect 547 1606 563 1640
rect 473 1568 563 1606
rect 621 1640 711 1656
rect 621 1606 637 1640
rect 695 1606 711 1640
rect 621 1568 711 1606
rect 769 1640 859 1656
rect 769 1606 785 1640
rect 843 1606 859 1640
rect 769 1568 859 1606
rect 917 1640 1007 1656
rect 917 1606 933 1640
rect 991 1606 1007 1640
rect 917 1568 1007 1606
rect 1065 1640 1155 1656
rect 1065 1606 1081 1640
rect 1139 1606 1155 1640
rect 1065 1568 1155 1606
rect 1213 1640 1303 1656
rect 1213 1606 1229 1640
rect 1287 1606 1303 1640
rect 1213 1568 1303 1606
rect 1361 1640 1451 1656
rect 1361 1606 1377 1640
rect 1435 1606 1451 1640
rect 1361 1568 1451 1606
rect 1509 1640 1599 1656
rect 1509 1606 1525 1640
rect 1583 1606 1599 1640
rect 1509 1568 1599 1606
rect 1657 1640 1747 1656
rect 1657 1606 1673 1640
rect 1731 1606 1747 1640
rect 1657 1568 1747 1606
rect 1805 1640 1895 1656
rect 1805 1606 1821 1640
rect 1879 1606 1895 1640
rect 1805 1568 1895 1606
rect 1953 1640 2043 1656
rect 1953 1606 1969 1640
rect 2027 1606 2043 1640
rect 1953 1568 2043 1606
rect 2101 1640 2191 1656
rect 2101 1606 2117 1640
rect 2175 1606 2191 1640
rect 2101 1568 2191 1606
rect 2249 1640 2339 1656
rect 2249 1606 2265 1640
rect 2323 1606 2339 1640
rect 2249 1568 2339 1606
rect 2397 1640 2487 1656
rect 2397 1606 2413 1640
rect 2471 1606 2487 1640
rect 2397 1568 2487 1606
rect 2545 1640 2635 1656
rect 2545 1606 2561 1640
rect 2619 1606 2635 1640
rect 2545 1568 2635 1606
rect 2693 1640 2783 1656
rect 2693 1606 2709 1640
rect 2767 1606 2783 1640
rect 2693 1568 2783 1606
rect 2841 1640 2931 1656
rect 2841 1606 2857 1640
rect 2915 1606 2931 1640
rect 2841 1568 2931 1606
rect 2989 1640 3079 1656
rect 2989 1606 3005 1640
rect 3063 1606 3079 1640
rect 2989 1568 3079 1606
rect 3137 1640 3227 1656
rect 3137 1606 3153 1640
rect 3211 1606 3227 1640
rect 3137 1568 3227 1606
rect 3285 1640 3375 1656
rect 3285 1606 3301 1640
rect 3359 1606 3375 1640
rect 3285 1568 3375 1606
rect 3433 1640 3523 1656
rect 3433 1606 3449 1640
rect 3507 1606 3523 1640
rect 3433 1568 3523 1606
rect 3581 1640 3671 1656
rect 3581 1606 3597 1640
rect 3655 1606 3671 1640
rect 3581 1568 3671 1606
rect -3671 630 -3581 668
rect -3671 596 -3655 630
rect -3597 596 -3581 630
rect -3671 580 -3581 596
rect -3523 630 -3433 668
rect -3523 596 -3507 630
rect -3449 596 -3433 630
rect -3523 580 -3433 596
rect -3375 630 -3285 668
rect -3375 596 -3359 630
rect -3301 596 -3285 630
rect -3375 580 -3285 596
rect -3227 630 -3137 668
rect -3227 596 -3211 630
rect -3153 596 -3137 630
rect -3227 580 -3137 596
rect -3079 630 -2989 668
rect -3079 596 -3063 630
rect -3005 596 -2989 630
rect -3079 580 -2989 596
rect -2931 630 -2841 668
rect -2931 596 -2915 630
rect -2857 596 -2841 630
rect -2931 580 -2841 596
rect -2783 630 -2693 668
rect -2783 596 -2767 630
rect -2709 596 -2693 630
rect -2783 580 -2693 596
rect -2635 630 -2545 668
rect -2635 596 -2619 630
rect -2561 596 -2545 630
rect -2635 580 -2545 596
rect -2487 630 -2397 668
rect -2487 596 -2471 630
rect -2413 596 -2397 630
rect -2487 580 -2397 596
rect -2339 630 -2249 668
rect -2339 596 -2323 630
rect -2265 596 -2249 630
rect -2339 580 -2249 596
rect -2191 630 -2101 668
rect -2191 596 -2175 630
rect -2117 596 -2101 630
rect -2191 580 -2101 596
rect -2043 630 -1953 668
rect -2043 596 -2027 630
rect -1969 596 -1953 630
rect -2043 580 -1953 596
rect -1895 630 -1805 668
rect -1895 596 -1879 630
rect -1821 596 -1805 630
rect -1895 580 -1805 596
rect -1747 630 -1657 668
rect -1747 596 -1731 630
rect -1673 596 -1657 630
rect -1747 580 -1657 596
rect -1599 630 -1509 668
rect -1599 596 -1583 630
rect -1525 596 -1509 630
rect -1599 580 -1509 596
rect -1451 630 -1361 668
rect -1451 596 -1435 630
rect -1377 596 -1361 630
rect -1451 580 -1361 596
rect -1303 630 -1213 668
rect -1303 596 -1287 630
rect -1229 596 -1213 630
rect -1303 580 -1213 596
rect -1155 630 -1065 668
rect -1155 596 -1139 630
rect -1081 596 -1065 630
rect -1155 580 -1065 596
rect -1007 630 -917 668
rect -1007 596 -991 630
rect -933 596 -917 630
rect -1007 580 -917 596
rect -859 630 -769 668
rect -859 596 -843 630
rect -785 596 -769 630
rect -859 580 -769 596
rect -711 630 -621 668
rect -711 596 -695 630
rect -637 596 -621 630
rect -711 580 -621 596
rect -563 630 -473 668
rect -563 596 -547 630
rect -489 596 -473 630
rect -563 580 -473 596
rect -415 630 -325 668
rect -415 596 -399 630
rect -341 596 -325 630
rect -415 580 -325 596
rect -267 630 -177 668
rect -267 596 -251 630
rect -193 596 -177 630
rect -267 580 -177 596
rect -119 630 -29 668
rect -119 596 -103 630
rect -45 596 -29 630
rect -119 580 -29 596
rect 29 630 119 668
rect 29 596 45 630
rect 103 596 119 630
rect 29 580 119 596
rect 177 630 267 668
rect 177 596 193 630
rect 251 596 267 630
rect 177 580 267 596
rect 325 630 415 668
rect 325 596 341 630
rect 399 596 415 630
rect 325 580 415 596
rect 473 630 563 668
rect 473 596 489 630
rect 547 596 563 630
rect 473 580 563 596
rect 621 630 711 668
rect 621 596 637 630
rect 695 596 711 630
rect 621 580 711 596
rect 769 630 859 668
rect 769 596 785 630
rect 843 596 859 630
rect 769 580 859 596
rect 917 630 1007 668
rect 917 596 933 630
rect 991 596 1007 630
rect 917 580 1007 596
rect 1065 630 1155 668
rect 1065 596 1081 630
rect 1139 596 1155 630
rect 1065 580 1155 596
rect 1213 630 1303 668
rect 1213 596 1229 630
rect 1287 596 1303 630
rect 1213 580 1303 596
rect 1361 630 1451 668
rect 1361 596 1377 630
rect 1435 596 1451 630
rect 1361 580 1451 596
rect 1509 630 1599 668
rect 1509 596 1525 630
rect 1583 596 1599 630
rect 1509 580 1599 596
rect 1657 630 1747 668
rect 1657 596 1673 630
rect 1731 596 1747 630
rect 1657 580 1747 596
rect 1805 630 1895 668
rect 1805 596 1821 630
rect 1879 596 1895 630
rect 1805 580 1895 596
rect 1953 630 2043 668
rect 1953 596 1969 630
rect 2027 596 2043 630
rect 1953 580 2043 596
rect 2101 630 2191 668
rect 2101 596 2117 630
rect 2175 596 2191 630
rect 2101 580 2191 596
rect 2249 630 2339 668
rect 2249 596 2265 630
rect 2323 596 2339 630
rect 2249 580 2339 596
rect 2397 630 2487 668
rect 2397 596 2413 630
rect 2471 596 2487 630
rect 2397 580 2487 596
rect 2545 630 2635 668
rect 2545 596 2561 630
rect 2619 596 2635 630
rect 2545 580 2635 596
rect 2693 630 2783 668
rect 2693 596 2709 630
rect 2767 596 2783 630
rect 2693 580 2783 596
rect 2841 630 2931 668
rect 2841 596 2857 630
rect 2915 596 2931 630
rect 2841 580 2931 596
rect 2989 630 3079 668
rect 2989 596 3005 630
rect 3063 596 3079 630
rect 2989 580 3079 596
rect 3137 630 3227 668
rect 3137 596 3153 630
rect 3211 596 3227 630
rect 3137 580 3227 596
rect 3285 630 3375 668
rect 3285 596 3301 630
rect 3359 596 3375 630
rect 3285 580 3375 596
rect 3433 630 3523 668
rect 3433 596 3449 630
rect 3507 596 3523 630
rect 3433 580 3523 596
rect 3581 630 3671 668
rect 3581 596 3597 630
rect 3655 596 3671 630
rect 3581 580 3671 596
rect -3671 522 -3581 538
rect -3671 488 -3655 522
rect -3597 488 -3581 522
rect -3671 450 -3581 488
rect -3523 522 -3433 538
rect -3523 488 -3507 522
rect -3449 488 -3433 522
rect -3523 450 -3433 488
rect -3375 522 -3285 538
rect -3375 488 -3359 522
rect -3301 488 -3285 522
rect -3375 450 -3285 488
rect -3227 522 -3137 538
rect -3227 488 -3211 522
rect -3153 488 -3137 522
rect -3227 450 -3137 488
rect -3079 522 -2989 538
rect -3079 488 -3063 522
rect -3005 488 -2989 522
rect -3079 450 -2989 488
rect -2931 522 -2841 538
rect -2931 488 -2915 522
rect -2857 488 -2841 522
rect -2931 450 -2841 488
rect -2783 522 -2693 538
rect -2783 488 -2767 522
rect -2709 488 -2693 522
rect -2783 450 -2693 488
rect -2635 522 -2545 538
rect -2635 488 -2619 522
rect -2561 488 -2545 522
rect -2635 450 -2545 488
rect -2487 522 -2397 538
rect -2487 488 -2471 522
rect -2413 488 -2397 522
rect -2487 450 -2397 488
rect -2339 522 -2249 538
rect -2339 488 -2323 522
rect -2265 488 -2249 522
rect -2339 450 -2249 488
rect -2191 522 -2101 538
rect -2191 488 -2175 522
rect -2117 488 -2101 522
rect -2191 450 -2101 488
rect -2043 522 -1953 538
rect -2043 488 -2027 522
rect -1969 488 -1953 522
rect -2043 450 -1953 488
rect -1895 522 -1805 538
rect -1895 488 -1879 522
rect -1821 488 -1805 522
rect -1895 450 -1805 488
rect -1747 522 -1657 538
rect -1747 488 -1731 522
rect -1673 488 -1657 522
rect -1747 450 -1657 488
rect -1599 522 -1509 538
rect -1599 488 -1583 522
rect -1525 488 -1509 522
rect -1599 450 -1509 488
rect -1451 522 -1361 538
rect -1451 488 -1435 522
rect -1377 488 -1361 522
rect -1451 450 -1361 488
rect -1303 522 -1213 538
rect -1303 488 -1287 522
rect -1229 488 -1213 522
rect -1303 450 -1213 488
rect -1155 522 -1065 538
rect -1155 488 -1139 522
rect -1081 488 -1065 522
rect -1155 450 -1065 488
rect -1007 522 -917 538
rect -1007 488 -991 522
rect -933 488 -917 522
rect -1007 450 -917 488
rect -859 522 -769 538
rect -859 488 -843 522
rect -785 488 -769 522
rect -859 450 -769 488
rect -711 522 -621 538
rect -711 488 -695 522
rect -637 488 -621 522
rect -711 450 -621 488
rect -563 522 -473 538
rect -563 488 -547 522
rect -489 488 -473 522
rect -563 450 -473 488
rect -415 522 -325 538
rect -415 488 -399 522
rect -341 488 -325 522
rect -415 450 -325 488
rect -267 522 -177 538
rect -267 488 -251 522
rect -193 488 -177 522
rect -267 450 -177 488
rect -119 522 -29 538
rect -119 488 -103 522
rect -45 488 -29 522
rect -119 450 -29 488
rect 29 522 119 538
rect 29 488 45 522
rect 103 488 119 522
rect 29 450 119 488
rect 177 522 267 538
rect 177 488 193 522
rect 251 488 267 522
rect 177 450 267 488
rect 325 522 415 538
rect 325 488 341 522
rect 399 488 415 522
rect 325 450 415 488
rect 473 522 563 538
rect 473 488 489 522
rect 547 488 563 522
rect 473 450 563 488
rect 621 522 711 538
rect 621 488 637 522
rect 695 488 711 522
rect 621 450 711 488
rect 769 522 859 538
rect 769 488 785 522
rect 843 488 859 522
rect 769 450 859 488
rect 917 522 1007 538
rect 917 488 933 522
rect 991 488 1007 522
rect 917 450 1007 488
rect 1065 522 1155 538
rect 1065 488 1081 522
rect 1139 488 1155 522
rect 1065 450 1155 488
rect 1213 522 1303 538
rect 1213 488 1229 522
rect 1287 488 1303 522
rect 1213 450 1303 488
rect 1361 522 1451 538
rect 1361 488 1377 522
rect 1435 488 1451 522
rect 1361 450 1451 488
rect 1509 522 1599 538
rect 1509 488 1525 522
rect 1583 488 1599 522
rect 1509 450 1599 488
rect 1657 522 1747 538
rect 1657 488 1673 522
rect 1731 488 1747 522
rect 1657 450 1747 488
rect 1805 522 1895 538
rect 1805 488 1821 522
rect 1879 488 1895 522
rect 1805 450 1895 488
rect 1953 522 2043 538
rect 1953 488 1969 522
rect 2027 488 2043 522
rect 1953 450 2043 488
rect 2101 522 2191 538
rect 2101 488 2117 522
rect 2175 488 2191 522
rect 2101 450 2191 488
rect 2249 522 2339 538
rect 2249 488 2265 522
rect 2323 488 2339 522
rect 2249 450 2339 488
rect 2397 522 2487 538
rect 2397 488 2413 522
rect 2471 488 2487 522
rect 2397 450 2487 488
rect 2545 522 2635 538
rect 2545 488 2561 522
rect 2619 488 2635 522
rect 2545 450 2635 488
rect 2693 522 2783 538
rect 2693 488 2709 522
rect 2767 488 2783 522
rect 2693 450 2783 488
rect 2841 522 2931 538
rect 2841 488 2857 522
rect 2915 488 2931 522
rect 2841 450 2931 488
rect 2989 522 3079 538
rect 2989 488 3005 522
rect 3063 488 3079 522
rect 2989 450 3079 488
rect 3137 522 3227 538
rect 3137 488 3153 522
rect 3211 488 3227 522
rect 3137 450 3227 488
rect 3285 522 3375 538
rect 3285 488 3301 522
rect 3359 488 3375 522
rect 3285 450 3375 488
rect 3433 522 3523 538
rect 3433 488 3449 522
rect 3507 488 3523 522
rect 3433 450 3523 488
rect 3581 522 3671 538
rect 3581 488 3597 522
rect 3655 488 3671 522
rect 3581 450 3671 488
rect -3671 -488 -3581 -450
rect -3671 -522 -3655 -488
rect -3597 -522 -3581 -488
rect -3671 -538 -3581 -522
rect -3523 -488 -3433 -450
rect -3523 -522 -3507 -488
rect -3449 -522 -3433 -488
rect -3523 -538 -3433 -522
rect -3375 -488 -3285 -450
rect -3375 -522 -3359 -488
rect -3301 -522 -3285 -488
rect -3375 -538 -3285 -522
rect -3227 -488 -3137 -450
rect -3227 -522 -3211 -488
rect -3153 -522 -3137 -488
rect -3227 -538 -3137 -522
rect -3079 -488 -2989 -450
rect -3079 -522 -3063 -488
rect -3005 -522 -2989 -488
rect -3079 -538 -2989 -522
rect -2931 -488 -2841 -450
rect -2931 -522 -2915 -488
rect -2857 -522 -2841 -488
rect -2931 -538 -2841 -522
rect -2783 -488 -2693 -450
rect -2783 -522 -2767 -488
rect -2709 -522 -2693 -488
rect -2783 -538 -2693 -522
rect -2635 -488 -2545 -450
rect -2635 -522 -2619 -488
rect -2561 -522 -2545 -488
rect -2635 -538 -2545 -522
rect -2487 -488 -2397 -450
rect -2487 -522 -2471 -488
rect -2413 -522 -2397 -488
rect -2487 -538 -2397 -522
rect -2339 -488 -2249 -450
rect -2339 -522 -2323 -488
rect -2265 -522 -2249 -488
rect -2339 -538 -2249 -522
rect -2191 -488 -2101 -450
rect -2191 -522 -2175 -488
rect -2117 -522 -2101 -488
rect -2191 -538 -2101 -522
rect -2043 -488 -1953 -450
rect -2043 -522 -2027 -488
rect -1969 -522 -1953 -488
rect -2043 -538 -1953 -522
rect -1895 -488 -1805 -450
rect -1895 -522 -1879 -488
rect -1821 -522 -1805 -488
rect -1895 -538 -1805 -522
rect -1747 -488 -1657 -450
rect -1747 -522 -1731 -488
rect -1673 -522 -1657 -488
rect -1747 -538 -1657 -522
rect -1599 -488 -1509 -450
rect -1599 -522 -1583 -488
rect -1525 -522 -1509 -488
rect -1599 -538 -1509 -522
rect -1451 -488 -1361 -450
rect -1451 -522 -1435 -488
rect -1377 -522 -1361 -488
rect -1451 -538 -1361 -522
rect -1303 -488 -1213 -450
rect -1303 -522 -1287 -488
rect -1229 -522 -1213 -488
rect -1303 -538 -1213 -522
rect -1155 -488 -1065 -450
rect -1155 -522 -1139 -488
rect -1081 -522 -1065 -488
rect -1155 -538 -1065 -522
rect -1007 -488 -917 -450
rect -1007 -522 -991 -488
rect -933 -522 -917 -488
rect -1007 -538 -917 -522
rect -859 -488 -769 -450
rect -859 -522 -843 -488
rect -785 -522 -769 -488
rect -859 -538 -769 -522
rect -711 -488 -621 -450
rect -711 -522 -695 -488
rect -637 -522 -621 -488
rect -711 -538 -621 -522
rect -563 -488 -473 -450
rect -563 -522 -547 -488
rect -489 -522 -473 -488
rect -563 -538 -473 -522
rect -415 -488 -325 -450
rect -415 -522 -399 -488
rect -341 -522 -325 -488
rect -415 -538 -325 -522
rect -267 -488 -177 -450
rect -267 -522 -251 -488
rect -193 -522 -177 -488
rect -267 -538 -177 -522
rect -119 -488 -29 -450
rect -119 -522 -103 -488
rect -45 -522 -29 -488
rect -119 -538 -29 -522
rect 29 -488 119 -450
rect 29 -522 45 -488
rect 103 -522 119 -488
rect 29 -538 119 -522
rect 177 -488 267 -450
rect 177 -522 193 -488
rect 251 -522 267 -488
rect 177 -538 267 -522
rect 325 -488 415 -450
rect 325 -522 341 -488
rect 399 -522 415 -488
rect 325 -538 415 -522
rect 473 -488 563 -450
rect 473 -522 489 -488
rect 547 -522 563 -488
rect 473 -538 563 -522
rect 621 -488 711 -450
rect 621 -522 637 -488
rect 695 -522 711 -488
rect 621 -538 711 -522
rect 769 -488 859 -450
rect 769 -522 785 -488
rect 843 -522 859 -488
rect 769 -538 859 -522
rect 917 -488 1007 -450
rect 917 -522 933 -488
rect 991 -522 1007 -488
rect 917 -538 1007 -522
rect 1065 -488 1155 -450
rect 1065 -522 1081 -488
rect 1139 -522 1155 -488
rect 1065 -538 1155 -522
rect 1213 -488 1303 -450
rect 1213 -522 1229 -488
rect 1287 -522 1303 -488
rect 1213 -538 1303 -522
rect 1361 -488 1451 -450
rect 1361 -522 1377 -488
rect 1435 -522 1451 -488
rect 1361 -538 1451 -522
rect 1509 -488 1599 -450
rect 1509 -522 1525 -488
rect 1583 -522 1599 -488
rect 1509 -538 1599 -522
rect 1657 -488 1747 -450
rect 1657 -522 1673 -488
rect 1731 -522 1747 -488
rect 1657 -538 1747 -522
rect 1805 -488 1895 -450
rect 1805 -522 1821 -488
rect 1879 -522 1895 -488
rect 1805 -538 1895 -522
rect 1953 -488 2043 -450
rect 1953 -522 1969 -488
rect 2027 -522 2043 -488
rect 1953 -538 2043 -522
rect 2101 -488 2191 -450
rect 2101 -522 2117 -488
rect 2175 -522 2191 -488
rect 2101 -538 2191 -522
rect 2249 -488 2339 -450
rect 2249 -522 2265 -488
rect 2323 -522 2339 -488
rect 2249 -538 2339 -522
rect 2397 -488 2487 -450
rect 2397 -522 2413 -488
rect 2471 -522 2487 -488
rect 2397 -538 2487 -522
rect 2545 -488 2635 -450
rect 2545 -522 2561 -488
rect 2619 -522 2635 -488
rect 2545 -538 2635 -522
rect 2693 -488 2783 -450
rect 2693 -522 2709 -488
rect 2767 -522 2783 -488
rect 2693 -538 2783 -522
rect 2841 -488 2931 -450
rect 2841 -522 2857 -488
rect 2915 -522 2931 -488
rect 2841 -538 2931 -522
rect 2989 -488 3079 -450
rect 2989 -522 3005 -488
rect 3063 -522 3079 -488
rect 2989 -538 3079 -522
rect 3137 -488 3227 -450
rect 3137 -522 3153 -488
rect 3211 -522 3227 -488
rect 3137 -538 3227 -522
rect 3285 -488 3375 -450
rect 3285 -522 3301 -488
rect 3359 -522 3375 -488
rect 3285 -538 3375 -522
rect 3433 -488 3523 -450
rect 3433 -522 3449 -488
rect 3507 -522 3523 -488
rect 3433 -538 3523 -522
rect 3581 -488 3671 -450
rect 3581 -522 3597 -488
rect 3655 -522 3671 -488
rect 3581 -538 3671 -522
rect -3671 -596 -3581 -580
rect -3671 -630 -3655 -596
rect -3597 -630 -3581 -596
rect -3671 -668 -3581 -630
rect -3523 -596 -3433 -580
rect -3523 -630 -3507 -596
rect -3449 -630 -3433 -596
rect -3523 -668 -3433 -630
rect -3375 -596 -3285 -580
rect -3375 -630 -3359 -596
rect -3301 -630 -3285 -596
rect -3375 -668 -3285 -630
rect -3227 -596 -3137 -580
rect -3227 -630 -3211 -596
rect -3153 -630 -3137 -596
rect -3227 -668 -3137 -630
rect -3079 -596 -2989 -580
rect -3079 -630 -3063 -596
rect -3005 -630 -2989 -596
rect -3079 -668 -2989 -630
rect -2931 -596 -2841 -580
rect -2931 -630 -2915 -596
rect -2857 -630 -2841 -596
rect -2931 -668 -2841 -630
rect -2783 -596 -2693 -580
rect -2783 -630 -2767 -596
rect -2709 -630 -2693 -596
rect -2783 -668 -2693 -630
rect -2635 -596 -2545 -580
rect -2635 -630 -2619 -596
rect -2561 -630 -2545 -596
rect -2635 -668 -2545 -630
rect -2487 -596 -2397 -580
rect -2487 -630 -2471 -596
rect -2413 -630 -2397 -596
rect -2487 -668 -2397 -630
rect -2339 -596 -2249 -580
rect -2339 -630 -2323 -596
rect -2265 -630 -2249 -596
rect -2339 -668 -2249 -630
rect -2191 -596 -2101 -580
rect -2191 -630 -2175 -596
rect -2117 -630 -2101 -596
rect -2191 -668 -2101 -630
rect -2043 -596 -1953 -580
rect -2043 -630 -2027 -596
rect -1969 -630 -1953 -596
rect -2043 -668 -1953 -630
rect -1895 -596 -1805 -580
rect -1895 -630 -1879 -596
rect -1821 -630 -1805 -596
rect -1895 -668 -1805 -630
rect -1747 -596 -1657 -580
rect -1747 -630 -1731 -596
rect -1673 -630 -1657 -596
rect -1747 -668 -1657 -630
rect -1599 -596 -1509 -580
rect -1599 -630 -1583 -596
rect -1525 -630 -1509 -596
rect -1599 -668 -1509 -630
rect -1451 -596 -1361 -580
rect -1451 -630 -1435 -596
rect -1377 -630 -1361 -596
rect -1451 -668 -1361 -630
rect -1303 -596 -1213 -580
rect -1303 -630 -1287 -596
rect -1229 -630 -1213 -596
rect -1303 -668 -1213 -630
rect -1155 -596 -1065 -580
rect -1155 -630 -1139 -596
rect -1081 -630 -1065 -596
rect -1155 -668 -1065 -630
rect -1007 -596 -917 -580
rect -1007 -630 -991 -596
rect -933 -630 -917 -596
rect -1007 -668 -917 -630
rect -859 -596 -769 -580
rect -859 -630 -843 -596
rect -785 -630 -769 -596
rect -859 -668 -769 -630
rect -711 -596 -621 -580
rect -711 -630 -695 -596
rect -637 -630 -621 -596
rect -711 -668 -621 -630
rect -563 -596 -473 -580
rect -563 -630 -547 -596
rect -489 -630 -473 -596
rect -563 -668 -473 -630
rect -415 -596 -325 -580
rect -415 -630 -399 -596
rect -341 -630 -325 -596
rect -415 -668 -325 -630
rect -267 -596 -177 -580
rect -267 -630 -251 -596
rect -193 -630 -177 -596
rect -267 -668 -177 -630
rect -119 -596 -29 -580
rect -119 -630 -103 -596
rect -45 -630 -29 -596
rect -119 -668 -29 -630
rect 29 -596 119 -580
rect 29 -630 45 -596
rect 103 -630 119 -596
rect 29 -668 119 -630
rect 177 -596 267 -580
rect 177 -630 193 -596
rect 251 -630 267 -596
rect 177 -668 267 -630
rect 325 -596 415 -580
rect 325 -630 341 -596
rect 399 -630 415 -596
rect 325 -668 415 -630
rect 473 -596 563 -580
rect 473 -630 489 -596
rect 547 -630 563 -596
rect 473 -668 563 -630
rect 621 -596 711 -580
rect 621 -630 637 -596
rect 695 -630 711 -596
rect 621 -668 711 -630
rect 769 -596 859 -580
rect 769 -630 785 -596
rect 843 -630 859 -596
rect 769 -668 859 -630
rect 917 -596 1007 -580
rect 917 -630 933 -596
rect 991 -630 1007 -596
rect 917 -668 1007 -630
rect 1065 -596 1155 -580
rect 1065 -630 1081 -596
rect 1139 -630 1155 -596
rect 1065 -668 1155 -630
rect 1213 -596 1303 -580
rect 1213 -630 1229 -596
rect 1287 -630 1303 -596
rect 1213 -668 1303 -630
rect 1361 -596 1451 -580
rect 1361 -630 1377 -596
rect 1435 -630 1451 -596
rect 1361 -668 1451 -630
rect 1509 -596 1599 -580
rect 1509 -630 1525 -596
rect 1583 -630 1599 -596
rect 1509 -668 1599 -630
rect 1657 -596 1747 -580
rect 1657 -630 1673 -596
rect 1731 -630 1747 -596
rect 1657 -668 1747 -630
rect 1805 -596 1895 -580
rect 1805 -630 1821 -596
rect 1879 -630 1895 -596
rect 1805 -668 1895 -630
rect 1953 -596 2043 -580
rect 1953 -630 1969 -596
rect 2027 -630 2043 -596
rect 1953 -668 2043 -630
rect 2101 -596 2191 -580
rect 2101 -630 2117 -596
rect 2175 -630 2191 -596
rect 2101 -668 2191 -630
rect 2249 -596 2339 -580
rect 2249 -630 2265 -596
rect 2323 -630 2339 -596
rect 2249 -668 2339 -630
rect 2397 -596 2487 -580
rect 2397 -630 2413 -596
rect 2471 -630 2487 -596
rect 2397 -668 2487 -630
rect 2545 -596 2635 -580
rect 2545 -630 2561 -596
rect 2619 -630 2635 -596
rect 2545 -668 2635 -630
rect 2693 -596 2783 -580
rect 2693 -630 2709 -596
rect 2767 -630 2783 -596
rect 2693 -668 2783 -630
rect 2841 -596 2931 -580
rect 2841 -630 2857 -596
rect 2915 -630 2931 -596
rect 2841 -668 2931 -630
rect 2989 -596 3079 -580
rect 2989 -630 3005 -596
rect 3063 -630 3079 -596
rect 2989 -668 3079 -630
rect 3137 -596 3227 -580
rect 3137 -630 3153 -596
rect 3211 -630 3227 -596
rect 3137 -668 3227 -630
rect 3285 -596 3375 -580
rect 3285 -630 3301 -596
rect 3359 -630 3375 -596
rect 3285 -668 3375 -630
rect 3433 -596 3523 -580
rect 3433 -630 3449 -596
rect 3507 -630 3523 -596
rect 3433 -668 3523 -630
rect 3581 -596 3671 -580
rect 3581 -630 3597 -596
rect 3655 -630 3671 -596
rect 3581 -668 3671 -630
rect -3671 -1606 -3581 -1568
rect -3671 -1640 -3655 -1606
rect -3597 -1640 -3581 -1606
rect -3671 -1656 -3581 -1640
rect -3523 -1606 -3433 -1568
rect -3523 -1640 -3507 -1606
rect -3449 -1640 -3433 -1606
rect -3523 -1656 -3433 -1640
rect -3375 -1606 -3285 -1568
rect -3375 -1640 -3359 -1606
rect -3301 -1640 -3285 -1606
rect -3375 -1656 -3285 -1640
rect -3227 -1606 -3137 -1568
rect -3227 -1640 -3211 -1606
rect -3153 -1640 -3137 -1606
rect -3227 -1656 -3137 -1640
rect -3079 -1606 -2989 -1568
rect -3079 -1640 -3063 -1606
rect -3005 -1640 -2989 -1606
rect -3079 -1656 -2989 -1640
rect -2931 -1606 -2841 -1568
rect -2931 -1640 -2915 -1606
rect -2857 -1640 -2841 -1606
rect -2931 -1656 -2841 -1640
rect -2783 -1606 -2693 -1568
rect -2783 -1640 -2767 -1606
rect -2709 -1640 -2693 -1606
rect -2783 -1656 -2693 -1640
rect -2635 -1606 -2545 -1568
rect -2635 -1640 -2619 -1606
rect -2561 -1640 -2545 -1606
rect -2635 -1656 -2545 -1640
rect -2487 -1606 -2397 -1568
rect -2487 -1640 -2471 -1606
rect -2413 -1640 -2397 -1606
rect -2487 -1656 -2397 -1640
rect -2339 -1606 -2249 -1568
rect -2339 -1640 -2323 -1606
rect -2265 -1640 -2249 -1606
rect -2339 -1656 -2249 -1640
rect -2191 -1606 -2101 -1568
rect -2191 -1640 -2175 -1606
rect -2117 -1640 -2101 -1606
rect -2191 -1656 -2101 -1640
rect -2043 -1606 -1953 -1568
rect -2043 -1640 -2027 -1606
rect -1969 -1640 -1953 -1606
rect -2043 -1656 -1953 -1640
rect -1895 -1606 -1805 -1568
rect -1895 -1640 -1879 -1606
rect -1821 -1640 -1805 -1606
rect -1895 -1656 -1805 -1640
rect -1747 -1606 -1657 -1568
rect -1747 -1640 -1731 -1606
rect -1673 -1640 -1657 -1606
rect -1747 -1656 -1657 -1640
rect -1599 -1606 -1509 -1568
rect -1599 -1640 -1583 -1606
rect -1525 -1640 -1509 -1606
rect -1599 -1656 -1509 -1640
rect -1451 -1606 -1361 -1568
rect -1451 -1640 -1435 -1606
rect -1377 -1640 -1361 -1606
rect -1451 -1656 -1361 -1640
rect -1303 -1606 -1213 -1568
rect -1303 -1640 -1287 -1606
rect -1229 -1640 -1213 -1606
rect -1303 -1656 -1213 -1640
rect -1155 -1606 -1065 -1568
rect -1155 -1640 -1139 -1606
rect -1081 -1640 -1065 -1606
rect -1155 -1656 -1065 -1640
rect -1007 -1606 -917 -1568
rect -1007 -1640 -991 -1606
rect -933 -1640 -917 -1606
rect -1007 -1656 -917 -1640
rect -859 -1606 -769 -1568
rect -859 -1640 -843 -1606
rect -785 -1640 -769 -1606
rect -859 -1656 -769 -1640
rect -711 -1606 -621 -1568
rect -711 -1640 -695 -1606
rect -637 -1640 -621 -1606
rect -711 -1656 -621 -1640
rect -563 -1606 -473 -1568
rect -563 -1640 -547 -1606
rect -489 -1640 -473 -1606
rect -563 -1656 -473 -1640
rect -415 -1606 -325 -1568
rect -415 -1640 -399 -1606
rect -341 -1640 -325 -1606
rect -415 -1656 -325 -1640
rect -267 -1606 -177 -1568
rect -267 -1640 -251 -1606
rect -193 -1640 -177 -1606
rect -267 -1656 -177 -1640
rect -119 -1606 -29 -1568
rect -119 -1640 -103 -1606
rect -45 -1640 -29 -1606
rect -119 -1656 -29 -1640
rect 29 -1606 119 -1568
rect 29 -1640 45 -1606
rect 103 -1640 119 -1606
rect 29 -1656 119 -1640
rect 177 -1606 267 -1568
rect 177 -1640 193 -1606
rect 251 -1640 267 -1606
rect 177 -1656 267 -1640
rect 325 -1606 415 -1568
rect 325 -1640 341 -1606
rect 399 -1640 415 -1606
rect 325 -1656 415 -1640
rect 473 -1606 563 -1568
rect 473 -1640 489 -1606
rect 547 -1640 563 -1606
rect 473 -1656 563 -1640
rect 621 -1606 711 -1568
rect 621 -1640 637 -1606
rect 695 -1640 711 -1606
rect 621 -1656 711 -1640
rect 769 -1606 859 -1568
rect 769 -1640 785 -1606
rect 843 -1640 859 -1606
rect 769 -1656 859 -1640
rect 917 -1606 1007 -1568
rect 917 -1640 933 -1606
rect 991 -1640 1007 -1606
rect 917 -1656 1007 -1640
rect 1065 -1606 1155 -1568
rect 1065 -1640 1081 -1606
rect 1139 -1640 1155 -1606
rect 1065 -1656 1155 -1640
rect 1213 -1606 1303 -1568
rect 1213 -1640 1229 -1606
rect 1287 -1640 1303 -1606
rect 1213 -1656 1303 -1640
rect 1361 -1606 1451 -1568
rect 1361 -1640 1377 -1606
rect 1435 -1640 1451 -1606
rect 1361 -1656 1451 -1640
rect 1509 -1606 1599 -1568
rect 1509 -1640 1525 -1606
rect 1583 -1640 1599 -1606
rect 1509 -1656 1599 -1640
rect 1657 -1606 1747 -1568
rect 1657 -1640 1673 -1606
rect 1731 -1640 1747 -1606
rect 1657 -1656 1747 -1640
rect 1805 -1606 1895 -1568
rect 1805 -1640 1821 -1606
rect 1879 -1640 1895 -1606
rect 1805 -1656 1895 -1640
rect 1953 -1606 2043 -1568
rect 1953 -1640 1969 -1606
rect 2027 -1640 2043 -1606
rect 1953 -1656 2043 -1640
rect 2101 -1606 2191 -1568
rect 2101 -1640 2117 -1606
rect 2175 -1640 2191 -1606
rect 2101 -1656 2191 -1640
rect 2249 -1606 2339 -1568
rect 2249 -1640 2265 -1606
rect 2323 -1640 2339 -1606
rect 2249 -1656 2339 -1640
rect 2397 -1606 2487 -1568
rect 2397 -1640 2413 -1606
rect 2471 -1640 2487 -1606
rect 2397 -1656 2487 -1640
rect 2545 -1606 2635 -1568
rect 2545 -1640 2561 -1606
rect 2619 -1640 2635 -1606
rect 2545 -1656 2635 -1640
rect 2693 -1606 2783 -1568
rect 2693 -1640 2709 -1606
rect 2767 -1640 2783 -1606
rect 2693 -1656 2783 -1640
rect 2841 -1606 2931 -1568
rect 2841 -1640 2857 -1606
rect 2915 -1640 2931 -1606
rect 2841 -1656 2931 -1640
rect 2989 -1606 3079 -1568
rect 2989 -1640 3005 -1606
rect 3063 -1640 3079 -1606
rect 2989 -1656 3079 -1640
rect 3137 -1606 3227 -1568
rect 3137 -1640 3153 -1606
rect 3211 -1640 3227 -1606
rect 3137 -1656 3227 -1640
rect 3285 -1606 3375 -1568
rect 3285 -1640 3301 -1606
rect 3359 -1640 3375 -1606
rect 3285 -1656 3375 -1640
rect 3433 -1606 3523 -1568
rect 3433 -1640 3449 -1606
rect 3507 -1640 3523 -1606
rect 3433 -1656 3523 -1640
rect 3581 -1606 3671 -1568
rect 3581 -1640 3597 -1606
rect 3655 -1640 3671 -1606
rect 3581 -1656 3671 -1640
<< polycont >>
rect -3655 1606 -3597 1640
rect -3507 1606 -3449 1640
rect -3359 1606 -3301 1640
rect -3211 1606 -3153 1640
rect -3063 1606 -3005 1640
rect -2915 1606 -2857 1640
rect -2767 1606 -2709 1640
rect -2619 1606 -2561 1640
rect -2471 1606 -2413 1640
rect -2323 1606 -2265 1640
rect -2175 1606 -2117 1640
rect -2027 1606 -1969 1640
rect -1879 1606 -1821 1640
rect -1731 1606 -1673 1640
rect -1583 1606 -1525 1640
rect -1435 1606 -1377 1640
rect -1287 1606 -1229 1640
rect -1139 1606 -1081 1640
rect -991 1606 -933 1640
rect -843 1606 -785 1640
rect -695 1606 -637 1640
rect -547 1606 -489 1640
rect -399 1606 -341 1640
rect -251 1606 -193 1640
rect -103 1606 -45 1640
rect 45 1606 103 1640
rect 193 1606 251 1640
rect 341 1606 399 1640
rect 489 1606 547 1640
rect 637 1606 695 1640
rect 785 1606 843 1640
rect 933 1606 991 1640
rect 1081 1606 1139 1640
rect 1229 1606 1287 1640
rect 1377 1606 1435 1640
rect 1525 1606 1583 1640
rect 1673 1606 1731 1640
rect 1821 1606 1879 1640
rect 1969 1606 2027 1640
rect 2117 1606 2175 1640
rect 2265 1606 2323 1640
rect 2413 1606 2471 1640
rect 2561 1606 2619 1640
rect 2709 1606 2767 1640
rect 2857 1606 2915 1640
rect 3005 1606 3063 1640
rect 3153 1606 3211 1640
rect 3301 1606 3359 1640
rect 3449 1606 3507 1640
rect 3597 1606 3655 1640
rect -3655 596 -3597 630
rect -3507 596 -3449 630
rect -3359 596 -3301 630
rect -3211 596 -3153 630
rect -3063 596 -3005 630
rect -2915 596 -2857 630
rect -2767 596 -2709 630
rect -2619 596 -2561 630
rect -2471 596 -2413 630
rect -2323 596 -2265 630
rect -2175 596 -2117 630
rect -2027 596 -1969 630
rect -1879 596 -1821 630
rect -1731 596 -1673 630
rect -1583 596 -1525 630
rect -1435 596 -1377 630
rect -1287 596 -1229 630
rect -1139 596 -1081 630
rect -991 596 -933 630
rect -843 596 -785 630
rect -695 596 -637 630
rect -547 596 -489 630
rect -399 596 -341 630
rect -251 596 -193 630
rect -103 596 -45 630
rect 45 596 103 630
rect 193 596 251 630
rect 341 596 399 630
rect 489 596 547 630
rect 637 596 695 630
rect 785 596 843 630
rect 933 596 991 630
rect 1081 596 1139 630
rect 1229 596 1287 630
rect 1377 596 1435 630
rect 1525 596 1583 630
rect 1673 596 1731 630
rect 1821 596 1879 630
rect 1969 596 2027 630
rect 2117 596 2175 630
rect 2265 596 2323 630
rect 2413 596 2471 630
rect 2561 596 2619 630
rect 2709 596 2767 630
rect 2857 596 2915 630
rect 3005 596 3063 630
rect 3153 596 3211 630
rect 3301 596 3359 630
rect 3449 596 3507 630
rect 3597 596 3655 630
rect -3655 488 -3597 522
rect -3507 488 -3449 522
rect -3359 488 -3301 522
rect -3211 488 -3153 522
rect -3063 488 -3005 522
rect -2915 488 -2857 522
rect -2767 488 -2709 522
rect -2619 488 -2561 522
rect -2471 488 -2413 522
rect -2323 488 -2265 522
rect -2175 488 -2117 522
rect -2027 488 -1969 522
rect -1879 488 -1821 522
rect -1731 488 -1673 522
rect -1583 488 -1525 522
rect -1435 488 -1377 522
rect -1287 488 -1229 522
rect -1139 488 -1081 522
rect -991 488 -933 522
rect -843 488 -785 522
rect -695 488 -637 522
rect -547 488 -489 522
rect -399 488 -341 522
rect -251 488 -193 522
rect -103 488 -45 522
rect 45 488 103 522
rect 193 488 251 522
rect 341 488 399 522
rect 489 488 547 522
rect 637 488 695 522
rect 785 488 843 522
rect 933 488 991 522
rect 1081 488 1139 522
rect 1229 488 1287 522
rect 1377 488 1435 522
rect 1525 488 1583 522
rect 1673 488 1731 522
rect 1821 488 1879 522
rect 1969 488 2027 522
rect 2117 488 2175 522
rect 2265 488 2323 522
rect 2413 488 2471 522
rect 2561 488 2619 522
rect 2709 488 2767 522
rect 2857 488 2915 522
rect 3005 488 3063 522
rect 3153 488 3211 522
rect 3301 488 3359 522
rect 3449 488 3507 522
rect 3597 488 3655 522
rect -3655 -522 -3597 -488
rect -3507 -522 -3449 -488
rect -3359 -522 -3301 -488
rect -3211 -522 -3153 -488
rect -3063 -522 -3005 -488
rect -2915 -522 -2857 -488
rect -2767 -522 -2709 -488
rect -2619 -522 -2561 -488
rect -2471 -522 -2413 -488
rect -2323 -522 -2265 -488
rect -2175 -522 -2117 -488
rect -2027 -522 -1969 -488
rect -1879 -522 -1821 -488
rect -1731 -522 -1673 -488
rect -1583 -522 -1525 -488
rect -1435 -522 -1377 -488
rect -1287 -522 -1229 -488
rect -1139 -522 -1081 -488
rect -991 -522 -933 -488
rect -843 -522 -785 -488
rect -695 -522 -637 -488
rect -547 -522 -489 -488
rect -399 -522 -341 -488
rect -251 -522 -193 -488
rect -103 -522 -45 -488
rect 45 -522 103 -488
rect 193 -522 251 -488
rect 341 -522 399 -488
rect 489 -522 547 -488
rect 637 -522 695 -488
rect 785 -522 843 -488
rect 933 -522 991 -488
rect 1081 -522 1139 -488
rect 1229 -522 1287 -488
rect 1377 -522 1435 -488
rect 1525 -522 1583 -488
rect 1673 -522 1731 -488
rect 1821 -522 1879 -488
rect 1969 -522 2027 -488
rect 2117 -522 2175 -488
rect 2265 -522 2323 -488
rect 2413 -522 2471 -488
rect 2561 -522 2619 -488
rect 2709 -522 2767 -488
rect 2857 -522 2915 -488
rect 3005 -522 3063 -488
rect 3153 -522 3211 -488
rect 3301 -522 3359 -488
rect 3449 -522 3507 -488
rect 3597 -522 3655 -488
rect -3655 -630 -3597 -596
rect -3507 -630 -3449 -596
rect -3359 -630 -3301 -596
rect -3211 -630 -3153 -596
rect -3063 -630 -3005 -596
rect -2915 -630 -2857 -596
rect -2767 -630 -2709 -596
rect -2619 -630 -2561 -596
rect -2471 -630 -2413 -596
rect -2323 -630 -2265 -596
rect -2175 -630 -2117 -596
rect -2027 -630 -1969 -596
rect -1879 -630 -1821 -596
rect -1731 -630 -1673 -596
rect -1583 -630 -1525 -596
rect -1435 -630 -1377 -596
rect -1287 -630 -1229 -596
rect -1139 -630 -1081 -596
rect -991 -630 -933 -596
rect -843 -630 -785 -596
rect -695 -630 -637 -596
rect -547 -630 -489 -596
rect -399 -630 -341 -596
rect -251 -630 -193 -596
rect -103 -630 -45 -596
rect 45 -630 103 -596
rect 193 -630 251 -596
rect 341 -630 399 -596
rect 489 -630 547 -596
rect 637 -630 695 -596
rect 785 -630 843 -596
rect 933 -630 991 -596
rect 1081 -630 1139 -596
rect 1229 -630 1287 -596
rect 1377 -630 1435 -596
rect 1525 -630 1583 -596
rect 1673 -630 1731 -596
rect 1821 -630 1879 -596
rect 1969 -630 2027 -596
rect 2117 -630 2175 -596
rect 2265 -630 2323 -596
rect 2413 -630 2471 -596
rect 2561 -630 2619 -596
rect 2709 -630 2767 -596
rect 2857 -630 2915 -596
rect 3005 -630 3063 -596
rect 3153 -630 3211 -596
rect 3301 -630 3359 -596
rect 3449 -630 3507 -596
rect 3597 -630 3655 -596
rect -3655 -1640 -3597 -1606
rect -3507 -1640 -3449 -1606
rect -3359 -1640 -3301 -1606
rect -3211 -1640 -3153 -1606
rect -3063 -1640 -3005 -1606
rect -2915 -1640 -2857 -1606
rect -2767 -1640 -2709 -1606
rect -2619 -1640 -2561 -1606
rect -2471 -1640 -2413 -1606
rect -2323 -1640 -2265 -1606
rect -2175 -1640 -2117 -1606
rect -2027 -1640 -1969 -1606
rect -1879 -1640 -1821 -1606
rect -1731 -1640 -1673 -1606
rect -1583 -1640 -1525 -1606
rect -1435 -1640 -1377 -1606
rect -1287 -1640 -1229 -1606
rect -1139 -1640 -1081 -1606
rect -991 -1640 -933 -1606
rect -843 -1640 -785 -1606
rect -695 -1640 -637 -1606
rect -547 -1640 -489 -1606
rect -399 -1640 -341 -1606
rect -251 -1640 -193 -1606
rect -103 -1640 -45 -1606
rect 45 -1640 103 -1606
rect 193 -1640 251 -1606
rect 341 -1640 399 -1606
rect 489 -1640 547 -1606
rect 637 -1640 695 -1606
rect 785 -1640 843 -1606
rect 933 -1640 991 -1606
rect 1081 -1640 1139 -1606
rect 1229 -1640 1287 -1606
rect 1377 -1640 1435 -1606
rect 1525 -1640 1583 -1606
rect 1673 -1640 1731 -1606
rect 1821 -1640 1879 -1606
rect 1969 -1640 2027 -1606
rect 2117 -1640 2175 -1606
rect 2265 -1640 2323 -1606
rect 2413 -1640 2471 -1606
rect 2561 -1640 2619 -1606
rect 2709 -1640 2767 -1606
rect 2857 -1640 2915 -1606
rect 3005 -1640 3063 -1606
rect 3153 -1640 3211 -1606
rect 3301 -1640 3359 -1606
rect 3449 -1640 3507 -1606
rect 3597 -1640 3655 -1606
<< locali >>
rect -3831 1708 -3735 1742
rect 3735 1708 3831 1742
rect -3831 1646 -3797 1708
rect 3797 1646 3831 1708
rect -3671 1606 -3655 1640
rect -3597 1606 -3581 1640
rect -3523 1606 -3507 1640
rect -3449 1606 -3433 1640
rect -3375 1606 -3359 1640
rect -3301 1606 -3285 1640
rect -3227 1606 -3211 1640
rect -3153 1606 -3137 1640
rect -3079 1606 -3063 1640
rect -3005 1606 -2989 1640
rect -2931 1606 -2915 1640
rect -2857 1606 -2841 1640
rect -2783 1606 -2767 1640
rect -2709 1606 -2693 1640
rect -2635 1606 -2619 1640
rect -2561 1606 -2545 1640
rect -2487 1606 -2471 1640
rect -2413 1606 -2397 1640
rect -2339 1606 -2323 1640
rect -2265 1606 -2249 1640
rect -2191 1606 -2175 1640
rect -2117 1606 -2101 1640
rect -2043 1606 -2027 1640
rect -1969 1606 -1953 1640
rect -1895 1606 -1879 1640
rect -1821 1606 -1805 1640
rect -1747 1606 -1731 1640
rect -1673 1606 -1657 1640
rect -1599 1606 -1583 1640
rect -1525 1606 -1509 1640
rect -1451 1606 -1435 1640
rect -1377 1606 -1361 1640
rect -1303 1606 -1287 1640
rect -1229 1606 -1213 1640
rect -1155 1606 -1139 1640
rect -1081 1606 -1065 1640
rect -1007 1606 -991 1640
rect -933 1606 -917 1640
rect -859 1606 -843 1640
rect -785 1606 -769 1640
rect -711 1606 -695 1640
rect -637 1606 -621 1640
rect -563 1606 -547 1640
rect -489 1606 -473 1640
rect -415 1606 -399 1640
rect -341 1606 -325 1640
rect -267 1606 -251 1640
rect -193 1606 -177 1640
rect -119 1606 -103 1640
rect -45 1606 -29 1640
rect 29 1606 45 1640
rect 103 1606 119 1640
rect 177 1606 193 1640
rect 251 1606 267 1640
rect 325 1606 341 1640
rect 399 1606 415 1640
rect 473 1606 489 1640
rect 547 1606 563 1640
rect 621 1606 637 1640
rect 695 1606 711 1640
rect 769 1606 785 1640
rect 843 1606 859 1640
rect 917 1606 933 1640
rect 991 1606 1007 1640
rect 1065 1606 1081 1640
rect 1139 1606 1155 1640
rect 1213 1606 1229 1640
rect 1287 1606 1303 1640
rect 1361 1606 1377 1640
rect 1435 1606 1451 1640
rect 1509 1606 1525 1640
rect 1583 1606 1599 1640
rect 1657 1606 1673 1640
rect 1731 1606 1747 1640
rect 1805 1606 1821 1640
rect 1879 1606 1895 1640
rect 1953 1606 1969 1640
rect 2027 1606 2043 1640
rect 2101 1606 2117 1640
rect 2175 1606 2191 1640
rect 2249 1606 2265 1640
rect 2323 1606 2339 1640
rect 2397 1606 2413 1640
rect 2471 1606 2487 1640
rect 2545 1606 2561 1640
rect 2619 1606 2635 1640
rect 2693 1606 2709 1640
rect 2767 1606 2783 1640
rect 2841 1606 2857 1640
rect 2915 1606 2931 1640
rect 2989 1606 3005 1640
rect 3063 1606 3079 1640
rect 3137 1606 3153 1640
rect 3211 1606 3227 1640
rect 3285 1606 3301 1640
rect 3359 1606 3375 1640
rect 3433 1606 3449 1640
rect 3507 1606 3523 1640
rect 3581 1606 3597 1640
rect 3655 1606 3671 1640
rect -3717 1556 -3683 1572
rect -3717 664 -3683 680
rect -3569 1556 -3535 1572
rect -3569 664 -3535 680
rect -3421 1556 -3387 1572
rect -3421 664 -3387 680
rect -3273 1556 -3239 1572
rect -3273 664 -3239 680
rect -3125 1556 -3091 1572
rect -3125 664 -3091 680
rect -2977 1556 -2943 1572
rect -2977 664 -2943 680
rect -2829 1556 -2795 1572
rect -2829 664 -2795 680
rect -2681 1556 -2647 1572
rect -2681 664 -2647 680
rect -2533 1556 -2499 1572
rect -2533 664 -2499 680
rect -2385 1556 -2351 1572
rect -2385 664 -2351 680
rect -2237 1556 -2203 1572
rect -2237 664 -2203 680
rect -2089 1556 -2055 1572
rect -2089 664 -2055 680
rect -1941 1556 -1907 1572
rect -1941 664 -1907 680
rect -1793 1556 -1759 1572
rect -1793 664 -1759 680
rect -1645 1556 -1611 1572
rect -1645 664 -1611 680
rect -1497 1556 -1463 1572
rect -1497 664 -1463 680
rect -1349 1556 -1315 1572
rect -1349 664 -1315 680
rect -1201 1556 -1167 1572
rect -1201 664 -1167 680
rect -1053 1556 -1019 1572
rect -1053 664 -1019 680
rect -905 1556 -871 1572
rect -905 664 -871 680
rect -757 1556 -723 1572
rect -757 664 -723 680
rect -609 1556 -575 1572
rect -609 664 -575 680
rect -461 1556 -427 1572
rect -461 664 -427 680
rect -313 1556 -279 1572
rect -313 664 -279 680
rect -165 1556 -131 1572
rect -165 664 -131 680
rect -17 1556 17 1572
rect -17 664 17 680
rect 131 1556 165 1572
rect 131 664 165 680
rect 279 1556 313 1572
rect 279 664 313 680
rect 427 1556 461 1572
rect 427 664 461 680
rect 575 1556 609 1572
rect 575 664 609 680
rect 723 1556 757 1572
rect 723 664 757 680
rect 871 1556 905 1572
rect 871 664 905 680
rect 1019 1556 1053 1572
rect 1019 664 1053 680
rect 1167 1556 1201 1572
rect 1167 664 1201 680
rect 1315 1556 1349 1572
rect 1315 664 1349 680
rect 1463 1556 1497 1572
rect 1463 664 1497 680
rect 1611 1556 1645 1572
rect 1611 664 1645 680
rect 1759 1556 1793 1572
rect 1759 664 1793 680
rect 1907 1556 1941 1572
rect 1907 664 1941 680
rect 2055 1556 2089 1572
rect 2055 664 2089 680
rect 2203 1556 2237 1572
rect 2203 664 2237 680
rect 2351 1556 2385 1572
rect 2351 664 2385 680
rect 2499 1556 2533 1572
rect 2499 664 2533 680
rect 2647 1556 2681 1572
rect 2647 664 2681 680
rect 2795 1556 2829 1572
rect 2795 664 2829 680
rect 2943 1556 2977 1572
rect 2943 664 2977 680
rect 3091 1556 3125 1572
rect 3091 664 3125 680
rect 3239 1556 3273 1572
rect 3239 664 3273 680
rect 3387 1556 3421 1572
rect 3387 664 3421 680
rect 3535 1556 3569 1572
rect 3535 664 3569 680
rect 3683 1556 3717 1572
rect 3683 664 3717 680
rect -3671 596 -3655 630
rect -3597 596 -3581 630
rect -3523 596 -3507 630
rect -3449 596 -3433 630
rect -3375 596 -3359 630
rect -3301 596 -3285 630
rect -3227 596 -3211 630
rect -3153 596 -3137 630
rect -3079 596 -3063 630
rect -3005 596 -2989 630
rect -2931 596 -2915 630
rect -2857 596 -2841 630
rect -2783 596 -2767 630
rect -2709 596 -2693 630
rect -2635 596 -2619 630
rect -2561 596 -2545 630
rect -2487 596 -2471 630
rect -2413 596 -2397 630
rect -2339 596 -2323 630
rect -2265 596 -2249 630
rect -2191 596 -2175 630
rect -2117 596 -2101 630
rect -2043 596 -2027 630
rect -1969 596 -1953 630
rect -1895 596 -1879 630
rect -1821 596 -1805 630
rect -1747 596 -1731 630
rect -1673 596 -1657 630
rect -1599 596 -1583 630
rect -1525 596 -1509 630
rect -1451 596 -1435 630
rect -1377 596 -1361 630
rect -1303 596 -1287 630
rect -1229 596 -1213 630
rect -1155 596 -1139 630
rect -1081 596 -1065 630
rect -1007 596 -991 630
rect -933 596 -917 630
rect -859 596 -843 630
rect -785 596 -769 630
rect -711 596 -695 630
rect -637 596 -621 630
rect -563 596 -547 630
rect -489 596 -473 630
rect -415 596 -399 630
rect -341 596 -325 630
rect -267 596 -251 630
rect -193 596 -177 630
rect -119 596 -103 630
rect -45 596 -29 630
rect 29 596 45 630
rect 103 596 119 630
rect 177 596 193 630
rect 251 596 267 630
rect 325 596 341 630
rect 399 596 415 630
rect 473 596 489 630
rect 547 596 563 630
rect 621 596 637 630
rect 695 596 711 630
rect 769 596 785 630
rect 843 596 859 630
rect 917 596 933 630
rect 991 596 1007 630
rect 1065 596 1081 630
rect 1139 596 1155 630
rect 1213 596 1229 630
rect 1287 596 1303 630
rect 1361 596 1377 630
rect 1435 596 1451 630
rect 1509 596 1525 630
rect 1583 596 1599 630
rect 1657 596 1673 630
rect 1731 596 1747 630
rect 1805 596 1821 630
rect 1879 596 1895 630
rect 1953 596 1969 630
rect 2027 596 2043 630
rect 2101 596 2117 630
rect 2175 596 2191 630
rect 2249 596 2265 630
rect 2323 596 2339 630
rect 2397 596 2413 630
rect 2471 596 2487 630
rect 2545 596 2561 630
rect 2619 596 2635 630
rect 2693 596 2709 630
rect 2767 596 2783 630
rect 2841 596 2857 630
rect 2915 596 2931 630
rect 2989 596 3005 630
rect 3063 596 3079 630
rect 3137 596 3153 630
rect 3211 596 3227 630
rect 3285 596 3301 630
rect 3359 596 3375 630
rect 3433 596 3449 630
rect 3507 596 3523 630
rect 3581 596 3597 630
rect 3655 596 3671 630
rect -3671 488 -3655 522
rect -3597 488 -3581 522
rect -3523 488 -3507 522
rect -3449 488 -3433 522
rect -3375 488 -3359 522
rect -3301 488 -3285 522
rect -3227 488 -3211 522
rect -3153 488 -3137 522
rect -3079 488 -3063 522
rect -3005 488 -2989 522
rect -2931 488 -2915 522
rect -2857 488 -2841 522
rect -2783 488 -2767 522
rect -2709 488 -2693 522
rect -2635 488 -2619 522
rect -2561 488 -2545 522
rect -2487 488 -2471 522
rect -2413 488 -2397 522
rect -2339 488 -2323 522
rect -2265 488 -2249 522
rect -2191 488 -2175 522
rect -2117 488 -2101 522
rect -2043 488 -2027 522
rect -1969 488 -1953 522
rect -1895 488 -1879 522
rect -1821 488 -1805 522
rect -1747 488 -1731 522
rect -1673 488 -1657 522
rect -1599 488 -1583 522
rect -1525 488 -1509 522
rect -1451 488 -1435 522
rect -1377 488 -1361 522
rect -1303 488 -1287 522
rect -1229 488 -1213 522
rect -1155 488 -1139 522
rect -1081 488 -1065 522
rect -1007 488 -991 522
rect -933 488 -917 522
rect -859 488 -843 522
rect -785 488 -769 522
rect -711 488 -695 522
rect -637 488 -621 522
rect -563 488 -547 522
rect -489 488 -473 522
rect -415 488 -399 522
rect -341 488 -325 522
rect -267 488 -251 522
rect -193 488 -177 522
rect -119 488 -103 522
rect -45 488 -29 522
rect 29 488 45 522
rect 103 488 119 522
rect 177 488 193 522
rect 251 488 267 522
rect 325 488 341 522
rect 399 488 415 522
rect 473 488 489 522
rect 547 488 563 522
rect 621 488 637 522
rect 695 488 711 522
rect 769 488 785 522
rect 843 488 859 522
rect 917 488 933 522
rect 991 488 1007 522
rect 1065 488 1081 522
rect 1139 488 1155 522
rect 1213 488 1229 522
rect 1287 488 1303 522
rect 1361 488 1377 522
rect 1435 488 1451 522
rect 1509 488 1525 522
rect 1583 488 1599 522
rect 1657 488 1673 522
rect 1731 488 1747 522
rect 1805 488 1821 522
rect 1879 488 1895 522
rect 1953 488 1969 522
rect 2027 488 2043 522
rect 2101 488 2117 522
rect 2175 488 2191 522
rect 2249 488 2265 522
rect 2323 488 2339 522
rect 2397 488 2413 522
rect 2471 488 2487 522
rect 2545 488 2561 522
rect 2619 488 2635 522
rect 2693 488 2709 522
rect 2767 488 2783 522
rect 2841 488 2857 522
rect 2915 488 2931 522
rect 2989 488 3005 522
rect 3063 488 3079 522
rect 3137 488 3153 522
rect 3211 488 3227 522
rect 3285 488 3301 522
rect 3359 488 3375 522
rect 3433 488 3449 522
rect 3507 488 3523 522
rect 3581 488 3597 522
rect 3655 488 3671 522
rect -3717 438 -3683 454
rect -3717 -454 -3683 -438
rect -3569 438 -3535 454
rect -3569 -454 -3535 -438
rect -3421 438 -3387 454
rect -3421 -454 -3387 -438
rect -3273 438 -3239 454
rect -3273 -454 -3239 -438
rect -3125 438 -3091 454
rect -3125 -454 -3091 -438
rect -2977 438 -2943 454
rect -2977 -454 -2943 -438
rect -2829 438 -2795 454
rect -2829 -454 -2795 -438
rect -2681 438 -2647 454
rect -2681 -454 -2647 -438
rect -2533 438 -2499 454
rect -2533 -454 -2499 -438
rect -2385 438 -2351 454
rect -2385 -454 -2351 -438
rect -2237 438 -2203 454
rect -2237 -454 -2203 -438
rect -2089 438 -2055 454
rect -2089 -454 -2055 -438
rect -1941 438 -1907 454
rect -1941 -454 -1907 -438
rect -1793 438 -1759 454
rect -1793 -454 -1759 -438
rect -1645 438 -1611 454
rect -1645 -454 -1611 -438
rect -1497 438 -1463 454
rect -1497 -454 -1463 -438
rect -1349 438 -1315 454
rect -1349 -454 -1315 -438
rect -1201 438 -1167 454
rect -1201 -454 -1167 -438
rect -1053 438 -1019 454
rect -1053 -454 -1019 -438
rect -905 438 -871 454
rect -905 -454 -871 -438
rect -757 438 -723 454
rect -757 -454 -723 -438
rect -609 438 -575 454
rect -609 -454 -575 -438
rect -461 438 -427 454
rect -461 -454 -427 -438
rect -313 438 -279 454
rect -313 -454 -279 -438
rect -165 438 -131 454
rect -165 -454 -131 -438
rect -17 438 17 454
rect -17 -454 17 -438
rect 131 438 165 454
rect 131 -454 165 -438
rect 279 438 313 454
rect 279 -454 313 -438
rect 427 438 461 454
rect 427 -454 461 -438
rect 575 438 609 454
rect 575 -454 609 -438
rect 723 438 757 454
rect 723 -454 757 -438
rect 871 438 905 454
rect 871 -454 905 -438
rect 1019 438 1053 454
rect 1019 -454 1053 -438
rect 1167 438 1201 454
rect 1167 -454 1201 -438
rect 1315 438 1349 454
rect 1315 -454 1349 -438
rect 1463 438 1497 454
rect 1463 -454 1497 -438
rect 1611 438 1645 454
rect 1611 -454 1645 -438
rect 1759 438 1793 454
rect 1759 -454 1793 -438
rect 1907 438 1941 454
rect 1907 -454 1941 -438
rect 2055 438 2089 454
rect 2055 -454 2089 -438
rect 2203 438 2237 454
rect 2203 -454 2237 -438
rect 2351 438 2385 454
rect 2351 -454 2385 -438
rect 2499 438 2533 454
rect 2499 -454 2533 -438
rect 2647 438 2681 454
rect 2647 -454 2681 -438
rect 2795 438 2829 454
rect 2795 -454 2829 -438
rect 2943 438 2977 454
rect 2943 -454 2977 -438
rect 3091 438 3125 454
rect 3091 -454 3125 -438
rect 3239 438 3273 454
rect 3239 -454 3273 -438
rect 3387 438 3421 454
rect 3387 -454 3421 -438
rect 3535 438 3569 454
rect 3535 -454 3569 -438
rect 3683 438 3717 454
rect 3683 -454 3717 -438
rect -3671 -522 -3655 -488
rect -3597 -522 -3581 -488
rect -3523 -522 -3507 -488
rect -3449 -522 -3433 -488
rect -3375 -522 -3359 -488
rect -3301 -522 -3285 -488
rect -3227 -522 -3211 -488
rect -3153 -522 -3137 -488
rect -3079 -522 -3063 -488
rect -3005 -522 -2989 -488
rect -2931 -522 -2915 -488
rect -2857 -522 -2841 -488
rect -2783 -522 -2767 -488
rect -2709 -522 -2693 -488
rect -2635 -522 -2619 -488
rect -2561 -522 -2545 -488
rect -2487 -522 -2471 -488
rect -2413 -522 -2397 -488
rect -2339 -522 -2323 -488
rect -2265 -522 -2249 -488
rect -2191 -522 -2175 -488
rect -2117 -522 -2101 -488
rect -2043 -522 -2027 -488
rect -1969 -522 -1953 -488
rect -1895 -522 -1879 -488
rect -1821 -522 -1805 -488
rect -1747 -522 -1731 -488
rect -1673 -522 -1657 -488
rect -1599 -522 -1583 -488
rect -1525 -522 -1509 -488
rect -1451 -522 -1435 -488
rect -1377 -522 -1361 -488
rect -1303 -522 -1287 -488
rect -1229 -522 -1213 -488
rect -1155 -522 -1139 -488
rect -1081 -522 -1065 -488
rect -1007 -522 -991 -488
rect -933 -522 -917 -488
rect -859 -522 -843 -488
rect -785 -522 -769 -488
rect -711 -522 -695 -488
rect -637 -522 -621 -488
rect -563 -522 -547 -488
rect -489 -522 -473 -488
rect -415 -522 -399 -488
rect -341 -522 -325 -488
rect -267 -522 -251 -488
rect -193 -522 -177 -488
rect -119 -522 -103 -488
rect -45 -522 -29 -488
rect 29 -522 45 -488
rect 103 -522 119 -488
rect 177 -522 193 -488
rect 251 -522 267 -488
rect 325 -522 341 -488
rect 399 -522 415 -488
rect 473 -522 489 -488
rect 547 -522 563 -488
rect 621 -522 637 -488
rect 695 -522 711 -488
rect 769 -522 785 -488
rect 843 -522 859 -488
rect 917 -522 933 -488
rect 991 -522 1007 -488
rect 1065 -522 1081 -488
rect 1139 -522 1155 -488
rect 1213 -522 1229 -488
rect 1287 -522 1303 -488
rect 1361 -522 1377 -488
rect 1435 -522 1451 -488
rect 1509 -522 1525 -488
rect 1583 -522 1599 -488
rect 1657 -522 1673 -488
rect 1731 -522 1747 -488
rect 1805 -522 1821 -488
rect 1879 -522 1895 -488
rect 1953 -522 1969 -488
rect 2027 -522 2043 -488
rect 2101 -522 2117 -488
rect 2175 -522 2191 -488
rect 2249 -522 2265 -488
rect 2323 -522 2339 -488
rect 2397 -522 2413 -488
rect 2471 -522 2487 -488
rect 2545 -522 2561 -488
rect 2619 -522 2635 -488
rect 2693 -522 2709 -488
rect 2767 -522 2783 -488
rect 2841 -522 2857 -488
rect 2915 -522 2931 -488
rect 2989 -522 3005 -488
rect 3063 -522 3079 -488
rect 3137 -522 3153 -488
rect 3211 -522 3227 -488
rect 3285 -522 3301 -488
rect 3359 -522 3375 -488
rect 3433 -522 3449 -488
rect 3507 -522 3523 -488
rect 3581 -522 3597 -488
rect 3655 -522 3671 -488
rect -3671 -630 -3655 -596
rect -3597 -630 -3581 -596
rect -3523 -630 -3507 -596
rect -3449 -630 -3433 -596
rect -3375 -630 -3359 -596
rect -3301 -630 -3285 -596
rect -3227 -630 -3211 -596
rect -3153 -630 -3137 -596
rect -3079 -630 -3063 -596
rect -3005 -630 -2989 -596
rect -2931 -630 -2915 -596
rect -2857 -630 -2841 -596
rect -2783 -630 -2767 -596
rect -2709 -630 -2693 -596
rect -2635 -630 -2619 -596
rect -2561 -630 -2545 -596
rect -2487 -630 -2471 -596
rect -2413 -630 -2397 -596
rect -2339 -630 -2323 -596
rect -2265 -630 -2249 -596
rect -2191 -630 -2175 -596
rect -2117 -630 -2101 -596
rect -2043 -630 -2027 -596
rect -1969 -630 -1953 -596
rect -1895 -630 -1879 -596
rect -1821 -630 -1805 -596
rect -1747 -630 -1731 -596
rect -1673 -630 -1657 -596
rect -1599 -630 -1583 -596
rect -1525 -630 -1509 -596
rect -1451 -630 -1435 -596
rect -1377 -630 -1361 -596
rect -1303 -630 -1287 -596
rect -1229 -630 -1213 -596
rect -1155 -630 -1139 -596
rect -1081 -630 -1065 -596
rect -1007 -630 -991 -596
rect -933 -630 -917 -596
rect -859 -630 -843 -596
rect -785 -630 -769 -596
rect -711 -630 -695 -596
rect -637 -630 -621 -596
rect -563 -630 -547 -596
rect -489 -630 -473 -596
rect -415 -630 -399 -596
rect -341 -630 -325 -596
rect -267 -630 -251 -596
rect -193 -630 -177 -596
rect -119 -630 -103 -596
rect -45 -630 -29 -596
rect 29 -630 45 -596
rect 103 -630 119 -596
rect 177 -630 193 -596
rect 251 -630 267 -596
rect 325 -630 341 -596
rect 399 -630 415 -596
rect 473 -630 489 -596
rect 547 -630 563 -596
rect 621 -630 637 -596
rect 695 -630 711 -596
rect 769 -630 785 -596
rect 843 -630 859 -596
rect 917 -630 933 -596
rect 991 -630 1007 -596
rect 1065 -630 1081 -596
rect 1139 -630 1155 -596
rect 1213 -630 1229 -596
rect 1287 -630 1303 -596
rect 1361 -630 1377 -596
rect 1435 -630 1451 -596
rect 1509 -630 1525 -596
rect 1583 -630 1599 -596
rect 1657 -630 1673 -596
rect 1731 -630 1747 -596
rect 1805 -630 1821 -596
rect 1879 -630 1895 -596
rect 1953 -630 1969 -596
rect 2027 -630 2043 -596
rect 2101 -630 2117 -596
rect 2175 -630 2191 -596
rect 2249 -630 2265 -596
rect 2323 -630 2339 -596
rect 2397 -630 2413 -596
rect 2471 -630 2487 -596
rect 2545 -630 2561 -596
rect 2619 -630 2635 -596
rect 2693 -630 2709 -596
rect 2767 -630 2783 -596
rect 2841 -630 2857 -596
rect 2915 -630 2931 -596
rect 2989 -630 3005 -596
rect 3063 -630 3079 -596
rect 3137 -630 3153 -596
rect 3211 -630 3227 -596
rect 3285 -630 3301 -596
rect 3359 -630 3375 -596
rect 3433 -630 3449 -596
rect 3507 -630 3523 -596
rect 3581 -630 3597 -596
rect 3655 -630 3671 -596
rect -3717 -680 -3683 -664
rect -3717 -1572 -3683 -1556
rect -3569 -680 -3535 -664
rect -3569 -1572 -3535 -1556
rect -3421 -680 -3387 -664
rect -3421 -1572 -3387 -1556
rect -3273 -680 -3239 -664
rect -3273 -1572 -3239 -1556
rect -3125 -680 -3091 -664
rect -3125 -1572 -3091 -1556
rect -2977 -680 -2943 -664
rect -2977 -1572 -2943 -1556
rect -2829 -680 -2795 -664
rect -2829 -1572 -2795 -1556
rect -2681 -680 -2647 -664
rect -2681 -1572 -2647 -1556
rect -2533 -680 -2499 -664
rect -2533 -1572 -2499 -1556
rect -2385 -680 -2351 -664
rect -2385 -1572 -2351 -1556
rect -2237 -680 -2203 -664
rect -2237 -1572 -2203 -1556
rect -2089 -680 -2055 -664
rect -2089 -1572 -2055 -1556
rect -1941 -680 -1907 -664
rect -1941 -1572 -1907 -1556
rect -1793 -680 -1759 -664
rect -1793 -1572 -1759 -1556
rect -1645 -680 -1611 -664
rect -1645 -1572 -1611 -1556
rect -1497 -680 -1463 -664
rect -1497 -1572 -1463 -1556
rect -1349 -680 -1315 -664
rect -1349 -1572 -1315 -1556
rect -1201 -680 -1167 -664
rect -1201 -1572 -1167 -1556
rect -1053 -680 -1019 -664
rect -1053 -1572 -1019 -1556
rect -905 -680 -871 -664
rect -905 -1572 -871 -1556
rect -757 -680 -723 -664
rect -757 -1572 -723 -1556
rect -609 -680 -575 -664
rect -609 -1572 -575 -1556
rect -461 -680 -427 -664
rect -461 -1572 -427 -1556
rect -313 -680 -279 -664
rect -313 -1572 -279 -1556
rect -165 -680 -131 -664
rect -165 -1572 -131 -1556
rect -17 -680 17 -664
rect -17 -1572 17 -1556
rect 131 -680 165 -664
rect 131 -1572 165 -1556
rect 279 -680 313 -664
rect 279 -1572 313 -1556
rect 427 -680 461 -664
rect 427 -1572 461 -1556
rect 575 -680 609 -664
rect 575 -1572 609 -1556
rect 723 -680 757 -664
rect 723 -1572 757 -1556
rect 871 -680 905 -664
rect 871 -1572 905 -1556
rect 1019 -680 1053 -664
rect 1019 -1572 1053 -1556
rect 1167 -680 1201 -664
rect 1167 -1572 1201 -1556
rect 1315 -680 1349 -664
rect 1315 -1572 1349 -1556
rect 1463 -680 1497 -664
rect 1463 -1572 1497 -1556
rect 1611 -680 1645 -664
rect 1611 -1572 1645 -1556
rect 1759 -680 1793 -664
rect 1759 -1572 1793 -1556
rect 1907 -680 1941 -664
rect 1907 -1572 1941 -1556
rect 2055 -680 2089 -664
rect 2055 -1572 2089 -1556
rect 2203 -680 2237 -664
rect 2203 -1572 2237 -1556
rect 2351 -680 2385 -664
rect 2351 -1572 2385 -1556
rect 2499 -680 2533 -664
rect 2499 -1572 2533 -1556
rect 2647 -680 2681 -664
rect 2647 -1572 2681 -1556
rect 2795 -680 2829 -664
rect 2795 -1572 2829 -1556
rect 2943 -680 2977 -664
rect 2943 -1572 2977 -1556
rect 3091 -680 3125 -664
rect 3091 -1572 3125 -1556
rect 3239 -680 3273 -664
rect 3239 -1572 3273 -1556
rect 3387 -680 3421 -664
rect 3387 -1572 3421 -1556
rect 3535 -680 3569 -664
rect 3535 -1572 3569 -1556
rect 3683 -680 3717 -664
rect 3683 -1572 3717 -1556
rect -3671 -1640 -3655 -1606
rect -3597 -1640 -3581 -1606
rect -3523 -1640 -3507 -1606
rect -3449 -1640 -3433 -1606
rect -3375 -1640 -3359 -1606
rect -3301 -1640 -3285 -1606
rect -3227 -1640 -3211 -1606
rect -3153 -1640 -3137 -1606
rect -3079 -1640 -3063 -1606
rect -3005 -1640 -2989 -1606
rect -2931 -1640 -2915 -1606
rect -2857 -1640 -2841 -1606
rect -2783 -1640 -2767 -1606
rect -2709 -1640 -2693 -1606
rect -2635 -1640 -2619 -1606
rect -2561 -1640 -2545 -1606
rect -2487 -1640 -2471 -1606
rect -2413 -1640 -2397 -1606
rect -2339 -1640 -2323 -1606
rect -2265 -1640 -2249 -1606
rect -2191 -1640 -2175 -1606
rect -2117 -1640 -2101 -1606
rect -2043 -1640 -2027 -1606
rect -1969 -1640 -1953 -1606
rect -1895 -1640 -1879 -1606
rect -1821 -1640 -1805 -1606
rect -1747 -1640 -1731 -1606
rect -1673 -1640 -1657 -1606
rect -1599 -1640 -1583 -1606
rect -1525 -1640 -1509 -1606
rect -1451 -1640 -1435 -1606
rect -1377 -1640 -1361 -1606
rect -1303 -1640 -1287 -1606
rect -1229 -1640 -1213 -1606
rect -1155 -1640 -1139 -1606
rect -1081 -1640 -1065 -1606
rect -1007 -1640 -991 -1606
rect -933 -1640 -917 -1606
rect -859 -1640 -843 -1606
rect -785 -1640 -769 -1606
rect -711 -1640 -695 -1606
rect -637 -1640 -621 -1606
rect -563 -1640 -547 -1606
rect -489 -1640 -473 -1606
rect -415 -1640 -399 -1606
rect -341 -1640 -325 -1606
rect -267 -1640 -251 -1606
rect -193 -1640 -177 -1606
rect -119 -1640 -103 -1606
rect -45 -1640 -29 -1606
rect 29 -1640 45 -1606
rect 103 -1640 119 -1606
rect 177 -1640 193 -1606
rect 251 -1640 267 -1606
rect 325 -1640 341 -1606
rect 399 -1640 415 -1606
rect 473 -1640 489 -1606
rect 547 -1640 563 -1606
rect 621 -1640 637 -1606
rect 695 -1640 711 -1606
rect 769 -1640 785 -1606
rect 843 -1640 859 -1606
rect 917 -1640 933 -1606
rect 991 -1640 1007 -1606
rect 1065 -1640 1081 -1606
rect 1139 -1640 1155 -1606
rect 1213 -1640 1229 -1606
rect 1287 -1640 1303 -1606
rect 1361 -1640 1377 -1606
rect 1435 -1640 1451 -1606
rect 1509 -1640 1525 -1606
rect 1583 -1640 1599 -1606
rect 1657 -1640 1673 -1606
rect 1731 -1640 1747 -1606
rect 1805 -1640 1821 -1606
rect 1879 -1640 1895 -1606
rect 1953 -1640 1969 -1606
rect 2027 -1640 2043 -1606
rect 2101 -1640 2117 -1606
rect 2175 -1640 2191 -1606
rect 2249 -1640 2265 -1606
rect 2323 -1640 2339 -1606
rect 2397 -1640 2413 -1606
rect 2471 -1640 2487 -1606
rect 2545 -1640 2561 -1606
rect 2619 -1640 2635 -1606
rect 2693 -1640 2709 -1606
rect 2767 -1640 2783 -1606
rect 2841 -1640 2857 -1606
rect 2915 -1640 2931 -1606
rect 2989 -1640 3005 -1606
rect 3063 -1640 3079 -1606
rect 3137 -1640 3153 -1606
rect 3211 -1640 3227 -1606
rect 3285 -1640 3301 -1606
rect 3359 -1640 3375 -1606
rect 3433 -1640 3449 -1606
rect 3507 -1640 3523 -1606
rect 3581 -1640 3597 -1606
rect 3655 -1640 3671 -1606
rect -3831 -1708 -3797 -1646
rect 3797 -1708 3831 -1646
rect -3831 -1742 -3735 -1708
rect 3735 -1742 3831 -1708
<< viali >>
rect -3655 1606 -3597 1640
rect -3507 1606 -3449 1640
rect -3359 1606 -3301 1640
rect -3211 1606 -3153 1640
rect -3063 1606 -3005 1640
rect -2915 1606 -2857 1640
rect -2767 1606 -2709 1640
rect -2619 1606 -2561 1640
rect -2471 1606 -2413 1640
rect -2323 1606 -2265 1640
rect -2175 1606 -2117 1640
rect -2027 1606 -1969 1640
rect -1879 1606 -1821 1640
rect -1731 1606 -1673 1640
rect -1583 1606 -1525 1640
rect -1435 1606 -1377 1640
rect -1287 1606 -1229 1640
rect -1139 1606 -1081 1640
rect -991 1606 -933 1640
rect -843 1606 -785 1640
rect -695 1606 -637 1640
rect -547 1606 -489 1640
rect -399 1606 -341 1640
rect -251 1606 -193 1640
rect -103 1606 -45 1640
rect 45 1606 103 1640
rect 193 1606 251 1640
rect 341 1606 399 1640
rect 489 1606 547 1640
rect 637 1606 695 1640
rect 785 1606 843 1640
rect 933 1606 991 1640
rect 1081 1606 1139 1640
rect 1229 1606 1287 1640
rect 1377 1606 1435 1640
rect 1525 1606 1583 1640
rect 1673 1606 1731 1640
rect 1821 1606 1879 1640
rect 1969 1606 2027 1640
rect 2117 1606 2175 1640
rect 2265 1606 2323 1640
rect 2413 1606 2471 1640
rect 2561 1606 2619 1640
rect 2709 1606 2767 1640
rect 2857 1606 2915 1640
rect 3005 1606 3063 1640
rect 3153 1606 3211 1640
rect 3301 1606 3359 1640
rect 3449 1606 3507 1640
rect 3597 1606 3655 1640
rect -3717 680 -3683 1556
rect -3569 680 -3535 1556
rect -3421 680 -3387 1556
rect -3273 680 -3239 1556
rect -3125 680 -3091 1556
rect -2977 680 -2943 1556
rect -2829 680 -2795 1556
rect -2681 680 -2647 1556
rect -2533 680 -2499 1556
rect -2385 680 -2351 1556
rect -2237 680 -2203 1556
rect -2089 680 -2055 1556
rect -1941 680 -1907 1556
rect -1793 680 -1759 1556
rect -1645 680 -1611 1556
rect -1497 680 -1463 1556
rect -1349 680 -1315 1556
rect -1201 680 -1167 1556
rect -1053 680 -1019 1556
rect -905 680 -871 1556
rect -757 680 -723 1556
rect -609 680 -575 1556
rect -461 680 -427 1556
rect -313 680 -279 1556
rect -165 680 -131 1556
rect -17 680 17 1556
rect 131 680 165 1556
rect 279 680 313 1556
rect 427 680 461 1556
rect 575 680 609 1556
rect 723 680 757 1556
rect 871 680 905 1556
rect 1019 680 1053 1556
rect 1167 680 1201 1556
rect 1315 680 1349 1556
rect 1463 680 1497 1556
rect 1611 680 1645 1556
rect 1759 680 1793 1556
rect 1907 680 1941 1556
rect 2055 680 2089 1556
rect 2203 680 2237 1556
rect 2351 680 2385 1556
rect 2499 680 2533 1556
rect 2647 680 2681 1556
rect 2795 680 2829 1556
rect 2943 680 2977 1556
rect 3091 680 3125 1556
rect 3239 680 3273 1556
rect 3387 680 3421 1556
rect 3535 680 3569 1556
rect 3683 680 3717 1556
rect -3655 596 -3597 630
rect -3507 596 -3449 630
rect -3359 596 -3301 630
rect -3211 596 -3153 630
rect -3063 596 -3005 630
rect -2915 596 -2857 630
rect -2767 596 -2709 630
rect -2619 596 -2561 630
rect -2471 596 -2413 630
rect -2323 596 -2265 630
rect -2175 596 -2117 630
rect -2027 596 -1969 630
rect -1879 596 -1821 630
rect -1731 596 -1673 630
rect -1583 596 -1525 630
rect -1435 596 -1377 630
rect -1287 596 -1229 630
rect -1139 596 -1081 630
rect -991 596 -933 630
rect -843 596 -785 630
rect -695 596 -637 630
rect -547 596 -489 630
rect -399 596 -341 630
rect -251 596 -193 630
rect -103 596 -45 630
rect 45 596 103 630
rect 193 596 251 630
rect 341 596 399 630
rect 489 596 547 630
rect 637 596 695 630
rect 785 596 843 630
rect 933 596 991 630
rect 1081 596 1139 630
rect 1229 596 1287 630
rect 1377 596 1435 630
rect 1525 596 1583 630
rect 1673 596 1731 630
rect 1821 596 1879 630
rect 1969 596 2027 630
rect 2117 596 2175 630
rect 2265 596 2323 630
rect 2413 596 2471 630
rect 2561 596 2619 630
rect 2709 596 2767 630
rect 2857 596 2915 630
rect 3005 596 3063 630
rect 3153 596 3211 630
rect 3301 596 3359 630
rect 3449 596 3507 630
rect 3597 596 3655 630
rect -3655 488 -3597 522
rect -3507 488 -3449 522
rect -3359 488 -3301 522
rect -3211 488 -3153 522
rect -3063 488 -3005 522
rect -2915 488 -2857 522
rect -2767 488 -2709 522
rect -2619 488 -2561 522
rect -2471 488 -2413 522
rect -2323 488 -2265 522
rect -2175 488 -2117 522
rect -2027 488 -1969 522
rect -1879 488 -1821 522
rect -1731 488 -1673 522
rect -1583 488 -1525 522
rect -1435 488 -1377 522
rect -1287 488 -1229 522
rect -1139 488 -1081 522
rect -991 488 -933 522
rect -843 488 -785 522
rect -695 488 -637 522
rect -547 488 -489 522
rect -399 488 -341 522
rect -251 488 -193 522
rect -103 488 -45 522
rect 45 488 103 522
rect 193 488 251 522
rect 341 488 399 522
rect 489 488 547 522
rect 637 488 695 522
rect 785 488 843 522
rect 933 488 991 522
rect 1081 488 1139 522
rect 1229 488 1287 522
rect 1377 488 1435 522
rect 1525 488 1583 522
rect 1673 488 1731 522
rect 1821 488 1879 522
rect 1969 488 2027 522
rect 2117 488 2175 522
rect 2265 488 2323 522
rect 2413 488 2471 522
rect 2561 488 2619 522
rect 2709 488 2767 522
rect 2857 488 2915 522
rect 3005 488 3063 522
rect 3153 488 3211 522
rect 3301 488 3359 522
rect 3449 488 3507 522
rect 3597 488 3655 522
rect -3717 -438 -3683 438
rect -3569 -438 -3535 438
rect -3421 -438 -3387 438
rect -3273 -438 -3239 438
rect -3125 -438 -3091 438
rect -2977 -438 -2943 438
rect -2829 -438 -2795 438
rect -2681 -438 -2647 438
rect -2533 -438 -2499 438
rect -2385 -438 -2351 438
rect -2237 -438 -2203 438
rect -2089 -438 -2055 438
rect -1941 -438 -1907 438
rect -1793 -438 -1759 438
rect -1645 -438 -1611 438
rect -1497 -438 -1463 438
rect -1349 -438 -1315 438
rect -1201 -438 -1167 438
rect -1053 -438 -1019 438
rect -905 -438 -871 438
rect -757 -438 -723 438
rect -609 -438 -575 438
rect -461 -438 -427 438
rect -313 -438 -279 438
rect -165 -438 -131 438
rect -17 -438 17 438
rect 131 -438 165 438
rect 279 -438 313 438
rect 427 -438 461 438
rect 575 -438 609 438
rect 723 -438 757 438
rect 871 -438 905 438
rect 1019 -438 1053 438
rect 1167 -438 1201 438
rect 1315 -438 1349 438
rect 1463 -438 1497 438
rect 1611 -438 1645 438
rect 1759 -438 1793 438
rect 1907 -438 1941 438
rect 2055 -438 2089 438
rect 2203 -438 2237 438
rect 2351 -438 2385 438
rect 2499 -438 2533 438
rect 2647 -438 2681 438
rect 2795 -438 2829 438
rect 2943 -438 2977 438
rect 3091 -438 3125 438
rect 3239 -438 3273 438
rect 3387 -438 3421 438
rect 3535 -438 3569 438
rect 3683 -438 3717 438
rect -3655 -522 -3597 -488
rect -3507 -522 -3449 -488
rect -3359 -522 -3301 -488
rect -3211 -522 -3153 -488
rect -3063 -522 -3005 -488
rect -2915 -522 -2857 -488
rect -2767 -522 -2709 -488
rect -2619 -522 -2561 -488
rect -2471 -522 -2413 -488
rect -2323 -522 -2265 -488
rect -2175 -522 -2117 -488
rect -2027 -522 -1969 -488
rect -1879 -522 -1821 -488
rect -1731 -522 -1673 -488
rect -1583 -522 -1525 -488
rect -1435 -522 -1377 -488
rect -1287 -522 -1229 -488
rect -1139 -522 -1081 -488
rect -991 -522 -933 -488
rect -843 -522 -785 -488
rect -695 -522 -637 -488
rect -547 -522 -489 -488
rect -399 -522 -341 -488
rect -251 -522 -193 -488
rect -103 -522 -45 -488
rect 45 -522 103 -488
rect 193 -522 251 -488
rect 341 -522 399 -488
rect 489 -522 547 -488
rect 637 -522 695 -488
rect 785 -522 843 -488
rect 933 -522 991 -488
rect 1081 -522 1139 -488
rect 1229 -522 1287 -488
rect 1377 -522 1435 -488
rect 1525 -522 1583 -488
rect 1673 -522 1731 -488
rect 1821 -522 1879 -488
rect 1969 -522 2027 -488
rect 2117 -522 2175 -488
rect 2265 -522 2323 -488
rect 2413 -522 2471 -488
rect 2561 -522 2619 -488
rect 2709 -522 2767 -488
rect 2857 -522 2915 -488
rect 3005 -522 3063 -488
rect 3153 -522 3211 -488
rect 3301 -522 3359 -488
rect 3449 -522 3507 -488
rect 3597 -522 3655 -488
rect -3655 -630 -3597 -596
rect -3507 -630 -3449 -596
rect -3359 -630 -3301 -596
rect -3211 -630 -3153 -596
rect -3063 -630 -3005 -596
rect -2915 -630 -2857 -596
rect -2767 -630 -2709 -596
rect -2619 -630 -2561 -596
rect -2471 -630 -2413 -596
rect -2323 -630 -2265 -596
rect -2175 -630 -2117 -596
rect -2027 -630 -1969 -596
rect -1879 -630 -1821 -596
rect -1731 -630 -1673 -596
rect -1583 -630 -1525 -596
rect -1435 -630 -1377 -596
rect -1287 -630 -1229 -596
rect -1139 -630 -1081 -596
rect -991 -630 -933 -596
rect -843 -630 -785 -596
rect -695 -630 -637 -596
rect -547 -630 -489 -596
rect -399 -630 -341 -596
rect -251 -630 -193 -596
rect -103 -630 -45 -596
rect 45 -630 103 -596
rect 193 -630 251 -596
rect 341 -630 399 -596
rect 489 -630 547 -596
rect 637 -630 695 -596
rect 785 -630 843 -596
rect 933 -630 991 -596
rect 1081 -630 1139 -596
rect 1229 -630 1287 -596
rect 1377 -630 1435 -596
rect 1525 -630 1583 -596
rect 1673 -630 1731 -596
rect 1821 -630 1879 -596
rect 1969 -630 2027 -596
rect 2117 -630 2175 -596
rect 2265 -630 2323 -596
rect 2413 -630 2471 -596
rect 2561 -630 2619 -596
rect 2709 -630 2767 -596
rect 2857 -630 2915 -596
rect 3005 -630 3063 -596
rect 3153 -630 3211 -596
rect 3301 -630 3359 -596
rect 3449 -630 3507 -596
rect 3597 -630 3655 -596
rect -3717 -1556 -3683 -680
rect -3569 -1556 -3535 -680
rect -3421 -1556 -3387 -680
rect -3273 -1556 -3239 -680
rect -3125 -1556 -3091 -680
rect -2977 -1556 -2943 -680
rect -2829 -1556 -2795 -680
rect -2681 -1556 -2647 -680
rect -2533 -1556 -2499 -680
rect -2385 -1556 -2351 -680
rect -2237 -1556 -2203 -680
rect -2089 -1556 -2055 -680
rect -1941 -1556 -1907 -680
rect -1793 -1556 -1759 -680
rect -1645 -1556 -1611 -680
rect -1497 -1556 -1463 -680
rect -1349 -1556 -1315 -680
rect -1201 -1556 -1167 -680
rect -1053 -1556 -1019 -680
rect -905 -1556 -871 -680
rect -757 -1556 -723 -680
rect -609 -1556 -575 -680
rect -461 -1556 -427 -680
rect -313 -1556 -279 -680
rect -165 -1556 -131 -680
rect -17 -1556 17 -680
rect 131 -1556 165 -680
rect 279 -1556 313 -680
rect 427 -1556 461 -680
rect 575 -1556 609 -680
rect 723 -1556 757 -680
rect 871 -1556 905 -680
rect 1019 -1556 1053 -680
rect 1167 -1556 1201 -680
rect 1315 -1556 1349 -680
rect 1463 -1556 1497 -680
rect 1611 -1556 1645 -680
rect 1759 -1556 1793 -680
rect 1907 -1556 1941 -680
rect 2055 -1556 2089 -680
rect 2203 -1556 2237 -680
rect 2351 -1556 2385 -680
rect 2499 -1556 2533 -680
rect 2647 -1556 2681 -680
rect 2795 -1556 2829 -680
rect 2943 -1556 2977 -680
rect 3091 -1556 3125 -680
rect 3239 -1556 3273 -680
rect 3387 -1556 3421 -680
rect 3535 -1556 3569 -680
rect 3683 -1556 3717 -680
rect -3655 -1640 -3597 -1606
rect -3507 -1640 -3449 -1606
rect -3359 -1640 -3301 -1606
rect -3211 -1640 -3153 -1606
rect -3063 -1640 -3005 -1606
rect -2915 -1640 -2857 -1606
rect -2767 -1640 -2709 -1606
rect -2619 -1640 -2561 -1606
rect -2471 -1640 -2413 -1606
rect -2323 -1640 -2265 -1606
rect -2175 -1640 -2117 -1606
rect -2027 -1640 -1969 -1606
rect -1879 -1640 -1821 -1606
rect -1731 -1640 -1673 -1606
rect -1583 -1640 -1525 -1606
rect -1435 -1640 -1377 -1606
rect -1287 -1640 -1229 -1606
rect -1139 -1640 -1081 -1606
rect -991 -1640 -933 -1606
rect -843 -1640 -785 -1606
rect -695 -1640 -637 -1606
rect -547 -1640 -489 -1606
rect -399 -1640 -341 -1606
rect -251 -1640 -193 -1606
rect -103 -1640 -45 -1606
rect 45 -1640 103 -1606
rect 193 -1640 251 -1606
rect 341 -1640 399 -1606
rect 489 -1640 547 -1606
rect 637 -1640 695 -1606
rect 785 -1640 843 -1606
rect 933 -1640 991 -1606
rect 1081 -1640 1139 -1606
rect 1229 -1640 1287 -1606
rect 1377 -1640 1435 -1606
rect 1525 -1640 1583 -1606
rect 1673 -1640 1731 -1606
rect 1821 -1640 1879 -1606
rect 1969 -1640 2027 -1606
rect 2117 -1640 2175 -1606
rect 2265 -1640 2323 -1606
rect 2413 -1640 2471 -1606
rect 2561 -1640 2619 -1606
rect 2709 -1640 2767 -1606
rect 2857 -1640 2915 -1606
rect 3005 -1640 3063 -1606
rect 3153 -1640 3211 -1606
rect 3301 -1640 3359 -1606
rect 3449 -1640 3507 -1606
rect 3597 -1640 3655 -1606
<< metal1 >>
rect -3667 1640 -3585 1646
rect -3667 1606 -3655 1640
rect -3597 1606 -3585 1640
rect -3667 1600 -3585 1606
rect -3519 1640 -3437 1646
rect -3519 1606 -3507 1640
rect -3449 1606 -3437 1640
rect -3519 1600 -3437 1606
rect -3371 1640 -3289 1646
rect -3371 1606 -3359 1640
rect -3301 1606 -3289 1640
rect -3371 1600 -3289 1606
rect -3223 1640 -3141 1646
rect -3223 1606 -3211 1640
rect -3153 1606 -3141 1640
rect -3223 1600 -3141 1606
rect -3075 1640 -2993 1646
rect -3075 1606 -3063 1640
rect -3005 1606 -2993 1640
rect -3075 1600 -2993 1606
rect -2927 1640 -2845 1646
rect -2927 1606 -2915 1640
rect -2857 1606 -2845 1640
rect -2927 1600 -2845 1606
rect -2779 1640 -2697 1646
rect -2779 1606 -2767 1640
rect -2709 1606 -2697 1640
rect -2779 1600 -2697 1606
rect -2631 1640 -2549 1646
rect -2631 1606 -2619 1640
rect -2561 1606 -2549 1640
rect -2631 1600 -2549 1606
rect -2483 1640 -2401 1646
rect -2483 1606 -2471 1640
rect -2413 1606 -2401 1640
rect -2483 1600 -2401 1606
rect -2335 1640 -2253 1646
rect -2335 1606 -2323 1640
rect -2265 1606 -2253 1640
rect -2335 1600 -2253 1606
rect -2187 1640 -2105 1646
rect -2187 1606 -2175 1640
rect -2117 1606 -2105 1640
rect -2187 1600 -2105 1606
rect -2039 1640 -1957 1646
rect -2039 1606 -2027 1640
rect -1969 1606 -1957 1640
rect -2039 1600 -1957 1606
rect -1891 1640 -1809 1646
rect -1891 1606 -1879 1640
rect -1821 1606 -1809 1640
rect -1891 1600 -1809 1606
rect -1743 1640 -1661 1646
rect -1743 1606 -1731 1640
rect -1673 1606 -1661 1640
rect -1743 1600 -1661 1606
rect -1595 1640 -1513 1646
rect -1595 1606 -1583 1640
rect -1525 1606 -1513 1640
rect -1595 1600 -1513 1606
rect -1447 1640 -1365 1646
rect -1447 1606 -1435 1640
rect -1377 1606 -1365 1640
rect -1447 1600 -1365 1606
rect -1299 1640 -1217 1646
rect -1299 1606 -1287 1640
rect -1229 1606 -1217 1640
rect -1299 1600 -1217 1606
rect -1151 1640 -1069 1646
rect -1151 1606 -1139 1640
rect -1081 1606 -1069 1640
rect -1151 1600 -1069 1606
rect -1003 1640 -921 1646
rect -1003 1606 -991 1640
rect -933 1606 -921 1640
rect -1003 1600 -921 1606
rect -855 1640 -773 1646
rect -855 1606 -843 1640
rect -785 1606 -773 1640
rect -855 1600 -773 1606
rect -707 1640 -625 1646
rect -707 1606 -695 1640
rect -637 1606 -625 1640
rect -707 1600 -625 1606
rect -559 1640 -477 1646
rect -559 1606 -547 1640
rect -489 1606 -477 1640
rect -559 1600 -477 1606
rect -411 1640 -329 1646
rect -411 1606 -399 1640
rect -341 1606 -329 1640
rect -411 1600 -329 1606
rect -263 1640 -181 1646
rect -263 1606 -251 1640
rect -193 1606 -181 1640
rect -263 1600 -181 1606
rect -115 1640 -33 1646
rect -115 1606 -103 1640
rect -45 1606 -33 1640
rect -115 1600 -33 1606
rect 33 1640 115 1646
rect 33 1606 45 1640
rect 103 1606 115 1640
rect 33 1600 115 1606
rect 181 1640 263 1646
rect 181 1606 193 1640
rect 251 1606 263 1640
rect 181 1600 263 1606
rect 329 1640 411 1646
rect 329 1606 341 1640
rect 399 1606 411 1640
rect 329 1600 411 1606
rect 477 1640 559 1646
rect 477 1606 489 1640
rect 547 1606 559 1640
rect 477 1600 559 1606
rect 625 1640 707 1646
rect 625 1606 637 1640
rect 695 1606 707 1640
rect 625 1600 707 1606
rect 773 1640 855 1646
rect 773 1606 785 1640
rect 843 1606 855 1640
rect 773 1600 855 1606
rect 921 1640 1003 1646
rect 921 1606 933 1640
rect 991 1606 1003 1640
rect 921 1600 1003 1606
rect 1069 1640 1151 1646
rect 1069 1606 1081 1640
rect 1139 1606 1151 1640
rect 1069 1600 1151 1606
rect 1217 1640 1299 1646
rect 1217 1606 1229 1640
rect 1287 1606 1299 1640
rect 1217 1600 1299 1606
rect 1365 1640 1447 1646
rect 1365 1606 1377 1640
rect 1435 1606 1447 1640
rect 1365 1600 1447 1606
rect 1513 1640 1595 1646
rect 1513 1606 1525 1640
rect 1583 1606 1595 1640
rect 1513 1600 1595 1606
rect 1661 1640 1743 1646
rect 1661 1606 1673 1640
rect 1731 1606 1743 1640
rect 1661 1600 1743 1606
rect 1809 1640 1891 1646
rect 1809 1606 1821 1640
rect 1879 1606 1891 1640
rect 1809 1600 1891 1606
rect 1957 1640 2039 1646
rect 1957 1606 1969 1640
rect 2027 1606 2039 1640
rect 1957 1600 2039 1606
rect 2105 1640 2187 1646
rect 2105 1606 2117 1640
rect 2175 1606 2187 1640
rect 2105 1600 2187 1606
rect 2253 1640 2335 1646
rect 2253 1606 2265 1640
rect 2323 1606 2335 1640
rect 2253 1600 2335 1606
rect 2401 1640 2483 1646
rect 2401 1606 2413 1640
rect 2471 1606 2483 1640
rect 2401 1600 2483 1606
rect 2549 1640 2631 1646
rect 2549 1606 2561 1640
rect 2619 1606 2631 1640
rect 2549 1600 2631 1606
rect 2697 1640 2779 1646
rect 2697 1606 2709 1640
rect 2767 1606 2779 1640
rect 2697 1600 2779 1606
rect 2845 1640 2927 1646
rect 2845 1606 2857 1640
rect 2915 1606 2927 1640
rect 2845 1600 2927 1606
rect 2993 1640 3075 1646
rect 2993 1606 3005 1640
rect 3063 1606 3075 1640
rect 2993 1600 3075 1606
rect 3141 1640 3223 1646
rect 3141 1606 3153 1640
rect 3211 1606 3223 1640
rect 3141 1600 3223 1606
rect 3289 1640 3371 1646
rect 3289 1606 3301 1640
rect 3359 1606 3371 1640
rect 3289 1600 3371 1606
rect 3437 1640 3519 1646
rect 3437 1606 3449 1640
rect 3507 1606 3519 1640
rect 3437 1600 3519 1606
rect 3585 1640 3667 1646
rect 3585 1606 3597 1640
rect 3655 1606 3667 1640
rect 3585 1600 3667 1606
rect -3723 1556 -3677 1568
rect -3723 680 -3717 1556
rect -3683 680 -3677 1556
rect -3723 668 -3677 680
rect -3575 1556 -3529 1568
rect -3575 680 -3569 1556
rect -3535 680 -3529 1556
rect -3575 668 -3529 680
rect -3427 1556 -3381 1568
rect -3427 680 -3421 1556
rect -3387 680 -3381 1556
rect -3427 668 -3381 680
rect -3279 1556 -3233 1568
rect -3279 680 -3273 1556
rect -3239 680 -3233 1556
rect -3279 668 -3233 680
rect -3131 1556 -3085 1568
rect -3131 680 -3125 1556
rect -3091 680 -3085 1556
rect -3131 668 -3085 680
rect -2983 1556 -2937 1568
rect -2983 680 -2977 1556
rect -2943 680 -2937 1556
rect -2983 668 -2937 680
rect -2835 1556 -2789 1568
rect -2835 680 -2829 1556
rect -2795 680 -2789 1556
rect -2835 668 -2789 680
rect -2687 1556 -2641 1568
rect -2687 680 -2681 1556
rect -2647 680 -2641 1556
rect -2687 668 -2641 680
rect -2539 1556 -2493 1568
rect -2539 680 -2533 1556
rect -2499 680 -2493 1556
rect -2539 668 -2493 680
rect -2391 1556 -2345 1568
rect -2391 680 -2385 1556
rect -2351 680 -2345 1556
rect -2391 668 -2345 680
rect -2243 1556 -2197 1568
rect -2243 680 -2237 1556
rect -2203 680 -2197 1556
rect -2243 668 -2197 680
rect -2095 1556 -2049 1568
rect -2095 680 -2089 1556
rect -2055 680 -2049 1556
rect -2095 668 -2049 680
rect -1947 1556 -1901 1568
rect -1947 680 -1941 1556
rect -1907 680 -1901 1556
rect -1947 668 -1901 680
rect -1799 1556 -1753 1568
rect -1799 680 -1793 1556
rect -1759 680 -1753 1556
rect -1799 668 -1753 680
rect -1651 1556 -1605 1568
rect -1651 680 -1645 1556
rect -1611 680 -1605 1556
rect -1651 668 -1605 680
rect -1503 1556 -1457 1568
rect -1503 680 -1497 1556
rect -1463 680 -1457 1556
rect -1503 668 -1457 680
rect -1355 1556 -1309 1568
rect -1355 680 -1349 1556
rect -1315 680 -1309 1556
rect -1355 668 -1309 680
rect -1207 1556 -1161 1568
rect -1207 680 -1201 1556
rect -1167 680 -1161 1556
rect -1207 668 -1161 680
rect -1059 1556 -1013 1568
rect -1059 680 -1053 1556
rect -1019 680 -1013 1556
rect -1059 668 -1013 680
rect -911 1556 -865 1568
rect -911 680 -905 1556
rect -871 680 -865 1556
rect -911 668 -865 680
rect -763 1556 -717 1568
rect -763 680 -757 1556
rect -723 680 -717 1556
rect -763 668 -717 680
rect -615 1556 -569 1568
rect -615 680 -609 1556
rect -575 680 -569 1556
rect -615 668 -569 680
rect -467 1556 -421 1568
rect -467 680 -461 1556
rect -427 680 -421 1556
rect -467 668 -421 680
rect -319 1556 -273 1568
rect -319 680 -313 1556
rect -279 680 -273 1556
rect -319 668 -273 680
rect -171 1556 -125 1568
rect -171 680 -165 1556
rect -131 680 -125 1556
rect -171 668 -125 680
rect -23 1556 23 1568
rect -23 680 -17 1556
rect 17 680 23 1556
rect -23 668 23 680
rect 125 1556 171 1568
rect 125 680 131 1556
rect 165 680 171 1556
rect 125 668 171 680
rect 273 1556 319 1568
rect 273 680 279 1556
rect 313 680 319 1556
rect 273 668 319 680
rect 421 1556 467 1568
rect 421 680 427 1556
rect 461 680 467 1556
rect 421 668 467 680
rect 569 1556 615 1568
rect 569 680 575 1556
rect 609 680 615 1556
rect 569 668 615 680
rect 717 1556 763 1568
rect 717 680 723 1556
rect 757 680 763 1556
rect 717 668 763 680
rect 865 1556 911 1568
rect 865 680 871 1556
rect 905 680 911 1556
rect 865 668 911 680
rect 1013 1556 1059 1568
rect 1013 680 1019 1556
rect 1053 680 1059 1556
rect 1013 668 1059 680
rect 1161 1556 1207 1568
rect 1161 680 1167 1556
rect 1201 680 1207 1556
rect 1161 668 1207 680
rect 1309 1556 1355 1568
rect 1309 680 1315 1556
rect 1349 680 1355 1556
rect 1309 668 1355 680
rect 1457 1556 1503 1568
rect 1457 680 1463 1556
rect 1497 680 1503 1556
rect 1457 668 1503 680
rect 1605 1556 1651 1568
rect 1605 680 1611 1556
rect 1645 680 1651 1556
rect 1605 668 1651 680
rect 1753 1556 1799 1568
rect 1753 680 1759 1556
rect 1793 680 1799 1556
rect 1753 668 1799 680
rect 1901 1556 1947 1568
rect 1901 680 1907 1556
rect 1941 680 1947 1556
rect 1901 668 1947 680
rect 2049 1556 2095 1568
rect 2049 680 2055 1556
rect 2089 680 2095 1556
rect 2049 668 2095 680
rect 2197 1556 2243 1568
rect 2197 680 2203 1556
rect 2237 680 2243 1556
rect 2197 668 2243 680
rect 2345 1556 2391 1568
rect 2345 680 2351 1556
rect 2385 680 2391 1556
rect 2345 668 2391 680
rect 2493 1556 2539 1568
rect 2493 680 2499 1556
rect 2533 680 2539 1556
rect 2493 668 2539 680
rect 2641 1556 2687 1568
rect 2641 680 2647 1556
rect 2681 680 2687 1556
rect 2641 668 2687 680
rect 2789 1556 2835 1568
rect 2789 680 2795 1556
rect 2829 680 2835 1556
rect 2789 668 2835 680
rect 2937 1556 2983 1568
rect 2937 680 2943 1556
rect 2977 680 2983 1556
rect 2937 668 2983 680
rect 3085 1556 3131 1568
rect 3085 680 3091 1556
rect 3125 680 3131 1556
rect 3085 668 3131 680
rect 3233 1556 3279 1568
rect 3233 680 3239 1556
rect 3273 680 3279 1556
rect 3233 668 3279 680
rect 3381 1556 3427 1568
rect 3381 680 3387 1556
rect 3421 680 3427 1556
rect 3381 668 3427 680
rect 3529 1556 3575 1568
rect 3529 680 3535 1556
rect 3569 680 3575 1556
rect 3529 668 3575 680
rect 3677 1556 3723 1568
rect 3677 680 3683 1556
rect 3717 680 3723 1556
rect 3677 668 3723 680
rect -3667 630 -3585 636
rect -3667 596 -3655 630
rect -3597 596 -3585 630
rect -3667 590 -3585 596
rect -3519 630 -3437 636
rect -3519 596 -3507 630
rect -3449 596 -3437 630
rect -3519 590 -3437 596
rect -3371 630 -3289 636
rect -3371 596 -3359 630
rect -3301 596 -3289 630
rect -3371 590 -3289 596
rect -3223 630 -3141 636
rect -3223 596 -3211 630
rect -3153 596 -3141 630
rect -3223 590 -3141 596
rect -3075 630 -2993 636
rect -3075 596 -3063 630
rect -3005 596 -2993 630
rect -3075 590 -2993 596
rect -2927 630 -2845 636
rect -2927 596 -2915 630
rect -2857 596 -2845 630
rect -2927 590 -2845 596
rect -2779 630 -2697 636
rect -2779 596 -2767 630
rect -2709 596 -2697 630
rect -2779 590 -2697 596
rect -2631 630 -2549 636
rect -2631 596 -2619 630
rect -2561 596 -2549 630
rect -2631 590 -2549 596
rect -2483 630 -2401 636
rect -2483 596 -2471 630
rect -2413 596 -2401 630
rect -2483 590 -2401 596
rect -2335 630 -2253 636
rect -2335 596 -2323 630
rect -2265 596 -2253 630
rect -2335 590 -2253 596
rect -2187 630 -2105 636
rect -2187 596 -2175 630
rect -2117 596 -2105 630
rect -2187 590 -2105 596
rect -2039 630 -1957 636
rect -2039 596 -2027 630
rect -1969 596 -1957 630
rect -2039 590 -1957 596
rect -1891 630 -1809 636
rect -1891 596 -1879 630
rect -1821 596 -1809 630
rect -1891 590 -1809 596
rect -1743 630 -1661 636
rect -1743 596 -1731 630
rect -1673 596 -1661 630
rect -1743 590 -1661 596
rect -1595 630 -1513 636
rect -1595 596 -1583 630
rect -1525 596 -1513 630
rect -1595 590 -1513 596
rect -1447 630 -1365 636
rect -1447 596 -1435 630
rect -1377 596 -1365 630
rect -1447 590 -1365 596
rect -1299 630 -1217 636
rect -1299 596 -1287 630
rect -1229 596 -1217 630
rect -1299 590 -1217 596
rect -1151 630 -1069 636
rect -1151 596 -1139 630
rect -1081 596 -1069 630
rect -1151 590 -1069 596
rect -1003 630 -921 636
rect -1003 596 -991 630
rect -933 596 -921 630
rect -1003 590 -921 596
rect -855 630 -773 636
rect -855 596 -843 630
rect -785 596 -773 630
rect -855 590 -773 596
rect -707 630 -625 636
rect -707 596 -695 630
rect -637 596 -625 630
rect -707 590 -625 596
rect -559 630 -477 636
rect -559 596 -547 630
rect -489 596 -477 630
rect -559 590 -477 596
rect -411 630 -329 636
rect -411 596 -399 630
rect -341 596 -329 630
rect -411 590 -329 596
rect -263 630 -181 636
rect -263 596 -251 630
rect -193 596 -181 630
rect -263 590 -181 596
rect -115 630 -33 636
rect -115 596 -103 630
rect -45 596 -33 630
rect -115 590 -33 596
rect 33 630 115 636
rect 33 596 45 630
rect 103 596 115 630
rect 33 590 115 596
rect 181 630 263 636
rect 181 596 193 630
rect 251 596 263 630
rect 181 590 263 596
rect 329 630 411 636
rect 329 596 341 630
rect 399 596 411 630
rect 329 590 411 596
rect 477 630 559 636
rect 477 596 489 630
rect 547 596 559 630
rect 477 590 559 596
rect 625 630 707 636
rect 625 596 637 630
rect 695 596 707 630
rect 625 590 707 596
rect 773 630 855 636
rect 773 596 785 630
rect 843 596 855 630
rect 773 590 855 596
rect 921 630 1003 636
rect 921 596 933 630
rect 991 596 1003 630
rect 921 590 1003 596
rect 1069 630 1151 636
rect 1069 596 1081 630
rect 1139 596 1151 630
rect 1069 590 1151 596
rect 1217 630 1299 636
rect 1217 596 1229 630
rect 1287 596 1299 630
rect 1217 590 1299 596
rect 1365 630 1447 636
rect 1365 596 1377 630
rect 1435 596 1447 630
rect 1365 590 1447 596
rect 1513 630 1595 636
rect 1513 596 1525 630
rect 1583 596 1595 630
rect 1513 590 1595 596
rect 1661 630 1743 636
rect 1661 596 1673 630
rect 1731 596 1743 630
rect 1661 590 1743 596
rect 1809 630 1891 636
rect 1809 596 1821 630
rect 1879 596 1891 630
rect 1809 590 1891 596
rect 1957 630 2039 636
rect 1957 596 1969 630
rect 2027 596 2039 630
rect 1957 590 2039 596
rect 2105 630 2187 636
rect 2105 596 2117 630
rect 2175 596 2187 630
rect 2105 590 2187 596
rect 2253 630 2335 636
rect 2253 596 2265 630
rect 2323 596 2335 630
rect 2253 590 2335 596
rect 2401 630 2483 636
rect 2401 596 2413 630
rect 2471 596 2483 630
rect 2401 590 2483 596
rect 2549 630 2631 636
rect 2549 596 2561 630
rect 2619 596 2631 630
rect 2549 590 2631 596
rect 2697 630 2779 636
rect 2697 596 2709 630
rect 2767 596 2779 630
rect 2697 590 2779 596
rect 2845 630 2927 636
rect 2845 596 2857 630
rect 2915 596 2927 630
rect 2845 590 2927 596
rect 2993 630 3075 636
rect 2993 596 3005 630
rect 3063 596 3075 630
rect 2993 590 3075 596
rect 3141 630 3223 636
rect 3141 596 3153 630
rect 3211 596 3223 630
rect 3141 590 3223 596
rect 3289 630 3371 636
rect 3289 596 3301 630
rect 3359 596 3371 630
rect 3289 590 3371 596
rect 3437 630 3519 636
rect 3437 596 3449 630
rect 3507 596 3519 630
rect 3437 590 3519 596
rect 3585 630 3667 636
rect 3585 596 3597 630
rect 3655 596 3667 630
rect 3585 590 3667 596
rect -3667 522 -3585 528
rect -3667 488 -3655 522
rect -3597 488 -3585 522
rect -3667 482 -3585 488
rect -3519 522 -3437 528
rect -3519 488 -3507 522
rect -3449 488 -3437 522
rect -3519 482 -3437 488
rect -3371 522 -3289 528
rect -3371 488 -3359 522
rect -3301 488 -3289 522
rect -3371 482 -3289 488
rect -3223 522 -3141 528
rect -3223 488 -3211 522
rect -3153 488 -3141 522
rect -3223 482 -3141 488
rect -3075 522 -2993 528
rect -3075 488 -3063 522
rect -3005 488 -2993 522
rect -3075 482 -2993 488
rect -2927 522 -2845 528
rect -2927 488 -2915 522
rect -2857 488 -2845 522
rect -2927 482 -2845 488
rect -2779 522 -2697 528
rect -2779 488 -2767 522
rect -2709 488 -2697 522
rect -2779 482 -2697 488
rect -2631 522 -2549 528
rect -2631 488 -2619 522
rect -2561 488 -2549 522
rect -2631 482 -2549 488
rect -2483 522 -2401 528
rect -2483 488 -2471 522
rect -2413 488 -2401 522
rect -2483 482 -2401 488
rect -2335 522 -2253 528
rect -2335 488 -2323 522
rect -2265 488 -2253 522
rect -2335 482 -2253 488
rect -2187 522 -2105 528
rect -2187 488 -2175 522
rect -2117 488 -2105 522
rect -2187 482 -2105 488
rect -2039 522 -1957 528
rect -2039 488 -2027 522
rect -1969 488 -1957 522
rect -2039 482 -1957 488
rect -1891 522 -1809 528
rect -1891 488 -1879 522
rect -1821 488 -1809 522
rect -1891 482 -1809 488
rect -1743 522 -1661 528
rect -1743 488 -1731 522
rect -1673 488 -1661 522
rect -1743 482 -1661 488
rect -1595 522 -1513 528
rect -1595 488 -1583 522
rect -1525 488 -1513 522
rect -1595 482 -1513 488
rect -1447 522 -1365 528
rect -1447 488 -1435 522
rect -1377 488 -1365 522
rect -1447 482 -1365 488
rect -1299 522 -1217 528
rect -1299 488 -1287 522
rect -1229 488 -1217 522
rect -1299 482 -1217 488
rect -1151 522 -1069 528
rect -1151 488 -1139 522
rect -1081 488 -1069 522
rect -1151 482 -1069 488
rect -1003 522 -921 528
rect -1003 488 -991 522
rect -933 488 -921 522
rect -1003 482 -921 488
rect -855 522 -773 528
rect -855 488 -843 522
rect -785 488 -773 522
rect -855 482 -773 488
rect -707 522 -625 528
rect -707 488 -695 522
rect -637 488 -625 522
rect -707 482 -625 488
rect -559 522 -477 528
rect -559 488 -547 522
rect -489 488 -477 522
rect -559 482 -477 488
rect -411 522 -329 528
rect -411 488 -399 522
rect -341 488 -329 522
rect -411 482 -329 488
rect -263 522 -181 528
rect -263 488 -251 522
rect -193 488 -181 522
rect -263 482 -181 488
rect -115 522 -33 528
rect -115 488 -103 522
rect -45 488 -33 522
rect -115 482 -33 488
rect 33 522 115 528
rect 33 488 45 522
rect 103 488 115 522
rect 33 482 115 488
rect 181 522 263 528
rect 181 488 193 522
rect 251 488 263 522
rect 181 482 263 488
rect 329 522 411 528
rect 329 488 341 522
rect 399 488 411 522
rect 329 482 411 488
rect 477 522 559 528
rect 477 488 489 522
rect 547 488 559 522
rect 477 482 559 488
rect 625 522 707 528
rect 625 488 637 522
rect 695 488 707 522
rect 625 482 707 488
rect 773 522 855 528
rect 773 488 785 522
rect 843 488 855 522
rect 773 482 855 488
rect 921 522 1003 528
rect 921 488 933 522
rect 991 488 1003 522
rect 921 482 1003 488
rect 1069 522 1151 528
rect 1069 488 1081 522
rect 1139 488 1151 522
rect 1069 482 1151 488
rect 1217 522 1299 528
rect 1217 488 1229 522
rect 1287 488 1299 522
rect 1217 482 1299 488
rect 1365 522 1447 528
rect 1365 488 1377 522
rect 1435 488 1447 522
rect 1365 482 1447 488
rect 1513 522 1595 528
rect 1513 488 1525 522
rect 1583 488 1595 522
rect 1513 482 1595 488
rect 1661 522 1743 528
rect 1661 488 1673 522
rect 1731 488 1743 522
rect 1661 482 1743 488
rect 1809 522 1891 528
rect 1809 488 1821 522
rect 1879 488 1891 522
rect 1809 482 1891 488
rect 1957 522 2039 528
rect 1957 488 1969 522
rect 2027 488 2039 522
rect 1957 482 2039 488
rect 2105 522 2187 528
rect 2105 488 2117 522
rect 2175 488 2187 522
rect 2105 482 2187 488
rect 2253 522 2335 528
rect 2253 488 2265 522
rect 2323 488 2335 522
rect 2253 482 2335 488
rect 2401 522 2483 528
rect 2401 488 2413 522
rect 2471 488 2483 522
rect 2401 482 2483 488
rect 2549 522 2631 528
rect 2549 488 2561 522
rect 2619 488 2631 522
rect 2549 482 2631 488
rect 2697 522 2779 528
rect 2697 488 2709 522
rect 2767 488 2779 522
rect 2697 482 2779 488
rect 2845 522 2927 528
rect 2845 488 2857 522
rect 2915 488 2927 522
rect 2845 482 2927 488
rect 2993 522 3075 528
rect 2993 488 3005 522
rect 3063 488 3075 522
rect 2993 482 3075 488
rect 3141 522 3223 528
rect 3141 488 3153 522
rect 3211 488 3223 522
rect 3141 482 3223 488
rect 3289 522 3371 528
rect 3289 488 3301 522
rect 3359 488 3371 522
rect 3289 482 3371 488
rect 3437 522 3519 528
rect 3437 488 3449 522
rect 3507 488 3519 522
rect 3437 482 3519 488
rect 3585 522 3667 528
rect 3585 488 3597 522
rect 3655 488 3667 522
rect 3585 482 3667 488
rect -3723 438 -3677 450
rect -3723 -438 -3717 438
rect -3683 -438 -3677 438
rect -3723 -450 -3677 -438
rect -3575 438 -3529 450
rect -3575 -438 -3569 438
rect -3535 -438 -3529 438
rect -3575 -450 -3529 -438
rect -3427 438 -3381 450
rect -3427 -438 -3421 438
rect -3387 -438 -3381 438
rect -3427 -450 -3381 -438
rect -3279 438 -3233 450
rect -3279 -438 -3273 438
rect -3239 -438 -3233 438
rect -3279 -450 -3233 -438
rect -3131 438 -3085 450
rect -3131 -438 -3125 438
rect -3091 -438 -3085 438
rect -3131 -450 -3085 -438
rect -2983 438 -2937 450
rect -2983 -438 -2977 438
rect -2943 -438 -2937 438
rect -2983 -450 -2937 -438
rect -2835 438 -2789 450
rect -2835 -438 -2829 438
rect -2795 -438 -2789 438
rect -2835 -450 -2789 -438
rect -2687 438 -2641 450
rect -2687 -438 -2681 438
rect -2647 -438 -2641 438
rect -2687 -450 -2641 -438
rect -2539 438 -2493 450
rect -2539 -438 -2533 438
rect -2499 -438 -2493 438
rect -2539 -450 -2493 -438
rect -2391 438 -2345 450
rect -2391 -438 -2385 438
rect -2351 -438 -2345 438
rect -2391 -450 -2345 -438
rect -2243 438 -2197 450
rect -2243 -438 -2237 438
rect -2203 -438 -2197 438
rect -2243 -450 -2197 -438
rect -2095 438 -2049 450
rect -2095 -438 -2089 438
rect -2055 -438 -2049 438
rect -2095 -450 -2049 -438
rect -1947 438 -1901 450
rect -1947 -438 -1941 438
rect -1907 -438 -1901 438
rect -1947 -450 -1901 -438
rect -1799 438 -1753 450
rect -1799 -438 -1793 438
rect -1759 -438 -1753 438
rect -1799 -450 -1753 -438
rect -1651 438 -1605 450
rect -1651 -438 -1645 438
rect -1611 -438 -1605 438
rect -1651 -450 -1605 -438
rect -1503 438 -1457 450
rect -1503 -438 -1497 438
rect -1463 -438 -1457 438
rect -1503 -450 -1457 -438
rect -1355 438 -1309 450
rect -1355 -438 -1349 438
rect -1315 -438 -1309 438
rect -1355 -450 -1309 -438
rect -1207 438 -1161 450
rect -1207 -438 -1201 438
rect -1167 -438 -1161 438
rect -1207 -450 -1161 -438
rect -1059 438 -1013 450
rect -1059 -438 -1053 438
rect -1019 -438 -1013 438
rect -1059 -450 -1013 -438
rect -911 438 -865 450
rect -911 -438 -905 438
rect -871 -438 -865 438
rect -911 -450 -865 -438
rect -763 438 -717 450
rect -763 -438 -757 438
rect -723 -438 -717 438
rect -763 -450 -717 -438
rect -615 438 -569 450
rect -615 -438 -609 438
rect -575 -438 -569 438
rect -615 -450 -569 -438
rect -467 438 -421 450
rect -467 -438 -461 438
rect -427 -438 -421 438
rect -467 -450 -421 -438
rect -319 438 -273 450
rect -319 -438 -313 438
rect -279 -438 -273 438
rect -319 -450 -273 -438
rect -171 438 -125 450
rect -171 -438 -165 438
rect -131 -438 -125 438
rect -171 -450 -125 -438
rect -23 438 23 450
rect -23 -438 -17 438
rect 17 -438 23 438
rect -23 -450 23 -438
rect 125 438 171 450
rect 125 -438 131 438
rect 165 -438 171 438
rect 125 -450 171 -438
rect 273 438 319 450
rect 273 -438 279 438
rect 313 -438 319 438
rect 273 -450 319 -438
rect 421 438 467 450
rect 421 -438 427 438
rect 461 -438 467 438
rect 421 -450 467 -438
rect 569 438 615 450
rect 569 -438 575 438
rect 609 -438 615 438
rect 569 -450 615 -438
rect 717 438 763 450
rect 717 -438 723 438
rect 757 -438 763 438
rect 717 -450 763 -438
rect 865 438 911 450
rect 865 -438 871 438
rect 905 -438 911 438
rect 865 -450 911 -438
rect 1013 438 1059 450
rect 1013 -438 1019 438
rect 1053 -438 1059 438
rect 1013 -450 1059 -438
rect 1161 438 1207 450
rect 1161 -438 1167 438
rect 1201 -438 1207 438
rect 1161 -450 1207 -438
rect 1309 438 1355 450
rect 1309 -438 1315 438
rect 1349 -438 1355 438
rect 1309 -450 1355 -438
rect 1457 438 1503 450
rect 1457 -438 1463 438
rect 1497 -438 1503 438
rect 1457 -450 1503 -438
rect 1605 438 1651 450
rect 1605 -438 1611 438
rect 1645 -438 1651 438
rect 1605 -450 1651 -438
rect 1753 438 1799 450
rect 1753 -438 1759 438
rect 1793 -438 1799 438
rect 1753 -450 1799 -438
rect 1901 438 1947 450
rect 1901 -438 1907 438
rect 1941 -438 1947 438
rect 1901 -450 1947 -438
rect 2049 438 2095 450
rect 2049 -438 2055 438
rect 2089 -438 2095 438
rect 2049 -450 2095 -438
rect 2197 438 2243 450
rect 2197 -438 2203 438
rect 2237 -438 2243 438
rect 2197 -450 2243 -438
rect 2345 438 2391 450
rect 2345 -438 2351 438
rect 2385 -438 2391 438
rect 2345 -450 2391 -438
rect 2493 438 2539 450
rect 2493 -438 2499 438
rect 2533 -438 2539 438
rect 2493 -450 2539 -438
rect 2641 438 2687 450
rect 2641 -438 2647 438
rect 2681 -438 2687 438
rect 2641 -450 2687 -438
rect 2789 438 2835 450
rect 2789 -438 2795 438
rect 2829 -438 2835 438
rect 2789 -450 2835 -438
rect 2937 438 2983 450
rect 2937 -438 2943 438
rect 2977 -438 2983 438
rect 2937 -450 2983 -438
rect 3085 438 3131 450
rect 3085 -438 3091 438
rect 3125 -438 3131 438
rect 3085 -450 3131 -438
rect 3233 438 3279 450
rect 3233 -438 3239 438
rect 3273 -438 3279 438
rect 3233 -450 3279 -438
rect 3381 438 3427 450
rect 3381 -438 3387 438
rect 3421 -438 3427 438
rect 3381 -450 3427 -438
rect 3529 438 3575 450
rect 3529 -438 3535 438
rect 3569 -438 3575 438
rect 3529 -450 3575 -438
rect 3677 438 3723 450
rect 3677 -438 3683 438
rect 3717 -438 3723 438
rect 3677 -450 3723 -438
rect -3667 -488 -3585 -482
rect -3667 -522 -3655 -488
rect -3597 -522 -3585 -488
rect -3667 -528 -3585 -522
rect -3519 -488 -3437 -482
rect -3519 -522 -3507 -488
rect -3449 -522 -3437 -488
rect -3519 -528 -3437 -522
rect -3371 -488 -3289 -482
rect -3371 -522 -3359 -488
rect -3301 -522 -3289 -488
rect -3371 -528 -3289 -522
rect -3223 -488 -3141 -482
rect -3223 -522 -3211 -488
rect -3153 -522 -3141 -488
rect -3223 -528 -3141 -522
rect -3075 -488 -2993 -482
rect -3075 -522 -3063 -488
rect -3005 -522 -2993 -488
rect -3075 -528 -2993 -522
rect -2927 -488 -2845 -482
rect -2927 -522 -2915 -488
rect -2857 -522 -2845 -488
rect -2927 -528 -2845 -522
rect -2779 -488 -2697 -482
rect -2779 -522 -2767 -488
rect -2709 -522 -2697 -488
rect -2779 -528 -2697 -522
rect -2631 -488 -2549 -482
rect -2631 -522 -2619 -488
rect -2561 -522 -2549 -488
rect -2631 -528 -2549 -522
rect -2483 -488 -2401 -482
rect -2483 -522 -2471 -488
rect -2413 -522 -2401 -488
rect -2483 -528 -2401 -522
rect -2335 -488 -2253 -482
rect -2335 -522 -2323 -488
rect -2265 -522 -2253 -488
rect -2335 -528 -2253 -522
rect -2187 -488 -2105 -482
rect -2187 -522 -2175 -488
rect -2117 -522 -2105 -488
rect -2187 -528 -2105 -522
rect -2039 -488 -1957 -482
rect -2039 -522 -2027 -488
rect -1969 -522 -1957 -488
rect -2039 -528 -1957 -522
rect -1891 -488 -1809 -482
rect -1891 -522 -1879 -488
rect -1821 -522 -1809 -488
rect -1891 -528 -1809 -522
rect -1743 -488 -1661 -482
rect -1743 -522 -1731 -488
rect -1673 -522 -1661 -488
rect -1743 -528 -1661 -522
rect -1595 -488 -1513 -482
rect -1595 -522 -1583 -488
rect -1525 -522 -1513 -488
rect -1595 -528 -1513 -522
rect -1447 -488 -1365 -482
rect -1447 -522 -1435 -488
rect -1377 -522 -1365 -488
rect -1447 -528 -1365 -522
rect -1299 -488 -1217 -482
rect -1299 -522 -1287 -488
rect -1229 -522 -1217 -488
rect -1299 -528 -1217 -522
rect -1151 -488 -1069 -482
rect -1151 -522 -1139 -488
rect -1081 -522 -1069 -488
rect -1151 -528 -1069 -522
rect -1003 -488 -921 -482
rect -1003 -522 -991 -488
rect -933 -522 -921 -488
rect -1003 -528 -921 -522
rect -855 -488 -773 -482
rect -855 -522 -843 -488
rect -785 -522 -773 -488
rect -855 -528 -773 -522
rect -707 -488 -625 -482
rect -707 -522 -695 -488
rect -637 -522 -625 -488
rect -707 -528 -625 -522
rect -559 -488 -477 -482
rect -559 -522 -547 -488
rect -489 -522 -477 -488
rect -559 -528 -477 -522
rect -411 -488 -329 -482
rect -411 -522 -399 -488
rect -341 -522 -329 -488
rect -411 -528 -329 -522
rect -263 -488 -181 -482
rect -263 -522 -251 -488
rect -193 -522 -181 -488
rect -263 -528 -181 -522
rect -115 -488 -33 -482
rect -115 -522 -103 -488
rect -45 -522 -33 -488
rect -115 -528 -33 -522
rect 33 -488 115 -482
rect 33 -522 45 -488
rect 103 -522 115 -488
rect 33 -528 115 -522
rect 181 -488 263 -482
rect 181 -522 193 -488
rect 251 -522 263 -488
rect 181 -528 263 -522
rect 329 -488 411 -482
rect 329 -522 341 -488
rect 399 -522 411 -488
rect 329 -528 411 -522
rect 477 -488 559 -482
rect 477 -522 489 -488
rect 547 -522 559 -488
rect 477 -528 559 -522
rect 625 -488 707 -482
rect 625 -522 637 -488
rect 695 -522 707 -488
rect 625 -528 707 -522
rect 773 -488 855 -482
rect 773 -522 785 -488
rect 843 -522 855 -488
rect 773 -528 855 -522
rect 921 -488 1003 -482
rect 921 -522 933 -488
rect 991 -522 1003 -488
rect 921 -528 1003 -522
rect 1069 -488 1151 -482
rect 1069 -522 1081 -488
rect 1139 -522 1151 -488
rect 1069 -528 1151 -522
rect 1217 -488 1299 -482
rect 1217 -522 1229 -488
rect 1287 -522 1299 -488
rect 1217 -528 1299 -522
rect 1365 -488 1447 -482
rect 1365 -522 1377 -488
rect 1435 -522 1447 -488
rect 1365 -528 1447 -522
rect 1513 -488 1595 -482
rect 1513 -522 1525 -488
rect 1583 -522 1595 -488
rect 1513 -528 1595 -522
rect 1661 -488 1743 -482
rect 1661 -522 1673 -488
rect 1731 -522 1743 -488
rect 1661 -528 1743 -522
rect 1809 -488 1891 -482
rect 1809 -522 1821 -488
rect 1879 -522 1891 -488
rect 1809 -528 1891 -522
rect 1957 -488 2039 -482
rect 1957 -522 1969 -488
rect 2027 -522 2039 -488
rect 1957 -528 2039 -522
rect 2105 -488 2187 -482
rect 2105 -522 2117 -488
rect 2175 -522 2187 -488
rect 2105 -528 2187 -522
rect 2253 -488 2335 -482
rect 2253 -522 2265 -488
rect 2323 -522 2335 -488
rect 2253 -528 2335 -522
rect 2401 -488 2483 -482
rect 2401 -522 2413 -488
rect 2471 -522 2483 -488
rect 2401 -528 2483 -522
rect 2549 -488 2631 -482
rect 2549 -522 2561 -488
rect 2619 -522 2631 -488
rect 2549 -528 2631 -522
rect 2697 -488 2779 -482
rect 2697 -522 2709 -488
rect 2767 -522 2779 -488
rect 2697 -528 2779 -522
rect 2845 -488 2927 -482
rect 2845 -522 2857 -488
rect 2915 -522 2927 -488
rect 2845 -528 2927 -522
rect 2993 -488 3075 -482
rect 2993 -522 3005 -488
rect 3063 -522 3075 -488
rect 2993 -528 3075 -522
rect 3141 -488 3223 -482
rect 3141 -522 3153 -488
rect 3211 -522 3223 -488
rect 3141 -528 3223 -522
rect 3289 -488 3371 -482
rect 3289 -522 3301 -488
rect 3359 -522 3371 -488
rect 3289 -528 3371 -522
rect 3437 -488 3519 -482
rect 3437 -522 3449 -488
rect 3507 -522 3519 -488
rect 3437 -528 3519 -522
rect 3585 -488 3667 -482
rect 3585 -522 3597 -488
rect 3655 -522 3667 -488
rect 3585 -528 3667 -522
rect -3667 -596 -3585 -590
rect -3667 -630 -3655 -596
rect -3597 -630 -3585 -596
rect -3667 -636 -3585 -630
rect -3519 -596 -3437 -590
rect -3519 -630 -3507 -596
rect -3449 -630 -3437 -596
rect -3519 -636 -3437 -630
rect -3371 -596 -3289 -590
rect -3371 -630 -3359 -596
rect -3301 -630 -3289 -596
rect -3371 -636 -3289 -630
rect -3223 -596 -3141 -590
rect -3223 -630 -3211 -596
rect -3153 -630 -3141 -596
rect -3223 -636 -3141 -630
rect -3075 -596 -2993 -590
rect -3075 -630 -3063 -596
rect -3005 -630 -2993 -596
rect -3075 -636 -2993 -630
rect -2927 -596 -2845 -590
rect -2927 -630 -2915 -596
rect -2857 -630 -2845 -596
rect -2927 -636 -2845 -630
rect -2779 -596 -2697 -590
rect -2779 -630 -2767 -596
rect -2709 -630 -2697 -596
rect -2779 -636 -2697 -630
rect -2631 -596 -2549 -590
rect -2631 -630 -2619 -596
rect -2561 -630 -2549 -596
rect -2631 -636 -2549 -630
rect -2483 -596 -2401 -590
rect -2483 -630 -2471 -596
rect -2413 -630 -2401 -596
rect -2483 -636 -2401 -630
rect -2335 -596 -2253 -590
rect -2335 -630 -2323 -596
rect -2265 -630 -2253 -596
rect -2335 -636 -2253 -630
rect -2187 -596 -2105 -590
rect -2187 -630 -2175 -596
rect -2117 -630 -2105 -596
rect -2187 -636 -2105 -630
rect -2039 -596 -1957 -590
rect -2039 -630 -2027 -596
rect -1969 -630 -1957 -596
rect -2039 -636 -1957 -630
rect -1891 -596 -1809 -590
rect -1891 -630 -1879 -596
rect -1821 -630 -1809 -596
rect -1891 -636 -1809 -630
rect -1743 -596 -1661 -590
rect -1743 -630 -1731 -596
rect -1673 -630 -1661 -596
rect -1743 -636 -1661 -630
rect -1595 -596 -1513 -590
rect -1595 -630 -1583 -596
rect -1525 -630 -1513 -596
rect -1595 -636 -1513 -630
rect -1447 -596 -1365 -590
rect -1447 -630 -1435 -596
rect -1377 -630 -1365 -596
rect -1447 -636 -1365 -630
rect -1299 -596 -1217 -590
rect -1299 -630 -1287 -596
rect -1229 -630 -1217 -596
rect -1299 -636 -1217 -630
rect -1151 -596 -1069 -590
rect -1151 -630 -1139 -596
rect -1081 -630 -1069 -596
rect -1151 -636 -1069 -630
rect -1003 -596 -921 -590
rect -1003 -630 -991 -596
rect -933 -630 -921 -596
rect -1003 -636 -921 -630
rect -855 -596 -773 -590
rect -855 -630 -843 -596
rect -785 -630 -773 -596
rect -855 -636 -773 -630
rect -707 -596 -625 -590
rect -707 -630 -695 -596
rect -637 -630 -625 -596
rect -707 -636 -625 -630
rect -559 -596 -477 -590
rect -559 -630 -547 -596
rect -489 -630 -477 -596
rect -559 -636 -477 -630
rect -411 -596 -329 -590
rect -411 -630 -399 -596
rect -341 -630 -329 -596
rect -411 -636 -329 -630
rect -263 -596 -181 -590
rect -263 -630 -251 -596
rect -193 -630 -181 -596
rect -263 -636 -181 -630
rect -115 -596 -33 -590
rect -115 -630 -103 -596
rect -45 -630 -33 -596
rect -115 -636 -33 -630
rect 33 -596 115 -590
rect 33 -630 45 -596
rect 103 -630 115 -596
rect 33 -636 115 -630
rect 181 -596 263 -590
rect 181 -630 193 -596
rect 251 -630 263 -596
rect 181 -636 263 -630
rect 329 -596 411 -590
rect 329 -630 341 -596
rect 399 -630 411 -596
rect 329 -636 411 -630
rect 477 -596 559 -590
rect 477 -630 489 -596
rect 547 -630 559 -596
rect 477 -636 559 -630
rect 625 -596 707 -590
rect 625 -630 637 -596
rect 695 -630 707 -596
rect 625 -636 707 -630
rect 773 -596 855 -590
rect 773 -630 785 -596
rect 843 -630 855 -596
rect 773 -636 855 -630
rect 921 -596 1003 -590
rect 921 -630 933 -596
rect 991 -630 1003 -596
rect 921 -636 1003 -630
rect 1069 -596 1151 -590
rect 1069 -630 1081 -596
rect 1139 -630 1151 -596
rect 1069 -636 1151 -630
rect 1217 -596 1299 -590
rect 1217 -630 1229 -596
rect 1287 -630 1299 -596
rect 1217 -636 1299 -630
rect 1365 -596 1447 -590
rect 1365 -630 1377 -596
rect 1435 -630 1447 -596
rect 1365 -636 1447 -630
rect 1513 -596 1595 -590
rect 1513 -630 1525 -596
rect 1583 -630 1595 -596
rect 1513 -636 1595 -630
rect 1661 -596 1743 -590
rect 1661 -630 1673 -596
rect 1731 -630 1743 -596
rect 1661 -636 1743 -630
rect 1809 -596 1891 -590
rect 1809 -630 1821 -596
rect 1879 -630 1891 -596
rect 1809 -636 1891 -630
rect 1957 -596 2039 -590
rect 1957 -630 1969 -596
rect 2027 -630 2039 -596
rect 1957 -636 2039 -630
rect 2105 -596 2187 -590
rect 2105 -630 2117 -596
rect 2175 -630 2187 -596
rect 2105 -636 2187 -630
rect 2253 -596 2335 -590
rect 2253 -630 2265 -596
rect 2323 -630 2335 -596
rect 2253 -636 2335 -630
rect 2401 -596 2483 -590
rect 2401 -630 2413 -596
rect 2471 -630 2483 -596
rect 2401 -636 2483 -630
rect 2549 -596 2631 -590
rect 2549 -630 2561 -596
rect 2619 -630 2631 -596
rect 2549 -636 2631 -630
rect 2697 -596 2779 -590
rect 2697 -630 2709 -596
rect 2767 -630 2779 -596
rect 2697 -636 2779 -630
rect 2845 -596 2927 -590
rect 2845 -630 2857 -596
rect 2915 -630 2927 -596
rect 2845 -636 2927 -630
rect 2993 -596 3075 -590
rect 2993 -630 3005 -596
rect 3063 -630 3075 -596
rect 2993 -636 3075 -630
rect 3141 -596 3223 -590
rect 3141 -630 3153 -596
rect 3211 -630 3223 -596
rect 3141 -636 3223 -630
rect 3289 -596 3371 -590
rect 3289 -630 3301 -596
rect 3359 -630 3371 -596
rect 3289 -636 3371 -630
rect 3437 -596 3519 -590
rect 3437 -630 3449 -596
rect 3507 -630 3519 -596
rect 3437 -636 3519 -630
rect 3585 -596 3667 -590
rect 3585 -630 3597 -596
rect 3655 -630 3667 -596
rect 3585 -636 3667 -630
rect -3723 -680 -3677 -668
rect -3723 -1556 -3717 -680
rect -3683 -1556 -3677 -680
rect -3723 -1568 -3677 -1556
rect -3575 -680 -3529 -668
rect -3575 -1556 -3569 -680
rect -3535 -1556 -3529 -680
rect -3575 -1568 -3529 -1556
rect -3427 -680 -3381 -668
rect -3427 -1556 -3421 -680
rect -3387 -1556 -3381 -680
rect -3427 -1568 -3381 -1556
rect -3279 -680 -3233 -668
rect -3279 -1556 -3273 -680
rect -3239 -1556 -3233 -680
rect -3279 -1568 -3233 -1556
rect -3131 -680 -3085 -668
rect -3131 -1556 -3125 -680
rect -3091 -1556 -3085 -680
rect -3131 -1568 -3085 -1556
rect -2983 -680 -2937 -668
rect -2983 -1556 -2977 -680
rect -2943 -1556 -2937 -680
rect -2983 -1568 -2937 -1556
rect -2835 -680 -2789 -668
rect -2835 -1556 -2829 -680
rect -2795 -1556 -2789 -680
rect -2835 -1568 -2789 -1556
rect -2687 -680 -2641 -668
rect -2687 -1556 -2681 -680
rect -2647 -1556 -2641 -680
rect -2687 -1568 -2641 -1556
rect -2539 -680 -2493 -668
rect -2539 -1556 -2533 -680
rect -2499 -1556 -2493 -680
rect -2539 -1568 -2493 -1556
rect -2391 -680 -2345 -668
rect -2391 -1556 -2385 -680
rect -2351 -1556 -2345 -680
rect -2391 -1568 -2345 -1556
rect -2243 -680 -2197 -668
rect -2243 -1556 -2237 -680
rect -2203 -1556 -2197 -680
rect -2243 -1568 -2197 -1556
rect -2095 -680 -2049 -668
rect -2095 -1556 -2089 -680
rect -2055 -1556 -2049 -680
rect -2095 -1568 -2049 -1556
rect -1947 -680 -1901 -668
rect -1947 -1556 -1941 -680
rect -1907 -1556 -1901 -680
rect -1947 -1568 -1901 -1556
rect -1799 -680 -1753 -668
rect -1799 -1556 -1793 -680
rect -1759 -1556 -1753 -680
rect -1799 -1568 -1753 -1556
rect -1651 -680 -1605 -668
rect -1651 -1556 -1645 -680
rect -1611 -1556 -1605 -680
rect -1651 -1568 -1605 -1556
rect -1503 -680 -1457 -668
rect -1503 -1556 -1497 -680
rect -1463 -1556 -1457 -680
rect -1503 -1568 -1457 -1556
rect -1355 -680 -1309 -668
rect -1355 -1556 -1349 -680
rect -1315 -1556 -1309 -680
rect -1355 -1568 -1309 -1556
rect -1207 -680 -1161 -668
rect -1207 -1556 -1201 -680
rect -1167 -1556 -1161 -680
rect -1207 -1568 -1161 -1556
rect -1059 -680 -1013 -668
rect -1059 -1556 -1053 -680
rect -1019 -1556 -1013 -680
rect -1059 -1568 -1013 -1556
rect -911 -680 -865 -668
rect -911 -1556 -905 -680
rect -871 -1556 -865 -680
rect -911 -1568 -865 -1556
rect -763 -680 -717 -668
rect -763 -1556 -757 -680
rect -723 -1556 -717 -680
rect -763 -1568 -717 -1556
rect -615 -680 -569 -668
rect -615 -1556 -609 -680
rect -575 -1556 -569 -680
rect -615 -1568 -569 -1556
rect -467 -680 -421 -668
rect -467 -1556 -461 -680
rect -427 -1556 -421 -680
rect -467 -1568 -421 -1556
rect -319 -680 -273 -668
rect -319 -1556 -313 -680
rect -279 -1556 -273 -680
rect -319 -1568 -273 -1556
rect -171 -680 -125 -668
rect -171 -1556 -165 -680
rect -131 -1556 -125 -680
rect -171 -1568 -125 -1556
rect -23 -680 23 -668
rect -23 -1556 -17 -680
rect 17 -1556 23 -680
rect -23 -1568 23 -1556
rect 125 -680 171 -668
rect 125 -1556 131 -680
rect 165 -1556 171 -680
rect 125 -1568 171 -1556
rect 273 -680 319 -668
rect 273 -1556 279 -680
rect 313 -1556 319 -680
rect 273 -1568 319 -1556
rect 421 -680 467 -668
rect 421 -1556 427 -680
rect 461 -1556 467 -680
rect 421 -1568 467 -1556
rect 569 -680 615 -668
rect 569 -1556 575 -680
rect 609 -1556 615 -680
rect 569 -1568 615 -1556
rect 717 -680 763 -668
rect 717 -1556 723 -680
rect 757 -1556 763 -680
rect 717 -1568 763 -1556
rect 865 -680 911 -668
rect 865 -1556 871 -680
rect 905 -1556 911 -680
rect 865 -1568 911 -1556
rect 1013 -680 1059 -668
rect 1013 -1556 1019 -680
rect 1053 -1556 1059 -680
rect 1013 -1568 1059 -1556
rect 1161 -680 1207 -668
rect 1161 -1556 1167 -680
rect 1201 -1556 1207 -680
rect 1161 -1568 1207 -1556
rect 1309 -680 1355 -668
rect 1309 -1556 1315 -680
rect 1349 -1556 1355 -680
rect 1309 -1568 1355 -1556
rect 1457 -680 1503 -668
rect 1457 -1556 1463 -680
rect 1497 -1556 1503 -680
rect 1457 -1568 1503 -1556
rect 1605 -680 1651 -668
rect 1605 -1556 1611 -680
rect 1645 -1556 1651 -680
rect 1605 -1568 1651 -1556
rect 1753 -680 1799 -668
rect 1753 -1556 1759 -680
rect 1793 -1556 1799 -680
rect 1753 -1568 1799 -1556
rect 1901 -680 1947 -668
rect 1901 -1556 1907 -680
rect 1941 -1556 1947 -680
rect 1901 -1568 1947 -1556
rect 2049 -680 2095 -668
rect 2049 -1556 2055 -680
rect 2089 -1556 2095 -680
rect 2049 -1568 2095 -1556
rect 2197 -680 2243 -668
rect 2197 -1556 2203 -680
rect 2237 -1556 2243 -680
rect 2197 -1568 2243 -1556
rect 2345 -680 2391 -668
rect 2345 -1556 2351 -680
rect 2385 -1556 2391 -680
rect 2345 -1568 2391 -1556
rect 2493 -680 2539 -668
rect 2493 -1556 2499 -680
rect 2533 -1556 2539 -680
rect 2493 -1568 2539 -1556
rect 2641 -680 2687 -668
rect 2641 -1556 2647 -680
rect 2681 -1556 2687 -680
rect 2641 -1568 2687 -1556
rect 2789 -680 2835 -668
rect 2789 -1556 2795 -680
rect 2829 -1556 2835 -680
rect 2789 -1568 2835 -1556
rect 2937 -680 2983 -668
rect 2937 -1556 2943 -680
rect 2977 -1556 2983 -680
rect 2937 -1568 2983 -1556
rect 3085 -680 3131 -668
rect 3085 -1556 3091 -680
rect 3125 -1556 3131 -680
rect 3085 -1568 3131 -1556
rect 3233 -680 3279 -668
rect 3233 -1556 3239 -680
rect 3273 -1556 3279 -680
rect 3233 -1568 3279 -1556
rect 3381 -680 3427 -668
rect 3381 -1556 3387 -680
rect 3421 -1556 3427 -680
rect 3381 -1568 3427 -1556
rect 3529 -680 3575 -668
rect 3529 -1556 3535 -680
rect 3569 -1556 3575 -680
rect 3529 -1568 3575 -1556
rect 3677 -680 3723 -668
rect 3677 -1556 3683 -680
rect 3717 -1556 3723 -680
rect 3677 -1568 3723 -1556
rect -3667 -1606 -3585 -1600
rect -3667 -1640 -3655 -1606
rect -3597 -1640 -3585 -1606
rect -3667 -1646 -3585 -1640
rect -3519 -1606 -3437 -1600
rect -3519 -1640 -3507 -1606
rect -3449 -1640 -3437 -1606
rect -3519 -1646 -3437 -1640
rect -3371 -1606 -3289 -1600
rect -3371 -1640 -3359 -1606
rect -3301 -1640 -3289 -1606
rect -3371 -1646 -3289 -1640
rect -3223 -1606 -3141 -1600
rect -3223 -1640 -3211 -1606
rect -3153 -1640 -3141 -1606
rect -3223 -1646 -3141 -1640
rect -3075 -1606 -2993 -1600
rect -3075 -1640 -3063 -1606
rect -3005 -1640 -2993 -1606
rect -3075 -1646 -2993 -1640
rect -2927 -1606 -2845 -1600
rect -2927 -1640 -2915 -1606
rect -2857 -1640 -2845 -1606
rect -2927 -1646 -2845 -1640
rect -2779 -1606 -2697 -1600
rect -2779 -1640 -2767 -1606
rect -2709 -1640 -2697 -1606
rect -2779 -1646 -2697 -1640
rect -2631 -1606 -2549 -1600
rect -2631 -1640 -2619 -1606
rect -2561 -1640 -2549 -1606
rect -2631 -1646 -2549 -1640
rect -2483 -1606 -2401 -1600
rect -2483 -1640 -2471 -1606
rect -2413 -1640 -2401 -1606
rect -2483 -1646 -2401 -1640
rect -2335 -1606 -2253 -1600
rect -2335 -1640 -2323 -1606
rect -2265 -1640 -2253 -1606
rect -2335 -1646 -2253 -1640
rect -2187 -1606 -2105 -1600
rect -2187 -1640 -2175 -1606
rect -2117 -1640 -2105 -1606
rect -2187 -1646 -2105 -1640
rect -2039 -1606 -1957 -1600
rect -2039 -1640 -2027 -1606
rect -1969 -1640 -1957 -1606
rect -2039 -1646 -1957 -1640
rect -1891 -1606 -1809 -1600
rect -1891 -1640 -1879 -1606
rect -1821 -1640 -1809 -1606
rect -1891 -1646 -1809 -1640
rect -1743 -1606 -1661 -1600
rect -1743 -1640 -1731 -1606
rect -1673 -1640 -1661 -1606
rect -1743 -1646 -1661 -1640
rect -1595 -1606 -1513 -1600
rect -1595 -1640 -1583 -1606
rect -1525 -1640 -1513 -1606
rect -1595 -1646 -1513 -1640
rect -1447 -1606 -1365 -1600
rect -1447 -1640 -1435 -1606
rect -1377 -1640 -1365 -1606
rect -1447 -1646 -1365 -1640
rect -1299 -1606 -1217 -1600
rect -1299 -1640 -1287 -1606
rect -1229 -1640 -1217 -1606
rect -1299 -1646 -1217 -1640
rect -1151 -1606 -1069 -1600
rect -1151 -1640 -1139 -1606
rect -1081 -1640 -1069 -1606
rect -1151 -1646 -1069 -1640
rect -1003 -1606 -921 -1600
rect -1003 -1640 -991 -1606
rect -933 -1640 -921 -1606
rect -1003 -1646 -921 -1640
rect -855 -1606 -773 -1600
rect -855 -1640 -843 -1606
rect -785 -1640 -773 -1606
rect -855 -1646 -773 -1640
rect -707 -1606 -625 -1600
rect -707 -1640 -695 -1606
rect -637 -1640 -625 -1606
rect -707 -1646 -625 -1640
rect -559 -1606 -477 -1600
rect -559 -1640 -547 -1606
rect -489 -1640 -477 -1606
rect -559 -1646 -477 -1640
rect -411 -1606 -329 -1600
rect -411 -1640 -399 -1606
rect -341 -1640 -329 -1606
rect -411 -1646 -329 -1640
rect -263 -1606 -181 -1600
rect -263 -1640 -251 -1606
rect -193 -1640 -181 -1606
rect -263 -1646 -181 -1640
rect -115 -1606 -33 -1600
rect -115 -1640 -103 -1606
rect -45 -1640 -33 -1606
rect -115 -1646 -33 -1640
rect 33 -1606 115 -1600
rect 33 -1640 45 -1606
rect 103 -1640 115 -1606
rect 33 -1646 115 -1640
rect 181 -1606 263 -1600
rect 181 -1640 193 -1606
rect 251 -1640 263 -1606
rect 181 -1646 263 -1640
rect 329 -1606 411 -1600
rect 329 -1640 341 -1606
rect 399 -1640 411 -1606
rect 329 -1646 411 -1640
rect 477 -1606 559 -1600
rect 477 -1640 489 -1606
rect 547 -1640 559 -1606
rect 477 -1646 559 -1640
rect 625 -1606 707 -1600
rect 625 -1640 637 -1606
rect 695 -1640 707 -1606
rect 625 -1646 707 -1640
rect 773 -1606 855 -1600
rect 773 -1640 785 -1606
rect 843 -1640 855 -1606
rect 773 -1646 855 -1640
rect 921 -1606 1003 -1600
rect 921 -1640 933 -1606
rect 991 -1640 1003 -1606
rect 921 -1646 1003 -1640
rect 1069 -1606 1151 -1600
rect 1069 -1640 1081 -1606
rect 1139 -1640 1151 -1606
rect 1069 -1646 1151 -1640
rect 1217 -1606 1299 -1600
rect 1217 -1640 1229 -1606
rect 1287 -1640 1299 -1606
rect 1217 -1646 1299 -1640
rect 1365 -1606 1447 -1600
rect 1365 -1640 1377 -1606
rect 1435 -1640 1447 -1606
rect 1365 -1646 1447 -1640
rect 1513 -1606 1595 -1600
rect 1513 -1640 1525 -1606
rect 1583 -1640 1595 -1606
rect 1513 -1646 1595 -1640
rect 1661 -1606 1743 -1600
rect 1661 -1640 1673 -1606
rect 1731 -1640 1743 -1606
rect 1661 -1646 1743 -1640
rect 1809 -1606 1891 -1600
rect 1809 -1640 1821 -1606
rect 1879 -1640 1891 -1606
rect 1809 -1646 1891 -1640
rect 1957 -1606 2039 -1600
rect 1957 -1640 1969 -1606
rect 2027 -1640 2039 -1606
rect 1957 -1646 2039 -1640
rect 2105 -1606 2187 -1600
rect 2105 -1640 2117 -1606
rect 2175 -1640 2187 -1606
rect 2105 -1646 2187 -1640
rect 2253 -1606 2335 -1600
rect 2253 -1640 2265 -1606
rect 2323 -1640 2335 -1606
rect 2253 -1646 2335 -1640
rect 2401 -1606 2483 -1600
rect 2401 -1640 2413 -1606
rect 2471 -1640 2483 -1606
rect 2401 -1646 2483 -1640
rect 2549 -1606 2631 -1600
rect 2549 -1640 2561 -1606
rect 2619 -1640 2631 -1606
rect 2549 -1646 2631 -1640
rect 2697 -1606 2779 -1600
rect 2697 -1640 2709 -1606
rect 2767 -1640 2779 -1606
rect 2697 -1646 2779 -1640
rect 2845 -1606 2927 -1600
rect 2845 -1640 2857 -1606
rect 2915 -1640 2927 -1606
rect 2845 -1646 2927 -1640
rect 2993 -1606 3075 -1600
rect 2993 -1640 3005 -1606
rect 3063 -1640 3075 -1606
rect 2993 -1646 3075 -1640
rect 3141 -1606 3223 -1600
rect 3141 -1640 3153 -1606
rect 3211 -1640 3223 -1606
rect 3141 -1646 3223 -1640
rect 3289 -1606 3371 -1600
rect 3289 -1640 3301 -1606
rect 3359 -1640 3371 -1606
rect 3289 -1646 3371 -1640
rect 3437 -1606 3519 -1600
rect 3437 -1640 3449 -1606
rect 3507 -1640 3519 -1606
rect 3437 -1646 3519 -1640
rect 3585 -1606 3667 -1600
rect 3585 -1640 3597 -1606
rect 3655 -1640 3667 -1606
rect 3585 -1646 3667 -1640
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -3814 -1725 3814 1725
string parameters w 4.5 l 0.45 m 3 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
