VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_id_programming
  CLASS BLOCK ;
  FOREIGN user_id_programming ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 35.000 ;
  PIN mask_rev[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 31.000 7.270 35.000 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 31.000 14.170 35.000 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 31.000 16.470 35.000 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 31.000 9.570 35.000 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 31.000 27.970 35.000 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 31.000 23.370 35.000 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.000 3.440 35.000 4.040 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.000 27.240 35.000 27.840 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.000 23.840 35.000 24.440 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.000 6.840 35.000 7.440 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 31.000 32.570 35.000 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.000 13.640 35.000 14.240 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 31.000 4.970 35.000 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 31.000 30.270 35.000 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 31.000 21.070 35.000 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.000 17.040 35.000 17.640 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END mask_rev[9]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.685 5.200 26.285 27.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.700 5.200 18.300 27.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.715 5.200 10.315 27.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 24.500 29.440 26.100 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 16.460 29.440 18.060 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 8.420 29.440 10.020 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 20.695 5.200 22.295 27.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 12.705 5.200 14.305 27.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 20.480 29.440 22.080 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 12.440 29.440 14.040 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 29.440 27.285 ;
      LAYER met1 ;
        RECT 2.370 5.200 32.590 27.440 ;
      LAYER met2 ;
        RECT 2.400 30.720 4.410 31.125 ;
        RECT 5.250 30.720 6.710 31.125 ;
        RECT 7.550 30.720 9.010 31.125 ;
        RECT 9.850 30.720 13.610 31.125 ;
        RECT 14.450 30.720 15.910 31.125 ;
        RECT 16.750 30.720 20.510 31.125 ;
        RECT 21.350 30.720 22.810 31.125 ;
        RECT 23.650 30.720 27.410 31.125 ;
        RECT 28.250 30.720 29.710 31.125 ;
        RECT 30.550 30.720 32.010 31.125 ;
        RECT 2.400 4.280 32.560 30.720 ;
        RECT 2.950 3.555 4.410 4.280 ;
        RECT 5.250 3.555 6.710 4.280 ;
        RECT 7.550 3.555 11.310 4.280 ;
        RECT 12.150 3.555 13.610 4.280 ;
        RECT 14.450 3.555 18.210 4.280 ;
        RECT 19.050 3.555 20.510 4.280 ;
        RECT 21.350 3.555 25.110 4.280 ;
        RECT 25.950 3.555 27.410 4.280 ;
        RECT 28.250 3.555 29.710 4.280 ;
        RECT 30.550 3.555 32.560 4.280 ;
      LAYER met3 ;
        RECT 4.400 30.240 31.000 31.105 ;
        RECT 4.000 28.240 31.000 30.240 ;
        RECT 4.400 26.840 30.600 28.240 ;
        RECT 4.000 24.840 31.000 26.840 ;
        RECT 4.000 23.440 30.600 24.840 ;
        RECT 4.000 21.440 31.000 23.440 ;
        RECT 4.400 20.040 31.000 21.440 ;
        RECT 4.000 18.040 31.000 20.040 ;
        RECT 4.400 16.640 30.600 18.040 ;
        RECT 4.000 14.640 31.000 16.640 ;
        RECT 4.000 13.240 30.600 14.640 ;
        RECT 4.000 11.240 31.000 13.240 ;
        RECT 4.400 9.840 31.000 11.240 ;
        RECT 4.000 7.840 31.000 9.840 ;
        RECT 4.400 6.440 30.600 7.840 ;
        RECT 4.000 4.440 31.000 6.440 ;
        RECT 4.000 3.575 30.600 4.440 ;
      LAYER met4 ;
        RECT 10.715 5.200 12.305 27.440 ;
        RECT 14.705 5.200 16.300 27.440 ;
        RECT 18.700 5.200 20.295 27.440 ;
  END
END user_id_programming
END LIBRARY

