.subckt sky130_fd_pr__diode_pd2nw_05v5 A C a=1 p=1
D A C  sky130_fd_pr__diode_pd2nw_05v5 area={a}
.ends
