magic
tech sky130A
magscale 1 2
timestamp 1607107346
<< obsli1 >>
rect 368 17 169556 12971
<< metal1 >>
rect 368 11920 169556 12016
rect 368 11376 169556 11472
<< obsm1 >>
rect 368 12072 169556 12980
rect 368 11528 169556 11864
rect 368 8 169556 11320
<< metal2 >>
rect 754 12200 810 13000
rect 1122 12200 1178 13000
rect 1490 12200 1546 13000
rect 1858 12200 1914 13000
rect 2226 12200 2282 13000
rect 2594 12200 2650 13000
rect 2962 12200 3018 13000
rect 3330 12200 3386 13000
rect 3698 12200 3754 13000
rect 4066 12200 4122 13000
rect 4434 12200 4490 13000
rect 4802 12200 4858 13000
rect 5170 12200 5226 13000
rect 5538 12200 5594 13000
rect 5906 12200 5962 13000
rect 6274 12200 6330 13000
rect 6642 12200 6698 13000
rect 7010 12200 7066 13000
rect 7378 12200 7434 13000
rect 7746 12200 7802 13000
rect 8114 12200 8170 13000
rect 8482 12200 8538 13000
rect 8850 12200 8906 13000
rect 9218 12200 9274 13000
rect 9586 12200 9642 13000
rect 9954 12200 10010 13000
rect 10322 12200 10378 13000
rect 10690 12200 10746 13000
rect 11058 12200 11114 13000
rect 11426 12200 11482 13000
rect 11794 12200 11850 13000
rect 12162 12200 12218 13000
rect 12530 12200 12586 13000
rect 12898 12200 12954 13000
rect 13266 12200 13322 13000
rect 13634 12200 13690 13000
rect 14002 12200 14058 13000
rect 14370 12200 14426 13000
rect 14738 12200 14794 13000
rect 15106 12200 15162 13000
rect 15474 12200 15530 13000
rect 15842 12200 15898 13000
rect 16210 12200 16266 13000
rect 16578 12200 16634 13000
rect 16946 12200 17002 13000
rect 17314 12200 17370 13000
rect 17682 12200 17738 13000
rect 18050 12200 18106 13000
rect 18418 12200 18474 13000
rect 18786 12200 18842 13000
rect 19154 12200 19210 13000
rect 19522 12200 19578 13000
rect 19890 12200 19946 13000
rect 20258 12200 20314 13000
rect 20626 12200 20682 13000
rect 20994 12200 21050 13000
rect 21362 12200 21418 13000
rect 21730 12200 21786 13000
rect 22098 12200 22154 13000
rect 22466 12200 22522 13000
rect 22834 12200 22890 13000
rect 23202 12200 23258 13000
rect 23570 12200 23626 13000
rect 23938 12200 23994 13000
rect 24306 12200 24362 13000
rect 24674 12200 24730 13000
rect 25042 12200 25098 13000
rect 25410 12200 25466 13000
rect 25778 12200 25834 13000
rect 26146 12200 26202 13000
rect 26514 12200 26570 13000
rect 26882 12200 26938 13000
rect 27250 12200 27306 13000
rect 27618 12200 27674 13000
rect 27986 12200 28042 13000
rect 28354 12200 28410 13000
rect 28722 12200 28778 13000
rect 29090 12200 29146 13000
rect 29458 12200 29514 13000
rect 29826 12200 29882 13000
rect 30194 12200 30250 13000
rect 30562 12200 30618 13000
rect 30930 12200 30986 13000
rect 31298 12200 31354 13000
rect 31666 12200 31722 13000
rect 32034 12200 32090 13000
rect 32402 12200 32458 13000
rect 32770 12200 32826 13000
rect 33138 12200 33194 13000
rect 33506 12200 33562 13000
rect 33874 12200 33930 13000
rect 34242 12200 34298 13000
rect 34610 12200 34666 13000
rect 34978 12200 35034 13000
rect 35346 12200 35402 13000
rect 35714 12200 35770 13000
rect 36082 12200 36138 13000
rect 36450 12200 36506 13000
rect 36818 12200 36874 13000
rect 37186 12200 37242 13000
rect 37554 12200 37610 13000
rect 37922 12200 37978 13000
rect 38290 12200 38346 13000
rect 38658 12200 38714 13000
rect 39026 12200 39082 13000
rect 39394 12200 39450 13000
rect 39762 12200 39818 13000
rect 40130 12200 40186 13000
rect 40498 12200 40554 13000
rect 40866 12200 40922 13000
rect 41234 12200 41290 13000
rect 41602 12200 41658 13000
rect 41970 12200 42026 13000
rect 42338 12200 42394 13000
rect 42706 12200 42762 13000
rect 43074 12200 43130 13000
rect 43442 12200 43498 13000
rect 43810 12200 43866 13000
rect 44178 12200 44234 13000
rect 44546 12200 44602 13000
rect 44914 12200 44970 13000
rect 45282 12200 45338 13000
rect 45650 12200 45706 13000
rect 46018 12200 46074 13000
rect 46386 12200 46442 13000
rect 46754 12200 46810 13000
rect 47122 12200 47178 13000
rect 47490 12200 47546 13000
rect 47858 12200 47914 13000
rect 48226 12200 48282 13000
rect 48594 12200 48650 13000
rect 48962 12200 49018 13000
rect 49330 12200 49386 13000
rect 49698 12200 49754 13000
rect 50066 12200 50122 13000
rect 50434 12200 50490 13000
rect 50802 12200 50858 13000
rect 51170 12200 51226 13000
rect 51538 12200 51594 13000
rect 51906 12200 51962 13000
rect 52274 12200 52330 13000
rect 52642 12200 52698 13000
rect 53010 12200 53066 13000
rect 53378 12200 53434 13000
rect 53746 12200 53802 13000
rect 54114 12200 54170 13000
rect 54482 12200 54538 13000
rect 54850 12200 54906 13000
rect 55218 12200 55274 13000
rect 55586 12200 55642 13000
rect 55954 12200 56010 13000
rect 56322 12200 56378 13000
rect 56690 12200 56746 13000
rect 57058 12200 57114 13000
rect 57426 12200 57482 13000
rect 57794 12200 57850 13000
rect 58162 12200 58218 13000
rect 58530 12200 58586 13000
rect 58898 12200 58954 13000
rect 59266 12200 59322 13000
rect 59634 12200 59690 13000
rect 60002 12200 60058 13000
rect 60370 12200 60426 13000
rect 60738 12200 60794 13000
rect 61106 12200 61162 13000
rect 61474 12200 61530 13000
rect 61842 12200 61898 13000
rect 62210 12200 62266 13000
rect 62578 12200 62634 13000
rect 62946 12200 63002 13000
rect 63314 12200 63370 13000
rect 63682 12200 63738 13000
rect 64050 12200 64106 13000
rect 64418 12200 64474 13000
rect 64786 12200 64842 13000
rect 65154 12200 65210 13000
rect 65522 12200 65578 13000
rect 65890 12200 65946 13000
rect 66258 12200 66314 13000
rect 66626 12200 66682 13000
rect 66994 12200 67050 13000
rect 67362 12200 67418 13000
rect 67730 12200 67786 13000
rect 68098 12200 68154 13000
rect 68466 12200 68522 13000
rect 68834 12200 68890 13000
rect 69202 12200 69258 13000
rect 69570 12200 69626 13000
rect 69938 12200 69994 13000
rect 70306 12200 70362 13000
rect 70674 12200 70730 13000
rect 71042 12200 71098 13000
rect 71410 12200 71466 13000
rect 71778 12200 71834 13000
rect 72146 12200 72202 13000
rect 72514 12200 72570 13000
rect 72882 12200 72938 13000
rect 73250 12200 73306 13000
rect 73618 12200 73674 13000
rect 73986 12200 74042 13000
rect 74354 12200 74410 13000
rect 74722 12200 74778 13000
rect 75090 12200 75146 13000
rect 75458 12200 75514 13000
rect 75826 12200 75882 13000
rect 76194 12200 76250 13000
rect 76562 12200 76618 13000
rect 76930 12200 76986 13000
rect 77298 12200 77354 13000
rect 77666 12200 77722 13000
rect 78034 12200 78090 13000
rect 78402 12200 78458 13000
rect 78770 12200 78826 13000
rect 79138 12200 79194 13000
rect 79506 12200 79562 13000
rect 79874 12200 79930 13000
rect 80242 12200 80298 13000
rect 80610 12200 80666 13000
rect 80978 12200 81034 13000
rect 81346 12200 81402 13000
rect 81714 12200 81770 13000
rect 82082 12200 82138 13000
rect 82450 12200 82506 13000
rect 82818 12200 82874 13000
rect 83186 12200 83242 13000
rect 83554 12200 83610 13000
rect 83922 12200 83978 13000
rect 84290 12200 84346 13000
rect 84658 12200 84714 13000
rect 85026 12200 85082 13000
rect 85394 12200 85450 13000
rect 85762 12200 85818 13000
rect 86130 12200 86186 13000
rect 86498 12200 86554 13000
rect 86866 12200 86922 13000
rect 87234 12200 87290 13000
rect 87602 12200 87658 13000
rect 87970 12200 88026 13000
rect 88338 12200 88394 13000
rect 88706 12200 88762 13000
rect 89074 12200 89130 13000
rect 89442 12200 89498 13000
rect 89810 12200 89866 13000
rect 90178 12200 90234 13000
rect 90546 12200 90602 13000
rect 90914 12200 90970 13000
rect 91282 12200 91338 13000
rect 91650 12200 91706 13000
rect 92018 12200 92074 13000
rect 92386 12200 92442 13000
rect 92754 12200 92810 13000
rect 93122 12200 93178 13000
rect 93490 12200 93546 13000
rect 93858 12200 93914 13000
rect 94226 12200 94282 13000
rect 94594 12200 94650 13000
rect 94962 12200 95018 13000
rect 95330 12200 95386 13000
rect 95698 12200 95754 13000
rect 96066 12200 96122 13000
rect 96434 12200 96490 13000
rect 96802 12200 96858 13000
rect 97170 12200 97226 13000
rect 97538 12200 97594 13000
rect 97906 12200 97962 13000
rect 98274 12200 98330 13000
rect 98642 12200 98698 13000
rect 99010 12200 99066 13000
rect 99378 12200 99434 13000
rect 99746 12200 99802 13000
rect 100114 12200 100170 13000
rect 100482 12200 100538 13000
rect 100850 12200 100906 13000
rect 101218 12200 101274 13000
rect 101586 12200 101642 13000
rect 101954 12200 102010 13000
rect 102322 12200 102378 13000
rect 102690 12200 102746 13000
rect 103058 12200 103114 13000
rect 103426 12200 103482 13000
rect 103794 12200 103850 13000
rect 104162 12200 104218 13000
rect 104530 12200 104586 13000
rect 104898 12200 104954 13000
rect 105266 12200 105322 13000
rect 105634 12200 105690 13000
rect 106002 12200 106058 13000
rect 106370 12200 106426 13000
rect 106738 12200 106794 13000
rect 107106 12200 107162 13000
rect 107474 12200 107530 13000
rect 107842 12200 107898 13000
rect 108210 12200 108266 13000
rect 108578 12200 108634 13000
rect 108946 12200 109002 13000
rect 109314 12200 109370 13000
rect 109682 12200 109738 13000
rect 110050 12200 110106 13000
rect 110418 12200 110474 13000
rect 110786 12200 110842 13000
rect 111154 12200 111210 13000
rect 111522 12200 111578 13000
rect 111890 12200 111946 13000
rect 112258 12200 112314 13000
rect 112626 12200 112682 13000
rect 112994 12200 113050 13000
rect 113362 12200 113418 13000
rect 113730 12200 113786 13000
rect 114098 12200 114154 13000
rect 114466 12200 114522 13000
rect 114834 12200 114890 13000
rect 115202 12200 115258 13000
rect 115570 12200 115626 13000
rect 115938 12200 115994 13000
rect 116306 12200 116362 13000
rect 116674 12200 116730 13000
rect 117042 12200 117098 13000
rect 117410 12200 117466 13000
rect 117778 12200 117834 13000
rect 118146 12200 118202 13000
rect 118514 12200 118570 13000
rect 118882 12200 118938 13000
rect 119250 12200 119306 13000
rect 119618 12200 119674 13000
rect 119986 12200 120042 13000
rect 120354 12200 120410 13000
rect 120722 12200 120778 13000
rect 121090 12200 121146 13000
rect 121458 12200 121514 13000
rect 121826 12200 121882 13000
rect 122194 12200 122250 13000
rect 122562 12200 122618 13000
rect 122930 12200 122986 13000
rect 123298 12200 123354 13000
rect 123666 12200 123722 13000
rect 124034 12200 124090 13000
rect 124402 12200 124458 13000
rect 124770 12200 124826 13000
rect 125138 12200 125194 13000
rect 125506 12200 125562 13000
rect 125874 12200 125930 13000
rect 126242 12200 126298 13000
rect 126610 12200 126666 13000
rect 126978 12200 127034 13000
rect 127346 12200 127402 13000
rect 127714 12200 127770 13000
rect 128082 12200 128138 13000
rect 128450 12200 128506 13000
rect 128818 12200 128874 13000
rect 129186 12200 129242 13000
rect 129554 12200 129610 13000
rect 129922 12200 129978 13000
rect 130290 12200 130346 13000
rect 130658 12200 130714 13000
rect 131026 12200 131082 13000
rect 131394 12200 131450 13000
rect 131762 12200 131818 13000
rect 132130 12200 132186 13000
rect 132498 12200 132554 13000
rect 132866 12200 132922 13000
rect 133234 12200 133290 13000
rect 133602 12200 133658 13000
rect 133970 12200 134026 13000
rect 134338 12200 134394 13000
rect 134706 12200 134762 13000
rect 135074 12200 135130 13000
rect 135442 12200 135498 13000
rect 135810 12200 135866 13000
rect 136178 12200 136234 13000
rect 136546 12200 136602 13000
rect 136914 12200 136970 13000
rect 137282 12200 137338 13000
rect 137650 12200 137706 13000
rect 138018 12200 138074 13000
rect 138386 12200 138442 13000
rect 138754 12200 138810 13000
rect 139122 12200 139178 13000
rect 139490 12200 139546 13000
rect 139858 12200 139914 13000
rect 140226 12200 140282 13000
rect 140594 12200 140650 13000
rect 140962 12200 141018 13000
rect 141330 12200 141386 13000
rect 141698 12200 141754 13000
rect 142066 12200 142122 13000
rect 142434 12200 142490 13000
rect 142802 12200 142858 13000
rect 143170 12200 143226 13000
rect 143538 12200 143594 13000
rect 143906 12200 143962 13000
rect 144274 12200 144330 13000
rect 144642 12200 144698 13000
rect 145010 12200 145066 13000
rect 145378 12200 145434 13000
rect 145746 12200 145802 13000
rect 146114 12200 146170 13000
rect 146482 12200 146538 13000
rect 146850 12200 146906 13000
rect 147218 12200 147274 13000
rect 147586 12200 147642 13000
rect 147954 12200 148010 13000
rect 148322 12200 148378 13000
rect 148690 12200 148746 13000
rect 149058 12200 149114 13000
rect 149426 12200 149482 13000
rect 149794 12200 149850 13000
rect 150162 12200 150218 13000
rect 150530 12200 150586 13000
rect 150898 12200 150954 13000
rect 151266 12200 151322 13000
rect 151634 12200 151690 13000
rect 152002 12200 152058 13000
rect 152370 12200 152426 13000
rect 152738 12200 152794 13000
rect 153106 12200 153162 13000
rect 153474 12200 153530 13000
rect 153842 12200 153898 13000
rect 154210 12200 154266 13000
rect 154578 12200 154634 13000
rect 154946 12200 155002 13000
rect 155314 12200 155370 13000
rect 155682 12200 155738 13000
rect 156050 12200 156106 13000
rect 156418 12200 156474 13000
rect 156786 12200 156842 13000
rect 157154 12200 157210 13000
rect 157522 12200 157578 13000
rect 157890 12200 157946 13000
rect 158258 12200 158314 13000
rect 158626 12200 158682 13000
rect 158994 12200 159050 13000
rect 159362 12200 159418 13000
rect 159730 12200 159786 13000
rect 160098 12200 160154 13000
rect 160466 12200 160522 13000
rect 160834 12200 160890 13000
rect 161202 12200 161258 13000
rect 161570 12200 161626 13000
rect 161938 12200 161994 13000
rect 162306 12200 162362 13000
rect 162674 12200 162730 13000
rect 163042 12200 163098 13000
rect 163410 12200 163466 13000
rect 163778 12200 163834 13000
rect 164146 12200 164202 13000
rect 164514 12200 164570 13000
rect 164882 12200 164938 13000
rect 570 0 626 800
rect 754 0 810 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 34058 0 34114 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 37002 0 37058 800
rect 37370 0 37426 800
rect 37738 0 37794 800
rect 38106 0 38162 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42522 0 42578 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43994 0 44050 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46202 0 46258 800
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47306 0 47362 800
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49146 0 49202 800
rect 49514 0 49570 800
rect 49882 0 49938 800
rect 50250 0 50306 800
rect 50618 0 50674 800
rect 50986 0 51042 800
rect 51354 0 51410 800
rect 51722 0 51778 800
rect 52090 0 52146 800
rect 52458 0 52514 800
rect 52826 0 52882 800
rect 53194 0 53250 800
rect 53562 0 53618 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54666 0 54722 800
rect 55034 0 55090 800
rect 55402 0 55458 800
rect 55770 0 55826 800
rect 56138 0 56194 800
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 57242 0 57298 800
rect 57610 0 57666 800
rect 57978 0 58034 800
rect 58346 0 58402 800
rect 58714 0 58770 800
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59818 0 59874 800
rect 60186 0 60242 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61290 0 61346 800
rect 61658 0 61714 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64602 0 64658 800
rect 64970 0 65026 800
rect 65338 0 65394 800
rect 65706 0 65762 800
rect 66074 0 66130 800
rect 66442 0 66498 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68282 0 68338 800
rect 68650 0 68706 800
rect 69018 0 69074 800
rect 69386 0 69442 800
rect 69754 0 69810 800
rect 70122 0 70178 800
rect 70490 0 70546 800
rect 70858 0 70914 800
rect 71226 0 71282 800
rect 71594 0 71650 800
rect 71962 0 72018 800
rect 72330 0 72386 800
rect 72698 0 72754 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73802 0 73858 800
rect 74170 0 74226 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75274 0 75330 800
rect 75642 0 75698 800
rect 76010 0 76066 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77114 0 77170 800
rect 77482 0 77538 800
rect 77850 0 77906 800
rect 78218 0 78274 800
rect 78586 0 78642 800
rect 78954 0 79010 800
rect 79322 0 79378 800
rect 79690 0 79746 800
rect 80058 0 80114 800
rect 80426 0 80482 800
rect 80794 0 80850 800
rect 81162 0 81218 800
rect 81530 0 81586 800
rect 81898 0 81954 800
rect 82266 0 82322 800
rect 82634 0 82690 800
rect 83002 0 83058 800
rect 83370 0 83426 800
rect 83738 0 83794 800
rect 84106 0 84162 800
rect 84474 0 84530 800
rect 84842 0 84898 800
rect 85210 0 85266 800
rect 85578 0 85634 800
rect 85946 0 86002 800
rect 86314 0 86370 800
rect 86682 0 86738 800
rect 87050 0 87106 800
rect 87418 0 87474 800
rect 87786 0 87842 800
rect 88154 0 88210 800
rect 88522 0 88578 800
rect 88890 0 88946 800
rect 89258 0 89314 800
rect 89626 0 89682 800
rect 89994 0 90050 800
rect 90362 0 90418 800
rect 90730 0 90786 800
rect 91098 0 91154 800
rect 91466 0 91522 800
rect 91834 0 91890 800
rect 92202 0 92258 800
rect 92570 0 92626 800
rect 92938 0 92994 800
rect 93306 0 93362 800
rect 93674 0 93730 800
rect 94042 0 94098 800
rect 94410 0 94466 800
rect 94778 0 94834 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96618 0 96674 800
rect 96986 0 97042 800
rect 97354 0 97410 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98458 0 98514 800
rect 98826 0 98882 800
rect 99194 0 99250 800
rect 99562 0 99618 800
rect 99930 0 99986 800
rect 100298 0 100354 800
rect 100666 0 100722 800
rect 101034 0 101090 800
rect 101402 0 101458 800
rect 101770 0 101826 800
rect 102138 0 102194 800
rect 102506 0 102562 800
rect 102874 0 102930 800
rect 103242 0 103298 800
rect 103610 0 103666 800
rect 103978 0 104034 800
rect 104346 0 104402 800
rect 104714 0 104770 800
rect 105082 0 105138 800
rect 105450 0 105506 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106554 0 106610 800
rect 106922 0 106978 800
rect 107290 0 107346 800
rect 107658 0 107714 800
rect 108026 0 108082 800
rect 108394 0 108450 800
rect 108762 0 108818 800
rect 109130 0 109186 800
rect 109498 0 109554 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 110970 0 111026 800
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 112074 0 112130 800
rect 112442 0 112498 800
rect 112810 0 112866 800
rect 113178 0 113234 800
rect 113546 0 113602 800
rect 113914 0 113970 800
rect 114282 0 114338 800
rect 114650 0 114706 800
rect 115018 0 115074 800
rect 115386 0 115442 800
rect 115754 0 115810 800
rect 116122 0 116178 800
rect 116490 0 116546 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117594 0 117650 800
rect 117962 0 118018 800
rect 118330 0 118386 800
rect 118698 0 118754 800
rect 119066 0 119122 800
rect 119434 0 119490 800
rect 119802 0 119858 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120906 0 120962 800
rect 121274 0 121330 800
rect 121642 0 121698 800
rect 122010 0 122066 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123850 0 123906 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126794 0 126850 800
rect 127162 0 127218 800
rect 127530 0 127586 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131578 0 131634 800
rect 131946 0 132002 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134154 0 134210 800
rect 134522 0 134578 800
rect 134890 0 134946 800
rect 135258 0 135314 800
rect 135626 0 135682 800
rect 135994 0 136050 800
rect 136362 0 136418 800
rect 136730 0 136786 800
rect 137098 0 137154 800
rect 137466 0 137522 800
rect 137834 0 137890 800
rect 138202 0 138258 800
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139306 0 139362 800
rect 139674 0 139730 800
rect 140042 0 140098 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141146 0 141202 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142618 0 142674 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143722 0 143778 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 145930 0 145986 800
rect 146298 0 146354 800
rect 146666 0 146722 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148874 0 148930 800
rect 149242 0 149298 800
rect 149610 0 149666 800
rect 149978 0 150034 800
rect 150346 0 150402 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151450 0 151506 800
rect 151818 0 151874 800
rect 152186 0 152242 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153658 0 153714 800
rect 154026 0 154082 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165802 0 165858 800
rect 166170 0 166226 800
rect 166538 0 166594 800
<< obsm2 >>
rect 572 12144 698 13025
rect 866 12144 1066 13025
rect 1234 12144 1434 13025
rect 1602 12144 1802 13025
rect 1970 12144 2170 13025
rect 2338 12144 2538 13025
rect 2706 12144 2906 13025
rect 3074 12144 3274 13025
rect 3442 12144 3642 13025
rect 3810 12144 4010 13025
rect 4178 12144 4378 13025
rect 4546 12144 4746 13025
rect 4914 12144 5114 13025
rect 5282 12144 5482 13025
rect 5650 12144 5850 13025
rect 6018 12144 6218 13025
rect 6386 12144 6586 13025
rect 6754 12144 6954 13025
rect 7122 12144 7322 13025
rect 7490 12144 7690 13025
rect 7858 12144 8058 13025
rect 8226 12144 8426 13025
rect 8594 12144 8794 13025
rect 8962 12144 9162 13025
rect 9330 12144 9530 13025
rect 9698 12144 9898 13025
rect 10066 12144 10266 13025
rect 10434 12144 10634 13025
rect 10802 12144 11002 13025
rect 11170 12144 11370 13025
rect 11538 12144 11738 13025
rect 11906 12144 12106 13025
rect 12274 12144 12474 13025
rect 12642 12144 12842 13025
rect 13010 12144 13210 13025
rect 13378 12144 13578 13025
rect 13746 12144 13946 13025
rect 14114 12144 14314 13025
rect 14482 12144 14682 13025
rect 14850 12144 15050 13025
rect 15218 12144 15418 13025
rect 15586 12144 15786 13025
rect 15954 12144 16154 13025
rect 16322 12144 16522 13025
rect 16690 12144 16890 13025
rect 17058 12144 17258 13025
rect 17426 12144 17626 13025
rect 17794 12144 17994 13025
rect 18162 12144 18362 13025
rect 18530 12144 18730 13025
rect 18898 12144 19098 13025
rect 19266 12144 19466 13025
rect 19634 12144 19834 13025
rect 20002 12144 20202 13025
rect 20370 12144 20570 13025
rect 20738 12144 20938 13025
rect 21106 12144 21306 13025
rect 21474 12144 21674 13025
rect 21842 12144 22042 13025
rect 22210 12144 22410 13025
rect 22578 12144 22778 13025
rect 22946 12144 23146 13025
rect 23314 12144 23514 13025
rect 23682 12144 23882 13025
rect 24050 12144 24250 13025
rect 24418 12144 24618 13025
rect 24786 12144 24986 13025
rect 25154 12144 25354 13025
rect 25522 12144 25722 13025
rect 25890 12144 26090 13025
rect 26258 12144 26458 13025
rect 26626 12144 26826 13025
rect 26994 12144 27194 13025
rect 27362 12144 27562 13025
rect 27730 12144 27930 13025
rect 28098 12144 28298 13025
rect 28466 12144 28666 13025
rect 28834 12144 29034 13025
rect 29202 12144 29402 13025
rect 29570 12144 29770 13025
rect 29938 12144 30138 13025
rect 30306 12144 30506 13025
rect 30674 12144 30874 13025
rect 31042 12144 31242 13025
rect 31410 12144 31610 13025
rect 31778 12144 31978 13025
rect 32146 12144 32346 13025
rect 32514 12144 32714 13025
rect 32882 12144 33082 13025
rect 33250 12144 33450 13025
rect 33618 12144 33818 13025
rect 33986 12144 34186 13025
rect 34354 12144 34554 13025
rect 34722 12144 34922 13025
rect 35090 12144 35290 13025
rect 35458 12144 35658 13025
rect 35826 12144 36026 13025
rect 36194 12144 36394 13025
rect 36562 12144 36762 13025
rect 36930 12144 37130 13025
rect 37298 12144 37498 13025
rect 37666 12144 37866 13025
rect 38034 12144 38234 13025
rect 38402 12144 38602 13025
rect 38770 12144 38970 13025
rect 39138 12144 39338 13025
rect 39506 12144 39706 13025
rect 39874 12144 40074 13025
rect 40242 12144 40442 13025
rect 40610 12144 40810 13025
rect 40978 12144 41178 13025
rect 41346 12144 41546 13025
rect 41714 12144 41914 13025
rect 42082 12144 42282 13025
rect 42450 12144 42650 13025
rect 42818 12144 43018 13025
rect 43186 12144 43386 13025
rect 43554 12144 43754 13025
rect 43922 12144 44122 13025
rect 44290 12144 44490 13025
rect 44658 12144 44858 13025
rect 45026 12144 45226 13025
rect 45394 12144 45594 13025
rect 45762 12144 45962 13025
rect 46130 12144 46330 13025
rect 46498 12144 46698 13025
rect 46866 12144 47066 13025
rect 47234 12144 47434 13025
rect 47602 12144 47802 13025
rect 47970 12144 48170 13025
rect 48338 12144 48538 13025
rect 48706 12144 48906 13025
rect 49074 12144 49274 13025
rect 49442 12144 49642 13025
rect 49810 12144 50010 13025
rect 50178 12144 50378 13025
rect 50546 12144 50746 13025
rect 50914 12144 51114 13025
rect 51282 12144 51482 13025
rect 51650 12144 51850 13025
rect 52018 12144 52218 13025
rect 52386 12144 52586 13025
rect 52754 12144 52954 13025
rect 53122 12144 53322 13025
rect 53490 12144 53690 13025
rect 53858 12144 54058 13025
rect 54226 12144 54426 13025
rect 54594 12144 54794 13025
rect 54962 12144 55162 13025
rect 55330 12144 55530 13025
rect 55698 12144 55898 13025
rect 56066 12144 56266 13025
rect 56434 12144 56634 13025
rect 56802 12144 57002 13025
rect 57170 12144 57370 13025
rect 57538 12144 57738 13025
rect 57906 12144 58106 13025
rect 58274 12144 58474 13025
rect 58642 12144 58842 13025
rect 59010 12144 59210 13025
rect 59378 12144 59578 13025
rect 59746 12144 59946 13025
rect 60114 12144 60314 13025
rect 60482 12144 60682 13025
rect 60850 12144 61050 13025
rect 61218 12144 61418 13025
rect 61586 12144 61786 13025
rect 61954 12144 62154 13025
rect 62322 12144 62522 13025
rect 62690 12144 62890 13025
rect 63058 12144 63258 13025
rect 63426 12144 63626 13025
rect 63794 12144 63994 13025
rect 64162 12144 64362 13025
rect 64530 12144 64730 13025
rect 64898 12144 65098 13025
rect 65266 12144 65466 13025
rect 65634 12144 65834 13025
rect 66002 12144 66202 13025
rect 66370 12144 66570 13025
rect 66738 12144 66938 13025
rect 67106 12144 67306 13025
rect 67474 12144 67674 13025
rect 67842 12144 68042 13025
rect 68210 12144 68410 13025
rect 68578 12144 68778 13025
rect 68946 12144 69146 13025
rect 69314 12144 69514 13025
rect 69682 12144 69882 13025
rect 70050 12144 70250 13025
rect 70418 12144 70618 13025
rect 70786 12144 70986 13025
rect 71154 12144 71354 13025
rect 71522 12144 71722 13025
rect 71890 12144 72090 13025
rect 72258 12144 72458 13025
rect 72626 12144 72826 13025
rect 72994 12144 73194 13025
rect 73362 12144 73562 13025
rect 73730 12144 73930 13025
rect 74098 12144 74298 13025
rect 74466 12144 74666 13025
rect 74834 12144 75034 13025
rect 75202 12144 75402 13025
rect 75570 12144 75770 13025
rect 75938 12144 76138 13025
rect 76306 12144 76506 13025
rect 76674 12144 76874 13025
rect 77042 12144 77242 13025
rect 77410 12144 77610 13025
rect 77778 12144 77978 13025
rect 78146 12144 78346 13025
rect 78514 12144 78714 13025
rect 78882 12144 79082 13025
rect 79250 12144 79450 13025
rect 79618 12144 79818 13025
rect 79986 12144 80186 13025
rect 80354 12144 80554 13025
rect 80722 12144 80922 13025
rect 81090 12144 81290 13025
rect 81458 12144 81658 13025
rect 81826 12144 82026 13025
rect 82194 12144 82394 13025
rect 82562 12144 82762 13025
rect 82930 12144 83130 13025
rect 83298 12144 83498 13025
rect 83666 12144 83866 13025
rect 84034 12144 84234 13025
rect 84402 12144 84602 13025
rect 84770 12144 84970 13025
rect 85138 12144 85338 13025
rect 85506 12144 85706 13025
rect 85874 12144 86074 13025
rect 86242 12144 86442 13025
rect 86610 12144 86810 13025
rect 86978 12144 87178 13025
rect 87346 12144 87546 13025
rect 87714 12144 87914 13025
rect 88082 12144 88282 13025
rect 88450 12144 88650 13025
rect 88818 12144 89018 13025
rect 89186 12144 89386 13025
rect 89554 12144 89754 13025
rect 89922 12144 90122 13025
rect 90290 12144 90490 13025
rect 90658 12144 90858 13025
rect 91026 12144 91226 13025
rect 91394 12144 91594 13025
rect 91762 12144 91962 13025
rect 92130 12144 92330 13025
rect 92498 12144 92698 13025
rect 92866 12144 93066 13025
rect 93234 12144 93434 13025
rect 93602 12144 93802 13025
rect 93970 12144 94170 13025
rect 94338 12144 94538 13025
rect 94706 12144 94906 13025
rect 95074 12144 95274 13025
rect 95442 12144 95642 13025
rect 95810 12144 96010 13025
rect 96178 12144 96378 13025
rect 96546 12144 96746 13025
rect 96914 12144 97114 13025
rect 97282 12144 97482 13025
rect 97650 12144 97850 13025
rect 98018 12144 98218 13025
rect 98386 12144 98586 13025
rect 98754 12144 98954 13025
rect 99122 12144 99322 13025
rect 99490 12144 99690 13025
rect 99858 12144 100058 13025
rect 100226 12144 100426 13025
rect 100594 12144 100794 13025
rect 100962 12144 101162 13025
rect 101330 12144 101530 13025
rect 101698 12144 101898 13025
rect 102066 12144 102266 13025
rect 102434 12144 102634 13025
rect 102802 12144 103002 13025
rect 103170 12144 103370 13025
rect 103538 12144 103738 13025
rect 103906 12144 104106 13025
rect 104274 12144 104474 13025
rect 104642 12144 104842 13025
rect 105010 12144 105210 13025
rect 105378 12144 105578 13025
rect 105746 12144 105946 13025
rect 106114 12144 106314 13025
rect 106482 12144 106682 13025
rect 106850 12144 107050 13025
rect 107218 12144 107418 13025
rect 107586 12144 107786 13025
rect 107954 12144 108154 13025
rect 108322 12144 108522 13025
rect 108690 12144 108890 13025
rect 109058 12144 109258 13025
rect 109426 12144 109626 13025
rect 109794 12144 109994 13025
rect 110162 12144 110362 13025
rect 110530 12144 110730 13025
rect 110898 12144 111098 13025
rect 111266 12144 111466 13025
rect 111634 12144 111834 13025
rect 112002 12144 112202 13025
rect 112370 12144 112570 13025
rect 112738 12144 112938 13025
rect 113106 12144 113306 13025
rect 113474 12144 113674 13025
rect 113842 12144 114042 13025
rect 114210 12144 114410 13025
rect 114578 12144 114778 13025
rect 114946 12144 115146 13025
rect 115314 12144 115514 13025
rect 115682 12144 115882 13025
rect 116050 12144 116250 13025
rect 116418 12144 116618 13025
rect 116786 12144 116986 13025
rect 117154 12144 117354 13025
rect 117522 12144 117722 13025
rect 117890 12144 118090 13025
rect 118258 12144 118458 13025
rect 118626 12144 118826 13025
rect 118994 12144 119194 13025
rect 119362 12144 119562 13025
rect 119730 12144 119930 13025
rect 120098 12144 120298 13025
rect 120466 12144 120666 13025
rect 120834 12144 121034 13025
rect 121202 12144 121402 13025
rect 121570 12144 121770 13025
rect 121938 12144 122138 13025
rect 122306 12144 122506 13025
rect 122674 12144 122874 13025
rect 123042 12144 123242 13025
rect 123410 12144 123610 13025
rect 123778 12144 123978 13025
rect 124146 12144 124346 13025
rect 124514 12144 124714 13025
rect 124882 12144 125082 13025
rect 125250 12144 125450 13025
rect 125618 12144 125818 13025
rect 125986 12144 126186 13025
rect 126354 12144 126554 13025
rect 126722 12144 126922 13025
rect 127090 12144 127290 13025
rect 127458 12144 127658 13025
rect 127826 12144 128026 13025
rect 128194 12144 128394 13025
rect 128562 12144 128762 13025
rect 128930 12144 129130 13025
rect 129298 12144 129498 13025
rect 129666 12144 129866 13025
rect 130034 12144 130234 13025
rect 130402 12144 130602 13025
rect 130770 12144 130970 13025
rect 131138 12144 131338 13025
rect 131506 12144 131706 13025
rect 131874 12144 132074 13025
rect 132242 12144 132442 13025
rect 132610 12144 132810 13025
rect 132978 12144 133178 13025
rect 133346 12144 133546 13025
rect 133714 12144 133914 13025
rect 134082 12144 134282 13025
rect 134450 12144 134650 13025
rect 134818 12144 135018 13025
rect 135186 12144 135386 13025
rect 135554 12144 135754 13025
rect 135922 12144 136122 13025
rect 136290 12144 136490 13025
rect 136658 12144 136858 13025
rect 137026 12144 137226 13025
rect 137394 12144 137594 13025
rect 137762 12144 137962 13025
rect 138130 12144 138330 13025
rect 138498 12144 138698 13025
rect 138866 12144 139066 13025
rect 139234 12144 139434 13025
rect 139602 12144 139802 13025
rect 139970 12144 140170 13025
rect 140338 12144 140538 13025
rect 140706 12144 140906 13025
rect 141074 12144 141274 13025
rect 141442 12144 141642 13025
rect 141810 12144 142010 13025
rect 142178 12144 142378 13025
rect 142546 12144 142746 13025
rect 142914 12144 143114 13025
rect 143282 12144 143482 13025
rect 143650 12144 143850 13025
rect 144018 12144 144218 13025
rect 144386 12144 144586 13025
rect 144754 12144 144954 13025
rect 145122 12144 145322 13025
rect 145490 12144 145690 13025
rect 145858 12144 146058 13025
rect 146226 12144 146426 13025
rect 146594 12144 146794 13025
rect 146962 12144 147162 13025
rect 147330 12144 147530 13025
rect 147698 12144 147898 13025
rect 148066 12144 148266 13025
rect 148434 12144 148634 13025
rect 148802 12144 149002 13025
rect 149170 12144 149370 13025
rect 149538 12144 149738 13025
rect 149906 12144 150106 13025
rect 150274 12144 150474 13025
rect 150642 12144 150842 13025
rect 151010 12144 151210 13025
rect 151378 12144 151578 13025
rect 151746 12144 151946 13025
rect 152114 12144 152314 13025
rect 152482 12144 152682 13025
rect 152850 12144 153050 13025
rect 153218 12144 153418 13025
rect 153586 12144 153786 13025
rect 153954 12144 154154 13025
rect 154322 12144 154522 13025
rect 154690 12144 154890 13025
rect 155058 12144 155258 13025
rect 155426 12144 155626 13025
rect 155794 12144 155994 13025
rect 156162 12144 156362 13025
rect 156530 12144 156730 13025
rect 156898 12144 157098 13025
rect 157266 12144 157466 13025
rect 157634 12144 157834 13025
rect 158002 12144 158202 13025
rect 158370 12144 158570 13025
rect 158738 12144 158938 13025
rect 159106 12144 159306 13025
rect 159474 12144 159674 13025
rect 159842 12144 160042 13025
rect 160210 12144 160410 13025
rect 160578 12144 160778 13025
rect 160946 12144 161146 13025
rect 161314 12144 161514 13025
rect 161682 12144 161882 13025
rect 162050 12144 162250 13025
rect 162418 12144 162618 13025
rect 162786 12144 162986 13025
rect 163154 12144 163354 13025
rect 163522 12144 163722 13025
rect 163890 12144 164090 13025
rect 164258 12144 164458 13025
rect 164626 12144 164826 13025
rect 164994 12144 167236 13025
rect 572 856 167236 12144
rect 682 2 698 856
rect 866 2 882 856
rect 1050 2 1250 856
rect 1418 2 1618 856
rect 1786 2 1986 856
rect 2154 2 2354 856
rect 2522 2 2722 856
rect 2890 2 3090 856
rect 3258 2 3458 856
rect 3626 2 3826 856
rect 3994 2 4194 856
rect 4362 2 4562 856
rect 4730 2 4930 856
rect 5098 2 5298 856
rect 5466 2 5666 856
rect 5834 2 6034 856
rect 6202 2 6402 856
rect 6570 2 6770 856
rect 6938 2 7138 856
rect 7306 2 7506 856
rect 7674 2 7874 856
rect 8042 2 8242 856
rect 8410 2 8610 856
rect 8778 2 8978 856
rect 9146 2 9346 856
rect 9514 2 9714 856
rect 9882 2 10082 856
rect 10250 2 10450 856
rect 10618 2 10818 856
rect 10986 2 11186 856
rect 11354 2 11554 856
rect 11722 2 11922 856
rect 12090 2 12290 856
rect 12458 2 12658 856
rect 12826 2 13026 856
rect 13194 2 13394 856
rect 13562 2 13762 856
rect 13930 2 14130 856
rect 14298 2 14498 856
rect 14666 2 14866 856
rect 15034 2 15234 856
rect 15402 2 15602 856
rect 15770 2 15970 856
rect 16138 2 16338 856
rect 16506 2 16706 856
rect 16874 2 17074 856
rect 17242 2 17442 856
rect 17610 2 17810 856
rect 17978 2 18178 856
rect 18346 2 18546 856
rect 18714 2 18914 856
rect 19082 2 19282 856
rect 19450 2 19650 856
rect 19818 2 20018 856
rect 20186 2 20386 856
rect 20554 2 20754 856
rect 20922 2 21122 856
rect 21290 2 21490 856
rect 21658 2 21858 856
rect 22026 2 22226 856
rect 22394 2 22594 856
rect 22762 2 22962 856
rect 23130 2 23330 856
rect 23498 2 23698 856
rect 23866 2 24066 856
rect 24234 2 24434 856
rect 24602 2 24802 856
rect 24970 2 25170 856
rect 25338 2 25538 856
rect 25706 2 25906 856
rect 26074 2 26274 856
rect 26442 2 26642 856
rect 26810 2 27010 856
rect 27178 2 27378 856
rect 27546 2 27746 856
rect 27914 2 28114 856
rect 28282 2 28482 856
rect 28650 2 28850 856
rect 29018 2 29218 856
rect 29386 2 29586 856
rect 29754 2 29954 856
rect 30122 2 30322 856
rect 30490 2 30690 856
rect 30858 2 31058 856
rect 31226 2 31426 856
rect 31594 2 31794 856
rect 31962 2 32162 856
rect 32330 2 32530 856
rect 32698 2 32898 856
rect 33066 2 33266 856
rect 33434 2 33634 856
rect 33802 2 34002 856
rect 34170 2 34370 856
rect 34538 2 34738 856
rect 34906 2 35106 856
rect 35274 2 35474 856
rect 35642 2 35842 856
rect 36010 2 36210 856
rect 36378 2 36578 856
rect 36746 2 36946 856
rect 37114 2 37314 856
rect 37482 2 37682 856
rect 37850 2 38050 856
rect 38218 2 38418 856
rect 38586 2 38786 856
rect 38954 2 39154 856
rect 39322 2 39522 856
rect 39690 2 39890 856
rect 40058 2 40258 856
rect 40426 2 40626 856
rect 40794 2 40994 856
rect 41162 2 41362 856
rect 41530 2 41730 856
rect 41898 2 42098 856
rect 42266 2 42466 856
rect 42634 2 42834 856
rect 43002 2 43202 856
rect 43370 2 43570 856
rect 43738 2 43938 856
rect 44106 2 44306 856
rect 44474 2 44674 856
rect 44842 2 45042 856
rect 45210 2 45410 856
rect 45578 2 45778 856
rect 45946 2 46146 856
rect 46314 2 46514 856
rect 46682 2 46882 856
rect 47050 2 47250 856
rect 47418 2 47618 856
rect 47786 2 47986 856
rect 48154 2 48354 856
rect 48522 2 48722 856
rect 48890 2 49090 856
rect 49258 2 49458 856
rect 49626 2 49826 856
rect 49994 2 50194 856
rect 50362 2 50562 856
rect 50730 2 50930 856
rect 51098 2 51298 856
rect 51466 2 51666 856
rect 51834 2 52034 856
rect 52202 2 52402 856
rect 52570 2 52770 856
rect 52938 2 53138 856
rect 53306 2 53506 856
rect 53674 2 53874 856
rect 54042 2 54242 856
rect 54410 2 54610 856
rect 54778 2 54978 856
rect 55146 2 55346 856
rect 55514 2 55714 856
rect 55882 2 56082 856
rect 56250 2 56450 856
rect 56618 2 56818 856
rect 56986 2 57186 856
rect 57354 2 57554 856
rect 57722 2 57922 856
rect 58090 2 58290 856
rect 58458 2 58658 856
rect 58826 2 59026 856
rect 59194 2 59394 856
rect 59562 2 59762 856
rect 59930 2 60130 856
rect 60298 2 60498 856
rect 60666 2 60866 856
rect 61034 2 61234 856
rect 61402 2 61602 856
rect 61770 2 61970 856
rect 62138 2 62338 856
rect 62506 2 62706 856
rect 62874 2 63074 856
rect 63242 2 63442 856
rect 63610 2 63810 856
rect 63978 2 64178 856
rect 64346 2 64546 856
rect 64714 2 64914 856
rect 65082 2 65282 856
rect 65450 2 65650 856
rect 65818 2 66018 856
rect 66186 2 66386 856
rect 66554 2 66754 856
rect 66922 2 67122 856
rect 67290 2 67490 856
rect 67658 2 67858 856
rect 68026 2 68226 856
rect 68394 2 68594 856
rect 68762 2 68962 856
rect 69130 2 69330 856
rect 69498 2 69698 856
rect 69866 2 70066 856
rect 70234 2 70434 856
rect 70602 2 70802 856
rect 70970 2 71170 856
rect 71338 2 71538 856
rect 71706 2 71906 856
rect 72074 2 72274 856
rect 72442 2 72642 856
rect 72810 2 73010 856
rect 73178 2 73378 856
rect 73546 2 73746 856
rect 73914 2 74114 856
rect 74282 2 74482 856
rect 74650 2 74850 856
rect 75018 2 75218 856
rect 75386 2 75586 856
rect 75754 2 75954 856
rect 76122 2 76322 856
rect 76490 2 76690 856
rect 76858 2 77058 856
rect 77226 2 77426 856
rect 77594 2 77794 856
rect 77962 2 78162 856
rect 78330 2 78530 856
rect 78698 2 78898 856
rect 79066 2 79266 856
rect 79434 2 79634 856
rect 79802 2 80002 856
rect 80170 2 80370 856
rect 80538 2 80738 856
rect 80906 2 81106 856
rect 81274 2 81474 856
rect 81642 2 81842 856
rect 82010 2 82210 856
rect 82378 2 82578 856
rect 82746 2 82946 856
rect 83114 2 83314 856
rect 83482 2 83682 856
rect 83850 2 84050 856
rect 84218 2 84418 856
rect 84586 2 84786 856
rect 84954 2 85154 856
rect 85322 2 85522 856
rect 85690 2 85890 856
rect 86058 2 86258 856
rect 86426 2 86626 856
rect 86794 2 86994 856
rect 87162 2 87362 856
rect 87530 2 87730 856
rect 87898 2 88098 856
rect 88266 2 88466 856
rect 88634 2 88834 856
rect 89002 2 89202 856
rect 89370 2 89570 856
rect 89738 2 89938 856
rect 90106 2 90306 856
rect 90474 2 90674 856
rect 90842 2 91042 856
rect 91210 2 91410 856
rect 91578 2 91778 856
rect 91946 2 92146 856
rect 92314 2 92514 856
rect 92682 2 92882 856
rect 93050 2 93250 856
rect 93418 2 93618 856
rect 93786 2 93986 856
rect 94154 2 94354 856
rect 94522 2 94722 856
rect 94890 2 95090 856
rect 95258 2 95458 856
rect 95626 2 95826 856
rect 95994 2 96194 856
rect 96362 2 96562 856
rect 96730 2 96930 856
rect 97098 2 97298 856
rect 97466 2 97666 856
rect 97834 2 98034 856
rect 98202 2 98402 856
rect 98570 2 98770 856
rect 98938 2 99138 856
rect 99306 2 99506 856
rect 99674 2 99874 856
rect 100042 2 100242 856
rect 100410 2 100610 856
rect 100778 2 100978 856
rect 101146 2 101346 856
rect 101514 2 101714 856
rect 101882 2 102082 856
rect 102250 2 102450 856
rect 102618 2 102818 856
rect 102986 2 103186 856
rect 103354 2 103554 856
rect 103722 2 103922 856
rect 104090 2 104290 856
rect 104458 2 104658 856
rect 104826 2 105026 856
rect 105194 2 105394 856
rect 105562 2 105762 856
rect 105930 2 106130 856
rect 106298 2 106498 856
rect 106666 2 106866 856
rect 107034 2 107234 856
rect 107402 2 107602 856
rect 107770 2 107970 856
rect 108138 2 108338 856
rect 108506 2 108706 856
rect 108874 2 109074 856
rect 109242 2 109442 856
rect 109610 2 109810 856
rect 109978 2 110178 856
rect 110346 2 110546 856
rect 110714 2 110914 856
rect 111082 2 111282 856
rect 111450 2 111650 856
rect 111818 2 112018 856
rect 112186 2 112386 856
rect 112554 2 112754 856
rect 112922 2 113122 856
rect 113290 2 113490 856
rect 113658 2 113858 856
rect 114026 2 114226 856
rect 114394 2 114594 856
rect 114762 2 114962 856
rect 115130 2 115330 856
rect 115498 2 115698 856
rect 115866 2 116066 856
rect 116234 2 116434 856
rect 116602 2 116802 856
rect 116970 2 117170 856
rect 117338 2 117538 856
rect 117706 2 117906 856
rect 118074 2 118274 856
rect 118442 2 118642 856
rect 118810 2 119010 856
rect 119178 2 119378 856
rect 119546 2 119746 856
rect 119914 2 120114 856
rect 120282 2 120482 856
rect 120650 2 120850 856
rect 121018 2 121218 856
rect 121386 2 121586 856
rect 121754 2 121954 856
rect 122122 2 122322 856
rect 122490 2 122690 856
rect 122858 2 123058 856
rect 123226 2 123426 856
rect 123594 2 123794 856
rect 123962 2 124162 856
rect 124330 2 124530 856
rect 124698 2 124898 856
rect 125066 2 125266 856
rect 125434 2 125634 856
rect 125802 2 126002 856
rect 126170 2 126370 856
rect 126538 2 126738 856
rect 126906 2 127106 856
rect 127274 2 127474 856
rect 127642 2 127842 856
rect 128010 2 128210 856
rect 128378 2 128578 856
rect 128746 2 128946 856
rect 129114 2 129314 856
rect 129482 2 129682 856
rect 129850 2 130050 856
rect 130218 2 130418 856
rect 130586 2 130786 856
rect 130954 2 131154 856
rect 131322 2 131522 856
rect 131690 2 131890 856
rect 132058 2 132258 856
rect 132426 2 132626 856
rect 132794 2 132994 856
rect 133162 2 133362 856
rect 133530 2 133730 856
rect 133898 2 134098 856
rect 134266 2 134466 856
rect 134634 2 134834 856
rect 135002 2 135202 856
rect 135370 2 135570 856
rect 135738 2 135938 856
rect 136106 2 136306 856
rect 136474 2 136674 856
rect 136842 2 137042 856
rect 137210 2 137410 856
rect 137578 2 137778 856
rect 137946 2 138146 856
rect 138314 2 138514 856
rect 138682 2 138882 856
rect 139050 2 139250 856
rect 139418 2 139618 856
rect 139786 2 139986 856
rect 140154 2 140354 856
rect 140522 2 140722 856
rect 140890 2 141090 856
rect 141258 2 141458 856
rect 141626 2 141826 856
rect 141994 2 142194 856
rect 142362 2 142562 856
rect 142730 2 142930 856
rect 143098 2 143298 856
rect 143466 2 143666 856
rect 143834 2 144034 856
rect 144202 2 144402 856
rect 144570 2 144770 856
rect 144938 2 145138 856
rect 145306 2 145506 856
rect 145674 2 145874 856
rect 146042 2 146242 856
rect 146410 2 146610 856
rect 146778 2 146978 856
rect 147146 2 147346 856
rect 147514 2 147714 856
rect 147882 2 148082 856
rect 148250 2 148450 856
rect 148618 2 148818 856
rect 148986 2 149186 856
rect 149354 2 149554 856
rect 149722 2 149922 856
rect 150090 2 150290 856
rect 150458 2 150658 856
rect 150826 2 151026 856
rect 151194 2 151394 856
rect 151562 2 151762 856
rect 151930 2 152130 856
rect 152298 2 152498 856
rect 152666 2 152866 856
rect 153034 2 153234 856
rect 153402 2 153602 856
rect 153770 2 153970 856
rect 154138 2 154338 856
rect 154506 2 154706 856
rect 154874 2 155074 856
rect 155242 2 155442 856
rect 155610 2 155810 856
rect 155978 2 156178 856
rect 156346 2 156546 856
rect 156714 2 156914 856
rect 157082 2 157282 856
rect 157450 2 157650 856
rect 157818 2 158018 856
rect 158186 2 158386 856
rect 158554 2 158754 856
rect 158922 2 159122 856
rect 159290 2 159490 856
rect 159658 2 159858 856
rect 160026 2 160226 856
rect 160394 2 160594 856
rect 160762 2 160962 856
rect 161130 2 161330 856
rect 161498 2 161698 856
rect 161866 2 162066 856
rect 162234 2 162434 856
rect 162602 2 162802 856
rect 162970 2 163170 856
rect 163338 2 163538 856
rect 163706 2 163906 856
rect 164074 2 164274 856
rect 164442 2 164642 856
rect 164810 2 165010 856
rect 165178 2 165378 856
rect 165546 2 165746 856
rect 165914 2 166114 856
rect 166282 2 166482 856
rect 166650 2 167236 856
<< metal3 >>
rect 0 11976 800 12096
rect 0 11432 800 11552
rect 0 10888 800 11008
rect 0 10344 800 10464
rect 0 9800 800 9920
rect 0 9256 800 9376
rect 0 8712 800 8832
rect 0 8168 800 8288
rect 0 7624 800 7744
rect 0 7080 800 7200
rect 0 6536 800 6656
rect 0 5992 800 6112
rect 0 5448 800 5568
rect 0 4904 800 5024
rect 0 4360 800 4480
rect 0 3816 800 3936
rect 0 3272 800 3392
rect 0 2728 800 2848
rect 0 2184 800 2304
rect 0 1640 800 1760
rect 0 1096 800 1216
<< obsm3 >>
rect 800 12176 166047 13021
rect 880 11896 166047 12176
rect 800 11632 166047 11896
rect 880 11352 166047 11632
rect 800 11088 166047 11352
rect 880 10808 166047 11088
rect 800 10544 166047 10808
rect 880 10264 166047 10544
rect 800 10000 166047 10264
rect 880 9720 166047 10000
rect 800 9456 166047 9720
rect 880 9176 166047 9456
rect 800 8912 166047 9176
rect 880 8632 166047 8912
rect 800 8368 166047 8632
rect 880 8088 166047 8368
rect 800 7824 166047 8088
rect 880 7544 166047 7824
rect 800 7280 166047 7544
rect 880 7000 166047 7280
rect 800 6736 166047 7000
rect 880 6456 166047 6736
rect 800 6192 166047 6456
rect 880 5912 166047 6192
rect 800 5648 166047 5912
rect 880 5368 166047 5648
rect 800 5104 166047 5368
rect 880 4824 166047 5104
rect 800 4560 166047 4824
rect 880 4280 166047 4560
rect 800 4016 166047 4280
rect 880 3736 166047 4016
rect 800 3472 166047 3736
rect 880 3192 166047 3472
rect 800 2928 166047 3192
rect 880 2648 166047 2928
rect 800 2384 166047 2648
rect 880 2104 166047 2384
rect 800 1840 166047 2104
rect 880 1560 166047 1840
rect 800 1296 166047 1560
rect 880 1016 166047 1296
rect 800 35 166047 1016
<< obsm4 >>
rect 5494 171 153213 13021
<< obsm5 >>
rect 368 180 169556 10582
<< labels >>
rlabel metal2 s 570 0 626 800 6 caravel_clk
port 1 nsew
rlabel metal2 s 938 0 994 800 6 caravel_clk2
port 2 nsew
rlabel metal3 s 0 1096 800 1216 6 caravel_rstn
port 3 nsew
rlabel metal2 s 754 12200 810 13000 6 la_data_in_core[0]
port 4 nsew
rlabel metal3 s 0 11976 800 12096 6 la_data_in_core[100]
port 5 nsew
rlabel metal2 s 1122 12200 1178 13000 6 la_data_in_core[101]
port 6 nsew
rlabel metal3 s 0 11432 800 11552 6 la_data_in_core[102]
port 7 nsew
rlabel metal2 s 1490 12200 1546 13000 6 la_data_in_core[103]
port 8 nsew
rlabel metal2 s 1858 12200 1914 13000 6 la_data_in_core[104]
port 9 nsew
rlabel metal3 s 0 10888 800 11008 6 la_data_in_core[105]
port 10 nsew
rlabel metal2 s 2226 12200 2282 13000 6 la_data_in_core[106]
port 11 nsew
rlabel metal3 s 0 10344 800 10464 6 la_data_in_core[107]
port 12 nsew
rlabel metal2 s 2594 12200 2650 13000 6 la_data_in_core[108]
port 13 nsew
rlabel metal2 s 2962 12200 3018 13000 6 la_data_in_core[109]
port 14 nsew
rlabel metal3 s 0 9800 800 9920 6 la_data_in_core[10]
port 15 nsew
rlabel metal2 s 3330 12200 3386 13000 6 la_data_in_core[110]
port 16 nsew
rlabel metal3 s 0 9256 800 9376 6 la_data_in_core[111]
port 17 nsew
rlabel metal2 s 3698 12200 3754 13000 6 la_data_in_core[112]
port 18 nsew
rlabel metal2 s 4066 12200 4122 13000 6 la_data_in_core[113]
port 19 nsew
rlabel metal3 s 0 8712 800 8832 6 la_data_in_core[114]
port 20 nsew
rlabel metal2 s 4434 12200 4490 13000 6 la_data_in_core[115]
port 21 nsew
rlabel metal3 s 0 8168 800 8288 6 la_data_in_core[116]
port 22 nsew
rlabel metal2 s 4802 12200 4858 13000 6 la_data_in_core[117]
port 23 nsew
rlabel metal2 s 5170 12200 5226 13000 6 la_data_in_core[118]
port 24 nsew
rlabel metal3 s 0 7624 800 7744 6 la_data_in_core[119]
port 25 nsew
rlabel metal2 s 5538 12200 5594 13000 6 la_data_in_core[11]
port 26 nsew
rlabel metal3 s 0 7080 800 7200 6 la_data_in_core[120]
port 27 nsew
rlabel metal2 s 5906 12200 5962 13000 6 la_data_in_core[121]
port 28 nsew
rlabel metal2 s 6274 12200 6330 13000 6 la_data_in_core[122]
port 29 nsew
rlabel metal3 s 0 6536 800 6656 6 la_data_in_core[123]
port 30 nsew
rlabel metal2 s 6642 12200 6698 13000 6 la_data_in_core[124]
port 31 nsew
rlabel metal3 s 0 5992 800 6112 6 la_data_in_core[125]
port 32 nsew
rlabel metal2 s 7010 12200 7066 13000 6 la_data_in_core[126]
port 33 nsew
rlabel metal2 s 7378 12200 7434 13000 6 la_data_in_core[127]
port 34 nsew
rlabel metal3 s 0 5448 800 5568 6 la_data_in_core[12]
port 35 nsew
rlabel metal2 s 7746 12200 7802 13000 6 la_data_in_core[13]
port 36 nsew
rlabel metal3 s 0 4904 800 5024 6 la_data_in_core[14]
port 37 nsew
rlabel metal2 s 8114 12200 8170 13000 6 la_data_in_core[15]
port 38 nsew
rlabel metal2 s 8482 12200 8538 13000 6 la_data_in_core[16]
port 39 nsew
rlabel metal3 s 0 4360 800 4480 6 la_data_in_core[17]
port 40 nsew
rlabel metal2 s 8850 12200 8906 13000 6 la_data_in_core[18]
port 41 nsew
rlabel metal3 s 0 3816 800 3936 6 la_data_in_core[19]
port 42 nsew
rlabel metal2 s 9218 12200 9274 13000 6 la_data_in_core[1]
port 43 nsew
rlabel metal2 s 9586 12200 9642 13000 6 la_data_in_core[20]
port 44 nsew
rlabel metal3 s 0 3272 800 3392 6 la_data_in_core[21]
port 45 nsew
rlabel metal2 s 9954 12200 10010 13000 6 la_data_in_core[22]
port 46 nsew
rlabel metal3 s 0 2728 800 2848 6 la_data_in_core[23]
port 47 nsew
rlabel metal2 s 10322 12200 10378 13000 6 la_data_in_core[24]
port 48 nsew
rlabel metal2 s 10690 12200 10746 13000 6 la_data_in_core[25]
port 49 nsew
rlabel metal3 s 0 2184 800 2304 6 la_data_in_core[26]
port 50 nsew
rlabel metal2 s 11058 12200 11114 13000 6 la_data_in_core[27]
port 51 nsew
rlabel metal3 s 0 1640 800 1760 6 la_data_in_core[28]
port 52 nsew
rlabel metal2 s 11426 12200 11482 13000 6 la_data_in_core[29]
port 53 nsew
rlabel metal2 s 11794 12200 11850 13000 6 la_data_in_core[2]
port 54 nsew
rlabel metal2 s 12162 12200 12218 13000 6 la_data_in_core[30]
port 55 nsew
rlabel metal2 s 12530 12200 12586 13000 6 la_data_in_core[31]
port 56 nsew
rlabel metal2 s 12898 12200 12954 13000 6 la_data_in_core[32]
port 57 nsew
rlabel metal2 s 13266 12200 13322 13000 6 la_data_in_core[33]
port 58 nsew
rlabel metal2 s 13634 12200 13690 13000 6 la_data_in_core[34]
port 59 nsew
rlabel metal2 s 14002 12200 14058 13000 6 la_data_in_core[35]
port 60 nsew
rlabel metal2 s 1306 0 1362 800 6 la_data_in_core[36]
port 61 nsew
rlabel metal2 s 14370 12200 14426 13000 6 la_data_in_core[37]
port 62 nsew
rlabel metal2 s 1674 0 1730 800 6 la_data_in_core[38]
port 63 nsew
rlabel metal2 s 14738 12200 14794 13000 6 la_data_in_core[39]
port 64 nsew
rlabel metal2 s 2042 0 2098 800 6 la_data_in_core[3]
port 65 nsew
rlabel metal2 s 15106 12200 15162 13000 6 la_data_in_core[40]
port 66 nsew
rlabel metal2 s 2410 0 2466 800 6 la_data_in_core[41]
port 67 nsew
rlabel metal2 s 15474 12200 15530 13000 6 la_data_in_core[42]
port 68 nsew
rlabel metal2 s 2778 0 2834 800 6 la_data_in_core[43]
port 69 nsew
rlabel metal2 s 15842 12200 15898 13000 6 la_data_in_core[44]
port 70 nsew
rlabel metal2 s 3146 0 3202 800 6 la_data_in_core[45]
port 71 nsew
rlabel metal2 s 16210 12200 16266 13000 6 la_data_in_core[46]
port 72 nsew
rlabel metal2 s 3514 0 3570 800 6 la_data_in_core[47]
port 73 nsew
rlabel metal2 s 16578 12200 16634 13000 6 la_data_in_core[48]
port 74 nsew
rlabel metal2 s 3882 0 3938 800 6 la_data_in_core[49]
port 75 nsew
rlabel metal2 s 16946 12200 17002 13000 6 la_data_in_core[4]
port 76 nsew
rlabel metal2 s 4250 0 4306 800 6 la_data_in_core[50]
port 77 nsew
rlabel metal2 s 17314 12200 17370 13000 6 la_data_in_core[51]
port 78 nsew
rlabel metal2 s 4618 0 4674 800 6 la_data_in_core[52]
port 79 nsew
rlabel metal2 s 17682 12200 17738 13000 6 la_data_in_core[53]
port 80 nsew
rlabel metal2 s 4986 0 5042 800 6 la_data_in_core[54]
port 81 nsew
rlabel metal2 s 18050 12200 18106 13000 6 la_data_in_core[55]
port 82 nsew
rlabel metal2 s 5354 0 5410 800 6 la_data_in_core[56]
port 83 nsew
rlabel metal2 s 18418 12200 18474 13000 6 la_data_in_core[57]
port 84 nsew
rlabel metal2 s 5722 0 5778 800 6 la_data_in_core[58]
port 85 nsew
rlabel metal2 s 18786 12200 18842 13000 6 la_data_in_core[59]
port 86 nsew
rlabel metal2 s 6090 0 6146 800 6 la_data_in_core[5]
port 87 nsew
rlabel metal2 s 19154 12200 19210 13000 6 la_data_in_core[60]
port 88 nsew
rlabel metal2 s 6458 0 6514 800 6 la_data_in_core[61]
port 89 nsew
rlabel metal2 s 19522 12200 19578 13000 6 la_data_in_core[62]
port 90 nsew
rlabel metal2 s 6826 0 6882 800 6 la_data_in_core[63]
port 91 nsew
rlabel metal2 s 19890 12200 19946 13000 6 la_data_in_core[64]
port 92 nsew
rlabel metal2 s 7194 0 7250 800 6 la_data_in_core[65]
port 93 nsew
rlabel metal2 s 20258 12200 20314 13000 6 la_data_in_core[66]
port 94 nsew
rlabel metal2 s 7562 0 7618 800 6 la_data_in_core[67]
port 95 nsew
rlabel metal2 s 20626 12200 20682 13000 6 la_data_in_core[68]
port 96 nsew
rlabel metal2 s 7930 0 7986 800 6 la_data_in_core[69]
port 97 nsew
rlabel metal2 s 20994 12200 21050 13000 6 la_data_in_core[6]
port 98 nsew
rlabel metal2 s 8298 0 8354 800 6 la_data_in_core[70]
port 99 nsew
rlabel metal2 s 21362 12200 21418 13000 6 la_data_in_core[71]
port 100 nsew
rlabel metal2 s 8666 0 8722 800 6 la_data_in_core[72]
port 101 nsew
rlabel metal2 s 21730 12200 21786 13000 6 la_data_in_core[73]
port 102 nsew
rlabel metal2 s 9034 0 9090 800 6 la_data_in_core[74]
port 103 nsew
rlabel metal2 s 22098 12200 22154 13000 6 la_data_in_core[75]
port 104 nsew
rlabel metal2 s 9402 0 9458 800 6 la_data_in_core[76]
port 105 nsew
rlabel metal2 s 22466 12200 22522 13000 6 la_data_in_core[77]
port 106 nsew
rlabel metal2 s 9770 0 9826 800 6 la_data_in_core[78]
port 107 nsew
rlabel metal2 s 22834 12200 22890 13000 6 la_data_in_core[79]
port 108 nsew
rlabel metal2 s 10138 0 10194 800 6 la_data_in_core[7]
port 109 nsew
rlabel metal2 s 23202 12200 23258 13000 6 la_data_in_core[80]
port 110 nsew
rlabel metal2 s 10506 0 10562 800 6 la_data_in_core[81]
port 111 nsew
rlabel metal2 s 23570 12200 23626 13000 6 la_data_in_core[82]
port 112 nsew
rlabel metal2 s 10874 0 10930 800 6 la_data_in_core[83]
port 113 nsew
rlabel metal2 s 23938 12200 23994 13000 6 la_data_in_core[84]
port 114 nsew
rlabel metal2 s 11242 0 11298 800 6 la_data_in_core[85]
port 115 nsew
rlabel metal2 s 24306 12200 24362 13000 6 la_data_in_core[86]
port 116 nsew
rlabel metal2 s 11610 0 11666 800 6 la_data_in_core[87]
port 117 nsew
rlabel metal2 s 24674 12200 24730 13000 6 la_data_in_core[88]
port 118 nsew
rlabel metal2 s 11978 0 12034 800 6 la_data_in_core[89]
port 119 nsew
rlabel metal2 s 25042 12200 25098 13000 6 la_data_in_core[8]
port 120 nsew
rlabel metal2 s 12346 0 12402 800 6 la_data_in_core[90]
port 121 nsew
rlabel metal2 s 25410 12200 25466 13000 6 la_data_in_core[91]
port 122 nsew
rlabel metal2 s 12714 0 12770 800 6 la_data_in_core[92]
port 123 nsew
rlabel metal2 s 25778 12200 25834 13000 6 la_data_in_core[93]
port 124 nsew
rlabel metal2 s 13082 0 13138 800 6 la_data_in_core[94]
port 125 nsew
rlabel metal2 s 26146 12200 26202 13000 6 la_data_in_core[95]
port 126 nsew
rlabel metal2 s 13450 0 13506 800 6 la_data_in_core[96]
port 127 nsew
rlabel metal2 s 26514 12200 26570 13000 6 la_data_in_core[97]
port 128 nsew
rlabel metal2 s 13818 0 13874 800 6 la_data_in_core[98]
port 129 nsew
rlabel metal2 s 26882 12200 26938 13000 6 la_data_in_core[99]
port 130 nsew
rlabel metal2 s 14186 0 14242 800 6 la_data_in_core[9]
port 131 nsew
rlabel metal2 s 14554 0 14610 800 6 la_data_in_mprj[0]
port 132 nsew
rlabel metal2 s 14922 0 14978 800 6 la_data_in_mprj[100]
port 133 nsew
rlabel metal2 s 15290 0 15346 800 6 la_data_in_mprj[101]
port 134 nsew
rlabel metal2 s 15658 0 15714 800 6 la_data_in_mprj[102]
port 135 nsew
rlabel metal2 s 16026 0 16082 800 6 la_data_in_mprj[103]
port 136 nsew
rlabel metal2 s 16394 0 16450 800 6 la_data_in_mprj[104]
port 137 nsew
rlabel metal2 s 16762 0 16818 800 6 la_data_in_mprj[105]
port 138 nsew
rlabel metal2 s 17130 0 17186 800 6 la_data_in_mprj[106]
port 139 nsew
rlabel metal2 s 17498 0 17554 800 6 la_data_in_mprj[107]
port 140 nsew
rlabel metal2 s 17866 0 17922 800 6 la_data_in_mprj[108]
port 141 nsew
rlabel metal2 s 18234 0 18290 800 6 la_data_in_mprj[109]
port 142 nsew
rlabel metal2 s 18602 0 18658 800 6 la_data_in_mprj[10]
port 143 nsew
rlabel metal2 s 18970 0 19026 800 6 la_data_in_mprj[110]
port 144 nsew
rlabel metal2 s 19338 0 19394 800 6 la_data_in_mprj[111]
port 145 nsew
rlabel metal2 s 19706 0 19762 800 6 la_data_in_mprj[112]
port 146 nsew
rlabel metal2 s 20074 0 20130 800 6 la_data_in_mprj[113]
port 147 nsew
rlabel metal2 s 20442 0 20498 800 6 la_data_in_mprj[114]
port 148 nsew
rlabel metal2 s 20810 0 20866 800 6 la_data_in_mprj[115]
port 149 nsew
rlabel metal2 s 21178 0 21234 800 6 la_data_in_mprj[116]
port 150 nsew
rlabel metal2 s 21546 0 21602 800 6 la_data_in_mprj[117]
port 151 nsew
rlabel metal2 s 21914 0 21970 800 6 la_data_in_mprj[118]
port 152 nsew
rlabel metal2 s 22282 0 22338 800 6 la_data_in_mprj[119]
port 153 nsew
rlabel metal2 s 22650 0 22706 800 6 la_data_in_mprj[11]
port 154 nsew
rlabel metal2 s 23018 0 23074 800 6 la_data_in_mprj[120]
port 155 nsew
rlabel metal2 s 23386 0 23442 800 6 la_data_in_mprj[121]
port 156 nsew
rlabel metal2 s 23754 0 23810 800 6 la_data_in_mprj[122]
port 157 nsew
rlabel metal2 s 24122 0 24178 800 6 la_data_in_mprj[123]
port 158 nsew
rlabel metal2 s 24490 0 24546 800 6 la_data_in_mprj[124]
port 159 nsew
rlabel metal2 s 24858 0 24914 800 6 la_data_in_mprj[125]
port 160 nsew
rlabel metal2 s 25226 0 25282 800 6 la_data_in_mprj[126]
port 161 nsew
rlabel metal2 s 25594 0 25650 800 6 la_data_in_mprj[127]
port 162 nsew
rlabel metal2 s 25962 0 26018 800 6 la_data_in_mprj[12]
port 163 nsew
rlabel metal2 s 26330 0 26386 800 6 la_data_in_mprj[13]
port 164 nsew
rlabel metal2 s 26698 0 26754 800 6 la_data_in_mprj[14]
port 165 nsew
rlabel metal2 s 27066 0 27122 800 6 la_data_in_mprj[15]
port 166 nsew
rlabel metal2 s 27434 0 27490 800 6 la_data_in_mprj[16]
port 167 nsew
rlabel metal2 s 27802 0 27858 800 6 la_data_in_mprj[17]
port 168 nsew
rlabel metal2 s 28170 0 28226 800 6 la_data_in_mprj[18]
port 169 nsew
rlabel metal2 s 28538 0 28594 800 6 la_data_in_mprj[19]
port 170 nsew
rlabel metal2 s 28906 0 28962 800 6 la_data_in_mprj[1]
port 171 nsew
rlabel metal2 s 29274 0 29330 800 6 la_data_in_mprj[20]
port 172 nsew
rlabel metal2 s 29642 0 29698 800 6 la_data_in_mprj[21]
port 173 nsew
rlabel metal2 s 30010 0 30066 800 6 la_data_in_mprj[22]
port 174 nsew
rlabel metal2 s 30378 0 30434 800 6 la_data_in_mprj[23]
port 175 nsew
rlabel metal2 s 30746 0 30802 800 6 la_data_in_mprj[24]
port 176 nsew
rlabel metal2 s 31114 0 31170 800 6 la_data_in_mprj[25]
port 177 nsew
rlabel metal2 s 31482 0 31538 800 6 la_data_in_mprj[26]
port 178 nsew
rlabel metal2 s 31850 0 31906 800 6 la_data_in_mprj[27]
port 179 nsew
rlabel metal2 s 32218 0 32274 800 6 la_data_in_mprj[28]
port 180 nsew
rlabel metal2 s 32586 0 32642 800 6 la_data_in_mprj[29]
port 181 nsew
rlabel metal2 s 32954 0 33010 800 6 la_data_in_mprj[2]
port 182 nsew
rlabel metal2 s 33322 0 33378 800 6 la_data_in_mprj[30]
port 183 nsew
rlabel metal2 s 33690 0 33746 800 6 la_data_in_mprj[31]
port 184 nsew
rlabel metal2 s 34058 0 34114 800 6 la_data_in_mprj[32]
port 185 nsew
rlabel metal2 s 34426 0 34482 800 6 la_data_in_mprj[33]
port 186 nsew
rlabel metal2 s 34794 0 34850 800 6 la_data_in_mprj[34]
port 187 nsew
rlabel metal2 s 35162 0 35218 800 6 la_data_in_mprj[35]
port 188 nsew
rlabel metal2 s 35530 0 35586 800 6 la_data_in_mprj[36]
port 189 nsew
rlabel metal2 s 35898 0 35954 800 6 la_data_in_mprj[37]
port 190 nsew
rlabel metal2 s 36266 0 36322 800 6 la_data_in_mprj[38]
port 191 nsew
rlabel metal2 s 36634 0 36690 800 6 la_data_in_mprj[39]
port 192 nsew
rlabel metal2 s 37002 0 37058 800 6 la_data_in_mprj[3]
port 193 nsew
rlabel metal2 s 37370 0 37426 800 6 la_data_in_mprj[40]
port 194 nsew
rlabel metal2 s 37738 0 37794 800 6 la_data_in_mprj[41]
port 195 nsew
rlabel metal2 s 38106 0 38162 800 6 la_data_in_mprj[42]
port 196 nsew
rlabel metal2 s 38474 0 38530 800 6 la_data_in_mprj[43]
port 197 nsew
rlabel metal2 s 38842 0 38898 800 6 la_data_in_mprj[44]
port 198 nsew
rlabel metal2 s 39210 0 39266 800 6 la_data_in_mprj[45]
port 199 nsew
rlabel metal2 s 39578 0 39634 800 6 la_data_in_mprj[46]
port 200 nsew
rlabel metal2 s 39946 0 40002 800 6 la_data_in_mprj[47]
port 201 nsew
rlabel metal2 s 27250 12200 27306 13000 6 la_data_in_mprj[48]
port 202 nsew
rlabel metal2 s 40314 0 40370 800 6 la_data_in_mprj[49]
port 203 nsew
rlabel metal2 s 27618 12200 27674 13000 6 la_data_in_mprj[4]
port 204 nsew
rlabel metal2 s 40682 0 40738 800 6 la_data_in_mprj[50]
port 205 nsew
rlabel metal2 s 27986 12200 28042 13000 6 la_data_in_mprj[51]
port 206 nsew
rlabel metal2 s 41050 0 41106 800 6 la_data_in_mprj[52]
port 207 nsew
rlabel metal2 s 28354 12200 28410 13000 6 la_data_in_mprj[53]
port 208 nsew
rlabel metal2 s 41418 0 41474 800 6 la_data_in_mprj[54]
port 209 nsew
rlabel metal2 s 28722 12200 28778 13000 6 la_data_in_mprj[55]
port 210 nsew
rlabel metal2 s 41786 0 41842 800 6 la_data_in_mprj[56]
port 211 nsew
rlabel metal2 s 29090 12200 29146 13000 6 la_data_in_mprj[57]
port 212 nsew
rlabel metal2 s 42154 0 42210 800 6 la_data_in_mprj[58]
port 213 nsew
rlabel metal2 s 29458 12200 29514 13000 6 la_data_in_mprj[59]
port 214 nsew
rlabel metal2 s 42522 0 42578 800 6 la_data_in_mprj[5]
port 215 nsew
rlabel metal2 s 29826 12200 29882 13000 6 la_data_in_mprj[60]
port 216 nsew
rlabel metal2 s 42890 0 42946 800 6 la_data_in_mprj[61]
port 217 nsew
rlabel metal2 s 30194 12200 30250 13000 6 la_data_in_mprj[62]
port 218 nsew
rlabel metal2 s 43258 0 43314 800 6 la_data_in_mprj[63]
port 219 nsew
rlabel metal2 s 30562 12200 30618 13000 6 la_data_in_mprj[64]
port 220 nsew
rlabel metal2 s 43626 0 43682 800 6 la_data_in_mprj[65]
port 221 nsew
rlabel metal2 s 30930 12200 30986 13000 6 la_data_in_mprj[66]
port 222 nsew
rlabel metal2 s 43994 0 44050 800 6 la_data_in_mprj[67]
port 223 nsew
rlabel metal2 s 31298 12200 31354 13000 6 la_data_in_mprj[68]
port 224 nsew
rlabel metal2 s 44362 0 44418 800 6 la_data_in_mprj[69]
port 225 nsew
rlabel metal2 s 31666 12200 31722 13000 6 la_data_in_mprj[6]
port 226 nsew
rlabel metal2 s 44730 0 44786 800 6 la_data_in_mprj[70]
port 227 nsew
rlabel metal2 s 32034 12200 32090 13000 6 la_data_in_mprj[71]
port 228 nsew
rlabel metal2 s 45098 0 45154 800 6 la_data_in_mprj[72]
port 229 nsew
rlabel metal2 s 32402 12200 32458 13000 6 la_data_in_mprj[73]
port 230 nsew
rlabel metal2 s 45466 0 45522 800 6 la_data_in_mprj[74]
port 231 nsew
rlabel metal2 s 32770 12200 32826 13000 6 la_data_in_mprj[75]
port 232 nsew
rlabel metal2 s 45834 0 45890 800 6 la_data_in_mprj[76]
port 233 nsew
rlabel metal2 s 33138 12200 33194 13000 6 la_data_in_mprj[77]
port 234 nsew
rlabel metal2 s 46202 0 46258 800 6 la_data_in_mprj[78]
port 235 nsew
rlabel metal2 s 33506 12200 33562 13000 6 la_data_in_mprj[79]
port 236 nsew
rlabel metal2 s 46570 0 46626 800 6 la_data_in_mprj[7]
port 237 nsew
rlabel metal2 s 33874 12200 33930 13000 6 la_data_in_mprj[80]
port 238 nsew
rlabel metal2 s 46938 0 46994 800 6 la_data_in_mprj[81]
port 239 nsew
rlabel metal2 s 34242 12200 34298 13000 6 la_data_in_mprj[82]
port 240 nsew
rlabel metal2 s 47306 0 47362 800 6 la_data_in_mprj[83]
port 241 nsew
rlabel metal2 s 34610 12200 34666 13000 6 la_data_in_mprj[84]
port 242 nsew
rlabel metal2 s 47674 0 47730 800 6 la_data_in_mprj[85]
port 243 nsew
rlabel metal2 s 34978 12200 35034 13000 6 la_data_in_mprj[86]
port 244 nsew
rlabel metal2 s 48042 0 48098 800 6 la_data_in_mprj[87]
port 245 nsew
rlabel metal2 s 35346 12200 35402 13000 6 la_data_in_mprj[88]
port 246 nsew
rlabel metal2 s 48410 0 48466 800 6 la_data_in_mprj[89]
port 247 nsew
rlabel metal2 s 35714 12200 35770 13000 6 la_data_in_mprj[8]
port 248 nsew
rlabel metal2 s 48778 0 48834 800 6 la_data_in_mprj[90]
port 249 nsew
rlabel metal2 s 36082 12200 36138 13000 6 la_data_in_mprj[91]
port 250 nsew
rlabel metal2 s 49146 0 49202 800 6 la_data_in_mprj[92]
port 251 nsew
rlabel metal2 s 36450 12200 36506 13000 6 la_data_in_mprj[93]
port 252 nsew
rlabel metal2 s 49514 0 49570 800 6 la_data_in_mprj[94]
port 253 nsew
rlabel metal2 s 36818 12200 36874 13000 6 la_data_in_mprj[95]
port 254 nsew
rlabel metal2 s 49882 0 49938 800 6 la_data_in_mprj[96]
port 255 nsew
rlabel metal2 s 37186 12200 37242 13000 6 la_data_in_mprj[97]
port 256 nsew
rlabel metal2 s 50250 0 50306 800 6 la_data_in_mprj[98]
port 257 nsew
rlabel metal2 s 37554 12200 37610 13000 6 la_data_in_mprj[99]
port 258 nsew
rlabel metal2 s 50618 0 50674 800 6 la_data_in_mprj[9]
port 259 nsew
rlabel metal2 s 37922 12200 37978 13000 6 la_data_out_core[0]
port 260 nsew
rlabel metal2 s 38290 12200 38346 13000 6 la_data_out_core[100]
port 261 nsew
rlabel metal2 s 38658 12200 38714 13000 6 la_data_out_core[101]
port 262 nsew
rlabel metal2 s 39026 12200 39082 13000 6 la_data_out_core[102]
port 263 nsew
rlabel metal2 s 39394 12200 39450 13000 6 la_data_out_core[103]
port 264 nsew
rlabel metal2 s 39762 12200 39818 13000 6 la_data_out_core[104]
port 265 nsew
rlabel metal2 s 40130 12200 40186 13000 6 la_data_out_core[105]
port 266 nsew
rlabel metal2 s 40498 12200 40554 13000 6 la_data_out_core[106]
port 267 nsew
rlabel metal2 s 40866 12200 40922 13000 6 la_data_out_core[107]
port 268 nsew
rlabel metal2 s 41234 12200 41290 13000 6 la_data_out_core[108]
port 269 nsew
rlabel metal2 s 41602 12200 41658 13000 6 la_data_out_core[109]
port 270 nsew
rlabel metal2 s 41970 12200 42026 13000 6 la_data_out_core[10]
port 271 nsew
rlabel metal2 s 42338 12200 42394 13000 6 la_data_out_core[110]
port 272 nsew
rlabel metal2 s 42706 12200 42762 13000 6 la_data_out_core[111]
port 273 nsew
rlabel metal2 s 43074 12200 43130 13000 6 la_data_out_core[112]
port 274 nsew
rlabel metal2 s 43442 12200 43498 13000 6 la_data_out_core[113]
port 275 nsew
rlabel metal2 s 43810 12200 43866 13000 6 la_data_out_core[114]
port 276 nsew
rlabel metal2 s 44178 12200 44234 13000 6 la_data_out_core[115]
port 277 nsew
rlabel metal2 s 44546 12200 44602 13000 6 la_data_out_core[116]
port 278 nsew
rlabel metal2 s 44914 12200 44970 13000 6 la_data_out_core[117]
port 279 nsew
rlabel metal2 s 45282 12200 45338 13000 6 la_data_out_core[118]
port 280 nsew
rlabel metal2 s 45650 12200 45706 13000 6 la_data_out_core[119]
port 281 nsew
rlabel metal2 s 46018 12200 46074 13000 6 la_data_out_core[11]
port 282 nsew
rlabel metal2 s 46386 12200 46442 13000 6 la_data_out_core[120]
port 283 nsew
rlabel metal2 s 46754 12200 46810 13000 6 la_data_out_core[121]
port 284 nsew
rlabel metal2 s 47122 12200 47178 13000 6 la_data_out_core[122]
port 285 nsew
rlabel metal2 s 47490 12200 47546 13000 6 la_data_out_core[123]
port 286 nsew
rlabel metal2 s 47858 12200 47914 13000 6 la_data_out_core[124]
port 287 nsew
rlabel metal2 s 48226 12200 48282 13000 6 la_data_out_core[125]
port 288 nsew
rlabel metal2 s 48594 12200 48650 13000 6 la_data_out_core[126]
port 289 nsew
rlabel metal2 s 48962 12200 49018 13000 6 la_data_out_core[127]
port 290 nsew
rlabel metal2 s 49330 12200 49386 13000 6 la_data_out_core[12]
port 291 nsew
rlabel metal2 s 49698 12200 49754 13000 6 la_data_out_core[13]
port 292 nsew
rlabel metal2 s 50066 12200 50122 13000 6 la_data_out_core[14]
port 293 nsew
rlabel metal2 s 50434 12200 50490 13000 6 la_data_out_core[15]
port 294 nsew
rlabel metal2 s 50802 12200 50858 13000 6 la_data_out_core[16]
port 295 nsew
rlabel metal2 s 51170 12200 51226 13000 6 la_data_out_core[17]
port 296 nsew
rlabel metal2 s 51538 12200 51594 13000 6 la_data_out_core[18]
port 297 nsew
rlabel metal2 s 51906 12200 51962 13000 6 la_data_out_core[19]
port 298 nsew
rlabel metal2 s 52274 12200 52330 13000 6 la_data_out_core[1]
port 299 nsew
rlabel metal2 s 52642 12200 52698 13000 6 la_data_out_core[20]
port 300 nsew
rlabel metal2 s 53010 12200 53066 13000 6 la_data_out_core[21]
port 301 nsew
rlabel metal2 s 53378 12200 53434 13000 6 la_data_out_core[22]
port 302 nsew
rlabel metal2 s 53746 12200 53802 13000 6 la_data_out_core[23]
port 303 nsew
rlabel metal2 s 54114 12200 54170 13000 6 la_data_out_core[24]
port 304 nsew
rlabel metal2 s 54482 12200 54538 13000 6 la_data_out_core[25]
port 305 nsew
rlabel metal2 s 54850 12200 54906 13000 6 la_data_out_core[26]
port 306 nsew
rlabel metal2 s 55218 12200 55274 13000 6 la_data_out_core[27]
port 307 nsew
rlabel metal2 s 55586 12200 55642 13000 6 la_data_out_core[28]
port 308 nsew
rlabel metal2 s 55954 12200 56010 13000 6 la_data_out_core[29]
port 309 nsew
rlabel metal2 s 56322 12200 56378 13000 6 la_data_out_core[2]
port 310 nsew
rlabel metal2 s 56690 12200 56746 13000 6 la_data_out_core[30]
port 311 nsew
rlabel metal2 s 57058 12200 57114 13000 6 la_data_out_core[31]
port 312 nsew
rlabel metal2 s 57426 12200 57482 13000 6 la_data_out_core[32]
port 313 nsew
rlabel metal2 s 57794 12200 57850 13000 6 la_data_out_core[33]
port 314 nsew
rlabel metal2 s 58162 12200 58218 13000 6 la_data_out_core[34]
port 315 nsew
rlabel metal2 s 58530 12200 58586 13000 6 la_data_out_core[35]
port 316 nsew
rlabel metal2 s 58898 12200 58954 13000 6 la_data_out_core[36]
port 317 nsew
rlabel metal2 s 59266 12200 59322 13000 6 la_data_out_core[37]
port 318 nsew
rlabel metal2 s 59634 12200 59690 13000 6 la_data_out_core[38]
port 319 nsew
rlabel metal2 s 60002 12200 60058 13000 6 la_data_out_core[39]
port 320 nsew
rlabel metal2 s 60370 12200 60426 13000 6 la_data_out_core[3]
port 321 nsew
rlabel metal2 s 60738 12200 60794 13000 6 la_data_out_core[40]
port 322 nsew
rlabel metal2 s 61106 12200 61162 13000 6 la_data_out_core[41]
port 323 nsew
rlabel metal2 s 61474 12200 61530 13000 6 la_data_out_core[42]
port 324 nsew
rlabel metal2 s 61842 12200 61898 13000 6 la_data_out_core[43]
port 325 nsew
rlabel metal2 s 62210 12200 62266 13000 6 la_data_out_core[44]
port 326 nsew
rlabel metal2 s 62578 12200 62634 13000 6 la_data_out_core[45]
port 327 nsew
rlabel metal2 s 62946 12200 63002 13000 6 la_data_out_core[46]
port 328 nsew
rlabel metal2 s 63314 12200 63370 13000 6 la_data_out_core[47]
port 329 nsew
rlabel metal2 s 63682 12200 63738 13000 6 la_data_out_core[48]
port 330 nsew
rlabel metal2 s 50986 0 51042 800 6 la_data_out_core[49]
port 331 nsew
rlabel metal2 s 64050 12200 64106 13000 6 la_data_out_core[4]
port 332 nsew
rlabel metal2 s 51354 0 51410 800 6 la_data_out_core[50]
port 333 nsew
rlabel metal2 s 64418 12200 64474 13000 6 la_data_out_core[51]
port 334 nsew
rlabel metal2 s 51722 0 51778 800 6 la_data_out_core[52]
port 335 nsew
rlabel metal2 s 64786 12200 64842 13000 6 la_data_out_core[53]
port 336 nsew
rlabel metal2 s 52090 0 52146 800 6 la_data_out_core[54]
port 337 nsew
rlabel metal2 s 65154 12200 65210 13000 6 la_data_out_core[55]
port 338 nsew
rlabel metal2 s 52458 0 52514 800 6 la_data_out_core[56]
port 339 nsew
rlabel metal2 s 65522 12200 65578 13000 6 la_data_out_core[57]
port 340 nsew
rlabel metal2 s 52826 0 52882 800 6 la_data_out_core[58]
port 341 nsew
rlabel metal2 s 65890 12200 65946 13000 6 la_data_out_core[59]
port 342 nsew
rlabel metal2 s 53194 0 53250 800 6 la_data_out_core[5]
port 343 nsew
rlabel metal2 s 66258 12200 66314 13000 6 la_data_out_core[60]
port 344 nsew
rlabel metal2 s 53562 0 53618 800 6 la_data_out_core[61]
port 345 nsew
rlabel metal2 s 66626 12200 66682 13000 6 la_data_out_core[62]
port 346 nsew
rlabel metal2 s 53930 0 53986 800 6 la_data_out_core[63]
port 347 nsew
rlabel metal2 s 66994 12200 67050 13000 6 la_data_out_core[64]
port 348 nsew
rlabel metal2 s 54298 0 54354 800 6 la_data_out_core[65]
port 349 nsew
rlabel metal2 s 67362 12200 67418 13000 6 la_data_out_core[66]
port 350 nsew
rlabel metal2 s 54666 0 54722 800 6 la_data_out_core[67]
port 351 nsew
rlabel metal2 s 67730 12200 67786 13000 6 la_data_out_core[68]
port 352 nsew
rlabel metal2 s 55034 0 55090 800 6 la_data_out_core[69]
port 353 nsew
rlabel metal2 s 68098 12200 68154 13000 6 la_data_out_core[6]
port 354 nsew
rlabel metal2 s 55402 0 55458 800 6 la_data_out_core[70]
port 355 nsew
rlabel metal2 s 68466 12200 68522 13000 6 la_data_out_core[71]
port 356 nsew
rlabel metal2 s 55770 0 55826 800 6 la_data_out_core[72]
port 357 nsew
rlabel metal2 s 68834 12200 68890 13000 6 la_data_out_core[73]
port 358 nsew
rlabel metal2 s 56138 0 56194 800 6 la_data_out_core[74]
port 359 nsew
rlabel metal2 s 69202 12200 69258 13000 6 la_data_out_core[75]
port 360 nsew
rlabel metal2 s 56506 0 56562 800 6 la_data_out_core[76]
port 361 nsew
rlabel metal2 s 69570 12200 69626 13000 6 la_data_out_core[77]
port 362 nsew
rlabel metal2 s 56874 0 56930 800 6 la_data_out_core[78]
port 363 nsew
rlabel metal2 s 69938 12200 69994 13000 6 la_data_out_core[79]
port 364 nsew
rlabel metal2 s 57242 0 57298 800 6 la_data_out_core[7]
port 365 nsew
rlabel metal2 s 70306 12200 70362 13000 6 la_data_out_core[80]
port 366 nsew
rlabel metal2 s 57610 0 57666 800 6 la_data_out_core[81]
port 367 nsew
rlabel metal2 s 70674 12200 70730 13000 6 la_data_out_core[82]
port 368 nsew
rlabel metal2 s 57978 0 58034 800 6 la_data_out_core[83]
port 369 nsew
rlabel metal2 s 71042 12200 71098 13000 6 la_data_out_core[84]
port 370 nsew
rlabel metal2 s 58346 0 58402 800 6 la_data_out_core[85]
port 371 nsew
rlabel metal2 s 71410 12200 71466 13000 6 la_data_out_core[86]
port 372 nsew
rlabel metal2 s 58714 0 58770 800 6 la_data_out_core[87]
port 373 nsew
rlabel metal2 s 71778 12200 71834 13000 6 la_data_out_core[88]
port 374 nsew
rlabel metal2 s 59082 0 59138 800 6 la_data_out_core[89]
port 375 nsew
rlabel metal2 s 72146 12200 72202 13000 6 la_data_out_core[8]
port 376 nsew
rlabel metal2 s 59450 0 59506 800 6 la_data_out_core[90]
port 377 nsew
rlabel metal2 s 72514 12200 72570 13000 6 la_data_out_core[91]
port 378 nsew
rlabel metal2 s 59818 0 59874 800 6 la_data_out_core[92]
port 379 nsew
rlabel metal2 s 72882 12200 72938 13000 6 la_data_out_core[93]
port 380 nsew
rlabel metal2 s 60186 0 60242 800 6 la_data_out_core[94]
port 381 nsew
rlabel metal2 s 73250 12200 73306 13000 6 la_data_out_core[95]
port 382 nsew
rlabel metal2 s 60554 0 60610 800 6 la_data_out_core[96]
port 383 nsew
rlabel metal2 s 73618 12200 73674 13000 6 la_data_out_core[97]
port 384 nsew
rlabel metal2 s 60922 0 60978 800 6 la_data_out_core[98]
port 385 nsew
rlabel metal2 s 73986 12200 74042 13000 6 la_data_out_core[99]
port 386 nsew
rlabel metal2 s 61290 0 61346 800 6 la_data_out_core[9]
port 387 nsew
rlabel metal2 s 61658 0 61714 800 6 la_data_out_mprj[0]
port 388 nsew
rlabel metal2 s 62026 0 62082 800 6 la_data_out_mprj[100]
port 389 nsew
rlabel metal2 s 62394 0 62450 800 6 la_data_out_mprj[101]
port 390 nsew
rlabel metal2 s 62762 0 62818 800 6 la_data_out_mprj[102]
port 391 nsew
rlabel metal2 s 63130 0 63186 800 6 la_data_out_mprj[103]
port 392 nsew
rlabel metal2 s 63498 0 63554 800 6 la_data_out_mprj[104]
port 393 nsew
rlabel metal2 s 63866 0 63922 800 6 la_data_out_mprj[105]
port 394 nsew
rlabel metal2 s 64234 0 64290 800 6 la_data_out_mprj[106]
port 395 nsew
rlabel metal2 s 64602 0 64658 800 6 la_data_out_mprj[107]
port 396 nsew
rlabel metal2 s 64970 0 65026 800 6 la_data_out_mprj[108]
port 397 nsew
rlabel metal2 s 65338 0 65394 800 6 la_data_out_mprj[109]
port 398 nsew
rlabel metal2 s 65706 0 65762 800 6 la_data_out_mprj[10]
port 399 nsew
rlabel metal2 s 66074 0 66130 800 6 la_data_out_mprj[110]
port 400 nsew
rlabel metal2 s 66442 0 66498 800 6 la_data_out_mprj[111]
port 401 nsew
rlabel metal2 s 66810 0 66866 800 6 la_data_out_mprj[112]
port 402 nsew
rlabel metal2 s 67178 0 67234 800 6 la_data_out_mprj[113]
port 403 nsew
rlabel metal2 s 67546 0 67602 800 6 la_data_out_mprj[114]
port 404 nsew
rlabel metal2 s 67914 0 67970 800 6 la_data_out_mprj[115]
port 405 nsew
rlabel metal2 s 68282 0 68338 800 6 la_data_out_mprj[116]
port 406 nsew
rlabel metal2 s 68650 0 68706 800 6 la_data_out_mprj[117]
port 407 nsew
rlabel metal2 s 69018 0 69074 800 6 la_data_out_mprj[118]
port 408 nsew
rlabel metal2 s 69386 0 69442 800 6 la_data_out_mprj[119]
port 409 nsew
rlabel metal2 s 69754 0 69810 800 6 la_data_out_mprj[11]
port 410 nsew
rlabel metal2 s 70122 0 70178 800 6 la_data_out_mprj[120]
port 411 nsew
rlabel metal2 s 70490 0 70546 800 6 la_data_out_mprj[121]
port 412 nsew
rlabel metal2 s 70858 0 70914 800 6 la_data_out_mprj[122]
port 413 nsew
rlabel metal2 s 71226 0 71282 800 6 la_data_out_mprj[123]
port 414 nsew
rlabel metal2 s 71594 0 71650 800 6 la_data_out_mprj[124]
port 415 nsew
rlabel metal2 s 71962 0 72018 800 6 la_data_out_mprj[125]
port 416 nsew
rlabel metal2 s 72330 0 72386 800 6 la_data_out_mprj[126]
port 417 nsew
rlabel metal2 s 72698 0 72754 800 6 la_data_out_mprj[127]
port 418 nsew
rlabel metal2 s 73066 0 73122 800 6 la_data_out_mprj[12]
port 419 nsew
rlabel metal2 s 73434 0 73490 800 6 la_data_out_mprj[13]
port 420 nsew
rlabel metal2 s 73802 0 73858 800 6 la_data_out_mprj[14]
port 421 nsew
rlabel metal2 s 74170 0 74226 800 6 la_data_out_mprj[15]
port 422 nsew
rlabel metal2 s 74538 0 74594 800 6 la_data_out_mprj[16]
port 423 nsew
rlabel metal2 s 74906 0 74962 800 6 la_data_out_mprj[17]
port 424 nsew
rlabel metal2 s 75274 0 75330 800 6 la_data_out_mprj[18]
port 425 nsew
rlabel metal2 s 75642 0 75698 800 6 la_data_out_mprj[19]
port 426 nsew
rlabel metal2 s 76010 0 76066 800 6 la_data_out_mprj[1]
port 427 nsew
rlabel metal2 s 76378 0 76434 800 6 la_data_out_mprj[20]
port 428 nsew
rlabel metal2 s 76746 0 76802 800 6 la_data_out_mprj[21]
port 429 nsew
rlabel metal2 s 77114 0 77170 800 6 la_data_out_mprj[22]
port 430 nsew
rlabel metal2 s 77482 0 77538 800 6 la_data_out_mprj[23]
port 431 nsew
rlabel metal2 s 77850 0 77906 800 6 la_data_out_mprj[24]
port 432 nsew
rlabel metal2 s 78218 0 78274 800 6 la_data_out_mprj[25]
port 433 nsew
rlabel metal2 s 78586 0 78642 800 6 la_data_out_mprj[26]
port 434 nsew
rlabel metal2 s 78954 0 79010 800 6 la_data_out_mprj[27]
port 435 nsew
rlabel metal2 s 79322 0 79378 800 6 la_data_out_mprj[28]
port 436 nsew
rlabel metal2 s 79690 0 79746 800 6 la_data_out_mprj[29]
port 437 nsew
rlabel metal2 s 80058 0 80114 800 6 la_data_out_mprj[2]
port 438 nsew
rlabel metal2 s 80426 0 80482 800 6 la_data_out_mprj[30]
port 439 nsew
rlabel metal2 s 80794 0 80850 800 6 la_data_out_mprj[31]
port 440 nsew
rlabel metal2 s 81162 0 81218 800 6 la_data_out_mprj[32]
port 441 nsew
rlabel metal2 s 81530 0 81586 800 6 la_data_out_mprj[33]
port 442 nsew
rlabel metal2 s 81898 0 81954 800 6 la_data_out_mprj[34]
port 443 nsew
rlabel metal2 s 82266 0 82322 800 6 la_data_out_mprj[35]
port 444 nsew
rlabel metal2 s 82634 0 82690 800 6 la_data_out_mprj[36]
port 445 nsew
rlabel metal2 s 83002 0 83058 800 6 la_data_out_mprj[37]
port 446 nsew
rlabel metal2 s 83370 0 83426 800 6 la_data_out_mprj[38]
port 447 nsew
rlabel metal2 s 83738 0 83794 800 6 la_data_out_mprj[39]
port 448 nsew
rlabel metal2 s 84106 0 84162 800 6 la_data_out_mprj[3]
port 449 nsew
rlabel metal2 s 84474 0 84530 800 6 la_data_out_mprj[40]
port 450 nsew
rlabel metal2 s 84842 0 84898 800 6 la_data_out_mprj[41]
port 451 nsew
rlabel metal2 s 85210 0 85266 800 6 la_data_out_mprj[42]
port 452 nsew
rlabel metal2 s 85578 0 85634 800 6 la_data_out_mprj[43]
port 453 nsew
rlabel metal2 s 85946 0 86002 800 6 la_data_out_mprj[44]
port 454 nsew
rlabel metal2 s 86314 0 86370 800 6 la_data_out_mprj[45]
port 455 nsew
rlabel metal2 s 86682 0 86738 800 6 la_data_out_mprj[46]
port 456 nsew
rlabel metal2 s 87050 0 87106 800 6 la_data_out_mprj[47]
port 457 nsew
rlabel metal2 s 74354 12200 74410 13000 6 la_data_out_mprj[48]
port 458 nsew
rlabel metal2 s 87418 0 87474 800 6 la_data_out_mprj[49]
port 459 nsew
rlabel metal2 s 74722 12200 74778 13000 6 la_data_out_mprj[4]
port 460 nsew
rlabel metal2 s 87786 0 87842 800 6 la_data_out_mprj[50]
port 461 nsew
rlabel metal2 s 75090 12200 75146 13000 6 la_data_out_mprj[51]
port 462 nsew
rlabel metal2 s 88154 0 88210 800 6 la_data_out_mprj[52]
port 463 nsew
rlabel metal2 s 75458 12200 75514 13000 6 la_data_out_mprj[53]
port 464 nsew
rlabel metal2 s 88522 0 88578 800 6 la_data_out_mprj[54]
port 465 nsew
rlabel metal2 s 75826 12200 75882 13000 6 la_data_out_mprj[55]
port 466 nsew
rlabel metal2 s 88890 0 88946 800 6 la_data_out_mprj[56]
port 467 nsew
rlabel metal2 s 76194 12200 76250 13000 6 la_data_out_mprj[57]
port 468 nsew
rlabel metal2 s 89258 0 89314 800 6 la_data_out_mprj[58]
port 469 nsew
rlabel metal2 s 76562 12200 76618 13000 6 la_data_out_mprj[59]
port 470 nsew
rlabel metal2 s 89626 0 89682 800 6 la_data_out_mprj[5]
port 471 nsew
rlabel metal2 s 76930 12200 76986 13000 6 la_data_out_mprj[60]
port 472 nsew
rlabel metal2 s 89994 0 90050 800 6 la_data_out_mprj[61]
port 473 nsew
rlabel metal2 s 77298 12200 77354 13000 6 la_data_out_mprj[62]
port 474 nsew
rlabel metal2 s 90362 0 90418 800 6 la_data_out_mprj[63]
port 475 nsew
rlabel metal2 s 77666 12200 77722 13000 6 la_data_out_mprj[64]
port 476 nsew
rlabel metal2 s 90730 0 90786 800 6 la_data_out_mprj[65]
port 477 nsew
rlabel metal2 s 78034 12200 78090 13000 6 la_data_out_mprj[66]
port 478 nsew
rlabel metal2 s 91098 0 91154 800 6 la_data_out_mprj[67]
port 479 nsew
rlabel metal2 s 78402 12200 78458 13000 6 la_data_out_mprj[68]
port 480 nsew
rlabel metal2 s 91466 0 91522 800 6 la_data_out_mprj[69]
port 481 nsew
rlabel metal2 s 78770 12200 78826 13000 6 la_data_out_mprj[6]
port 482 nsew
rlabel metal2 s 91834 0 91890 800 6 la_data_out_mprj[70]
port 483 nsew
rlabel metal2 s 79138 12200 79194 13000 6 la_data_out_mprj[71]
port 484 nsew
rlabel metal2 s 92202 0 92258 800 6 la_data_out_mprj[72]
port 485 nsew
rlabel metal2 s 79506 12200 79562 13000 6 la_data_out_mprj[73]
port 486 nsew
rlabel metal2 s 92570 0 92626 800 6 la_data_out_mprj[74]
port 487 nsew
rlabel metal2 s 79874 12200 79930 13000 6 la_data_out_mprj[75]
port 488 nsew
rlabel metal2 s 92938 0 92994 800 6 la_data_out_mprj[76]
port 489 nsew
rlabel metal2 s 80242 12200 80298 13000 6 la_data_out_mprj[77]
port 490 nsew
rlabel metal2 s 93306 0 93362 800 6 la_data_out_mprj[78]
port 491 nsew
rlabel metal2 s 80610 12200 80666 13000 6 la_data_out_mprj[79]
port 492 nsew
rlabel metal2 s 93674 0 93730 800 6 la_data_out_mprj[7]
port 493 nsew
rlabel metal2 s 80978 12200 81034 13000 6 la_data_out_mprj[80]
port 494 nsew
rlabel metal2 s 94042 0 94098 800 6 la_data_out_mprj[81]
port 495 nsew
rlabel metal2 s 81346 12200 81402 13000 6 la_data_out_mprj[82]
port 496 nsew
rlabel metal2 s 94410 0 94466 800 6 la_data_out_mprj[83]
port 497 nsew
rlabel metal2 s 81714 12200 81770 13000 6 la_data_out_mprj[84]
port 498 nsew
rlabel metal2 s 94778 0 94834 800 6 la_data_out_mprj[85]
port 499 nsew
rlabel metal2 s 82082 12200 82138 13000 6 la_data_out_mprj[86]
port 500 nsew
rlabel metal2 s 95146 0 95202 800 6 la_data_out_mprj[87]
port 501 nsew
rlabel metal2 s 82450 12200 82506 13000 6 la_data_out_mprj[88]
port 502 nsew
rlabel metal2 s 95514 0 95570 800 6 la_data_out_mprj[89]
port 503 nsew
rlabel metal2 s 82818 12200 82874 13000 6 la_data_out_mprj[8]
port 504 nsew
rlabel metal2 s 95882 0 95938 800 6 la_data_out_mprj[90]
port 505 nsew
rlabel metal2 s 83186 12200 83242 13000 6 la_data_out_mprj[91]
port 506 nsew
rlabel metal2 s 96250 0 96306 800 6 la_data_out_mprj[92]
port 507 nsew
rlabel metal2 s 83554 12200 83610 13000 6 la_data_out_mprj[93]
port 508 nsew
rlabel metal2 s 96618 0 96674 800 6 la_data_out_mprj[94]
port 509 nsew
rlabel metal2 s 83922 12200 83978 13000 6 la_data_out_mprj[95]
port 510 nsew
rlabel metal2 s 96986 0 97042 800 6 la_data_out_mprj[96]
port 511 nsew
rlabel metal2 s 84290 12200 84346 13000 6 la_data_out_mprj[97]
port 512 nsew
rlabel metal2 s 97354 0 97410 800 6 la_data_out_mprj[98]
port 513 nsew
rlabel metal2 s 84658 12200 84714 13000 6 la_data_out_mprj[99]
port 514 nsew
rlabel metal2 s 97722 0 97778 800 6 la_data_out_mprj[9]
port 515 nsew
rlabel metal2 s 85026 12200 85082 13000 6 la_oen_core[0]
port 516 nsew
rlabel metal2 s 85394 12200 85450 13000 6 la_oen_core[100]
port 517 nsew
rlabel metal2 s 85762 12200 85818 13000 6 la_oen_core[101]
port 518 nsew
rlabel metal2 s 86130 12200 86186 13000 6 la_oen_core[102]
port 519 nsew
rlabel metal2 s 86498 12200 86554 13000 6 la_oen_core[103]
port 520 nsew
rlabel metal2 s 86866 12200 86922 13000 6 la_oen_core[104]
port 521 nsew
rlabel metal2 s 87234 12200 87290 13000 6 la_oen_core[105]
port 522 nsew
rlabel metal2 s 87602 12200 87658 13000 6 la_oen_core[106]
port 523 nsew
rlabel metal2 s 87970 12200 88026 13000 6 la_oen_core[107]
port 524 nsew
rlabel metal2 s 88338 12200 88394 13000 6 la_oen_core[108]
port 525 nsew
rlabel metal2 s 88706 12200 88762 13000 6 la_oen_core[109]
port 526 nsew
rlabel metal2 s 89074 12200 89130 13000 6 la_oen_core[10]
port 527 nsew
rlabel metal2 s 89442 12200 89498 13000 6 la_oen_core[110]
port 528 nsew
rlabel metal2 s 89810 12200 89866 13000 6 la_oen_core[111]
port 529 nsew
rlabel metal2 s 90178 12200 90234 13000 6 la_oen_core[112]
port 530 nsew
rlabel metal2 s 90546 12200 90602 13000 6 la_oen_core[113]
port 531 nsew
rlabel metal2 s 90914 12200 90970 13000 6 la_oen_core[114]
port 532 nsew
rlabel metal2 s 91282 12200 91338 13000 6 la_oen_core[115]
port 533 nsew
rlabel metal2 s 91650 12200 91706 13000 6 la_oen_core[116]
port 534 nsew
rlabel metal2 s 92018 12200 92074 13000 6 la_oen_core[117]
port 535 nsew
rlabel metal2 s 92386 12200 92442 13000 6 la_oen_core[118]
port 536 nsew
rlabel metal2 s 92754 12200 92810 13000 6 la_oen_core[119]
port 537 nsew
rlabel metal2 s 93122 12200 93178 13000 6 la_oen_core[11]
port 538 nsew
rlabel metal2 s 93490 12200 93546 13000 6 la_oen_core[120]
port 539 nsew
rlabel metal2 s 93858 12200 93914 13000 6 la_oen_core[121]
port 540 nsew
rlabel metal2 s 94226 12200 94282 13000 6 la_oen_core[122]
port 541 nsew
rlabel metal2 s 94594 12200 94650 13000 6 la_oen_core[123]
port 542 nsew
rlabel metal2 s 94962 12200 95018 13000 6 la_oen_core[124]
port 543 nsew
rlabel metal2 s 95330 12200 95386 13000 6 la_oen_core[125]
port 544 nsew
rlabel metal2 s 95698 12200 95754 13000 6 la_oen_core[126]
port 545 nsew
rlabel metal2 s 96066 12200 96122 13000 6 la_oen_core[127]
port 546 nsew
rlabel metal2 s 96434 12200 96490 13000 6 la_oen_core[12]
port 547 nsew
rlabel metal2 s 96802 12200 96858 13000 6 la_oen_core[13]
port 548 nsew
rlabel metal2 s 97170 12200 97226 13000 6 la_oen_core[14]
port 549 nsew
rlabel metal2 s 97538 12200 97594 13000 6 la_oen_core[15]
port 550 nsew
rlabel metal2 s 97906 12200 97962 13000 6 la_oen_core[16]
port 551 nsew
rlabel metal2 s 98274 12200 98330 13000 6 la_oen_core[17]
port 552 nsew
rlabel metal2 s 98642 12200 98698 13000 6 la_oen_core[18]
port 553 nsew
rlabel metal2 s 99010 12200 99066 13000 6 la_oen_core[19]
port 554 nsew
rlabel metal2 s 99378 12200 99434 13000 6 la_oen_core[1]
port 555 nsew
rlabel metal2 s 99746 12200 99802 13000 6 la_oen_core[20]
port 556 nsew
rlabel metal2 s 100114 12200 100170 13000 6 la_oen_core[21]
port 557 nsew
rlabel metal2 s 100482 12200 100538 13000 6 la_oen_core[22]
port 558 nsew
rlabel metal2 s 100850 12200 100906 13000 6 la_oen_core[23]
port 559 nsew
rlabel metal2 s 101218 12200 101274 13000 6 la_oen_core[24]
port 560 nsew
rlabel metal2 s 101586 12200 101642 13000 6 la_oen_core[25]
port 561 nsew
rlabel metal2 s 101954 12200 102010 13000 6 la_oen_core[26]
port 562 nsew
rlabel metal2 s 102322 12200 102378 13000 6 la_oen_core[27]
port 563 nsew
rlabel metal2 s 102690 12200 102746 13000 6 la_oen_core[28]
port 564 nsew
rlabel metal2 s 103058 12200 103114 13000 6 la_oen_core[29]
port 565 nsew
rlabel metal2 s 103426 12200 103482 13000 6 la_oen_core[2]
port 566 nsew
rlabel metal2 s 103794 12200 103850 13000 6 la_oen_core[30]
port 567 nsew
rlabel metal2 s 104162 12200 104218 13000 6 la_oen_core[31]
port 568 nsew
rlabel metal2 s 104530 12200 104586 13000 6 la_oen_core[32]
port 569 nsew
rlabel metal2 s 104898 12200 104954 13000 6 la_oen_core[33]
port 570 nsew
rlabel metal2 s 105266 12200 105322 13000 6 la_oen_core[34]
port 571 nsew
rlabel metal2 s 105634 12200 105690 13000 6 la_oen_core[35]
port 572 nsew
rlabel metal2 s 106002 12200 106058 13000 6 la_oen_core[36]
port 573 nsew
rlabel metal2 s 106370 12200 106426 13000 6 la_oen_core[37]
port 574 nsew
rlabel metal2 s 106738 12200 106794 13000 6 la_oen_core[38]
port 575 nsew
rlabel metal2 s 107106 12200 107162 13000 6 la_oen_core[39]
port 576 nsew
rlabel metal2 s 107474 12200 107530 13000 6 la_oen_core[3]
port 577 nsew
rlabel metal2 s 107842 12200 107898 13000 6 la_oen_core[40]
port 578 nsew
rlabel metal2 s 108210 12200 108266 13000 6 la_oen_core[41]
port 579 nsew
rlabel metal2 s 108578 12200 108634 13000 6 la_oen_core[42]
port 580 nsew
rlabel metal2 s 108946 12200 109002 13000 6 la_oen_core[43]
port 581 nsew
rlabel metal2 s 109314 12200 109370 13000 6 la_oen_core[44]
port 582 nsew
rlabel metal2 s 109682 12200 109738 13000 6 la_oen_core[45]
port 583 nsew
rlabel metal2 s 110050 12200 110106 13000 6 la_oen_core[46]
port 584 nsew
rlabel metal2 s 110418 12200 110474 13000 6 la_oen_core[47]
port 585 nsew
rlabel metal2 s 110786 12200 110842 13000 6 la_oen_core[48]
port 586 nsew
rlabel metal2 s 98090 0 98146 800 6 la_oen_core[49]
port 587 nsew
rlabel metal2 s 111154 12200 111210 13000 6 la_oen_core[4]
port 588 nsew
rlabel metal2 s 98458 0 98514 800 6 la_oen_core[50]
port 589 nsew
rlabel metal2 s 111522 12200 111578 13000 6 la_oen_core[51]
port 590 nsew
rlabel metal2 s 98826 0 98882 800 6 la_oen_core[52]
port 591 nsew
rlabel metal2 s 111890 12200 111946 13000 6 la_oen_core[53]
port 592 nsew
rlabel metal2 s 99194 0 99250 800 6 la_oen_core[54]
port 593 nsew
rlabel metal2 s 112258 12200 112314 13000 6 la_oen_core[55]
port 594 nsew
rlabel metal2 s 99562 0 99618 800 6 la_oen_core[56]
port 595 nsew
rlabel metal2 s 112626 12200 112682 13000 6 la_oen_core[57]
port 596 nsew
rlabel metal2 s 99930 0 99986 800 6 la_oen_core[58]
port 597 nsew
rlabel metal2 s 112994 12200 113050 13000 6 la_oen_core[59]
port 598 nsew
rlabel metal2 s 100298 0 100354 800 6 la_oen_core[5]
port 599 nsew
rlabel metal2 s 113362 12200 113418 13000 6 la_oen_core[60]
port 600 nsew
rlabel metal2 s 100666 0 100722 800 6 la_oen_core[61]
port 601 nsew
rlabel metal2 s 113730 12200 113786 13000 6 la_oen_core[62]
port 602 nsew
rlabel metal2 s 101034 0 101090 800 6 la_oen_core[63]
port 603 nsew
rlabel metal2 s 114098 12200 114154 13000 6 la_oen_core[64]
port 604 nsew
rlabel metal2 s 101402 0 101458 800 6 la_oen_core[65]
port 605 nsew
rlabel metal2 s 114466 12200 114522 13000 6 la_oen_core[66]
port 606 nsew
rlabel metal2 s 101770 0 101826 800 6 la_oen_core[67]
port 607 nsew
rlabel metal2 s 114834 12200 114890 13000 6 la_oen_core[68]
port 608 nsew
rlabel metal2 s 102138 0 102194 800 6 la_oen_core[69]
port 609 nsew
rlabel metal2 s 115202 12200 115258 13000 6 la_oen_core[6]
port 610 nsew
rlabel metal2 s 102506 0 102562 800 6 la_oen_core[70]
port 611 nsew
rlabel metal2 s 115570 12200 115626 13000 6 la_oen_core[71]
port 612 nsew
rlabel metal2 s 102874 0 102930 800 6 la_oen_core[72]
port 613 nsew
rlabel metal2 s 115938 12200 115994 13000 6 la_oen_core[73]
port 614 nsew
rlabel metal2 s 103242 0 103298 800 6 la_oen_core[74]
port 615 nsew
rlabel metal2 s 116306 12200 116362 13000 6 la_oen_core[75]
port 616 nsew
rlabel metal2 s 103610 0 103666 800 6 la_oen_core[76]
port 617 nsew
rlabel metal2 s 116674 12200 116730 13000 6 la_oen_core[77]
port 618 nsew
rlabel metal2 s 103978 0 104034 800 6 la_oen_core[78]
port 619 nsew
rlabel metal2 s 117042 12200 117098 13000 6 la_oen_core[79]
port 620 nsew
rlabel metal2 s 104346 0 104402 800 6 la_oen_core[7]
port 621 nsew
rlabel metal2 s 117410 12200 117466 13000 6 la_oen_core[80]
port 622 nsew
rlabel metal2 s 104714 0 104770 800 6 la_oen_core[81]
port 623 nsew
rlabel metal2 s 117778 12200 117834 13000 6 la_oen_core[82]
port 624 nsew
rlabel metal2 s 105082 0 105138 800 6 la_oen_core[83]
port 625 nsew
rlabel metal2 s 118146 12200 118202 13000 6 la_oen_core[84]
port 626 nsew
rlabel metal2 s 105450 0 105506 800 6 la_oen_core[85]
port 627 nsew
rlabel metal2 s 118514 12200 118570 13000 6 la_oen_core[86]
port 628 nsew
rlabel metal2 s 105818 0 105874 800 6 la_oen_core[87]
port 629 nsew
rlabel metal2 s 118882 12200 118938 13000 6 la_oen_core[88]
port 630 nsew
rlabel metal2 s 106186 0 106242 800 6 la_oen_core[89]
port 631 nsew
rlabel metal2 s 119250 12200 119306 13000 6 la_oen_core[8]
port 632 nsew
rlabel metal2 s 106554 0 106610 800 6 la_oen_core[90]
port 633 nsew
rlabel metal2 s 119618 12200 119674 13000 6 la_oen_core[91]
port 634 nsew
rlabel metal2 s 106922 0 106978 800 6 la_oen_core[92]
port 635 nsew
rlabel metal2 s 119986 12200 120042 13000 6 la_oen_core[93]
port 636 nsew
rlabel metal2 s 107290 0 107346 800 6 la_oen_core[94]
port 637 nsew
rlabel metal2 s 120354 12200 120410 13000 6 la_oen_core[95]
port 638 nsew
rlabel metal2 s 107658 0 107714 800 6 la_oen_core[96]
port 639 nsew
rlabel metal2 s 120722 12200 120778 13000 6 la_oen_core[97]
port 640 nsew
rlabel metal2 s 108026 0 108082 800 6 la_oen_core[98]
port 641 nsew
rlabel metal2 s 121090 12200 121146 13000 6 la_oen_core[99]
port 642 nsew
rlabel metal2 s 108394 0 108450 800 6 la_oen_core[9]
port 643 nsew
rlabel metal2 s 108762 0 108818 800 6 la_oen_mprj[0]
port 644 nsew
rlabel metal2 s 109130 0 109186 800 6 la_oen_mprj[100]
port 645 nsew
rlabel metal2 s 109498 0 109554 800 6 la_oen_mprj[101]
port 646 nsew
rlabel metal2 s 109866 0 109922 800 6 la_oen_mprj[102]
port 647 nsew
rlabel metal2 s 110234 0 110290 800 6 la_oen_mprj[103]
port 648 nsew
rlabel metal2 s 110602 0 110658 800 6 la_oen_mprj[104]
port 649 nsew
rlabel metal2 s 110970 0 111026 800 6 la_oen_mprj[105]
port 650 nsew
rlabel metal2 s 111338 0 111394 800 6 la_oen_mprj[106]
port 651 nsew
rlabel metal2 s 111706 0 111762 800 6 la_oen_mprj[107]
port 652 nsew
rlabel metal2 s 112074 0 112130 800 6 la_oen_mprj[108]
port 653 nsew
rlabel metal2 s 112442 0 112498 800 6 la_oen_mprj[109]
port 654 nsew
rlabel metal2 s 112810 0 112866 800 6 la_oen_mprj[10]
port 655 nsew
rlabel metal2 s 113178 0 113234 800 6 la_oen_mprj[110]
port 656 nsew
rlabel metal2 s 113546 0 113602 800 6 la_oen_mprj[111]
port 657 nsew
rlabel metal2 s 113914 0 113970 800 6 la_oen_mprj[112]
port 658 nsew
rlabel metal2 s 114282 0 114338 800 6 la_oen_mprj[113]
port 659 nsew
rlabel metal2 s 114650 0 114706 800 6 la_oen_mprj[114]
port 660 nsew
rlabel metal2 s 115018 0 115074 800 6 la_oen_mprj[115]
port 661 nsew
rlabel metal2 s 115386 0 115442 800 6 la_oen_mprj[116]
port 662 nsew
rlabel metal2 s 115754 0 115810 800 6 la_oen_mprj[117]
port 663 nsew
rlabel metal2 s 116122 0 116178 800 6 la_oen_mprj[118]
port 664 nsew
rlabel metal2 s 116490 0 116546 800 6 la_oen_mprj[119]
port 665 nsew
rlabel metal2 s 116858 0 116914 800 6 la_oen_mprj[11]
port 666 nsew
rlabel metal2 s 117226 0 117282 800 6 la_oen_mprj[120]
port 667 nsew
rlabel metal2 s 117594 0 117650 800 6 la_oen_mprj[121]
port 668 nsew
rlabel metal2 s 117962 0 118018 800 6 la_oen_mprj[122]
port 669 nsew
rlabel metal2 s 118330 0 118386 800 6 la_oen_mprj[123]
port 670 nsew
rlabel metal2 s 118698 0 118754 800 6 la_oen_mprj[124]
port 671 nsew
rlabel metal2 s 119066 0 119122 800 6 la_oen_mprj[125]
port 672 nsew
rlabel metal2 s 119434 0 119490 800 6 la_oen_mprj[126]
port 673 nsew
rlabel metal2 s 119802 0 119858 800 6 la_oen_mprj[127]
port 674 nsew
rlabel metal2 s 120170 0 120226 800 6 la_oen_mprj[12]
port 675 nsew
rlabel metal2 s 120538 0 120594 800 6 la_oen_mprj[13]
port 676 nsew
rlabel metal2 s 120906 0 120962 800 6 la_oen_mprj[14]
port 677 nsew
rlabel metal2 s 121274 0 121330 800 6 la_oen_mprj[15]
port 678 nsew
rlabel metal2 s 121642 0 121698 800 6 la_oen_mprj[16]
port 679 nsew
rlabel metal2 s 122010 0 122066 800 6 la_oen_mprj[17]
port 680 nsew
rlabel metal2 s 122378 0 122434 800 6 la_oen_mprj[18]
port 681 nsew
rlabel metal2 s 122746 0 122802 800 6 la_oen_mprj[19]
port 682 nsew
rlabel metal2 s 123114 0 123170 800 6 la_oen_mprj[1]
port 683 nsew
rlabel metal2 s 123482 0 123538 800 6 la_oen_mprj[20]
port 684 nsew
rlabel metal2 s 123850 0 123906 800 6 la_oen_mprj[21]
port 685 nsew
rlabel metal2 s 124218 0 124274 800 6 la_oen_mprj[22]
port 686 nsew
rlabel metal2 s 124586 0 124642 800 6 la_oen_mprj[23]
port 687 nsew
rlabel metal2 s 124954 0 125010 800 6 la_oen_mprj[24]
port 688 nsew
rlabel metal2 s 125322 0 125378 800 6 la_oen_mprj[25]
port 689 nsew
rlabel metal2 s 125690 0 125746 800 6 la_oen_mprj[26]
port 690 nsew
rlabel metal2 s 126058 0 126114 800 6 la_oen_mprj[27]
port 691 nsew
rlabel metal2 s 126426 0 126482 800 6 la_oen_mprj[28]
port 692 nsew
rlabel metal2 s 126794 0 126850 800 6 la_oen_mprj[29]
port 693 nsew
rlabel metal2 s 127162 0 127218 800 6 la_oen_mprj[2]
port 694 nsew
rlabel metal2 s 127530 0 127586 800 6 la_oen_mprj[30]
port 695 nsew
rlabel metal2 s 127898 0 127954 800 6 la_oen_mprj[31]
port 696 nsew
rlabel metal2 s 128266 0 128322 800 6 la_oen_mprj[32]
port 697 nsew
rlabel metal2 s 128634 0 128690 800 6 la_oen_mprj[33]
port 698 nsew
rlabel metal2 s 129002 0 129058 800 6 la_oen_mprj[34]
port 699 nsew
rlabel metal2 s 129370 0 129426 800 6 la_oen_mprj[35]
port 700 nsew
rlabel metal2 s 129738 0 129794 800 6 la_oen_mprj[36]
port 701 nsew
rlabel metal2 s 130106 0 130162 800 6 la_oen_mprj[37]
port 702 nsew
rlabel metal2 s 130474 0 130530 800 6 la_oen_mprj[38]
port 703 nsew
rlabel metal2 s 130842 0 130898 800 6 la_oen_mprj[39]
port 704 nsew
rlabel metal2 s 131210 0 131266 800 6 la_oen_mprj[3]
port 705 nsew
rlabel metal2 s 131578 0 131634 800 6 la_oen_mprj[40]
port 706 nsew
rlabel metal2 s 131946 0 132002 800 6 la_oen_mprj[41]
port 707 nsew
rlabel metal2 s 132314 0 132370 800 6 la_oen_mprj[42]
port 708 nsew
rlabel metal2 s 132682 0 132738 800 6 la_oen_mprj[43]
port 709 nsew
rlabel metal2 s 133050 0 133106 800 6 la_oen_mprj[44]
port 710 nsew
rlabel metal2 s 133418 0 133474 800 6 la_oen_mprj[45]
port 711 nsew
rlabel metal2 s 133786 0 133842 800 6 la_oen_mprj[46]
port 712 nsew
rlabel metal2 s 134154 0 134210 800 6 la_oen_mprj[47]
port 713 nsew
rlabel metal2 s 121458 12200 121514 13000 6 la_oen_mprj[48]
port 714 nsew
rlabel metal2 s 134522 0 134578 800 6 la_oen_mprj[49]
port 715 nsew
rlabel metal2 s 121826 12200 121882 13000 6 la_oen_mprj[4]
port 716 nsew
rlabel metal2 s 134890 0 134946 800 6 la_oen_mprj[50]
port 717 nsew
rlabel metal2 s 122194 12200 122250 13000 6 la_oen_mprj[51]
port 718 nsew
rlabel metal2 s 135258 0 135314 800 6 la_oen_mprj[52]
port 719 nsew
rlabel metal2 s 122562 12200 122618 13000 6 la_oen_mprj[53]
port 720 nsew
rlabel metal2 s 135626 0 135682 800 6 la_oen_mprj[54]
port 721 nsew
rlabel metal2 s 122930 12200 122986 13000 6 la_oen_mprj[55]
port 722 nsew
rlabel metal2 s 135994 0 136050 800 6 la_oen_mprj[56]
port 723 nsew
rlabel metal2 s 123298 12200 123354 13000 6 la_oen_mprj[57]
port 724 nsew
rlabel metal2 s 136362 0 136418 800 6 la_oen_mprj[58]
port 725 nsew
rlabel metal2 s 123666 12200 123722 13000 6 la_oen_mprj[59]
port 726 nsew
rlabel metal2 s 136730 0 136786 800 6 la_oen_mprj[5]
port 727 nsew
rlabel metal2 s 124034 12200 124090 13000 6 la_oen_mprj[60]
port 728 nsew
rlabel metal2 s 137098 0 137154 800 6 la_oen_mprj[61]
port 729 nsew
rlabel metal2 s 124402 12200 124458 13000 6 la_oen_mprj[62]
port 730 nsew
rlabel metal2 s 137466 0 137522 800 6 la_oen_mprj[63]
port 731 nsew
rlabel metal2 s 124770 12200 124826 13000 6 la_oen_mprj[64]
port 732 nsew
rlabel metal2 s 137834 0 137890 800 6 la_oen_mprj[65]
port 733 nsew
rlabel metal2 s 125138 12200 125194 13000 6 la_oen_mprj[66]
port 734 nsew
rlabel metal2 s 138202 0 138258 800 6 la_oen_mprj[67]
port 735 nsew
rlabel metal2 s 125506 12200 125562 13000 6 la_oen_mprj[68]
port 736 nsew
rlabel metal2 s 138570 0 138626 800 6 la_oen_mprj[69]
port 737 nsew
rlabel metal2 s 125874 12200 125930 13000 6 la_oen_mprj[6]
port 738 nsew
rlabel metal2 s 138938 0 138994 800 6 la_oen_mprj[70]
port 739 nsew
rlabel metal2 s 126242 12200 126298 13000 6 la_oen_mprj[71]
port 740 nsew
rlabel metal2 s 139306 0 139362 800 6 la_oen_mprj[72]
port 741 nsew
rlabel metal2 s 126610 12200 126666 13000 6 la_oen_mprj[73]
port 742 nsew
rlabel metal2 s 139674 0 139730 800 6 la_oen_mprj[74]
port 743 nsew
rlabel metal2 s 126978 12200 127034 13000 6 la_oen_mprj[75]
port 744 nsew
rlabel metal2 s 140042 0 140098 800 6 la_oen_mprj[76]
port 745 nsew
rlabel metal2 s 127346 12200 127402 13000 6 la_oen_mprj[77]
port 746 nsew
rlabel metal2 s 140410 0 140466 800 6 la_oen_mprj[78]
port 747 nsew
rlabel metal2 s 127714 12200 127770 13000 6 la_oen_mprj[79]
port 748 nsew
rlabel metal2 s 140778 0 140834 800 6 la_oen_mprj[7]
port 749 nsew
rlabel metal2 s 128082 12200 128138 13000 6 la_oen_mprj[80]
port 750 nsew
rlabel metal2 s 141146 0 141202 800 6 la_oen_mprj[81]
port 751 nsew
rlabel metal2 s 128450 12200 128506 13000 6 la_oen_mprj[82]
port 752 nsew
rlabel metal2 s 141514 0 141570 800 6 la_oen_mprj[83]
port 753 nsew
rlabel metal2 s 128818 12200 128874 13000 6 la_oen_mprj[84]
port 754 nsew
rlabel metal2 s 141882 0 141938 800 6 la_oen_mprj[85]
port 755 nsew
rlabel metal2 s 129186 12200 129242 13000 6 la_oen_mprj[86]
port 756 nsew
rlabel metal2 s 142250 0 142306 800 6 la_oen_mprj[87]
port 757 nsew
rlabel metal2 s 129554 12200 129610 13000 6 la_oen_mprj[88]
port 758 nsew
rlabel metal2 s 142618 0 142674 800 6 la_oen_mprj[89]
port 759 nsew
rlabel metal2 s 129922 12200 129978 13000 6 la_oen_mprj[8]
port 760 nsew
rlabel metal2 s 142986 0 143042 800 6 la_oen_mprj[90]
port 761 nsew
rlabel metal2 s 130290 12200 130346 13000 6 la_oen_mprj[91]
port 762 nsew
rlabel metal2 s 143354 0 143410 800 6 la_oen_mprj[92]
port 763 nsew
rlabel metal2 s 130658 12200 130714 13000 6 la_oen_mprj[93]
port 764 nsew
rlabel metal2 s 143722 0 143778 800 6 la_oen_mprj[94]
port 765 nsew
rlabel metal2 s 131026 12200 131082 13000 6 la_oen_mprj[95]
port 766 nsew
rlabel metal2 s 144090 0 144146 800 6 la_oen_mprj[96]
port 767 nsew
rlabel metal2 s 131394 12200 131450 13000 6 la_oen_mprj[97]
port 768 nsew
rlabel metal2 s 144458 0 144514 800 6 la_oen_mprj[98]
port 769 nsew
rlabel metal2 s 131762 12200 131818 13000 6 la_oen_mprj[99]
port 770 nsew
rlabel metal2 s 144826 0 144882 800 6 la_oen_mprj[9]
port 771 nsew
rlabel metal2 s 132130 12200 132186 13000 6 mprj_adr_o_core[0]
port 772 nsew
rlabel metal2 s 145194 0 145250 800 6 mprj_adr_o_core[10]
port 773 nsew
rlabel metal2 s 132498 12200 132554 13000 6 mprj_adr_o_core[11]
port 774 nsew
rlabel metal2 s 145562 0 145618 800 6 mprj_adr_o_core[12]
port 775 nsew
rlabel metal2 s 132866 12200 132922 13000 6 mprj_adr_o_core[13]
port 776 nsew
rlabel metal2 s 145930 0 145986 800 6 mprj_adr_o_core[14]
port 777 nsew
rlabel metal2 s 133234 12200 133290 13000 6 mprj_adr_o_core[15]
port 778 nsew
rlabel metal2 s 146298 0 146354 800 6 mprj_adr_o_core[16]
port 779 nsew
rlabel metal2 s 133602 12200 133658 13000 6 mprj_adr_o_core[17]
port 780 nsew
rlabel metal2 s 146666 0 146722 800 6 mprj_adr_o_core[18]
port 781 nsew
rlabel metal2 s 133970 12200 134026 13000 6 mprj_adr_o_core[19]
port 782 nsew
rlabel metal2 s 147034 0 147090 800 6 mprj_adr_o_core[1]
port 783 nsew
rlabel metal2 s 134338 12200 134394 13000 6 mprj_adr_o_core[20]
port 784 nsew
rlabel metal2 s 147402 0 147458 800 6 mprj_adr_o_core[21]
port 785 nsew
rlabel metal2 s 134706 12200 134762 13000 6 mprj_adr_o_core[22]
port 786 nsew
rlabel metal2 s 147770 0 147826 800 6 mprj_adr_o_core[23]
port 787 nsew
rlabel metal2 s 135074 12200 135130 13000 6 mprj_adr_o_core[24]
port 788 nsew
rlabel metal2 s 148138 0 148194 800 6 mprj_adr_o_core[25]
port 789 nsew
rlabel metal2 s 135442 12200 135498 13000 6 mprj_adr_o_core[26]
port 790 nsew
rlabel metal2 s 148506 0 148562 800 6 mprj_adr_o_core[27]
port 791 nsew
rlabel metal2 s 135810 12200 135866 13000 6 mprj_adr_o_core[28]
port 792 nsew
rlabel metal2 s 148874 0 148930 800 6 mprj_adr_o_core[29]
port 793 nsew
rlabel metal2 s 136178 12200 136234 13000 6 mprj_adr_o_core[2]
port 794 nsew
rlabel metal2 s 149242 0 149298 800 6 mprj_adr_o_core[30]
port 795 nsew
rlabel metal2 s 136546 12200 136602 13000 6 mprj_adr_o_core[31]
port 796 nsew
rlabel metal2 s 149610 0 149666 800 6 mprj_adr_o_core[3]
port 797 nsew
rlabel metal2 s 136914 12200 136970 13000 6 mprj_adr_o_core[4]
port 798 nsew
rlabel metal2 s 149978 0 150034 800 6 mprj_adr_o_core[5]
port 799 nsew
rlabel metal2 s 137282 12200 137338 13000 6 mprj_adr_o_core[6]
port 800 nsew
rlabel metal2 s 150346 0 150402 800 6 mprj_adr_o_core[7]
port 801 nsew
rlabel metal2 s 137650 12200 137706 13000 6 mprj_adr_o_core[8]
port 802 nsew
rlabel metal2 s 150714 0 150770 800 6 mprj_adr_o_core[9]
port 803 nsew
rlabel metal2 s 138018 12200 138074 13000 6 mprj_adr_o_user[0]
port 804 nsew
rlabel metal2 s 138386 12200 138442 13000 6 mprj_adr_o_user[10]
port 805 nsew
rlabel metal2 s 138754 12200 138810 13000 6 mprj_adr_o_user[11]
port 806 nsew
rlabel metal2 s 139122 12200 139178 13000 6 mprj_adr_o_user[12]
port 807 nsew
rlabel metal2 s 139490 12200 139546 13000 6 mprj_adr_o_user[13]
port 808 nsew
rlabel metal2 s 139858 12200 139914 13000 6 mprj_adr_o_user[14]
port 809 nsew
rlabel metal2 s 140226 12200 140282 13000 6 mprj_adr_o_user[15]
port 810 nsew
rlabel metal2 s 140594 12200 140650 13000 6 mprj_adr_o_user[16]
port 811 nsew
rlabel metal2 s 140962 12200 141018 13000 6 mprj_adr_o_user[17]
port 812 nsew
rlabel metal2 s 141330 12200 141386 13000 6 mprj_adr_o_user[18]
port 813 nsew
rlabel metal2 s 141698 12200 141754 13000 6 mprj_adr_o_user[19]
port 814 nsew
rlabel metal2 s 142066 12200 142122 13000 6 mprj_adr_o_user[1]
port 815 nsew
rlabel metal2 s 142434 12200 142490 13000 6 mprj_adr_o_user[20]
port 816 nsew
rlabel metal2 s 142802 12200 142858 13000 6 mprj_adr_o_user[21]
port 817 nsew
rlabel metal2 s 143170 12200 143226 13000 6 mprj_adr_o_user[22]
port 818 nsew
rlabel metal2 s 143538 12200 143594 13000 6 mprj_adr_o_user[23]
port 819 nsew
rlabel metal2 s 143906 12200 143962 13000 6 mprj_adr_o_user[24]
port 820 nsew
rlabel metal2 s 144274 12200 144330 13000 6 mprj_adr_o_user[25]
port 821 nsew
rlabel metal2 s 144642 12200 144698 13000 6 mprj_adr_o_user[26]
port 822 nsew
rlabel metal2 s 145010 12200 145066 13000 6 mprj_adr_o_user[27]
port 823 nsew
rlabel metal2 s 145378 12200 145434 13000 6 mprj_adr_o_user[28]
port 824 nsew
rlabel metal2 s 145746 12200 145802 13000 6 mprj_adr_o_user[29]
port 825 nsew
rlabel metal2 s 146114 12200 146170 13000 6 mprj_adr_o_user[2]
port 826 nsew
rlabel metal2 s 146482 12200 146538 13000 6 mprj_adr_o_user[30]
port 827 nsew
rlabel metal2 s 146850 12200 146906 13000 6 mprj_adr_o_user[31]
port 828 nsew
rlabel metal2 s 147218 12200 147274 13000 6 mprj_adr_o_user[3]
port 829 nsew
rlabel metal2 s 147586 12200 147642 13000 6 mprj_adr_o_user[4]
port 830 nsew
rlabel metal2 s 147954 12200 148010 13000 6 mprj_adr_o_user[5]
port 831 nsew
rlabel metal2 s 148322 12200 148378 13000 6 mprj_adr_o_user[6]
port 832 nsew
rlabel metal2 s 148690 12200 148746 13000 6 mprj_adr_o_user[7]
port 833 nsew
rlabel metal2 s 149058 12200 149114 13000 6 mprj_adr_o_user[8]
port 834 nsew
rlabel metal2 s 149426 12200 149482 13000 6 mprj_adr_o_user[9]
port 835 nsew
rlabel metal2 s 151082 0 151138 800 6 mprj_cyc_o_core
port 836 nsew
rlabel metal2 s 149794 12200 149850 13000 6 mprj_cyc_o_user
port 837 nsew
rlabel metal2 s 151450 0 151506 800 6 mprj_dat_o_core[0]
port 838 nsew
rlabel metal2 s 151818 0 151874 800 6 mprj_dat_o_core[10]
port 839 nsew
rlabel metal2 s 152186 0 152242 800 6 mprj_dat_o_core[11]
port 840 nsew
rlabel metal2 s 152554 0 152610 800 6 mprj_dat_o_core[12]
port 841 nsew
rlabel metal2 s 152922 0 152978 800 6 mprj_dat_o_core[13]
port 842 nsew
rlabel metal2 s 153290 0 153346 800 6 mprj_dat_o_core[14]
port 843 nsew
rlabel metal2 s 153658 0 153714 800 6 mprj_dat_o_core[15]
port 844 nsew
rlabel metal2 s 154026 0 154082 800 6 mprj_dat_o_core[16]
port 845 nsew
rlabel metal2 s 154394 0 154450 800 6 mprj_dat_o_core[17]
port 846 nsew
rlabel metal2 s 154762 0 154818 800 6 mprj_dat_o_core[18]
port 847 nsew
rlabel metal2 s 155130 0 155186 800 6 mprj_dat_o_core[19]
port 848 nsew
rlabel metal2 s 155498 0 155554 800 6 mprj_dat_o_core[1]
port 849 nsew
rlabel metal2 s 155866 0 155922 800 6 mprj_dat_o_core[20]
port 850 nsew
rlabel metal2 s 156234 0 156290 800 6 mprj_dat_o_core[21]
port 851 nsew
rlabel metal2 s 156602 0 156658 800 6 mprj_dat_o_core[22]
port 852 nsew
rlabel metal2 s 156970 0 157026 800 6 mprj_dat_o_core[23]
port 853 nsew
rlabel metal2 s 157338 0 157394 800 6 mprj_dat_o_core[24]
port 854 nsew
rlabel metal2 s 157706 0 157762 800 6 mprj_dat_o_core[25]
port 855 nsew
rlabel metal2 s 158074 0 158130 800 6 mprj_dat_o_core[26]
port 856 nsew
rlabel metal2 s 158442 0 158498 800 6 mprj_dat_o_core[27]
port 857 nsew
rlabel metal2 s 158810 0 158866 800 6 mprj_dat_o_core[28]
port 858 nsew
rlabel metal2 s 159178 0 159234 800 6 mprj_dat_o_core[29]
port 859 nsew
rlabel metal2 s 159546 0 159602 800 6 mprj_dat_o_core[2]
port 860 nsew
rlabel metal2 s 159914 0 159970 800 6 mprj_dat_o_core[30]
port 861 nsew
rlabel metal2 s 160282 0 160338 800 6 mprj_dat_o_core[31]
port 862 nsew
rlabel metal2 s 160650 0 160706 800 6 mprj_dat_o_core[3]
port 863 nsew
rlabel metal2 s 161018 0 161074 800 6 mprj_dat_o_core[4]
port 864 nsew
rlabel metal2 s 161386 0 161442 800 6 mprj_dat_o_core[5]
port 865 nsew
rlabel metal2 s 161754 0 161810 800 6 mprj_dat_o_core[6]
port 866 nsew
rlabel metal2 s 162122 0 162178 800 6 mprj_dat_o_core[7]
port 867 nsew
rlabel metal2 s 162490 0 162546 800 6 mprj_dat_o_core[8]
port 868 nsew
rlabel metal2 s 162858 0 162914 800 6 mprj_dat_o_core[9]
port 869 nsew
rlabel metal2 s 150162 12200 150218 13000 6 mprj_dat_o_user[0]
port 870 nsew
rlabel metal2 s 150530 12200 150586 13000 6 mprj_dat_o_user[10]
port 871 nsew
rlabel metal2 s 150898 12200 150954 13000 6 mprj_dat_o_user[11]
port 872 nsew
rlabel metal2 s 151266 12200 151322 13000 6 mprj_dat_o_user[12]
port 873 nsew
rlabel metal2 s 151634 12200 151690 13000 6 mprj_dat_o_user[13]
port 874 nsew
rlabel metal2 s 152002 12200 152058 13000 6 mprj_dat_o_user[14]
port 875 nsew
rlabel metal2 s 152370 12200 152426 13000 6 mprj_dat_o_user[15]
port 876 nsew
rlabel metal2 s 152738 12200 152794 13000 6 mprj_dat_o_user[16]
port 877 nsew
rlabel metal2 s 153106 12200 153162 13000 6 mprj_dat_o_user[17]
port 878 nsew
rlabel metal2 s 153474 12200 153530 13000 6 mprj_dat_o_user[18]
port 879 nsew
rlabel metal2 s 153842 12200 153898 13000 6 mprj_dat_o_user[19]
port 880 nsew
rlabel metal2 s 154210 12200 154266 13000 6 mprj_dat_o_user[1]
port 881 nsew
rlabel metal2 s 154578 12200 154634 13000 6 mprj_dat_o_user[20]
port 882 nsew
rlabel metal2 s 154946 12200 155002 13000 6 mprj_dat_o_user[21]
port 883 nsew
rlabel metal2 s 155314 12200 155370 13000 6 mprj_dat_o_user[22]
port 884 nsew
rlabel metal2 s 155682 12200 155738 13000 6 mprj_dat_o_user[23]
port 885 nsew
rlabel metal2 s 156050 12200 156106 13000 6 mprj_dat_o_user[24]
port 886 nsew
rlabel metal2 s 156418 12200 156474 13000 6 mprj_dat_o_user[25]
port 887 nsew
rlabel metal2 s 156786 12200 156842 13000 6 mprj_dat_o_user[26]
port 888 nsew
rlabel metal2 s 157154 12200 157210 13000 6 mprj_dat_o_user[27]
port 889 nsew
rlabel metal2 s 157522 12200 157578 13000 6 mprj_dat_o_user[28]
port 890 nsew
rlabel metal2 s 157890 12200 157946 13000 6 mprj_dat_o_user[29]
port 891 nsew
rlabel metal2 s 158258 12200 158314 13000 6 mprj_dat_o_user[2]
port 892 nsew
rlabel metal2 s 158626 12200 158682 13000 6 mprj_dat_o_user[30]
port 893 nsew
rlabel metal2 s 158994 12200 159050 13000 6 mprj_dat_o_user[31]
port 894 nsew
rlabel metal2 s 159362 12200 159418 13000 6 mprj_dat_o_user[3]
port 895 nsew
rlabel metal2 s 159730 12200 159786 13000 6 mprj_dat_o_user[4]
port 896 nsew
rlabel metal2 s 160098 12200 160154 13000 6 mprj_dat_o_user[5]
port 897 nsew
rlabel metal2 s 160466 12200 160522 13000 6 mprj_dat_o_user[6]
port 898 nsew
rlabel metal2 s 160834 12200 160890 13000 6 mprj_dat_o_user[7]
port 899 nsew
rlabel metal2 s 161202 12200 161258 13000 6 mprj_dat_o_user[8]
port 900 nsew
rlabel metal2 s 161570 12200 161626 13000 6 mprj_dat_o_user[9]
port 901 nsew
rlabel metal2 s 163226 0 163282 800 6 mprj_sel_o_core[0]
port 902 nsew
rlabel metal2 s 163594 0 163650 800 6 mprj_sel_o_core[1]
port 903 nsew
rlabel metal2 s 163962 0 164018 800 6 mprj_sel_o_core[2]
port 904 nsew
rlabel metal2 s 164330 0 164386 800 6 mprj_sel_o_core[3]
port 905 nsew
rlabel metal2 s 161938 12200 161994 13000 6 mprj_sel_o_user[0]
port 906 nsew
rlabel metal2 s 162306 12200 162362 13000 6 mprj_sel_o_user[1]
port 907 nsew
rlabel metal2 s 162674 12200 162730 13000 6 mprj_sel_o_user[2]
port 908 nsew
rlabel metal2 s 163042 12200 163098 13000 6 mprj_sel_o_user[3]
port 909 nsew
rlabel metal2 s 164698 0 164754 800 6 mprj_stb_o_core
port 910 nsew
rlabel metal2 s 163410 12200 163466 13000 6 mprj_stb_o_user
port 911 nsew
rlabel metal2 s 165066 0 165122 800 6 mprj_we_o_core
port 912 nsew
rlabel metal2 s 163778 12200 163834 13000 6 mprj_we_o_user
port 913 nsew
rlabel metal2 s 165434 0 165490 800 6 user1_vcc_powergood
port 914 nsew
rlabel metal2 s 165802 0 165858 800 6 user1_vdd_powergood
port 915 nsew
rlabel metal2 s 166170 0 166226 800 6 user2_vcc_powergood
port 916 nsew
rlabel metal2 s 166538 0 166594 800 6 user2_vdd_powergood
port 917 nsew
rlabel metal2 s 164146 12200 164202 13000 6 user_clock
port 918 nsew
rlabel metal2 s 164514 12200 164570 13000 6 user_clock2
port 919 nsew
rlabel metal2 s 164882 12200 164938 13000 6 user_reset
port 920 nsew
rlabel metal2 s 754 0 810 800 6 user_resetn
port 921 nsew
rlabel metal1 s 368 11376 169556 11472 6 VPWR
port 922 nsew power default
rlabel metal1 s 368 11920 169556 12016 6 VGND
port 923 nsew ground default
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 169594 13025
string LEFview TRUE
<< end >>

