* NGSPICE file created from gpio_control_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

.subckt gpio_control_block mgmt_gpio_in mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en
+ pad_gpio_ana_pol pad_gpio_ana_sel pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover
+ pad_gpio_ib_mode_sel pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel
+ pad_gpio_vtrip_sel resetn serial_clock serial_data_in serial_data_out user_gpio_in
+ user_gpio_oeb user_gpio_out zero vccd vssd1 vccd1
XFILLER_9_55 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_062_ _064_/A vssd1 vssd1 vccd vccd _062_/X sky130_fd_sc_hd__buf_2
XFILLER_13_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_8
X_045_ _044_/A vssd1 vssd1 vccd vccd _045_/X sky130_fd_sc_hd__buf_2
XFILLER_15_7 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_36 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_061_ _064_/A vssd1 vssd1 vccd vccd _061_/X sky130_fd_sc_hd__buf_2
X_044_ _044_/A vssd1 vssd1 vccd vccd _044_/X sky130_fd_sc_hd__buf_2
X_060_ _064_/A vssd1 vssd1 vccd vccd _060_/X sky130_fd_sc_hd__buf_2
X_043_ _044_/A vssd1 vssd1 vccd vccd _043_/X sky130_fd_sc_hd__buf_2
XFILLER_15_45 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_042_ _041_/X vssd1 vssd1 vccd vccd _044_/A sky130_fd_sc_hd__buf_2
XFILLER_9_26 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_041_ _065_/A vssd1 vssd1 vccd vccd _041_/X sky130_fd_sc_hd__buf_2
XFILLER_15_36 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_49 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_040_ _081_/A resetn vssd1 vssd1 vccd vccd _065_/A sky130_fd_sc_hd__or2_4
XFILLER_1_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_099_ _081_/A _098_/Q _052_/X vssd1 vssd1 vccd vccd _099_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
Xconst_source vssd1 vssd1 vccd vccd one zero sky130_fd_sc_hd__conb_1
XFILLER_4_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_098_ _081_/A _084_/D _054_/X vssd1 vssd1 vccd vccd _098_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_63 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__tapvpwrvgnd_1_0 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_097_ _081_/A serial_data_in _055_/X vssd1 vssd1 vccd vccd _084_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_10_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_096_ _081_/X _105_/D _056_/X vssd1 vssd1 vccd vccd pad_gpio_ana_pol sky130_fd_sc_hd__dfrtp_4
XFILLER_1_7 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_079_ pad_gpio_in vssd1 vssd1 vccd vccd _079_/Y sky130_fd_sc_hd__inv_2
XPHY_4 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_40 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_095_ _081_/X _103_/Q _057_/X vssd1 vssd1 vccd vccd pad_gpio_ana_sel sky130_fd_sc_hd__dfrtp_4
X_078_ _084_/Q _076_/X _077_/Y _072_/Y user_gpio_out vssd1 vssd1 vccd vccd pad_gpio_out
+ sky130_fd_sc_hd__a32o_4
XFILLER_16_63 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_094_ _081_/X _102_/Q _058_/X vssd1 vssd1 vccd vccd pad_gpio_ana_en sky130_fd_sc_hd__dfrtp_4
X_077_ pad_gpio_dm[0] _075_/X vssd1 vssd1 vccd vccd _077_/Y sky130_fd_sc_hd__nand2_4
XPHY_6 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_32 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_093_ _081_/X serial_data_out _060_/X vssd1 vssd1 vccd vccd pad_gpio_dm[2] sky130_fd_sc_hd__dfstp_4
XFILLER_8_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_6
X_076_ mgmt_gpio_out _075_/X vssd1 vssd1 vccd vccd _076_/X sky130_fd_sc_hd__or2_4
XFILLER_16_32 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_8
XPHY_7 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_059_ _041_/X vssd1 vssd1 vccd vccd _064_/A sky130_fd_sc_hd__buf_2
XFILLER_13_11 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
Xgpio_in_buf _079_/Y gpio_in_buf/TE vssd1 vssd1 vccd vccd user_gpio_in sky130_fd_sc_hd__einvp_8
X_092_ _081_/X _109_/D _061_/X vssd1 vssd1 vccd vccd pad_gpio_dm[1] sky130_fd_sc_hd__dfstp_4
X_058_ _055_/A vssd1 vssd1 vccd vccd _058_/X sky130_fd_sc_hd__buf_2
X_075_ mgmt_gpio_oeb _075_/B pad_gpio_dm[1] vssd1 vssd1 vccd vccd _075_/X sky130_fd_sc_hd__and3_4
XPHY_8 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_44 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_091_ _081_/X _107_/Q _062_/X vssd1 vssd1 vccd vccd pad_gpio_dm[0] sky130_fd_sc_hd__dfrtp_4
X_074_ pad_gpio_dm[2] vssd1 vssd1 vccd vccd _075_/B sky130_fd_sc_hd__inv_2
X_057_ _055_/A vssd1 vssd1 vccd vccd _057_/X sky130_fd_sc_hd__buf_2
XPHY_9 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_36 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_109_ _081_/A _109_/D _082_/X vssd1 vssd1 vccd vccd serial_data_out sky130_fd_sc_hd__dfrtp_4
X_090_ _081_/X _098_/Q _063_/X vssd1 vssd1 vccd vccd _090_/Q sky130_fd_sc_hd__dfstp_4
X_073_ _090_/Q mgmt_gpio_oeb _084_/Q user_gpio_oeb _072_/Y vssd1 vssd1 vccd vccd pad_gpio_outenb
+ sky130_fd_sc_hd__a32o_4
X_056_ _055_/A vssd1 vssd1 vccd vccd _056_/X sky130_fd_sc_hd__buf_2
XFILLER_7_26 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_108_ _106_/CLK _107_/Q _044_/A vssd1 vssd1 vccd vccd _109_/D sky130_fd_sc_hd__dfrtp_4
X_072_ _084_/Q vssd1 vssd1 vccd vccd _072_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_59 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_25 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_6
X_055_ _055_/A vssd1 vssd1 vccd vccd _055_/X sky130_fd_sc_hd__buf_2
XFILLER_16_6 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_serial_clock clkbuf_0_serial_clock/X vssd1 vssd1 vccd vccd _081_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_107_ _081_/A _087_/D _043_/X vssd1 vssd1 vccd vccd _107_/Q sky130_fd_sc_hd__dfrtp_4
X_071_ pad_gpio_inenb vssd1 vssd1 vccd vccd _071_/X sky130_fd_sc_hd__buf_2
X_054_ _055_/A vssd1 vssd1 vccd vccd _054_/X sky130_fd_sc_hd__buf_2
X_106_ _106_/CLK _086_/D _044_/X vssd1 vssd1 vccd vccd _087_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_8_9 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_070_ _070_/A vssd1 vssd1 vccd vccd _070_/X sky130_fd_sc_hd__buf_2
X_053_ _041_/X vssd1 vssd1 vccd vccd _055_/A sky130_fd_sc_hd__buf_2
XFILLER_2_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_105_ _106_/CLK _105_/D _045_/X vssd1 vssd1 vccd vccd _086_/D sky130_fd_sc_hd__dfrtp_4
X_052_ _052_/A vssd1 vssd1 vccd vccd _052_/X sky130_fd_sc_hd__buf_2
X_104_ _106_/CLK _103_/Q _046_/X vssd1 vssd1 vccd vccd _105_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_12_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_30 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_051_ _052_/A vssd1 vssd1 vccd vccd _051_/X sky130_fd_sc_hd__buf_2
XFILLER_16_18 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_103_ _106_/CLK _102_/Q _048_/X vssd1 vssd1 vccd vccd _103_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_50 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_30 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_8
X_102_ _106_/CLK _089_/D _049_/X vssd1 vssd1 vccd vccd _102_/Q sky130_fd_sc_hd__dfrtp_4
X_050_ _052_/A vssd1 vssd1 vccd vccd _050_/X sky130_fd_sc_hd__buf_2
Xgpio_logic_high vssd1 vssd1 vccd1 vccd1 gpio_in_buf/TE gpio_logic_high/LO sky130_fd_sc_hd__conb_1
XFILLER_5_32 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XPHY_51 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_11 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_101_ _106_/CLK _100_/Q _050_/X vssd1 vssd1 vccd vccd _089_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_10_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XPHY_52 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_32 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_100_ _081_/A _099_/Q _051_/X vssd1 vssd1 vccd vccd _100_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_31 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_089_ _081_/X _089_/D _064_/X vssd1 vssd1 vccd vccd pad_gpio_ib_mode_sel sky130_fd_sc_hd__dfrtp_4
Xclkbuf_1_0_0_serial_clock clkbuf_0_serial_clock/X vssd1 vssd1 vccd vccd _106_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XPHY_33 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_serial_clock serial_clock vssd1 vssd1 vccd vccd clkbuf_0_serial_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XPHY_11 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_088_ _081_/X _100_/Q _066_/X vssd1 vssd1 vccd vccd pad_gpio_inenb sky130_fd_sc_hd__dfrtp_4
XFILLER_5_37 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_12 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_087_ _081_/X _087_/D _067_/X vssd1 vssd1 vccd vccd pad_gpio_vtrip_sel sky130_fd_sc_hd__dfrtp_4
XPHY_24 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_086_ _081_/X _086_/D _068_/X vssd1 vssd1 vccd vccd pad_gpio_slow_sel sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_49 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_069_ _070_/A vssd1 vssd1 vccd vccd _069_/X sky130_fd_sc_hd__buf_2
XPHY_25 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_085_ _081_/X _099_/Q _069_/X vssd1 vssd1 vccd vccd pad_gpio_holdover sky130_fd_sc_hd__dfrtp_4
X_068_ _070_/A vssd1 vssd1 vccd vccd _068_/X sky130_fd_sc_hd__buf_2
XPHY_48 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_067_ _070_/A vssd1 vssd1 vccd vccd _067_/X sky130_fd_sc_hd__buf_2
X_084_ _081_/X _084_/D _070_/X vssd1 vssd1 vccd vccd _084_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_63 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_18 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_4
XPHY_27 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_0 pad_gpio_inenb vssd1 vssd1 vccd vccd sky130_fd_sc_hd__diode_2
XPHY_38 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_30 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_083_ pad_gpio_in _071_/X vssd1 vssd1 vccd vccd mgmt_gpio_in sky130_fd_sc_hd__ebufn_2
X_049_ _052_/A vssd1 vssd1 vccd vccd _049_/X sky130_fd_sc_hd__buf_2
X_066_ _070_/A vssd1 vssd1 vccd vccd _066_/X sky130_fd_sc_hd__buf_2
XPHY_28 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_065_ _065_/A vssd1 vssd1 vccd vccd _070_/A sky130_fd_sc_hd__buf_2
XFILLER_12_62 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_2
X_082_ _041_/X vssd1 vssd1 vccd vccd _082_/X sky130_fd_sc_hd__buf_2
XFILLER_15_3 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_63 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__fill_1
X_048_ _052_/A vssd1 vssd1 vccd vccd _048_/X sky130_fd_sc_hd__buf_2
XPHY_29 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_081_ _081_/A _081_/B vssd1 vssd1 vccd vccd _081_/X sky130_fd_sc_hd__and2_4
XFILLER_12_52 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_6
X_064_ _064_/A vssd1 vssd1 vccd vccd _064_/X sky130_fd_sc_hd__buf_2
X_047_ _041_/X vssd1 vssd1 vccd vccd _052_/A sky130_fd_sc_hd__buf_2
XPHY_19 vssd1 vssd1 vccd vccd sky130_fd_sc_hd__decap_3
X_080_ resetn vssd1 vssd1 vccd vccd _081_/B sky130_fd_sc_hd__inv_2
X_063_ _064_/A vssd1 vssd1 vccd vccd _063_/X sky130_fd_sc_hd__buf_2
X_046_ _044_/A vssd1 vssd1 vccd vccd _046_/X sky130_fd_sc_hd__buf_2
.ends

