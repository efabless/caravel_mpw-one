VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_pll
  CLASS BLOCK ;
  FOREIGN digital_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 85.000 ;
  PIN clockp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 81.000 30.270 85.000 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 81.000 41.770 85.000 ;
    END
  END dco
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 81.000 55.570 85.000 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 17.040 75.000 17.640 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END div[4]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 81.000 69.370 85.000 ;
    END
  END enable
  PIN ext_trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 81.000 34.870 85.000 ;
    END
  END ext_trim[0]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END ext_trim[10]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END ext_trim[11]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 81.000 16.470 85.000 ;
    END
  END ext_trim[12]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 81.000 23.370 85.000 ;
    END
  END ext_trim[13]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END ext_trim[14]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END ext_trim[15]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 44.240 75.000 44.840 ;
    END
  END ext_trim[16]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END ext_trim[17]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 6.840 75.000 7.440 ;
    END
  END ext_trim[18]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 81.000 62.470 85.000 ;
    END
  END ext_trim[19]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END ext_trim[1]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END ext_trim[20]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END ext_trim[21]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 64.640 75.000 65.240 ;
    END
  END ext_trim[22]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 81.000 9.570 85.000 ;
    END
  END ext_trim[23]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 81.000 2.670 85.000 ;
    END
  END ext_trim[24]
  PIN ext_trim[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END ext_trim[25]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END ext_trim[2]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 81.000 48.670 85.000 ;
    END
  END ext_trim[3]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END ext_trim[4]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END ext_trim[5]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END ext_trim[6]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 54.440 75.000 55.040 ;
    END
  END ext_trim[7]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 23.840 75.000 24.440 ;
    END
  END ext_trim[8]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 74.840 75.000 75.440 ;
    END
  END ext_trim[9]
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 34.040 75.000 34.640 ;
    END
  END osc
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END resetb
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 61.040 5.200 62.640 79.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 79.120 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 41.040 5.200 42.640 79.120 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 69.460 78.965 ;
      LAYER met1 ;
        RECT 2.370 5.200 69.460 79.120 ;
      LAYER met2 ;
        RECT 2.950 80.720 9.010 81.000 ;
        RECT 9.850 80.720 15.910 81.000 ;
        RECT 16.750 80.720 22.810 81.000 ;
        RECT 23.650 80.720 29.710 81.000 ;
        RECT 30.550 80.720 34.310 81.000 ;
        RECT 35.150 80.720 41.210 81.000 ;
        RECT 42.050 80.720 48.110 81.000 ;
        RECT 48.950 80.720 55.010 81.000 ;
        RECT 55.850 80.720 61.910 81.000 ;
        RECT 62.750 80.720 68.810 81.000 ;
        RECT 2.400 4.280 69.370 80.720 ;
        RECT 2.950 4.000 6.710 4.280 ;
        RECT 7.550 4.000 13.610 4.280 ;
        RECT 14.450 4.000 20.510 4.280 ;
        RECT 21.350 4.000 27.410 4.280 ;
        RECT 28.250 4.000 34.310 4.280 ;
        RECT 35.150 4.000 41.210 4.280 ;
        RECT 42.050 4.000 48.110 4.280 ;
        RECT 48.950 4.000 55.010 4.280 ;
        RECT 55.850 4.000 61.910 4.280 ;
        RECT 62.750 4.000 68.810 4.280 ;
      LAYER met3 ;
        RECT 4.000 75.840 71.000 79.045 ;
        RECT 4.000 74.440 70.600 75.840 ;
        RECT 4.000 72.440 71.000 74.440 ;
        RECT 4.400 71.040 71.000 72.440 ;
        RECT 4.000 65.640 71.000 71.040 ;
        RECT 4.000 64.240 70.600 65.640 ;
        RECT 4.000 62.240 71.000 64.240 ;
        RECT 4.400 60.840 71.000 62.240 ;
        RECT 4.000 55.440 71.000 60.840 ;
        RECT 4.000 54.040 70.600 55.440 ;
        RECT 4.000 52.040 71.000 54.040 ;
        RECT 4.400 50.640 71.000 52.040 ;
        RECT 4.000 45.240 71.000 50.640 ;
        RECT 4.000 43.840 70.600 45.240 ;
        RECT 4.000 41.840 71.000 43.840 ;
        RECT 4.400 40.440 71.000 41.840 ;
        RECT 4.000 35.040 71.000 40.440 ;
        RECT 4.000 33.640 70.600 35.040 ;
        RECT 4.000 31.640 71.000 33.640 ;
        RECT 4.400 30.240 71.000 31.640 ;
        RECT 4.000 24.840 71.000 30.240 ;
        RECT 4.000 23.440 70.600 24.840 ;
        RECT 4.000 21.440 71.000 23.440 ;
        RECT 4.400 20.040 71.000 21.440 ;
        RECT 4.000 18.040 71.000 20.040 ;
        RECT 4.000 16.640 70.600 18.040 ;
        RECT 4.000 11.240 71.000 16.640 ;
        RECT 4.400 9.840 71.000 11.240 ;
        RECT 4.000 7.840 71.000 9.840 ;
        RECT 4.000 6.440 70.600 7.840 ;
        RECT 4.000 5.275 71.000 6.440 ;
  END
END digital_pll
END LIBRARY

