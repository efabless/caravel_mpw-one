magic
tech sky130A
magscale 1 2
timestamp 1625004077
<< metal1 >>
rect 585778 996412 585784 996464
rect 585836 996452 585842 996464
rect 674742 996452 674748 996464
rect 585836 996424 674748 996452
rect 585836 996412 585842 996424
rect 674742 996412 674748 996424
rect 674800 996412 674806 996464
rect 42242 996344 42248 996396
rect 42300 996384 42306 996396
rect 339494 996384 339500 996396
rect 42300 996356 339500 996384
rect 42300 996344 42306 996356
rect 339494 996344 339500 996356
rect 339552 996384 339558 996396
rect 673546 996384 673552 996396
rect 339552 996356 673552 996384
rect 339552 996344 339558 996356
rect 673546 996344 673552 996356
rect 673604 996344 673610 996396
rect 44910 990088 44916 990140
rect 44968 990128 44974 990140
rect 673638 990128 673644 990140
rect 44968 990100 673644 990128
rect 44968 990088 44974 990100
rect 673638 990088 673644 990100
rect 673696 990088 673702 990140
rect 42334 990020 42340 990072
rect 42392 990060 42398 990072
rect 673454 990060 673460 990072
rect 42392 990032 673460 990060
rect 42392 990020 42398 990032
rect 673454 990020 673460 990032
rect 673512 990020 673518 990072
rect 42426 861160 42432 861212
rect 42484 861200 42490 861212
rect 44174 861200 44180 861212
rect 42484 861172 44180 861200
rect 42484 861160 42490 861172
rect 44174 861160 44180 861172
rect 44232 861160 44238 861212
rect 673546 859120 673552 859172
rect 673604 859160 673610 859172
rect 675386 859160 675392 859172
rect 673604 859132 675392 859160
rect 673604 859120 673610 859132
rect 675386 859120 675392 859132
rect 675444 859120 675450 859172
rect 673638 856060 673644 856112
rect 673696 856100 673702 856112
rect 675386 856100 675392 856112
rect 673696 856072 675392 856100
rect 673696 856060 673702 856072
rect 675386 856060 675392 856072
rect 675444 856060 675450 856112
rect 673730 855380 673736 855432
rect 673788 855420 673794 855432
rect 675386 855420 675392 855432
rect 673788 855392 675392 855420
rect 673788 855380 673794 855392
rect 675386 855380 675392 855392
rect 675444 855380 675450 855432
rect 673454 849668 673460 849720
rect 673512 849708 673518 849720
rect 675386 849708 675392 849720
rect 673512 849680 675392 849708
rect 673512 849668 673518 849680
rect 675386 849668 675392 849680
rect 675444 849668 675450 849720
rect 675294 803768 675300 803820
rect 675352 803808 675358 803820
rect 677594 803808 677600 803820
rect 675352 803780 677600 803808
rect 675352 803768 675358 803780
rect 677594 803768 677600 803780
rect 677652 803768 677658 803820
rect 42242 800980 42248 801032
rect 42300 801020 42306 801032
rect 42610 801020 42616 801032
rect 42300 800992 42616 801020
rect 42300 800980 42306 800992
rect 42610 800980 42616 800992
rect 42668 800980 42674 801032
rect 41782 798532 41788 798584
rect 41840 798572 41846 798584
rect 42334 798572 42340 798584
rect 41840 798544 42340 798572
rect 41840 798532 41846 798544
rect 42334 798532 42340 798544
rect 42392 798532 42398 798584
rect 41782 792072 41788 792124
rect 41840 792112 41846 792124
rect 42426 792112 42432 792124
rect 41840 792084 42432 792112
rect 41840 792072 41846 792084
rect 42426 792072 42432 792084
rect 42484 792072 42490 792124
rect 41782 789080 41788 789132
rect 41840 789120 41846 789132
rect 42610 789120 42616 789132
rect 41840 789092 42616 789120
rect 41840 789080 41846 789092
rect 42610 789080 42616 789092
rect 42668 789080 42674 789132
rect 42242 787992 42248 788044
rect 42300 788032 42306 788044
rect 42426 788032 42432 788044
rect 42300 788004 42432 788032
rect 42300 787992 42306 788004
rect 42426 787992 42432 788004
rect 42484 787992 42490 788044
rect 673730 773304 673736 773356
rect 673788 773344 673794 773356
rect 675202 773344 675208 773356
rect 673788 773316 675208 773344
rect 673788 773304 673794 773316
rect 675202 773304 675208 773316
rect 675260 773344 675266 773356
rect 675386 773344 675392 773356
rect 675260 773316 675392 773344
rect 675260 773304 675266 773316
rect 675386 773304 675392 773316
rect 675444 773304 675450 773356
rect 673546 772760 673552 772812
rect 673604 772800 673610 772812
rect 675386 772800 675392 772812
rect 673604 772772 675392 772800
rect 673604 772760 673610 772772
rect 675386 772760 675392 772772
rect 675444 772760 675450 772812
rect 673638 769632 673644 769684
rect 673696 769672 673702 769684
rect 673914 769672 673920 769684
rect 673696 769644 673920 769672
rect 673696 769632 673702 769644
rect 673914 769632 673920 769644
rect 673972 769672 673978 769684
rect 675386 769672 675392 769684
rect 673972 769644 675392 769672
rect 673972 769632 673978 769644
rect 675386 769632 675392 769644
rect 675444 769632 675450 769684
rect 673730 769088 673736 769140
rect 673788 769128 673794 769140
rect 675202 769128 675208 769140
rect 673788 769100 675208 769128
rect 673788 769088 673794 769100
rect 675202 769088 675208 769100
rect 675260 769128 675266 769140
rect 675386 769128 675392 769140
rect 675260 769100 675392 769128
rect 675260 769088 675266 769100
rect 675386 769088 675392 769100
rect 675444 769088 675450 769140
rect 675202 767592 675208 767644
rect 675260 767632 675266 767644
rect 675386 767632 675392 767644
rect 675260 767604 675392 767632
rect 675260 767592 675266 767604
rect 675386 767592 675392 767604
rect 675444 767592 675450 767644
rect 673454 761268 673460 761320
rect 673512 761308 673518 761320
rect 674006 761308 674012 761320
rect 673512 761280 674012 761308
rect 673512 761268 673518 761280
rect 674006 761268 674012 761280
rect 674064 761308 674070 761320
rect 675386 761308 675392 761320
rect 674064 761280 675392 761308
rect 674064 761268 674070 761280
rect 675386 761268 675392 761280
rect 675444 761268 675450 761320
rect 675202 760180 675208 760232
rect 675260 760220 675266 760232
rect 675386 760220 675392 760232
rect 675260 760192 675392 760220
rect 675260 760180 675266 760192
rect 675386 760180 675392 760192
rect 675444 760180 675450 760232
rect 41782 756236 41788 756288
rect 41840 756276 41846 756288
rect 42334 756276 42340 756288
rect 41840 756248 42340 756276
rect 41840 756236 41846 756248
rect 42334 756236 42340 756248
rect 42392 756276 42398 756288
rect 42610 756276 42616 756288
rect 42392 756248 42616 756276
rect 42392 756236 42398 756248
rect 42610 756236 42616 756248
rect 42668 756236 42674 756288
rect 41782 748280 41788 748332
rect 41840 748320 41846 748332
rect 42518 748320 42524 748332
rect 41840 748292 42524 748320
rect 41840 748280 41846 748292
rect 42518 748280 42524 748292
rect 42576 748280 42582 748332
rect 41782 744812 41788 744864
rect 41840 744852 41846 744864
rect 42426 744852 42432 744864
rect 41840 744824 42432 744852
rect 41840 744812 41846 744824
rect 42426 744812 42432 744824
rect 42484 744852 42490 744864
rect 42702 744852 42708 744864
rect 42484 744824 42708 744852
rect 42484 744812 42490 744824
rect 42702 744812 42708 744824
rect 42760 744812 42766 744864
rect 673730 728560 673736 728612
rect 673788 728600 673794 728612
rect 675386 728600 675392 728612
rect 673788 728572 675392 728600
rect 673788 728560 673794 728572
rect 675386 728560 675392 728572
rect 675444 728560 675450 728612
rect 673546 728356 673552 728408
rect 673604 728396 673610 728408
rect 675386 728396 675392 728408
rect 673604 728368 675392 728396
rect 673604 728356 673610 728368
rect 675386 728356 675392 728368
rect 675444 728356 675450 728408
rect 673914 725228 673920 725280
rect 673972 725268 673978 725280
rect 675386 725268 675392 725280
rect 673972 725240 675392 725268
rect 673972 725228 673978 725240
rect 675386 725228 675392 725240
rect 675444 725228 675450 725280
rect 673454 724004 673460 724056
rect 673512 724044 673518 724056
rect 675386 724044 675392 724056
rect 673512 724016 675392 724044
rect 673512 724004 673518 724016
rect 675386 724004 675392 724016
rect 675444 724004 675450 724056
rect 673638 717816 673644 717868
rect 673696 717856 673702 717868
rect 674006 717856 674012 717868
rect 673696 717828 674012 717856
rect 673696 717816 673702 717828
rect 674006 717816 674012 717828
rect 674064 717856 674070 717868
rect 675386 717856 675392 717868
rect 674064 717828 675392 717856
rect 674064 717816 674070 717828
rect 675386 717816 675392 717828
rect 675444 717816 675450 717868
rect 41782 713056 41788 713108
rect 41840 713096 41846 713108
rect 42610 713096 42616 713108
rect 41840 713068 42616 713096
rect 41840 713056 41846 713068
rect 42610 713056 42616 713068
rect 42668 713056 42674 713108
rect 41782 704760 41788 704812
rect 41840 704800 41846 704812
rect 42518 704800 42524 704812
rect 41840 704772 42524 704800
rect 41840 704760 41846 704772
rect 42518 704760 42524 704772
rect 42576 704760 42582 704812
rect 41782 701632 41788 701684
rect 41840 701672 41846 701684
rect 42426 701672 42432 701684
rect 41840 701644 42432 701672
rect 41840 701632 41846 701644
rect 42426 701632 42432 701644
rect 42484 701632 42490 701684
rect 673454 684292 673460 684344
rect 673512 684332 673518 684344
rect 675294 684332 675300 684344
rect 673512 684304 675300 684332
rect 673512 684292 673518 684304
rect 675294 684292 675300 684304
rect 675352 684292 675358 684344
rect 673546 683068 673552 683120
rect 673604 683108 673610 683120
rect 673730 683108 673736 683120
rect 673604 683080 673736 683108
rect 673604 683068 673610 683080
rect 673730 683068 673736 683080
rect 673788 683108 673794 683120
rect 675386 683108 675392 683120
rect 673788 683080 675392 683108
rect 673788 683068 673794 683080
rect 675386 683068 675392 683080
rect 675444 683068 675450 683120
rect 673546 680416 673552 680468
rect 673604 680456 673610 680468
rect 673914 680456 673920 680468
rect 673604 680428 673920 680456
rect 673604 680416 673610 680428
rect 673914 680416 673920 680428
rect 673972 680456 673978 680468
rect 675386 680456 675392 680468
rect 673972 680428 675392 680456
rect 673972 680416 673978 680428
rect 675386 680416 675392 680428
rect 675444 680416 675450 680468
rect 673822 680076 673828 680128
rect 673880 680116 673886 680128
rect 675386 680116 675392 680128
rect 673880 680088 675392 680116
rect 673880 680076 673886 680088
rect 675386 680076 675392 680088
rect 675444 680076 675450 680128
rect 675202 678784 675208 678836
rect 675260 678824 675266 678836
rect 675386 678824 675392 678836
rect 675260 678796 675392 678824
rect 675260 678784 675266 678796
rect 675386 678784 675392 678796
rect 675444 678784 675450 678836
rect 673638 673616 673644 673668
rect 673696 673656 673702 673668
rect 674006 673656 674012 673668
rect 673696 673628 674012 673656
rect 673696 673616 673702 673628
rect 674006 673616 674012 673628
rect 674064 673656 674070 673668
rect 675386 673656 675392 673668
rect 674064 673628 675392 673656
rect 674064 673616 674070 673628
rect 675386 673616 675392 673628
rect 675444 673616 675450 673668
rect 41782 668720 41788 668772
rect 41840 668760 41846 668772
rect 42610 668760 42616 668772
rect 41840 668732 42616 668760
rect 41840 668720 41846 668732
rect 42610 668720 42616 668732
rect 42668 668720 42674 668772
rect 41782 661308 41788 661360
rect 41840 661348 41846 661360
rect 42518 661348 42524 661360
rect 41840 661320 42524 661348
rect 41840 661308 41846 661320
rect 42518 661308 42524 661320
rect 42576 661308 42582 661360
rect 41782 659268 41788 659320
rect 41840 659308 41846 659320
rect 42426 659308 42432 659320
rect 41840 659280 42432 659308
rect 41840 659268 41846 659280
rect 42426 659268 42432 659280
rect 42484 659308 42490 659320
rect 42702 659308 42708 659320
rect 42484 659280 42708 659308
rect 42484 659268 42490 659280
rect 42702 659268 42708 659280
rect 42760 659268 42766 659320
rect 673822 640092 673828 640144
rect 673880 640132 673886 640144
rect 675294 640132 675300 640144
rect 673880 640104 675300 640132
rect 673880 640092 673886 640104
rect 675294 640092 675300 640104
rect 675352 640092 675358 640144
rect 673638 638868 673644 638920
rect 673696 638908 673702 638920
rect 675386 638908 675392 638920
rect 673696 638880 675392 638908
rect 673696 638868 673702 638880
rect 675386 638868 675392 638880
rect 675444 638868 675450 638920
rect 673546 636284 673552 636336
rect 673604 636324 673610 636336
rect 675386 636324 675392 636336
rect 673604 636296 675392 636324
rect 673604 636284 673610 636296
rect 675386 636284 675392 636296
rect 675444 636284 675450 636336
rect 673730 635740 673736 635792
rect 673788 635780 673794 635792
rect 675294 635780 675300 635792
rect 673788 635752 675300 635780
rect 673788 635740 673794 635752
rect 675294 635740 675300 635752
rect 675352 635740 675358 635792
rect 675202 634584 675208 634636
rect 675260 634624 675266 634636
rect 675386 634624 675392 634636
rect 675260 634596 675392 634624
rect 675260 634584 675266 634596
rect 675386 634584 675392 634596
rect 675444 634584 675450 634636
rect 673454 629416 673460 629468
rect 673512 629456 673518 629468
rect 674006 629456 674012 629468
rect 673512 629428 674012 629456
rect 673512 629416 673518 629428
rect 674006 629416 674012 629428
rect 674064 629456 674070 629468
rect 675386 629456 675392 629468
rect 674064 629428 675392 629456
rect 674064 629416 674070 629428
rect 675386 629416 675392 629428
rect 675444 629416 675450 629468
rect 41782 625472 41788 625524
rect 41840 625512 41846 625524
rect 42610 625512 42616 625524
rect 41840 625484 42616 625512
rect 41840 625472 41846 625484
rect 42610 625472 42616 625484
rect 42668 625472 42674 625524
rect 41782 618128 41788 618180
rect 41840 618168 41846 618180
rect 42518 618168 42524 618180
rect 41840 618140 42524 618168
rect 41840 618128 41846 618140
rect 42518 618128 42524 618140
rect 42576 618128 42582 618180
rect 41782 615000 41788 615052
rect 41840 615040 41846 615052
rect 42702 615040 42708 615052
rect 41840 615012 42708 615040
rect 41840 615000 41846 615012
rect 42260 614712 42288 615012
rect 42702 615000 42708 615012
rect 42760 615000 42766 615052
rect 42242 614660 42248 614712
rect 42300 614660 42306 614712
rect 673730 596096 673736 596148
rect 673788 596136 673794 596148
rect 675202 596136 675208 596148
rect 673788 596108 675208 596136
rect 673788 596096 673794 596108
rect 675202 596096 675208 596108
rect 675260 596136 675266 596148
rect 675386 596136 675392 596148
rect 675260 596108 675392 596136
rect 675260 596096 675266 596108
rect 675386 596096 675392 596108
rect 675444 596096 675450 596148
rect 673638 595144 673644 595196
rect 673696 595184 673702 595196
rect 675386 595184 675392 595196
rect 673696 595156 675392 595184
rect 673696 595144 673702 595156
rect 675386 595144 675392 595156
rect 675444 595144 675450 595196
rect 673546 591880 673552 591932
rect 673604 591920 673610 591932
rect 675386 591920 675392 591932
rect 673604 591892 675392 591920
rect 673604 591880 673610 591892
rect 675386 591880 675392 591892
rect 675444 591880 675450 591932
rect 673730 590792 673736 590844
rect 673788 590832 673794 590844
rect 675202 590832 675208 590844
rect 673788 590804 675208 590832
rect 673788 590792 673794 590804
rect 675202 590792 675208 590804
rect 675260 590832 675266 590844
rect 675386 590832 675392 590844
rect 675260 590804 675392 590832
rect 675260 590792 675266 590804
rect 675386 590792 675392 590804
rect 675444 590792 675450 590844
rect 673454 584128 673460 584180
rect 673512 584168 673518 584180
rect 673914 584168 673920 584180
rect 673512 584140 673920 584168
rect 673512 584128 673518 584140
rect 673914 584128 673920 584140
rect 673972 584168 673978 584180
rect 675386 584168 675392 584180
rect 673972 584140 675392 584168
rect 673972 584128 673978 584140
rect 675386 584128 675392 584140
rect 675444 584128 675450 584180
rect 41782 583244 41788 583296
rect 41840 583284 41846 583296
rect 42610 583284 42616 583296
rect 41840 583256 42616 583284
rect 41840 583244 41846 583256
rect 42610 583244 42616 583256
rect 42668 583244 42674 583296
rect 41782 576512 41788 576564
rect 41840 576552 41846 576564
rect 42242 576552 42248 576564
rect 41840 576524 42248 576552
rect 41840 576512 41846 576524
rect 42242 576512 42248 576524
rect 42300 576552 42306 576564
rect 42426 576552 42432 576564
rect 42300 576524 42432 576552
rect 42300 576512 42306 576524
rect 42426 576512 42432 576524
rect 42484 576512 42490 576564
rect 41782 575900 41788 575952
rect 41840 575940 41846 575952
rect 42518 575940 42524 575952
rect 41840 575912 42524 575940
rect 41840 575900 41846 575912
rect 42518 575900 42524 575912
rect 42576 575900 42582 575952
rect 41782 571820 41788 571872
rect 41840 571860 41846 571872
rect 42426 571860 42432 571872
rect 41840 571832 42432 571860
rect 41840 571820 41846 571832
rect 42426 571820 42432 571832
rect 42484 571820 42490 571872
rect 673730 551488 673736 551540
rect 673788 551528 673794 551540
rect 675202 551528 675208 551540
rect 673788 551500 675208 551528
rect 673788 551488 673794 551500
rect 675202 551488 675208 551500
rect 675260 551488 675266 551540
rect 673638 551352 673644 551404
rect 673696 551392 673702 551404
rect 675386 551392 675392 551404
rect 673696 551364 675392 551392
rect 673696 551352 673702 551364
rect 675386 551352 675392 551364
rect 675444 551352 675450 551404
rect 673546 548224 673552 548276
rect 673604 548264 673610 548276
rect 675386 548264 675392 548276
rect 673604 548236 675392 548264
rect 673604 548224 673610 548236
rect 675386 548224 675392 548236
rect 675444 548224 675450 548276
rect 673454 547000 673460 547052
rect 673512 547040 673518 547052
rect 675202 547040 675208 547052
rect 673512 547012 675208 547040
rect 673512 547000 673518 547012
rect 675202 547000 675208 547012
rect 675260 547040 675266 547052
rect 675386 547040 675392 547052
rect 675260 547012 675392 547040
rect 675260 547000 675266 547012
rect 675386 547000 675392 547012
rect 675444 547000 675450 547052
rect 673914 540880 673920 540932
rect 673972 540920 673978 540932
rect 675386 540920 675392 540932
rect 673972 540892 675392 540920
rect 673972 540880 673978 540892
rect 675386 540880 675392 540892
rect 675444 540880 675450 540932
rect 41782 540064 41788 540116
rect 41840 540104 41846 540116
rect 42610 540104 42616 540116
rect 41840 540076 42616 540104
rect 41840 540064 41846 540076
rect 42610 540064 42616 540076
rect 42668 540064 42674 540116
rect 41782 531768 41788 531820
rect 41840 531808 41846 531820
rect 42518 531808 42524 531820
rect 41840 531780 42524 531808
rect 41840 531768 41846 531780
rect 42518 531768 42524 531780
rect 42576 531808 42582 531820
rect 42702 531808 42708 531820
rect 42576 531780 42708 531808
rect 42576 531768 42582 531780
rect 42702 531768 42708 531780
rect 42760 531768 42766 531820
rect 41782 528640 41788 528692
rect 41840 528680 41846 528692
rect 42426 528680 42432 528692
rect 41840 528652 42432 528680
rect 41840 528640 41846 528652
rect 42426 528640 42432 528652
rect 42484 528640 42490 528692
rect 675294 499468 675300 499520
rect 675352 499508 675358 499520
rect 676122 499508 676128 499520
rect 675352 499480 676128 499508
rect 675352 499468 675358 499480
rect 676122 499468 676128 499480
rect 676180 499468 676186 499520
rect 676122 494844 676128 494896
rect 676180 494884 676186 494896
rect 677962 494884 677968 494896
rect 676180 494856 677968 494884
rect 676180 494844 676186 494856
rect 677962 494844 677968 494856
rect 678020 494844 678026 494896
rect 674006 422220 674012 422272
rect 674064 422260 674070 422272
rect 674742 422260 674748 422272
rect 674064 422232 674748 422260
rect 674064 422220 674070 422232
rect 674742 422220 674748 422232
rect 674800 422220 674806 422272
rect 674006 419160 674012 419212
rect 674064 419200 674070 419212
rect 677502 419200 677508 419212
rect 674064 419172 677508 419200
rect 674064 419160 674070 419172
rect 677502 419160 677508 419172
rect 677560 419160 677566 419212
rect 41782 411272 41788 411324
rect 41840 411312 41846 411324
rect 42518 411312 42524 411324
rect 41840 411284 42524 411312
rect 41840 411272 41846 411284
rect 42518 411272 42524 411284
rect 42576 411272 42582 411324
rect 41782 404880 41788 404932
rect 41840 404920 41846 404932
rect 42702 404920 42708 404932
rect 41840 404892 42708 404920
rect 41840 404880 41846 404892
rect 42702 404880 42708 404892
rect 42760 404880 42766 404932
rect 41782 401888 41788 401940
rect 41840 401928 41846 401940
rect 42426 401928 42432 401940
rect 41840 401900 42432 401928
rect 41840 401888 41846 401900
rect 42426 401888 42432 401900
rect 42484 401888 42490 401940
rect 673914 376116 673920 376168
rect 673972 376156 673978 376168
rect 675386 376156 675392 376168
rect 673972 376128 675392 376156
rect 673972 376116 673978 376128
rect 675386 376116 675392 376128
rect 675444 376116 675450 376168
rect 673730 373056 673736 373108
rect 673788 373096 673794 373108
rect 675386 373096 675392 373108
rect 673788 373068 675392 373096
rect 673788 373056 673794 373068
rect 675386 373056 675392 373068
rect 675444 373056 675450 373108
rect 673546 372784 673552 372836
rect 673604 372824 673610 372836
rect 675386 372824 675392 372836
rect 673604 372796 675392 372824
rect 673604 372784 673610 372796
rect 675386 372784 675392 372796
rect 675444 372784 675450 372836
rect 41782 369044 41788 369096
rect 41840 369084 41846 369096
rect 42518 369084 42524 369096
rect 41840 369056 42524 369084
rect 41840 369044 41846 369056
rect 42518 369044 42524 369056
rect 42576 369044 42582 369096
rect 674006 365712 674012 365764
rect 674064 365752 674070 365764
rect 675386 365752 675392 365764
rect 674064 365724 675392 365752
rect 674064 365712 674070 365724
rect 675386 365712 675392 365724
rect 675444 365712 675450 365764
rect 41782 361292 41788 361344
rect 41840 361332 41846 361344
rect 42610 361332 42616 361344
rect 41840 361304 42616 361332
rect 41840 361292 41846 361304
rect 42610 361292 42616 361304
rect 42668 361292 42674 361344
rect 41782 357620 41788 357672
rect 41840 357660 41846 357672
rect 42426 357660 42432 357672
rect 41840 357632 42432 357660
rect 41840 357620 41846 357632
rect 42426 357620 42432 357632
rect 42484 357660 42490 357672
rect 42702 357660 42708 357672
rect 42484 357632 42708 357660
rect 42484 357620 42490 357632
rect 42702 357620 42708 357632
rect 42760 357620 42766 357672
rect 673730 333956 673736 334008
rect 673788 333996 673794 334008
rect 675202 333996 675208 334008
rect 673788 333968 675208 333996
rect 673788 333956 673794 333968
rect 675202 333956 675208 333968
rect 675260 333956 675266 334008
rect 673546 333072 673552 333124
rect 673604 333112 673610 333124
rect 675294 333112 675300 333124
rect 673604 333084 675300 333112
rect 673604 333072 673610 333084
rect 675294 333072 675300 333084
rect 675352 333072 675358 333124
rect 673454 331916 673460 331968
rect 673512 331956 673518 331968
rect 673914 331956 673920 331968
rect 673512 331928 673920 331956
rect 673512 331916 673518 331928
rect 673914 331916 673920 331928
rect 673972 331956 673978 331968
rect 675386 331956 675392 331968
rect 673972 331928 675392 331956
rect 673972 331916 673978 331928
rect 675386 331916 675392 331928
rect 675444 331916 675450 331968
rect 673546 328856 673552 328908
rect 673604 328896 673610 328908
rect 675202 328896 675208 328908
rect 673604 328868 675208 328896
rect 673604 328856 673610 328868
rect 675202 328856 675208 328868
rect 675260 328896 675266 328908
rect 675386 328896 675392 328908
rect 675260 328868 675392 328896
rect 675260 328856 675266 328868
rect 675386 328856 675392 328868
rect 675444 328856 675450 328908
rect 673730 328244 673736 328296
rect 673788 328284 673794 328296
rect 675386 328284 675392 328296
rect 673788 328256 675392 328284
rect 673788 328244 673794 328256
rect 675386 328244 675392 328256
rect 675444 328244 675450 328296
rect 41782 325660 41788 325712
rect 41840 325700 41846 325712
rect 42518 325700 42524 325712
rect 41840 325672 42524 325700
rect 41840 325660 41846 325672
rect 42518 325660 42524 325672
rect 42576 325660 42582 325712
rect 673638 322464 673644 322516
rect 673696 322504 673702 322516
rect 674006 322504 674012 322516
rect 673696 322476 674012 322504
rect 673696 322464 673702 322476
rect 674006 322464 674012 322476
rect 674064 322504 674070 322516
rect 675386 322504 675392 322516
rect 674064 322476 675392 322504
rect 674064 322464 674070 322476
rect 675386 322464 675392 322476
rect 675444 322464 675450 322516
rect 41782 317364 41788 317416
rect 41840 317404 41846 317416
rect 42610 317404 42616 317416
rect 41840 317376 42616 317404
rect 41840 317364 41846 317376
rect 42610 317364 42616 317376
rect 42668 317364 42674 317416
rect 41782 314236 41788 314288
rect 41840 314276 41846 314288
rect 42518 314276 42524 314288
rect 41840 314248 42524 314276
rect 41840 314236 41846 314248
rect 42518 314236 42524 314248
rect 42576 314276 42582 314288
rect 42702 314276 42708 314288
rect 42576 314248 42708 314276
rect 42576 314236 42582 314248
rect 42702 314236 42708 314248
rect 42760 314236 42766 314288
rect 42242 313080 42248 313132
rect 42300 313120 42306 313132
rect 42300 313092 42380 313120
rect 42300 313080 42306 313092
rect 42352 312928 42380 313092
rect 42334 312876 42340 312928
rect 42392 312876 42398 312928
rect 673730 289280 673736 289332
rect 673788 289320 673794 289332
rect 675386 289320 675392 289332
rect 673788 289292 675392 289320
rect 673788 289280 673794 289292
rect 675386 289280 675392 289292
rect 675444 289280 675450 289332
rect 673454 288736 673460 288788
rect 673512 288776 673518 288788
rect 675386 288776 675392 288788
rect 673512 288748 675392 288776
rect 673512 288736 673518 288748
rect 675386 288736 675392 288748
rect 675444 288736 675450 288788
rect 673546 285268 673552 285320
rect 673604 285308 673610 285320
rect 675386 285308 675392 285320
rect 673604 285280 675392 285308
rect 673604 285268 673610 285280
rect 675386 285268 675392 285280
rect 675444 285268 675450 285320
rect 42334 284112 42340 284164
rect 42392 284112 42398 284164
rect 42352 283960 42380 284112
rect 673730 284044 673736 284096
rect 673788 284084 673794 284096
rect 675386 284084 675392 284096
rect 673788 284056 675392 284084
rect 673788 284044 673794 284056
rect 675386 284044 675392 284056
rect 675444 284044 675450 284096
rect 42334 283908 42340 283960
rect 42392 283908 42398 283960
rect 41782 281528 41788 281580
rect 41840 281568 41846 281580
rect 42426 281568 42432 281580
rect 41840 281540 42432 281568
rect 41840 281528 41846 281540
rect 42426 281528 42432 281540
rect 42484 281568 42490 281580
rect 42702 281568 42708 281580
rect 42484 281540 42708 281568
rect 42484 281528 42490 281540
rect 42702 281528 42708 281540
rect 42760 281528 42766 281580
rect 673638 277312 673644 277364
rect 673696 277352 673702 277364
rect 675386 277352 675392 277364
rect 673696 277324 675392 277352
rect 673696 277312 673702 277324
rect 675386 277312 675392 277324
rect 675444 277312 675450 277364
rect 41782 274660 41788 274712
rect 41840 274700 41846 274712
rect 42610 274700 42616 274712
rect 41840 274672 42616 274700
rect 41840 274660 41846 274672
rect 42610 274660 42616 274672
rect 42668 274660 42674 274712
rect 41782 272076 41788 272128
rect 41840 272116 41846 272128
rect 42518 272116 42524 272128
rect 41840 272088 42524 272116
rect 41840 272076 41846 272088
rect 42518 272076 42524 272088
rect 42576 272076 42582 272128
rect 673730 244604 673736 244656
rect 673788 244644 673794 244656
rect 675386 244644 675392 244656
rect 673788 244616 675392 244644
rect 673788 244604 673794 244616
rect 675386 244604 675392 244616
rect 675444 244604 675450 244656
rect 673454 243720 673460 243772
rect 673512 243760 673518 243772
rect 675386 243760 675392 243772
rect 673512 243732 675392 243760
rect 673512 243720 673518 243732
rect 675386 243720 675392 243732
rect 675444 243720 675450 243772
rect 673546 240252 673552 240304
rect 673604 240292 673610 240304
rect 675386 240292 675392 240304
rect 673604 240264 675392 240292
rect 673604 240252 673610 240264
rect 675386 240252 675392 240264
rect 675444 240252 675450 240304
rect 673730 239640 673736 239692
rect 673788 239680 673794 239692
rect 675386 239680 675392 239692
rect 673788 239652 675392 239680
rect 673788 239640 673794 239652
rect 675386 239640 675392 239652
rect 675444 239640 675450 239692
rect 41782 238280 41788 238332
rect 41840 238320 41846 238332
rect 42426 238320 42432 238332
rect 41840 238292 42432 238320
rect 41840 238280 41846 238292
rect 42426 238280 42432 238292
rect 42484 238320 42490 238332
rect 42702 238320 42708 238332
rect 42484 238292 42708 238320
rect 42484 238280 42490 238292
rect 42702 238280 42708 238292
rect 42760 238280 42766 238332
rect 673638 233860 673644 233912
rect 673696 233900 673702 233912
rect 675386 233900 675392 233912
rect 673696 233872 675392 233900
rect 673696 233860 673702 233872
rect 675386 233860 675392 233872
rect 675444 233860 675450 233912
rect 41782 231888 41788 231940
rect 41840 231928 41846 231940
rect 42610 231928 42616 231940
rect 41840 231900 42616 231928
rect 41840 231888 41846 231900
rect 42610 231888 42616 231900
rect 42668 231888 42674 231940
rect 41782 228828 41788 228880
rect 41840 228868 41846 228880
rect 42518 228868 42524 228880
rect 41840 228840 42524 228868
rect 41840 228828 41846 228840
rect 42518 228828 42524 228840
rect 42576 228828 42582 228880
rect 673730 200404 673736 200456
rect 673788 200444 673794 200456
rect 675386 200444 675392 200456
rect 673788 200416 675392 200444
rect 673788 200404 673794 200416
rect 675386 200404 675392 200416
rect 675444 200404 675450 200456
rect 673454 199112 673460 199164
rect 673512 199152 673518 199164
rect 675386 199152 675392 199164
rect 673512 199124 675392 199152
rect 673512 199112 673518 199124
rect 675386 199112 675392 199124
rect 675444 199112 675450 199164
rect 673546 197004 673552 197056
rect 673604 197044 673610 197056
rect 675386 197044 675392 197056
rect 673604 197016 675392 197044
rect 673604 197004 673610 197016
rect 675386 197004 675392 197016
rect 675444 197004 675450 197056
rect 673730 195780 673736 195832
rect 673788 195820 673794 195832
rect 675386 195820 675392 195832
rect 673788 195792 675392 195820
rect 673788 195780 673794 195792
rect 675386 195780 675392 195792
rect 675444 195780 675450 195832
rect 41782 195100 41788 195152
rect 41840 195140 41846 195152
rect 42426 195140 42432 195152
rect 41840 195112 42432 195140
rect 41840 195100 41846 195112
rect 42426 195100 42432 195112
rect 42484 195100 42490 195152
rect 673638 189252 673644 189304
rect 673696 189292 673702 189304
rect 675386 189292 675392 189304
rect 673696 189264 675392 189292
rect 673696 189252 673702 189264
rect 675386 189252 675392 189264
rect 675444 189252 675450 189304
rect 41782 188708 41788 188760
rect 41840 188748 41846 188760
rect 42518 188748 42524 188760
rect 41840 188720 42524 188748
rect 41840 188708 41846 188720
rect 42518 188708 42524 188720
rect 42576 188748 42582 188760
rect 42794 188748 42800 188760
rect 42576 188720 42800 188748
rect 42576 188708 42582 188720
rect 42794 188708 42800 188720
rect 42852 188708 42858 188760
rect 41782 185648 41788 185700
rect 41840 185688 41846 185700
rect 42702 185688 42708 185700
rect 41840 185660 42708 185688
rect 41840 185648 41846 185660
rect 42702 185648 42708 185660
rect 42760 185648 42766 185700
rect 42242 184356 42248 184408
rect 42300 184396 42306 184408
rect 42702 184396 42708 184408
rect 42300 184368 42708 184396
rect 42300 184356 42306 184368
rect 42702 184356 42708 184368
rect 42760 184356 42766 184408
rect 673730 156272 673736 156324
rect 673788 156312 673794 156324
rect 675386 156312 675392 156324
rect 673788 156284 675392 156312
rect 673788 156272 673794 156284
rect 675386 156272 675392 156284
rect 675444 156272 675450 156324
rect 673454 155932 673460 155984
rect 673512 155972 673518 155984
rect 673914 155972 673920 155984
rect 673512 155944 673920 155972
rect 673512 155932 673518 155944
rect 673914 155932 673920 155944
rect 673972 155972 673978 155984
rect 675386 155972 675392 155984
rect 673972 155944 675392 155972
rect 673972 155932 673978 155944
rect 675386 155932 675392 155944
rect 675444 155932 675450 155984
rect 673546 152804 673552 152856
rect 673604 152844 673610 152856
rect 675386 152844 675392 152856
rect 673604 152816 675392 152844
rect 673604 152804 673610 152816
rect 675386 152804 675392 152816
rect 675444 152804 675450 152856
rect 673822 151716 673828 151768
rect 673880 151756 673886 151768
rect 675294 151756 675300 151768
rect 673880 151728 675300 151756
rect 673880 151716 673886 151728
rect 675294 151716 675300 151728
rect 675352 151716 675358 151768
rect 673730 144508 673736 144560
rect 673788 144548 673794 144560
rect 675386 144548 675392 144560
rect 673788 144520 675392 144548
rect 673788 144508 673794 144520
rect 675386 144508 675392 144520
rect 675444 144508 675450 144560
rect 42518 121456 42524 121508
rect 42576 121496 42582 121508
rect 44174 121496 44180 121508
rect 42576 121468 44180 121496
rect 42576 121456 42582 121468
rect 44174 121456 44180 121468
rect 44232 121456 44238 121508
rect 673822 111800 673828 111852
rect 673880 111840 673886 111852
rect 675386 111840 675392 111852
rect 673880 111812 675392 111840
rect 673880 111800 673886 111812
rect 675386 111800 675392 111812
rect 675444 111800 675450 111852
rect 673454 111528 673460 111580
rect 673512 111568 673518 111580
rect 673914 111568 673920 111580
rect 673512 111540 673920 111568
rect 673512 111528 673518 111540
rect 673914 111528 673920 111540
rect 673972 111568 673978 111580
rect 675386 111568 675392 111580
rect 673972 111540 675392 111568
rect 673972 111528 673978 111540
rect 675386 111528 675392 111540
rect 675444 111528 675450 111580
rect 673546 108400 673552 108452
rect 673604 108440 673610 108452
rect 675386 108440 675392 108452
rect 673604 108412 675392 108440
rect 673604 108400 673610 108412
rect 675386 108400 675392 108412
rect 675444 108400 675450 108452
rect 673638 107312 673644 107364
rect 673696 107352 673702 107364
rect 675294 107352 675300 107364
rect 673696 107324 675300 107352
rect 673696 107312 673702 107324
rect 675294 107312 675300 107324
rect 675352 107312 675358 107364
rect 42426 106020 42432 106072
rect 42484 106060 42490 106072
rect 44174 106060 44180 106072
rect 42484 106032 44180 106060
rect 42484 106020 42490 106032
rect 44174 106020 44180 106032
rect 44232 106020 44238 106072
rect 44818 46928 44824 46980
rect 44876 46928 44882 46980
rect 673638 46968 673644 46980
rect 200868 46940 297772 46968
rect 44836 46900 44864 46928
rect 200868 46912 200896 46940
rect 143534 46900 143540 46912
rect 44836 46872 143540 46900
rect 143534 46860 143540 46872
rect 143592 46860 143598 46912
rect 200850 46860 200856 46912
rect 200908 46860 200914 46912
rect 240888 46900 240916 46940
rect 297744 46912 297772 46940
rect 309428 46940 352604 46968
rect 309428 46912 309456 46940
rect 352576 46912 352604 46940
rect 364260 46940 407436 46968
rect 364260 46912 364288 46940
rect 407408 46912 407436 46940
rect 419092 46940 462176 46968
rect 419092 46912 419120 46940
rect 462148 46912 462176 46940
rect 473832 46940 517008 46968
rect 473832 46912 473860 46940
rect 516980 46912 517008 46940
rect 527468 46940 673644 46968
rect 527468 46912 527496 46940
rect 673638 46928 673644 46940
rect 673696 46928 673702 46980
rect 256234 46900 256240 46912
rect 240888 46872 256240 46900
rect 256234 46860 256240 46872
rect 256292 46860 256298 46912
rect 297726 46860 297732 46912
rect 297784 46860 297790 46912
rect 309410 46860 309416 46912
rect 309468 46860 309474 46912
rect 352558 46860 352564 46912
rect 352616 46860 352622 46912
rect 364242 46860 364248 46912
rect 364300 46860 364306 46912
rect 407390 46860 407396 46912
rect 407448 46860 407454 46912
rect 419074 46860 419080 46912
rect 419132 46860 419138 46912
rect 462130 46860 462136 46912
rect 462188 46860 462194 46912
rect 473814 46860 473820 46912
rect 473872 46860 473878 46912
rect 516962 46860 516968 46912
rect 517020 46860 517026 46912
rect 527450 46860 527456 46912
rect 527508 46860 527514 46912
rect 42242 45636 42248 45688
rect 42300 45676 42306 45688
rect 140958 45676 140964 45688
rect 42300 45648 140964 45676
rect 42300 45636 42306 45648
rect 140958 45636 140964 45648
rect 141016 45636 141022 45688
rect 42334 45568 42340 45620
rect 42392 45608 42398 45620
rect 143626 45608 143632 45620
rect 42392 45580 143632 45608
rect 42392 45568 42398 45580
rect 143626 45568 143632 45580
rect 143684 45568 143690 45620
rect 186682 45568 186688 45620
rect 186740 45608 186746 45620
rect 194686 45608 194692 45620
rect 186740 45580 194692 45608
rect 186740 45568 186746 45580
rect 194686 45568 194692 45580
rect 194744 45568 194750 45620
rect 523770 45568 523776 45620
rect 523828 45608 523834 45620
rect 673546 45608 673552 45620
rect 523828 45580 673552 45608
rect 523828 45568 523834 45580
rect 673546 45568 673552 45580
rect 673604 45568 673610 45620
rect 44910 45500 44916 45552
rect 44968 45540 44974 45552
rect 195974 45540 195980 45552
rect 44968 45512 195980 45540
rect 44968 45500 44974 45512
rect 195974 45500 195980 45512
rect 196032 45500 196038 45552
rect 518710 45500 518716 45552
rect 518768 45540 518774 45552
rect 673730 45540 673736 45552
rect 518768 45512 673736 45540
rect 518768 45500 518774 45512
rect 673730 45500 673736 45512
rect 673788 45500 673794 45552
rect 349982 44412 349988 44464
rect 350040 44452 350046 44464
rect 359366 44452 359372 44464
rect 350040 44424 359372 44452
rect 350040 44412 350046 44424
rect 359366 44412 359372 44424
rect 359424 44452 359430 44464
rect 414198 44452 414204 44464
rect 359424 44424 414204 44452
rect 359424 44412 359430 44424
rect 414198 44412 414204 44424
rect 414256 44412 414262 44464
rect 188522 44344 188528 44396
rect 188580 44384 188586 44396
rect 192846 44384 192852 44396
rect 188580 44356 192852 44384
rect 188580 44344 188586 44356
rect 192846 44344 192852 44356
rect 192904 44384 192910 44396
rect 297082 44384 297088 44396
rect 192904 44356 201540 44384
rect 192904 44344 192910 44356
rect 201512 44328 201540 44356
rect 284266 44356 297088 44384
rect 195974 44276 195980 44328
rect 196032 44316 196038 44328
rect 196032 44288 199792 44316
rect 196032 44276 196038 44288
rect 143626 44140 143632 44192
rect 143684 44180 143690 44192
rect 145098 44180 145104 44192
rect 143684 44152 145104 44180
rect 143684 44140 143690 44152
rect 145098 44140 145104 44152
rect 145156 44180 145162 44192
rect 195330 44180 195336 44192
rect 145156 44152 195336 44180
rect 145156 44140 145162 44152
rect 195330 44140 195336 44152
rect 195388 44180 195394 44192
rect 199654 44180 199660 44192
rect 195388 44152 199660 44180
rect 195388 44140 195394 44152
rect 199654 44140 199660 44152
rect 199712 44140 199718 44192
rect 199764 44180 199792 44288
rect 201494 44276 201500 44328
rect 201552 44316 201558 44328
rect 284266 44316 284294 44356
rect 297082 44344 297088 44356
rect 297140 44384 297146 44396
rect 299566 44384 299572 44396
rect 297140 44356 299572 44384
rect 297140 44344 297146 44356
rect 299566 44344 299572 44356
rect 299624 44384 299630 44396
rect 305730 44384 305736 44396
rect 299624 44356 305736 44384
rect 299624 44344 299630 44356
rect 305730 44344 305736 44356
rect 305788 44384 305794 44396
rect 305788 44356 322934 44384
rect 305788 44344 305794 44356
rect 201552 44288 284294 44316
rect 201552 44276 201558 44288
rect 295242 44276 295248 44328
rect 295300 44316 295306 44328
rect 303246 44316 303252 44328
rect 295300 44288 303252 44316
rect 295300 44276 295306 44288
rect 303246 44276 303252 44288
rect 303304 44276 303310 44328
rect 322906 44316 322934 44356
rect 468938 44344 468944 44396
rect 468996 44384 469002 44396
rect 523770 44384 523776 44396
rect 468996 44356 523776 44384
rect 468996 44344 469002 44356
rect 523770 44344 523776 44356
rect 523828 44344 523834 44396
rect 351914 44316 351920 44328
rect 303586 44288 303936 44316
rect 322906 44288 351920 44316
rect 199838 44208 199844 44260
rect 199896 44248 199902 44260
rect 303586 44248 303614 44288
rect 303908 44260 303936 44288
rect 351914 44276 351920 44288
rect 351972 44316 351978 44328
rect 354398 44316 354404 44328
rect 351972 44288 354404 44316
rect 351972 44276 351978 44288
rect 354398 44276 354404 44288
rect 354456 44316 354462 44328
rect 360562 44316 360568 44328
rect 354456 44288 360568 44316
rect 354456 44276 354462 44288
rect 360562 44276 360568 44288
rect 360620 44276 360626 44328
rect 363046 44316 363052 44328
rect 361546 44288 363052 44316
rect 199896 44220 303614 44248
rect 199896 44208 199902 44220
rect 303890 44208 303896 44260
rect 303948 44248 303954 44260
rect 308214 44248 308220 44260
rect 303948 44220 308220 44248
rect 303948 44208 303954 44220
rect 308214 44208 308220 44220
rect 308272 44248 308278 44260
rect 358722 44248 358728 44260
rect 308272 44220 358728 44248
rect 308272 44208 308278 44220
rect 358722 44208 358728 44220
rect 358780 44248 358786 44260
rect 361546 44248 361574 44288
rect 363046 44276 363052 44288
rect 363104 44316 363110 44328
rect 413554 44316 413560 44328
rect 363104 44288 413560 44316
rect 363104 44276 363110 44288
rect 413554 44276 413560 44288
rect 413612 44316 413618 44328
rect 417878 44316 417884 44328
rect 413612 44288 417884 44316
rect 413612 44276 413618 44288
rect 417878 44276 417884 44288
rect 417936 44316 417942 44328
rect 468294 44316 468300 44328
rect 417936 44288 468300 44316
rect 417936 44276 417942 44288
rect 468294 44276 468300 44288
rect 468352 44316 468358 44328
rect 472618 44316 472624 44328
rect 468352 44288 472624 44316
rect 468352 44276 468358 44288
rect 472618 44276 472624 44288
rect 472676 44316 472682 44328
rect 472676 44288 523172 44316
rect 472676 44276 472682 44288
rect 406746 44248 406752 44260
rect 358780 44220 361574 44248
rect 380866 44220 406752 44248
rect 358780 44208 358786 44220
rect 304534 44180 304540 44192
rect 199764 44152 304540 44180
rect 304534 44140 304540 44152
rect 304592 44180 304598 44192
rect 349982 44180 349988 44192
rect 304592 44152 349988 44180
rect 304592 44140 304598 44152
rect 349982 44140 349988 44152
rect 350040 44140 350046 44192
rect 350074 44140 350080 44192
rect 350132 44180 350138 44192
rect 358078 44180 358084 44192
rect 350132 44152 358084 44180
rect 350132 44140 350138 44152
rect 358078 44140 358084 44152
rect 358136 44140 358142 44192
rect 360562 44140 360568 44192
rect 360620 44180 360626 44192
rect 380866 44180 380894 44220
rect 406746 44208 406752 44220
rect 406804 44248 406810 44260
rect 461486 44248 461492 44260
rect 406804 44220 461492 44248
rect 406804 44208 406810 44220
rect 461486 44208 461492 44220
rect 461544 44248 461550 44260
rect 516318 44248 516324 44260
rect 461544 44220 516324 44248
rect 461544 44208 461550 44220
rect 516318 44208 516324 44220
rect 516376 44248 516382 44260
rect 518710 44248 518716 44260
rect 516376 44220 518716 44248
rect 516376 44208 516382 44220
rect 518710 44208 518716 44220
rect 518768 44208 518774 44260
rect 523144 44192 523172 44288
rect 360620 44152 380894 44180
rect 360620 44140 360626 44152
rect 414198 44140 414204 44192
rect 414256 44180 414262 44192
rect 468938 44180 468944 44192
rect 414256 44152 468944 44180
rect 414256 44140 414262 44152
rect 468938 44140 468944 44152
rect 468996 44140 469002 44192
rect 523126 44140 523132 44192
rect 523184 44180 523190 44192
rect 527450 44180 527456 44192
rect 523184 44152 527456 44180
rect 523184 44140 523190 44152
rect 527450 44140 527456 44152
rect 527508 44140 527514 44192
rect 579890 42712 579896 42764
rect 579948 42752 579954 42764
rect 673454 42752 673460 42764
rect 579948 42724 673460 42752
rect 579948 42712 579954 42724
rect 673454 42712 673460 42724
rect 673512 42712 673518 42764
rect 189258 41896 189264 41948
rect 189316 41936 189322 41948
rect 191098 41936 191104 41948
rect 189316 41908 191104 41936
rect 189316 41896 189322 41908
rect 191098 41896 191104 41908
rect 191156 41936 191162 41948
rect 192294 41936 192300 41948
rect 191156 41908 192300 41936
rect 191156 41896 191162 41908
rect 192294 41896 192300 41908
rect 192352 41936 192358 41948
rect 193582 41936 193588 41948
rect 192352 41908 193588 41936
rect 192352 41896 192358 41908
rect 193582 41896 193588 41908
rect 193640 41936 193646 41948
rect 196434 41936 196440 41948
rect 193640 41908 196440 41936
rect 193640 41896 193646 41908
rect 196434 41896 196440 41908
rect 196492 41896 196498 41948
rect 198458 41896 198464 41948
rect 198516 41936 198522 41948
rect 200114 41936 200120 41948
rect 198516 41908 200120 41936
rect 198516 41896 198522 41908
rect 200114 41896 200120 41908
rect 200172 41896 200178 41948
rect 297910 41896 297916 41948
rect 297968 41936 297974 41948
rect 300670 41936 300676 41948
rect 297968 41908 300676 41936
rect 297968 41896 297974 41908
rect 300670 41896 300676 41908
rect 300728 41896 300734 41948
rect 302234 41896 302240 41948
rect 302292 41936 302298 41948
rect 305270 41936 305276 41948
rect 302292 41908 305276 41936
rect 302292 41896 302298 41908
rect 305270 41896 305276 41908
rect 305328 41936 305334 41948
rect 306558 41936 306564 41948
rect 305328 41908 306564 41936
rect 305328 41896 305334 41908
rect 306558 41896 306564 41908
rect 306616 41936 306622 41948
rect 308674 41936 308680 41948
rect 306616 41908 308680 41936
rect 306616 41896 306622 41908
rect 308674 41896 308680 41908
rect 308732 41896 308738 41948
rect 352650 41896 352656 41948
rect 352708 41936 352714 41948
rect 355502 41936 355508 41948
rect 352708 41908 355508 41936
rect 352708 41896 352714 41908
rect 355502 41896 355508 41908
rect 355560 41896 355566 41948
rect 356974 41896 356980 41948
rect 357032 41936 357038 41948
rect 359826 41936 359832 41948
rect 357032 41908 359832 41936
rect 357032 41896 357038 41908
rect 359826 41896 359832 41908
rect 359884 41936 359890 41948
rect 361114 41936 361120 41948
rect 359884 41908 361120 41936
rect 359884 41896 359890 41908
rect 361114 41896 361120 41908
rect 361172 41936 361178 41948
rect 363506 41936 363512 41948
rect 361172 41908 363512 41936
rect 361172 41896 361178 41908
rect 363506 41896 363512 41908
rect 363564 41896 363570 41948
rect 407482 41896 407488 41948
rect 407540 41936 407546 41948
rect 410242 41936 410248 41948
rect 407540 41908 410248 41936
rect 407540 41896 407546 41908
rect 410242 41896 410248 41908
rect 410300 41936 410306 41948
rect 411530 41936 411536 41948
rect 410300 41908 411536 41936
rect 410300 41896 410306 41908
rect 411530 41896 411536 41908
rect 411588 41936 411594 41948
rect 414566 41936 414572 41948
rect 411588 41908 414572 41936
rect 411588 41896 411594 41908
rect 414566 41896 414572 41908
rect 414624 41936 414630 41948
rect 415854 41936 415860 41948
rect 414624 41908 415860 41936
rect 414624 41896 414630 41908
rect 415854 41896 415860 41908
rect 415912 41936 415918 41948
rect 418246 41936 418252 41948
rect 415912 41908 418252 41936
rect 415912 41896 415918 41908
rect 418246 41896 418252 41908
rect 418304 41896 418310 41948
rect 462314 41896 462320 41948
rect 462372 41936 462378 41948
rect 465074 41936 465080 41948
rect 462372 41908 465080 41936
rect 462372 41896 462378 41908
rect 465074 41896 465080 41908
rect 465132 41936 465138 41948
rect 466362 41936 466368 41948
rect 465132 41908 466368 41936
rect 465132 41896 465138 41908
rect 466362 41896 466368 41908
rect 466420 41936 466426 41948
rect 469398 41936 469404 41948
rect 466420 41908 469404 41936
rect 466420 41896 466426 41908
rect 469398 41896 469404 41908
rect 469456 41936 469462 41948
rect 470686 41936 470692 41948
rect 469456 41908 470692 41936
rect 469456 41896 469462 41908
rect 470686 41896 470692 41908
rect 470744 41936 470750 41948
rect 473078 41936 473084 41948
rect 470744 41908 473084 41936
rect 470744 41896 470750 41908
rect 473078 41896 473084 41908
rect 473136 41896 473142 41948
rect 517054 41896 517060 41948
rect 517112 41936 517118 41948
rect 519906 41936 519912 41948
rect 517112 41908 519912 41936
rect 517112 41896 517118 41908
rect 519906 41896 519912 41908
rect 519964 41936 519970 41948
rect 521194 41936 521200 41948
rect 519964 41908 521200 41936
rect 519964 41896 519970 41908
rect 521194 41896 521200 41908
rect 521252 41936 521258 41948
rect 524230 41936 524236 41948
rect 521252 41908 524236 41936
rect 521252 41896 521258 41908
rect 524230 41896 524236 41908
rect 524288 41936 524294 41948
rect 525518 41936 525524 41948
rect 524288 41908 525524 41936
rect 524288 41896 524294 41908
rect 525518 41896 525524 41908
rect 525576 41936 525582 41948
rect 527910 41936 527916 41948
rect 525576 41908 527916 41936
rect 525576 41896 525582 41908
rect 527910 41896 527916 41908
rect 527968 41896 527974 41948
rect 146294 41828 146300 41880
rect 146352 41868 146358 41880
rect 568850 41868 568856 41880
rect 146352 41840 568856 41868
rect 146352 41828 146358 41840
rect 568850 41828 568856 41840
rect 568908 41868 568914 41880
rect 579890 41868 579896 41880
rect 568908 41840 579896 41868
rect 568908 41828 568914 41840
rect 579890 41828 579896 41840
rect 579948 41828 579954 41880
rect 198918 41800 198924 41812
rect 168346 41772 198924 41800
rect 93762 41488 93768 41540
rect 93820 41528 93826 41540
rect 168346 41528 168374 41772
rect 198918 41760 198924 41772
rect 198976 41800 198982 41812
rect 307754 41800 307760 41812
rect 198976 41772 307760 41800
rect 198976 41760 198982 41772
rect 307754 41760 307760 41772
rect 307812 41800 307818 41812
rect 362494 41800 362500 41812
rect 307812 41772 362500 41800
rect 307812 41760 307818 41772
rect 362494 41760 362500 41772
rect 362552 41800 362558 41812
rect 362552 41772 380894 41800
rect 362552 41760 362558 41772
rect 93820 41500 168374 41528
rect 380866 41528 380894 41772
rect 409322 41760 409328 41812
rect 409380 41800 409386 41812
rect 412358 41800 412364 41812
rect 409380 41772 412364 41800
rect 409380 41760 409386 41772
rect 412358 41760 412364 41772
rect 412416 41800 412422 41812
rect 415210 41800 415216 41812
rect 412416 41772 415216 41800
rect 412416 41760 412422 41772
rect 415210 41760 415216 41772
rect 415268 41760 415274 41812
rect 417326 41800 417332 41812
rect 417252 41772 417332 41800
rect 417252 41528 417280 41772
rect 417326 41760 417332 41772
rect 417384 41760 417390 41812
rect 464154 41760 464160 41812
rect 464212 41800 464218 41812
rect 467190 41800 467196 41812
rect 464212 41772 467196 41800
rect 464212 41760 464218 41772
rect 467190 41760 467196 41772
rect 467248 41800 467254 41812
rect 470042 41800 470048 41812
rect 467248 41772 470048 41800
rect 467248 41760 467254 41772
rect 470042 41760 470048 41772
rect 470100 41760 470106 41812
rect 472158 41800 472164 41812
rect 472084 41772 472164 41800
rect 472084 41528 472112 41772
rect 472158 41760 472164 41772
rect 472216 41760 472222 41812
rect 526714 41800 526720 41812
rect 516106 41772 526720 41800
rect 516106 41528 516134 41772
rect 526714 41760 526720 41772
rect 526772 41760 526778 41812
rect 380866 41500 516134 41528
rect 93820 41488 93826 41500
rect 135162 40196 135168 40248
rect 135220 40236 135226 40248
rect 143534 40236 143540 40248
rect 135220 40208 143540 40236
rect 135220 40196 135226 40208
rect 143534 40196 143540 40208
rect 143592 40196 143598 40248
rect 140990 40060 140996 40112
rect 141048 40100 141054 40112
rect 143066 40100 143072 40112
rect 141048 40072 143072 40100
rect 141048 40060 141054 40072
rect 142586 39950 142614 40072
rect 143066 40060 143072 40072
rect 143124 40100 143130 40112
rect 144546 40100 144552 40112
rect 143124 40072 144552 40100
rect 143124 40060 143130 40072
rect 144546 40060 144552 40072
rect 144604 40100 144610 40112
rect 146294 40100 146300 40112
rect 144604 40072 146300 40100
rect 144604 40060 144610 40072
rect 146294 40060 146300 40072
rect 146352 40060 146358 40112
<< via1 >>
rect 585784 996412 585836 996464
rect 674748 996412 674800 996464
rect 42248 996344 42300 996396
rect 339500 996344 339552 996396
rect 673552 996344 673604 996396
rect 44916 990088 44968 990140
rect 673644 990088 673696 990140
rect 42340 990020 42392 990072
rect 673460 990020 673512 990072
rect 42432 861160 42484 861212
rect 44180 861160 44232 861212
rect 673552 859120 673604 859172
rect 675392 859120 675444 859172
rect 673644 856060 673696 856112
rect 675392 856060 675444 856112
rect 673736 855380 673788 855432
rect 675392 855380 675444 855432
rect 673460 849668 673512 849720
rect 675392 849668 675444 849720
rect 675300 803768 675352 803820
rect 677600 803768 677652 803820
rect 42248 800980 42300 801032
rect 42616 800980 42668 801032
rect 41788 798532 41840 798584
rect 42340 798532 42392 798584
rect 41788 792072 41840 792124
rect 42432 792072 42484 792124
rect 41788 789080 41840 789132
rect 42616 789080 42668 789132
rect 42248 787992 42300 788044
rect 42432 787992 42484 788044
rect 673736 773304 673788 773356
rect 675208 773304 675260 773356
rect 675392 773304 675444 773356
rect 673552 772760 673604 772812
rect 675392 772760 675444 772812
rect 673644 769632 673696 769684
rect 673920 769632 673972 769684
rect 675392 769632 675444 769684
rect 673736 769088 673788 769140
rect 675208 769088 675260 769140
rect 675392 769088 675444 769140
rect 675208 767592 675260 767644
rect 675392 767592 675444 767644
rect 673460 761268 673512 761320
rect 674012 761268 674064 761320
rect 675392 761268 675444 761320
rect 675208 760180 675260 760232
rect 675392 760180 675444 760232
rect 41788 756236 41840 756288
rect 42340 756236 42392 756288
rect 42616 756236 42668 756288
rect 41788 748280 41840 748332
rect 42524 748280 42576 748332
rect 41788 744812 41840 744864
rect 42432 744812 42484 744864
rect 42708 744812 42760 744864
rect 673736 728560 673788 728612
rect 675392 728560 675444 728612
rect 673552 728356 673604 728408
rect 675392 728356 675444 728408
rect 673920 725228 673972 725280
rect 675392 725228 675444 725280
rect 673460 724004 673512 724056
rect 675392 724004 675444 724056
rect 673644 717816 673696 717868
rect 674012 717816 674064 717868
rect 675392 717816 675444 717868
rect 41788 713056 41840 713108
rect 42616 713056 42668 713108
rect 41788 704760 41840 704812
rect 42524 704760 42576 704812
rect 41788 701632 41840 701684
rect 42432 701632 42484 701684
rect 673460 684292 673512 684344
rect 675300 684292 675352 684344
rect 673552 683068 673604 683120
rect 673736 683068 673788 683120
rect 675392 683068 675444 683120
rect 673552 680416 673604 680468
rect 673920 680416 673972 680468
rect 675392 680416 675444 680468
rect 673828 680076 673880 680128
rect 675392 680076 675444 680128
rect 675208 678784 675260 678836
rect 675392 678784 675444 678836
rect 673644 673616 673696 673668
rect 674012 673616 674064 673668
rect 675392 673616 675444 673668
rect 41788 668720 41840 668772
rect 42616 668720 42668 668772
rect 41788 661308 41840 661360
rect 42524 661308 42576 661360
rect 41788 659268 41840 659320
rect 42432 659268 42484 659320
rect 42708 659268 42760 659320
rect 673828 640092 673880 640144
rect 675300 640092 675352 640144
rect 673644 638868 673696 638920
rect 675392 638868 675444 638920
rect 673552 636284 673604 636336
rect 675392 636284 675444 636336
rect 673736 635740 673788 635792
rect 675300 635740 675352 635792
rect 675208 634584 675260 634636
rect 675392 634584 675444 634636
rect 673460 629416 673512 629468
rect 674012 629416 674064 629468
rect 675392 629416 675444 629468
rect 41788 625472 41840 625524
rect 42616 625472 42668 625524
rect 41788 618128 41840 618180
rect 42524 618128 42576 618180
rect 41788 615000 41840 615052
rect 42708 615000 42760 615052
rect 42248 614660 42300 614712
rect 673736 596096 673788 596148
rect 675208 596096 675260 596148
rect 675392 596096 675444 596148
rect 673644 595144 673696 595196
rect 675392 595144 675444 595196
rect 673552 591880 673604 591932
rect 675392 591880 675444 591932
rect 673736 590792 673788 590844
rect 675208 590792 675260 590844
rect 675392 590792 675444 590844
rect 673460 584128 673512 584180
rect 673920 584128 673972 584180
rect 675392 584128 675444 584180
rect 41788 583244 41840 583296
rect 42616 583244 42668 583296
rect 41788 576512 41840 576564
rect 42248 576512 42300 576564
rect 42432 576512 42484 576564
rect 41788 575900 41840 575952
rect 42524 575900 42576 575952
rect 41788 571820 41840 571872
rect 42432 571820 42484 571872
rect 673736 551488 673788 551540
rect 675208 551488 675260 551540
rect 673644 551352 673696 551404
rect 675392 551352 675444 551404
rect 673552 548224 673604 548276
rect 675392 548224 675444 548276
rect 673460 547000 673512 547052
rect 675208 547000 675260 547052
rect 675392 547000 675444 547052
rect 673920 540880 673972 540932
rect 675392 540880 675444 540932
rect 41788 540064 41840 540116
rect 42616 540064 42668 540116
rect 41788 531768 41840 531820
rect 42524 531768 42576 531820
rect 42708 531768 42760 531820
rect 41788 528640 41840 528692
rect 42432 528640 42484 528692
rect 675300 499468 675352 499520
rect 676128 499468 676180 499520
rect 676128 494844 676180 494896
rect 677968 494844 678020 494896
rect 674012 422220 674064 422272
rect 674748 422220 674800 422272
rect 674012 419160 674064 419212
rect 677508 419160 677560 419212
rect 41788 411272 41840 411324
rect 42524 411272 42576 411324
rect 41788 404880 41840 404932
rect 42708 404880 42760 404932
rect 41788 401888 41840 401940
rect 42432 401888 42484 401940
rect 673920 376116 673972 376168
rect 675392 376116 675444 376168
rect 673736 373056 673788 373108
rect 675392 373056 675444 373108
rect 673552 372784 673604 372836
rect 675392 372784 675444 372836
rect 41788 369044 41840 369096
rect 42524 369044 42576 369096
rect 674012 365712 674064 365764
rect 675392 365712 675444 365764
rect 41788 361292 41840 361344
rect 42616 361292 42668 361344
rect 41788 357620 41840 357672
rect 42432 357620 42484 357672
rect 42708 357620 42760 357672
rect 673736 333956 673788 334008
rect 675208 333956 675260 334008
rect 673552 333072 673604 333124
rect 675300 333072 675352 333124
rect 673460 331916 673512 331968
rect 673920 331916 673972 331968
rect 675392 331916 675444 331968
rect 673552 328856 673604 328908
rect 675208 328856 675260 328908
rect 675392 328856 675444 328908
rect 673736 328244 673788 328296
rect 675392 328244 675444 328296
rect 41788 325660 41840 325712
rect 42524 325660 42576 325712
rect 673644 322464 673696 322516
rect 674012 322464 674064 322516
rect 675392 322464 675444 322516
rect 41788 317364 41840 317416
rect 42616 317364 42668 317416
rect 41788 314236 41840 314288
rect 42524 314236 42576 314288
rect 42708 314236 42760 314288
rect 42248 313080 42300 313132
rect 42340 312876 42392 312928
rect 673736 289280 673788 289332
rect 675392 289280 675444 289332
rect 673460 288736 673512 288788
rect 675392 288736 675444 288788
rect 673552 285268 673604 285320
rect 675392 285268 675444 285320
rect 42340 284112 42392 284164
rect 673736 284044 673788 284096
rect 675392 284044 675444 284096
rect 42340 283908 42392 283960
rect 41788 281528 41840 281580
rect 42432 281528 42484 281580
rect 42708 281528 42760 281580
rect 673644 277312 673696 277364
rect 675392 277312 675444 277364
rect 41788 274660 41840 274712
rect 42616 274660 42668 274712
rect 41788 272076 41840 272128
rect 42524 272076 42576 272128
rect 673736 244604 673788 244656
rect 675392 244604 675444 244656
rect 673460 243720 673512 243772
rect 675392 243720 675444 243772
rect 673552 240252 673604 240304
rect 675392 240252 675444 240304
rect 673736 239640 673788 239692
rect 675392 239640 675444 239692
rect 41788 238280 41840 238332
rect 42432 238280 42484 238332
rect 42708 238280 42760 238332
rect 673644 233860 673696 233912
rect 675392 233860 675444 233912
rect 41788 231888 41840 231940
rect 42616 231888 42668 231940
rect 41788 228828 41840 228880
rect 42524 228828 42576 228880
rect 673736 200404 673788 200456
rect 675392 200404 675444 200456
rect 673460 199112 673512 199164
rect 675392 199112 675444 199164
rect 673552 197004 673604 197056
rect 675392 197004 675444 197056
rect 673736 195780 673788 195832
rect 675392 195780 675444 195832
rect 41788 195100 41840 195152
rect 42432 195100 42484 195152
rect 673644 189252 673696 189304
rect 675392 189252 675444 189304
rect 41788 188708 41840 188760
rect 42524 188708 42576 188760
rect 42800 188708 42852 188760
rect 41788 185648 41840 185700
rect 42708 185648 42760 185700
rect 42248 184356 42300 184408
rect 42708 184356 42760 184408
rect 673736 156272 673788 156324
rect 675392 156272 675444 156324
rect 673460 155932 673512 155984
rect 673920 155932 673972 155984
rect 675392 155932 675444 155984
rect 673552 152804 673604 152856
rect 675392 152804 675444 152856
rect 673828 151716 673880 151768
rect 675300 151716 675352 151768
rect 673736 144508 673788 144560
rect 675392 144508 675444 144560
rect 42524 121456 42576 121508
rect 44180 121456 44232 121508
rect 673828 111800 673880 111852
rect 675392 111800 675444 111852
rect 673460 111528 673512 111580
rect 673920 111528 673972 111580
rect 675392 111528 675444 111580
rect 673552 108400 673604 108452
rect 675392 108400 675444 108452
rect 673644 107312 673696 107364
rect 675300 107312 675352 107364
rect 42432 106020 42484 106072
rect 44180 106020 44232 106072
rect 44824 46928 44876 46980
rect 143540 46860 143592 46912
rect 200856 46860 200908 46912
rect 673644 46928 673696 46980
rect 256240 46860 256292 46912
rect 297732 46860 297784 46912
rect 309416 46860 309468 46912
rect 352564 46860 352616 46912
rect 364248 46860 364300 46912
rect 407396 46860 407448 46912
rect 419080 46860 419132 46912
rect 462136 46860 462188 46912
rect 473820 46860 473872 46912
rect 516968 46860 517020 46912
rect 527456 46860 527508 46912
rect 42248 45636 42300 45688
rect 140964 45636 141016 45688
rect 42340 45568 42392 45620
rect 143632 45568 143684 45620
rect 186688 45568 186740 45620
rect 194692 45568 194744 45620
rect 523776 45568 523828 45620
rect 673552 45568 673604 45620
rect 44916 45500 44968 45552
rect 195980 45500 196032 45552
rect 518716 45500 518768 45552
rect 673736 45500 673788 45552
rect 349988 44412 350040 44464
rect 359372 44412 359424 44464
rect 414204 44412 414256 44464
rect 188528 44344 188580 44396
rect 192852 44344 192904 44396
rect 195980 44276 196032 44328
rect 143632 44140 143684 44192
rect 145104 44140 145156 44192
rect 195336 44140 195388 44192
rect 199660 44140 199712 44192
rect 201500 44276 201552 44328
rect 297088 44344 297140 44396
rect 299572 44344 299624 44396
rect 305736 44344 305788 44396
rect 295248 44276 295300 44328
rect 303252 44276 303304 44328
rect 468944 44344 468996 44396
rect 523776 44344 523828 44396
rect 199844 44208 199896 44260
rect 351920 44276 351972 44328
rect 354404 44276 354456 44328
rect 360568 44276 360620 44328
rect 303896 44208 303948 44260
rect 308220 44208 308272 44260
rect 358728 44208 358780 44260
rect 363052 44276 363104 44328
rect 413560 44276 413612 44328
rect 417884 44276 417936 44328
rect 468300 44276 468352 44328
rect 472624 44276 472676 44328
rect 304540 44140 304592 44192
rect 349988 44140 350040 44192
rect 350080 44140 350132 44192
rect 358084 44140 358136 44192
rect 360568 44140 360620 44192
rect 406752 44208 406804 44260
rect 461492 44208 461544 44260
rect 516324 44208 516376 44260
rect 518716 44208 518768 44260
rect 414204 44140 414256 44192
rect 468944 44140 468996 44192
rect 523132 44140 523184 44192
rect 527456 44140 527508 44192
rect 579896 42712 579948 42764
rect 673460 42712 673512 42764
rect 189264 41896 189316 41948
rect 191104 41896 191156 41948
rect 192300 41896 192352 41948
rect 193588 41896 193640 41948
rect 196440 41896 196492 41948
rect 198464 41896 198516 41948
rect 200120 41896 200172 41948
rect 297916 41896 297968 41948
rect 300676 41896 300728 41948
rect 302240 41896 302292 41948
rect 305276 41896 305328 41948
rect 306564 41896 306616 41948
rect 308680 41896 308732 41948
rect 352656 41896 352708 41948
rect 355508 41896 355560 41948
rect 356980 41896 357032 41948
rect 359832 41896 359884 41948
rect 361120 41896 361172 41948
rect 363512 41896 363564 41948
rect 407488 41896 407540 41948
rect 410248 41896 410300 41948
rect 411536 41896 411588 41948
rect 414572 41896 414624 41948
rect 415860 41896 415912 41948
rect 418252 41896 418304 41948
rect 462320 41896 462372 41948
rect 465080 41896 465132 41948
rect 466368 41896 466420 41948
rect 469404 41896 469456 41948
rect 470692 41896 470744 41948
rect 473084 41896 473136 41948
rect 517060 41896 517112 41948
rect 519912 41896 519964 41948
rect 521200 41896 521252 41948
rect 524236 41896 524288 41948
rect 525524 41896 525576 41948
rect 527916 41896 527968 41948
rect 146300 41828 146352 41880
rect 568856 41828 568908 41880
rect 579896 41828 579948 41880
rect 93768 41488 93820 41540
rect 198924 41760 198976 41812
rect 307760 41760 307812 41812
rect 362500 41760 362552 41812
rect 409328 41760 409380 41812
rect 412364 41760 412416 41812
rect 415216 41760 415268 41812
rect 417332 41760 417384 41812
rect 464160 41760 464212 41812
rect 467196 41760 467248 41812
rect 470048 41760 470100 41812
rect 472164 41760 472216 41812
rect 526720 41760 526772 41812
rect 135168 40196 135220 40248
rect 143540 40196 143592 40248
rect 140996 40060 141048 40112
rect 143072 40060 143124 40112
rect 144552 40060 144604 40112
rect 146300 40060 146352 40112
<< metal2 >>
rect 229499 997600 234279 998010
rect 239478 997600 244258 1002732
rect 280899 997600 285679 998010
rect 290878 997600 295658 1002732
rect 585782 997520 585838 997529
rect 585782 997455 585838 997464
rect 339498 997112 339554 997121
rect 339498 997047 339554 997056
rect 339512 996402 339540 997047
rect 585796 996470 585824 997455
rect 585784 996464 585836 996470
rect 585784 996406 585836 996412
rect 674748 996464 674800 996470
rect 674748 996406 674800 996412
rect 42248 996396 42300 996402
rect 42248 996338 42300 996344
rect 339500 996396 339552 996402
rect 339500 996338 339552 996344
rect 673552 996396 673604 996402
rect 673552 996338 673604 996344
rect 42260 801038 42288 996338
rect 44916 990140 44968 990146
rect 44916 990082 44968 990088
rect 42340 990072 42392 990078
rect 42340 990014 42392 990020
rect 42248 801032 42300 801038
rect 42248 800974 42300 800980
rect 41722 800875 42288 800903
rect 41713 800217 42193 800273
rect 41722 799054 41828 799082
rect 41800 798590 41828 799054
rect 41788 798584 41840 798590
rect 41788 798526 41840 798532
rect 41713 798377 42193 798433
rect 41713 797733 42193 797789
rect 41713 796537 42193 796593
rect 41713 795893 42193 795949
rect 41713 795341 42193 795397
rect 41713 794697 42193 794753
rect 41713 794053 42193 794109
rect 41713 793501 42193 793557
rect 42260 793098 42288 800875
rect 42352 798590 42380 990014
rect 44928 902534 44956 990082
rect 673460 990072 673512 990078
rect 673460 990014 673512 990020
rect 44836 902506 44956 902534
rect 44836 885873 44864 902506
rect 44178 885864 44234 885873
rect 44178 885799 44234 885808
rect 44822 885864 44878 885873
rect 44822 885799 44878 885808
rect 44192 871049 44220 885799
rect 44178 871040 44234 871049
rect 44178 870975 44234 870984
rect 44192 861218 44220 870975
rect 42432 861212 42484 861218
rect 42432 861154 42484 861160
rect 44180 861212 44232 861218
rect 44180 861154 44232 861160
rect 42340 798584 42392 798590
rect 42340 798526 42392 798532
rect 41800 793070 42288 793098
rect 41800 792899 41828 793070
rect 41722 792871 41828 792899
rect 41722 792254 42288 792282
rect 41788 792124 41840 792130
rect 41788 792066 41840 792072
rect 41800 791602 41828 792066
rect 41722 791574 41828 791602
rect 41713 791017 42193 791073
rect 41713 790373 42193 790429
rect 41713 789729 42193 789785
rect 41713 789177 42193 789233
rect 41788 789132 41840 789138
rect 41788 789074 41840 789080
rect 41800 788575 41828 789074
rect 41722 788547 41828 788575
rect 42260 788066 42288 792254
rect 41892 788050 42288 788066
rect 41892 788044 42300 788050
rect 41892 788038 42248 788044
rect 41892 787930 41920 788038
rect 42248 787986 42300 787992
rect 42260 787955 42288 787986
rect 41722 787902 41920 787930
rect 41713 787337 42193 787393
rect 41713 786693 42193 786749
rect 41713 786049 42193 786105
rect 41713 785497 42193 785553
rect 41722 757675 42288 757703
rect 41713 757017 42193 757073
rect 41788 756288 41840 756294
rect 41788 756230 41840 756236
rect 41800 755863 41828 756230
rect 41722 755835 41828 755863
rect 41713 755177 42193 755233
rect 41713 754533 42193 754589
rect 41713 753337 42193 753393
rect 41713 752693 42193 752749
rect 41713 752141 42193 752197
rect 41713 751497 42193 751553
rect 41713 750853 42193 750909
rect 41713 750301 42193 750357
rect 42260 749850 42288 757675
rect 42352 756294 42380 798526
rect 42444 792130 42472 861154
rect 673472 849726 673500 990014
rect 673564 859178 673592 996338
rect 673644 990140 673696 990146
rect 673644 990082 673696 990088
rect 673552 859172 673604 859178
rect 673552 859114 673604 859120
rect 673460 849720 673512 849726
rect 673460 849662 673512 849668
rect 42616 801032 42668 801038
rect 42616 800974 42668 800980
rect 42432 792124 42484 792130
rect 42432 792066 42484 792072
rect 42444 792010 42472 792066
rect 42444 791982 42564 792010
rect 42432 788044 42484 788050
rect 42432 787986 42484 787992
rect 42340 756288 42392 756294
rect 42340 756230 42392 756236
rect 41800 749822 42288 749850
rect 41800 749714 41828 749822
rect 41722 749686 41828 749714
rect 42444 749578 42472 787986
rect 41800 749550 42472 749578
rect 41800 749034 41828 749550
rect 41722 749006 41828 749034
rect 41722 748383 41828 748411
rect 41800 748338 41828 748383
rect 41788 748332 41840 748338
rect 41788 748274 41840 748280
rect 41713 747817 42193 747873
rect 41713 747173 42193 747229
rect 41713 746529 42193 746585
rect 41713 745977 42193 746033
rect 41722 745334 41828 745362
rect 41800 744870 41828 745334
rect 41788 744864 41840 744870
rect 41788 744806 41840 744812
rect 42260 744731 42288 749550
rect 42536 748338 42564 791982
rect 42628 789138 42656 800974
rect 42616 789132 42668 789138
rect 42616 789074 42668 789080
rect 42628 786614 42656 789074
rect 42628 786586 42748 786614
rect 42616 756288 42668 756294
rect 42616 756230 42668 756236
rect 42524 748332 42576 748338
rect 42524 748274 42576 748280
rect 42432 744864 42484 744870
rect 42432 744806 42484 744812
rect 41722 744703 42288 744731
rect 41713 744137 42193 744193
rect 41713 743493 42193 743549
rect 41713 742849 42193 742905
rect 41713 742297 42193 742353
rect 42260 728654 42288 744703
rect 42260 728626 42380 728654
rect 41722 714462 41920 714490
rect 41892 714218 41920 714462
rect 41892 714190 42288 714218
rect 41713 713817 42193 713873
rect 41788 713108 41840 713114
rect 41788 713050 41840 713056
rect 41800 712663 41828 713050
rect 41722 712635 41828 712663
rect 41713 711977 42193 712033
rect 41713 711333 42193 711389
rect 41713 710137 42193 710193
rect 41713 709493 42193 709549
rect 41713 708941 42193 708997
rect 41713 708297 42193 708353
rect 41713 707653 42193 707709
rect 41713 707101 42193 707157
rect 42260 706499 42288 714190
rect 41722 706471 42288 706499
rect 42352 705855 42380 728626
rect 41722 705827 42380 705855
rect 41722 705183 41828 705211
rect 41800 704818 41828 705183
rect 41788 704812 41840 704818
rect 41788 704754 41840 704760
rect 41713 704617 42193 704673
rect 41713 703973 42193 704029
rect 41713 703329 42193 703385
rect 41713 702777 42193 702833
rect 41722 702147 41828 702175
rect 41800 701690 41828 702147
rect 41788 701684 41840 701690
rect 41788 701626 41840 701632
rect 41722 701503 41920 701531
rect 41892 701434 41920 701503
rect 42260 701434 42288 705827
rect 42444 701690 42472 744806
rect 42536 704818 42564 748274
rect 42628 713114 42656 756230
rect 42720 744870 42748 786586
rect 673472 761326 673500 849662
rect 673564 772818 673592 859114
rect 673656 856118 673684 990082
rect 673644 856112 673696 856118
rect 673644 856054 673696 856060
rect 673552 772812 673604 772818
rect 673552 772754 673604 772760
rect 673460 761320 673512 761326
rect 673460 761262 673512 761268
rect 42708 744864 42760 744870
rect 42708 744806 42760 744812
rect 673564 728414 673592 772754
rect 673656 769690 673684 856054
rect 673736 855432 673788 855438
rect 673736 855374 673788 855380
rect 673748 773362 673776 855374
rect 673736 773356 673788 773362
rect 673736 773298 673788 773304
rect 673644 769684 673696 769690
rect 673644 769626 673696 769632
rect 673920 769684 673972 769690
rect 673920 769626 673972 769632
rect 673736 769140 673788 769146
rect 673736 769082 673788 769088
rect 673748 728618 673776 769082
rect 673736 728612 673788 728618
rect 673736 728554 673788 728560
rect 673552 728408 673604 728414
rect 673552 728350 673604 728356
rect 673460 724056 673512 724062
rect 673460 723998 673512 724004
rect 42616 713108 42668 713114
rect 42616 713050 42668 713056
rect 42524 704812 42576 704818
rect 42524 704754 42576 704760
rect 42432 701684 42484 701690
rect 42432 701626 42484 701632
rect 41892 701406 42288 701434
rect 41713 700937 42193 700993
rect 41713 700293 42193 700349
rect 41713 699649 42193 699705
rect 41713 699097 42193 699153
rect 42260 690014 42288 701406
rect 42260 689986 42380 690014
rect 41722 671078 41828 671106
rect 41800 670694 41828 671078
rect 41800 670666 42288 670694
rect 41713 670417 42193 670473
rect 41722 669235 41828 669263
rect 41800 668778 41828 669235
rect 41788 668772 41840 668778
rect 41788 668714 41840 668720
rect 41713 668577 42193 668633
rect 41713 667933 42193 667989
rect 41713 666737 42193 666793
rect 41713 666093 42193 666149
rect 41713 665541 42193 665597
rect 41713 664897 42193 664953
rect 41713 664253 42193 664309
rect 41713 663701 42193 663757
rect 42260 663626 42288 670666
rect 41892 663598 42288 663626
rect 41892 663082 41920 663598
rect 41722 663054 41920 663082
rect 42352 662538 42380 689986
rect 41892 662510 42380 662538
rect 41892 662455 41920 662510
rect 41722 662427 41920 662455
rect 41722 661783 41828 661811
rect 41800 661366 41828 661783
rect 41788 661360 41840 661366
rect 41788 661302 41840 661308
rect 41713 661217 42193 661273
rect 41713 660573 42193 660629
rect 41713 659929 42193 659985
rect 41713 659377 42193 659433
rect 41788 659320 41840 659326
rect 41788 659262 41840 659268
rect 41800 658775 41828 659262
rect 41722 658747 41828 658775
rect 42260 658131 42288 662510
rect 42444 659326 42472 701626
rect 42536 661366 42564 704754
rect 42628 668778 42656 713050
rect 673472 684350 673500 723998
rect 673460 684344 673512 684350
rect 673460 684286 673512 684292
rect 673564 683126 673592 728350
rect 673932 725286 673960 769626
rect 674012 761320 674064 761326
rect 674012 761262 674064 761268
rect 673920 725280 673972 725286
rect 673920 725222 673972 725228
rect 673644 717868 673696 717874
rect 673644 717810 673696 717816
rect 673552 683120 673604 683126
rect 673552 683062 673604 683068
rect 673552 680468 673604 680474
rect 673552 680410 673604 680416
rect 42616 668772 42668 668778
rect 42616 668714 42668 668720
rect 42524 661360 42576 661366
rect 42524 661302 42576 661308
rect 42432 659320 42484 659326
rect 42432 659262 42484 659268
rect 41722 658103 42288 658131
rect 41713 657537 42193 657593
rect 41713 656893 42193 656949
rect 41713 656249 42193 656305
rect 41713 655697 42193 655753
rect 42260 651374 42288 658103
rect 42260 651346 42380 651374
rect 41722 627875 42288 627903
rect 41713 627217 42193 627273
rect 41722 626062 41828 626090
rect 41800 625530 41828 626062
rect 41788 625524 41840 625530
rect 41788 625466 41840 625472
rect 41713 625377 42193 625433
rect 41713 624733 42193 624789
rect 41713 623537 42193 623593
rect 41713 622893 42193 622949
rect 41713 622341 42193 622397
rect 41713 621697 42193 621753
rect 41713 621053 42193 621109
rect 41713 620501 42193 620557
rect 42260 620378 42288 627875
rect 41892 620350 42288 620378
rect 41892 619899 41920 620350
rect 41722 619871 41920 619899
rect 41722 619227 41920 619255
rect 41892 619154 41920 619227
rect 42352 619154 42380 651346
rect 41892 619126 42380 619154
rect 41722 618582 41828 618610
rect 41800 618186 41828 618582
rect 41788 618180 41840 618186
rect 41788 618122 41840 618128
rect 41713 618017 42193 618073
rect 41713 617373 42193 617429
rect 41713 616729 42193 616785
rect 41713 616177 42193 616233
rect 41722 615547 41828 615575
rect 41800 615058 41828 615547
rect 41788 615052 41840 615058
rect 41788 614994 41840 615000
rect 41722 614910 41828 614938
rect 41800 614802 41828 614910
rect 42260 614802 42288 619126
rect 42536 618186 42564 661302
rect 42628 625530 42656 668714
rect 42708 659320 42760 659326
rect 42708 659262 42760 659268
rect 42616 625524 42668 625530
rect 42616 625466 42668 625472
rect 42524 618180 42576 618186
rect 42524 618122 42576 618128
rect 41800 614774 42380 614802
rect 42248 614712 42300 614718
rect 42248 614654 42300 614660
rect 41713 614337 42193 614393
rect 41713 613693 42193 613749
rect 41713 613049 42193 613105
rect 41713 612497 42193 612553
rect 42260 584882 42288 614654
rect 42352 604454 42380 614774
rect 42352 604426 42472 604454
rect 42260 584854 42380 584882
rect 41722 584675 42288 584703
rect 41713 584017 42193 584073
rect 41788 583296 41840 583302
rect 41788 583238 41840 583244
rect 41800 582842 41828 583238
rect 41722 582814 41828 582842
rect 41713 582177 42193 582233
rect 41713 581533 42193 581589
rect 41713 580337 42193 580393
rect 41713 579693 42193 579749
rect 41713 579141 42193 579197
rect 41713 578497 42193 578553
rect 41713 577853 42193 577909
rect 41713 577301 42193 577357
rect 42260 576858 42288 584675
rect 41892 576830 42288 576858
rect 41892 576722 41920 576830
rect 41722 576694 41920 576722
rect 41788 576564 41840 576570
rect 41788 576506 41840 576512
rect 42248 576564 42300 576570
rect 42248 576506 42300 576512
rect 41800 576042 41828 576506
rect 41722 576014 41828 576042
rect 41788 575952 41840 575958
rect 41788 575894 41840 575900
rect 41800 575411 41828 575894
rect 41722 575383 41828 575411
rect 41713 574817 42193 574873
rect 41713 574173 42193 574229
rect 41713 573529 42193 573585
rect 41713 572977 42193 573033
rect 41722 572342 41828 572370
rect 41800 571878 41828 572342
rect 41788 571872 41840 571878
rect 41788 571814 41840 571820
rect 42260 571731 42288 576506
rect 42352 574094 42380 584854
rect 42444 576570 42472 604426
rect 42432 576564 42484 576570
rect 42432 576506 42484 576512
rect 42536 575958 42564 618122
rect 42628 583302 42656 625466
rect 42720 615058 42748 659262
rect 673564 636342 673592 680410
rect 673656 673674 673684 717810
rect 673736 683120 673788 683126
rect 673736 683062 673788 683068
rect 673644 673668 673696 673674
rect 673644 673610 673696 673616
rect 673748 643094 673776 683062
rect 673932 680474 673960 725222
rect 674024 717874 674052 761262
rect 674012 717868 674064 717874
rect 674012 717810 674064 717816
rect 673920 680468 673972 680474
rect 673920 680410 673972 680416
rect 673828 680128 673880 680134
rect 673828 680070 673880 680076
rect 673656 643066 673776 643094
rect 673656 638926 673684 643066
rect 673840 640150 673868 680070
rect 674012 673668 674064 673674
rect 674012 673610 674064 673616
rect 673828 640144 673880 640150
rect 673828 640086 673880 640092
rect 673644 638920 673696 638926
rect 673644 638862 673696 638868
rect 673552 636336 673604 636342
rect 673552 636278 673604 636284
rect 673460 629468 673512 629474
rect 673460 629410 673512 629416
rect 42708 615052 42760 615058
rect 42708 614994 42760 615000
rect 673472 584186 673500 629410
rect 673564 591938 673592 636278
rect 673656 595202 673684 638862
rect 673736 635792 673788 635798
rect 673736 635734 673788 635740
rect 673748 596154 673776 635734
rect 674024 629474 674052 673610
rect 674012 629468 674064 629474
rect 674012 629410 674064 629416
rect 673736 596148 673788 596154
rect 673736 596090 673788 596096
rect 673644 595196 673696 595202
rect 673644 595138 673696 595144
rect 673552 591932 673604 591938
rect 673552 591874 673604 591880
rect 673460 584180 673512 584186
rect 673460 584122 673512 584128
rect 42616 583296 42668 583302
rect 42616 583238 42668 583244
rect 42524 575952 42576 575958
rect 42524 575894 42576 575900
rect 42352 574066 42472 574094
rect 42444 571878 42472 574066
rect 42432 571872 42484 571878
rect 42432 571814 42484 571820
rect 41722 571703 42380 571731
rect 41713 571137 42193 571193
rect 41713 570493 42193 570549
rect 41713 569849 42193 569905
rect 41713 569297 42193 569353
rect 41722 541470 41828 541498
rect 41800 541362 41828 541470
rect 41800 541334 42288 541362
rect 41713 540817 42193 540873
rect 41788 540116 41840 540122
rect 41788 540058 41840 540064
rect 41800 539663 41828 540058
rect 41722 539635 41828 539663
rect 41713 538977 42193 539033
rect 41713 538333 42193 538389
rect 41713 537137 42193 537193
rect 41713 536493 42193 536549
rect 41713 535941 42193 535997
rect 41713 535297 42193 535353
rect 41713 534653 42193 534709
rect 41713 534101 42193 534157
rect 42260 533610 42288 541334
rect 41892 533582 42288 533610
rect 41892 533474 41920 533582
rect 41722 533446 41920 533474
rect 42352 532855 42380 571703
rect 41722 532827 42380 532855
rect 41722 532183 41828 532211
rect 41800 531826 41828 532183
rect 41788 531820 41840 531826
rect 41788 531762 41840 531768
rect 41713 531617 42193 531673
rect 41713 530973 42193 531029
rect 41713 530329 42193 530385
rect 41713 529777 42193 529833
rect 41722 529147 41828 529175
rect 41800 528698 41828 529147
rect 41788 528692 41840 528698
rect 41788 528634 41840 528640
rect 41722 528503 41920 528531
rect 41892 528442 41920 528503
rect 42260 528442 42288 532827
rect 42444 528698 42472 571814
rect 42536 531826 42564 575894
rect 42628 540122 42656 583238
rect 673564 548282 673592 591874
rect 673656 551410 673684 595138
rect 673736 590844 673788 590850
rect 673736 590786 673788 590792
rect 673748 551546 673776 590786
rect 673920 584180 673972 584186
rect 673920 584122 673972 584128
rect 673736 551540 673788 551546
rect 673736 551482 673788 551488
rect 673644 551404 673696 551410
rect 673644 551346 673696 551352
rect 673552 548276 673604 548282
rect 673552 548218 673604 548224
rect 673460 547052 673512 547058
rect 673460 546994 673512 547000
rect 42616 540116 42668 540122
rect 42616 540058 42668 540064
rect 42524 531820 42576 531826
rect 42524 531762 42576 531768
rect 42432 528692 42484 528698
rect 42432 528634 42484 528640
rect 41892 528414 42288 528442
rect 41713 527937 42193 527993
rect 41713 527293 42193 527349
rect 41713 526649 42193 526705
rect 41713 526097 42193 526153
rect 42260 419534 42288 528414
rect 42260 419506 42380 419534
rect 41722 413675 42288 413703
rect 41713 413017 42193 413073
rect 41722 411862 41828 411890
rect 41800 411330 41828 411862
rect 41788 411324 41840 411330
rect 41788 411266 41840 411272
rect 41713 411177 42193 411233
rect 41713 410533 42193 410589
rect 41713 409337 42193 409393
rect 41713 408693 42193 408749
rect 41713 408141 42193 408197
rect 41713 407497 42193 407553
rect 41713 406853 42193 406909
rect 41713 406301 42193 406357
rect 42260 405770 42288 413675
rect 41892 405742 42288 405770
rect 41892 405699 41920 405742
rect 41722 405671 41920 405699
rect 42352 405498 42380 419506
rect 41800 405470 42380 405498
rect 41800 405055 41828 405470
rect 41722 405027 41828 405055
rect 41788 404932 41840 404938
rect 41788 404874 41840 404880
rect 41800 404410 41828 404874
rect 41722 404382 41828 404410
rect 41713 403817 42193 403873
rect 41713 403173 42193 403229
rect 41713 402529 42193 402585
rect 41713 401977 42193 402033
rect 41788 401940 41840 401946
rect 41788 401882 41840 401888
rect 41800 401375 41828 401882
rect 41722 401347 41828 401375
rect 42260 400738 42288 405470
rect 42444 401946 42472 528634
rect 42628 419534 42656 540058
rect 42708 531820 42760 531826
rect 42708 531762 42760 531768
rect 42536 419506 42656 419534
rect 42536 411330 42564 419506
rect 42524 411324 42576 411330
rect 42524 411266 42576 411272
rect 42432 401940 42484 401946
rect 42432 401882 42484 401888
rect 41722 400710 42288 400738
rect 41713 400137 42193 400193
rect 41713 399493 42193 399549
rect 41713 398849 42193 398905
rect 41713 398297 42193 398353
rect 42260 380894 42288 400710
rect 42260 380866 42380 380894
rect 41722 370475 42288 370503
rect 41713 369817 42193 369873
rect 41788 369096 41840 369102
rect 41788 369038 41840 369044
rect 41800 368642 41828 369038
rect 41722 368614 41828 368642
rect 41713 367977 42193 368033
rect 41713 367333 42193 367389
rect 41713 366137 42193 366193
rect 41713 365493 42193 365549
rect 41713 364941 42193 364997
rect 41713 364297 42193 364353
rect 41713 363653 42193 363709
rect 41713 363101 42193 363157
rect 42260 362658 42288 370475
rect 41800 362630 42288 362658
rect 41800 362522 41828 362630
rect 41722 362494 41828 362522
rect 41722 361814 41828 361842
rect 41800 361574 41828 361814
rect 42352 361574 42380 380866
rect 41800 361546 42380 361574
rect 41788 361344 41840 361350
rect 41788 361286 41840 361292
rect 41800 361211 41828 361286
rect 41722 361183 41828 361211
rect 41713 360617 42193 360673
rect 41713 359973 42193 360029
rect 41713 359329 42193 359385
rect 41713 358777 42193 358833
rect 41722 358142 41828 358170
rect 41800 357678 41828 358142
rect 41788 357672 41840 357678
rect 41788 357614 41840 357620
rect 42260 357531 42288 361546
rect 42444 357678 42472 401882
rect 42536 369102 42564 411266
rect 42720 404938 42748 531762
rect 42708 404932 42760 404938
rect 42708 404874 42760 404880
rect 42720 400214 42748 404874
rect 42628 400186 42748 400214
rect 42524 369096 42576 369102
rect 42524 369038 42576 369044
rect 42432 357672 42484 357678
rect 42432 357614 42484 357620
rect 41722 357503 42380 357531
rect 41713 356937 42193 356993
rect 41713 356293 42193 356349
rect 41713 355649 42193 355705
rect 41713 355097 42193 355153
rect 41722 327075 42288 327103
rect 41713 326417 42193 326473
rect 41788 325712 41840 325718
rect 41788 325654 41840 325660
rect 41800 325258 41828 325654
rect 41722 325230 41828 325258
rect 41713 324577 42193 324633
rect 41713 323933 42193 323989
rect 41713 322737 42193 322793
rect 41713 322093 42193 322149
rect 41713 321541 42193 321597
rect 41713 320897 42193 320953
rect 41713 320253 42193 320309
rect 41713 319701 42193 319757
rect 42260 319099 42288 327075
rect 41722 319071 42288 319099
rect 41722 318430 41920 318458
rect 41892 318322 41920 318430
rect 42352 318322 42380 357503
rect 42536 325718 42564 369038
rect 42628 361350 42656 400186
rect 673472 380894 673500 546994
rect 673932 540938 673960 584122
rect 673920 540932 673972 540938
rect 673920 540874 673972 540880
rect 674760 422278 674788 996406
rect 677600 954121 678010 958901
rect 677600 944142 682732 948922
rect 675407 862647 675887 862703
rect 675407 862095 675887 862151
rect 675407 861451 675887 861507
rect 675407 860807 675887 860863
rect 675312 860254 675418 860282
rect 675312 855973 675340 860254
rect 675404 859178 675432 859639
rect 675392 859172 675444 859178
rect 675392 859114 675444 859120
rect 675407 858967 675887 859023
rect 675407 858415 675887 858471
rect 675407 857771 675887 857827
rect 675407 857127 675887 857183
rect 675404 856118 675432 856596
rect 675392 856112 675444 856118
rect 675392 856054 675444 856060
rect 675312 855959 675418 855973
rect 675312 855945 675432 855959
rect 675404 855438 675432 855945
rect 675392 855432 675444 855438
rect 675392 855374 675444 855380
rect 675312 855301 675418 855329
rect 675312 847325 675340 855301
rect 675407 854643 675887 854699
rect 675407 854091 675887 854147
rect 675407 853447 675887 853503
rect 675407 852803 675887 852859
rect 675407 852251 675887 852307
rect 675407 851607 675887 851663
rect 675407 850411 675887 850467
rect 675407 849767 675887 849823
rect 675392 849720 675444 849726
rect 675392 849662 675444 849668
rect 675404 849151 675432 849662
rect 675407 847927 675887 847983
rect 675312 847297 675418 847325
rect 677598 803856 677654 803865
rect 675300 803820 675352 803826
rect 677598 803791 677600 803800
rect 675300 803762 675352 803768
rect 677652 803791 677654 803800
rect 677600 803762 677652 803768
rect 675208 773356 675260 773362
rect 675208 773298 675260 773304
rect 675220 769146 675248 773298
rect 675208 769140 675260 769146
rect 675208 769082 675260 769088
rect 675208 767644 675260 767650
rect 675208 767586 675260 767592
rect 675220 760238 675248 767586
rect 675208 760232 675260 760238
rect 675208 760174 675260 760180
rect 675312 739694 675340 803762
rect 675407 775247 675887 775303
rect 675407 774695 675887 774751
rect 675407 774051 675887 774107
rect 675407 773407 675887 773463
rect 675392 773356 675444 773362
rect 675392 773298 675444 773304
rect 675404 772883 675432 773298
rect 675392 772812 675444 772818
rect 675392 772754 675444 772760
rect 675404 772239 675432 772754
rect 675407 771567 675887 771623
rect 675407 771015 675887 771071
rect 675407 770371 675887 770427
rect 675407 769727 675887 769783
rect 675392 769684 675444 769690
rect 675392 769626 675444 769632
rect 675404 769203 675432 769626
rect 675392 769140 675444 769146
rect 675392 769082 675444 769088
rect 675404 768559 675432 769082
rect 675404 767650 675432 767924
rect 675392 767644 675444 767650
rect 675392 767586 675444 767592
rect 675407 767243 675887 767299
rect 675407 766691 675887 766747
rect 675407 766047 675887 766103
rect 675407 765403 675887 765459
rect 675407 764851 675887 764907
rect 675407 764207 675887 764263
rect 675407 763011 675887 763067
rect 675407 762367 675887 762423
rect 675404 761326 675432 761751
rect 675392 761320 675444 761326
rect 675392 761262 675444 761268
rect 675407 760527 675887 760583
rect 675392 760232 675444 760238
rect 675392 760174 675444 760180
rect 675404 759900 675432 760174
rect 675128 739666 675340 739694
rect 675128 709334 675156 739666
rect 675407 730847 675887 730903
rect 675407 730295 675887 730351
rect 675407 729651 675887 729707
rect 675407 729007 675887 729063
rect 675392 728612 675444 728618
rect 675392 728554 675444 728560
rect 675404 728498 675432 728554
rect 675312 728484 675432 728498
rect 675312 728470 675418 728484
rect 675312 724690 675340 728470
rect 675392 728408 675444 728414
rect 675392 728350 675444 728356
rect 675404 727839 675432 728350
rect 675407 727167 675887 727223
rect 675407 726615 675887 726671
rect 675407 725971 675887 726027
rect 675407 725327 675887 725383
rect 675392 725280 675444 725286
rect 675392 725222 675444 725228
rect 675404 724812 675432 725222
rect 675312 724662 675432 724690
rect 675404 724062 675432 724662
rect 675392 724056 675444 724062
rect 675392 723998 675444 724004
rect 675220 723501 675418 723529
rect 675220 715525 675248 723501
rect 675407 722843 675887 722899
rect 675407 722291 675887 722347
rect 675407 721647 675887 721703
rect 675407 721003 675887 721059
rect 675407 720451 675887 720507
rect 675407 719807 675887 719863
rect 675407 718611 675887 718667
rect 675407 717967 675887 718023
rect 675392 717868 675444 717874
rect 675392 717810 675444 717816
rect 675404 717332 675432 717810
rect 675407 716127 675887 716183
rect 675220 715497 675418 715525
rect 675128 709306 675340 709334
rect 675312 690014 675340 709306
rect 675128 689986 675340 690014
rect 675128 670694 675156 689986
rect 675407 686647 675887 686703
rect 675407 686095 675887 686151
rect 675407 685451 675887 685507
rect 675407 684807 675887 684863
rect 675312 684350 675340 684381
rect 675300 684344 675352 684350
rect 675352 684292 675418 684298
rect 675300 684286 675418 684292
rect 675312 684270 675418 684286
rect 675312 680354 675340 684270
rect 675404 683126 675432 683639
rect 675392 683120 675444 683126
rect 675392 683062 675444 683068
rect 675407 682967 675887 683023
rect 675407 682415 675887 682471
rect 675407 681771 675887 681827
rect 675407 681127 675887 681183
rect 675404 680474 675432 680612
rect 675392 680468 675444 680474
rect 675392 680410 675444 680416
rect 675312 680326 675432 680354
rect 675404 680134 675432 680326
rect 675392 680128 675444 680134
rect 675392 680070 675444 680076
rect 675404 679932 675432 680070
rect 675404 678842 675432 679315
rect 675208 678836 675260 678842
rect 675208 678778 675260 678784
rect 675392 678836 675444 678842
rect 675392 678778 675444 678784
rect 675220 671325 675248 678778
rect 675407 678643 675887 678699
rect 675407 678091 675887 678147
rect 675407 677447 675887 677503
rect 675407 676803 675887 676859
rect 675407 676251 675887 676307
rect 675407 675607 675887 675663
rect 675407 674411 675887 674467
rect 675407 673767 675887 673823
rect 675392 673668 675444 673674
rect 675392 673610 675444 673616
rect 675404 673132 675432 673610
rect 675407 671927 675887 671983
rect 675220 671297 675418 671325
rect 675128 670666 675340 670694
rect 675312 651374 675340 670666
rect 675128 651346 675340 651374
rect 675128 623774 675156 651346
rect 675407 642447 675887 642503
rect 675407 641895 675887 641951
rect 675407 641251 675887 641307
rect 675407 640607 675887 640663
rect 675312 640150 675340 640181
rect 675300 640144 675352 640150
rect 675352 640092 675418 640098
rect 675300 640086 675418 640092
rect 675312 640070 675418 640086
rect 675312 635882 675340 640070
rect 675404 638926 675432 639439
rect 675392 638920 675444 638926
rect 675392 638862 675444 638868
rect 675407 638767 675887 638823
rect 675407 638215 675887 638271
rect 675407 637571 675887 637627
rect 675407 636927 675887 636983
rect 675404 636342 675432 636412
rect 675392 636336 675444 636342
rect 675392 636278 675444 636284
rect 675312 635854 675432 635882
rect 675312 635798 675340 635854
rect 675300 635792 675352 635798
rect 675300 635734 675352 635740
rect 675404 635732 675432 635854
rect 675404 634642 675432 635115
rect 675208 634636 675260 634642
rect 675208 634578 675260 634584
rect 675392 634636 675444 634642
rect 675392 634578 675444 634584
rect 675220 627125 675248 634578
rect 675407 634443 675887 634499
rect 675407 633891 675887 633947
rect 675407 633247 675887 633303
rect 675407 632603 675887 632659
rect 675407 632051 675887 632107
rect 675407 631407 675887 631463
rect 675407 630211 675887 630267
rect 675407 629567 675887 629623
rect 675392 629468 675444 629474
rect 675392 629410 675444 629416
rect 675404 628932 675432 629410
rect 675407 627727 675887 627783
rect 675220 627097 675418 627125
rect 675128 623746 675340 623774
rect 675208 596148 675260 596154
rect 675208 596090 675260 596096
rect 675220 590850 675248 596090
rect 675208 590844 675260 590850
rect 675208 590786 675260 590792
rect 675312 590322 675340 623746
rect 675407 598047 675887 598103
rect 675407 597495 675887 597551
rect 675407 596851 675887 596907
rect 675407 596207 675887 596263
rect 675392 596148 675444 596154
rect 675392 596090 675444 596096
rect 675404 595683 675432 596090
rect 675392 595196 675444 595202
rect 675392 595138 675444 595144
rect 675404 595039 675432 595138
rect 675407 594367 675887 594423
rect 675407 593815 675887 593871
rect 675407 593171 675887 593227
rect 675407 592527 675887 592583
rect 675404 591938 675432 592003
rect 675392 591932 675444 591938
rect 675392 591874 675444 591880
rect 675404 590850 675432 591359
rect 675392 590844 675444 590850
rect 675392 590786 675444 590792
rect 675128 590294 675340 590322
rect 675128 535454 675156 590294
rect 675404 590186 675432 590716
rect 675312 590158 675432 590186
rect 675312 583250 675340 590158
rect 675407 590043 675887 590099
rect 675407 589491 675887 589547
rect 675407 588847 675887 588903
rect 675407 588203 675887 588259
rect 675407 587651 675887 587707
rect 675407 587007 675887 587063
rect 675407 585811 675887 585867
rect 675407 585167 675887 585223
rect 675404 584186 675432 584551
rect 675392 584180 675444 584186
rect 675392 584122 675444 584128
rect 675407 583327 675887 583383
rect 675312 583222 675432 583250
rect 675404 582692 675432 583222
rect 675407 553847 675887 553903
rect 675407 553295 675887 553351
rect 675407 552651 675887 552707
rect 675407 552007 675887 552063
rect 675220 551546 675248 551580
rect 675208 551540 675260 551546
rect 675260 551488 675418 551497
rect 675208 551482 675418 551488
rect 675220 551469 675418 551482
rect 675220 547058 675248 551469
rect 675392 551404 675444 551410
rect 675392 551346 675444 551352
rect 675404 550839 675432 551346
rect 675407 550167 675887 550223
rect 675407 549615 675887 549671
rect 675407 548971 675887 549027
rect 675407 548327 675887 548383
rect 675392 548276 675444 548282
rect 675392 548218 675444 548224
rect 675404 547803 675432 548218
rect 675404 547058 675432 547159
rect 675208 547052 675260 547058
rect 675208 546994 675260 547000
rect 675392 547052 675444 547058
rect 675392 546994 675444 547000
rect 675312 546502 675418 546530
rect 675312 539050 675340 546502
rect 675407 545843 675887 545899
rect 675407 545291 675887 545347
rect 675407 544647 675887 544703
rect 675407 544003 675887 544059
rect 675407 543451 675887 543507
rect 675407 542807 675887 542863
rect 675407 541611 675887 541667
rect 675407 540967 675887 541023
rect 675392 540932 675444 540938
rect 675392 540874 675444 540880
rect 675404 540351 675432 540874
rect 675407 539127 675887 539183
rect 675312 539022 675432 539050
rect 675404 538492 675432 539022
rect 675128 535426 675340 535454
rect 675312 499526 675340 535426
rect 675300 499520 675352 499526
rect 675300 499462 675352 499468
rect 676128 499520 676180 499526
rect 676128 499462 676180 499468
rect 676140 494902 676168 499462
rect 676128 494896 676180 494902
rect 677968 494896 678020 494902
rect 676128 494838 676180 494844
rect 677966 494864 677968 494873
rect 678020 494864 678022 494873
rect 677966 494799 678022 494808
rect 674012 422272 674064 422278
rect 674012 422214 674064 422220
rect 674748 422272 674800 422278
rect 674748 422214 674800 422220
rect 674024 419937 674052 422214
rect 674010 419928 674066 419937
rect 674010 419863 674066 419872
rect 674010 419248 674066 419257
rect 674010 419183 674012 419192
rect 674064 419183 674066 419192
rect 677508 419212 677560 419218
rect 674012 419154 674064 419160
rect 677508 419154 677560 419160
rect 677520 418441 677548 419154
rect 677506 418432 677562 418441
rect 677506 418367 677562 418376
rect 673472 380866 673592 380894
rect 673564 372842 673592 380866
rect 675407 379647 675887 379703
rect 675407 379095 675887 379151
rect 675407 378451 675887 378507
rect 675407 377807 675887 377863
rect 675312 377269 675418 377297
rect 673920 376168 673972 376174
rect 673920 376110 673972 376116
rect 673736 373108 673788 373114
rect 673736 373050 673788 373056
rect 673552 372836 673604 372842
rect 673552 372778 673604 372784
rect 42616 361344 42668 361350
rect 42616 361286 42668 361292
rect 42524 325712 42576 325718
rect 42524 325654 42576 325660
rect 42536 322934 42564 325654
rect 41892 318294 42380 318322
rect 42444 322906 42564 322934
rect 41722 317783 41828 317811
rect 41800 317422 41828 317783
rect 41788 317416 41840 317422
rect 41788 317358 41840 317364
rect 41713 317217 42193 317273
rect 41713 316573 42193 316629
rect 41713 315929 42193 315985
rect 41713 315377 42193 315433
rect 41722 314758 41828 314786
rect 41800 314294 41828 314758
rect 41788 314288 41840 314294
rect 41788 314230 41840 314236
rect 41722 314078 41920 314106
rect 41892 313970 41920 314078
rect 42260 313970 42288 318294
rect 41892 313942 42288 313970
rect 41713 313537 42193 313593
rect 42260 313138 42288 313942
rect 42248 313132 42300 313138
rect 42248 313074 42300 313080
rect 42444 313018 42472 322906
rect 42628 317422 42656 361286
rect 42708 357672 42760 357678
rect 42708 357614 42760 357620
rect 42616 317416 42668 317422
rect 42616 317358 42668 317364
rect 42524 314288 42576 314294
rect 42524 314230 42576 314236
rect 42260 312990 42472 313018
rect 41713 312893 42193 312949
rect 41713 312249 42193 312305
rect 41713 311697 42193 311753
rect 42260 284050 42288 312990
rect 42340 312928 42392 312934
rect 42340 312870 42392 312876
rect 42352 284170 42380 312870
rect 42340 284164 42392 284170
rect 42340 284106 42392 284112
rect 42260 284022 42472 284050
rect 42340 283960 42392 283966
rect 41722 283886 42288 283914
rect 42340 283902 42392 283908
rect 41713 283217 42193 283273
rect 41722 282035 41828 282063
rect 41800 281586 41828 282035
rect 41788 281580 41840 281586
rect 41788 281522 41840 281528
rect 41713 281377 42193 281433
rect 41713 280733 42193 280789
rect 41713 279537 42193 279593
rect 41713 278893 42193 278949
rect 41713 278341 42193 278397
rect 41713 277697 42193 277753
rect 41713 277053 42193 277109
rect 41713 276501 42193 276557
rect 42260 276026 42288 283886
rect 41800 275998 42288 276026
rect 41800 275890 41828 275998
rect 41722 275862 41828 275890
rect 42352 275346 42380 283902
rect 42444 281586 42472 284022
rect 42432 281580 42484 281586
rect 42432 281522 42484 281528
rect 41800 275318 42380 275346
rect 41800 275255 41828 275318
rect 41722 275227 41828 275255
rect 41788 274712 41840 274718
rect 41788 274654 41840 274660
rect 41800 274611 41828 274654
rect 41722 274583 41828 274611
rect 41713 274017 42193 274073
rect 41713 273373 42193 273429
rect 41713 272729 42193 272785
rect 41713 272177 42193 272233
rect 41788 272128 41840 272134
rect 41788 272070 41840 272076
rect 41800 271575 41828 272070
rect 41722 271547 41828 271575
rect 42260 270931 42288 275318
rect 42536 272134 42564 314230
rect 42628 274718 42656 317358
rect 42720 314294 42748 357614
rect 673564 333130 673592 372778
rect 673748 334014 673776 373050
rect 673736 334008 673788 334014
rect 673736 333950 673788 333956
rect 673552 333124 673604 333130
rect 673552 333066 673604 333072
rect 673932 331974 673960 376110
rect 675312 372858 675340 377269
rect 675404 376174 675432 376652
rect 675392 376168 675444 376174
rect 675392 376110 675444 376116
rect 675407 375967 675887 376023
rect 675407 375415 675887 375471
rect 675407 374771 675887 374827
rect 675407 374127 675887 374183
rect 675404 373114 675432 373603
rect 675392 373108 675444 373114
rect 675392 373050 675444 373056
rect 675404 372858 675432 372980
rect 675312 372842 675432 372858
rect 675312 372836 675444 372842
rect 675312 372830 675392 372836
rect 675392 372778 675444 372784
rect 675312 372286 675418 372314
rect 674012 365764 674064 365770
rect 674012 365706 674064 365712
rect 673460 331968 673512 331974
rect 673460 331910 673512 331916
rect 673920 331968 673972 331974
rect 673920 331910 673972 331916
rect 42708 314288 42760 314294
rect 42708 314230 42760 314236
rect 673472 288794 673500 331910
rect 673552 328908 673604 328914
rect 673552 328850 673604 328856
rect 673460 288788 673512 288794
rect 673460 288730 673512 288736
rect 42708 281580 42760 281586
rect 42708 281522 42760 281528
rect 42616 274712 42668 274718
rect 42616 274654 42668 274660
rect 42524 272128 42576 272134
rect 42524 272070 42576 272076
rect 41722 270903 42288 270931
rect 41713 270337 42193 270393
rect 41713 269693 42193 269749
rect 41713 269049 42193 269105
rect 41713 268497 42193 268553
rect 42260 264974 42288 270903
rect 42260 264946 42380 264974
rect 41722 240675 42288 240703
rect 41713 240017 42193 240073
rect 41722 238835 41828 238863
rect 41800 238338 41828 238835
rect 41788 238332 41840 238338
rect 41788 238274 41840 238280
rect 41713 238177 42193 238233
rect 41713 236337 42193 236393
rect 41713 235141 42193 235197
rect 41713 234497 42193 234553
rect 41713 233853 42193 233909
rect 41713 233301 42193 233357
rect 42260 232778 42288 240675
rect 41800 232750 42288 232778
rect 41800 232699 41828 232750
rect 41722 232671 41828 232699
rect 42352 232506 42380 264946
rect 42432 238332 42484 238338
rect 42432 238274 42484 238280
rect 41800 232478 42380 232506
rect 41800 232055 41828 232478
rect 41722 232027 41828 232055
rect 41788 231940 41840 231946
rect 41788 231882 41840 231888
rect 41800 231418 41828 231882
rect 41722 231390 41828 231418
rect 41713 230817 42193 230873
rect 41713 230173 42193 230229
rect 41713 229529 42193 229585
rect 41713 228977 42193 229033
rect 41788 228880 41840 228886
rect 41788 228822 41840 228828
rect 41800 228375 41828 228822
rect 41722 228347 41828 228375
rect 42260 227882 42288 232478
rect 41800 227854 42288 227882
rect 41800 227746 41828 227854
rect 41722 227718 41828 227746
rect 41713 227137 42193 227193
rect 41713 226493 42193 226549
rect 42260 226334 42288 227854
rect 42260 226306 42380 226334
rect 41713 225849 42193 225905
rect 41713 225297 42193 225353
rect 41722 197475 42288 197503
rect 41713 196817 42193 196873
rect 41722 195622 41828 195650
rect 41800 195158 41828 195622
rect 41788 195152 41840 195158
rect 41788 195094 41840 195100
rect 41713 194977 42193 195033
rect 41713 193137 42193 193193
rect 41713 191941 42193 191997
rect 41713 191297 42193 191353
rect 41713 190653 42193 190709
rect 41713 190101 42193 190157
rect 42260 189530 42288 197475
rect 41708 189502 42288 189530
rect 41708 189485 41736 189502
rect 42352 188986 42380 226306
rect 42444 195158 42472 238274
rect 42536 228886 42564 272070
rect 42628 231946 42656 274654
rect 42720 238338 42748 281522
rect 673472 243778 673500 288730
rect 673564 285326 673592 328850
rect 673736 328296 673788 328302
rect 673736 328238 673788 328244
rect 673644 322516 673696 322522
rect 673644 322458 673696 322464
rect 673552 285320 673604 285326
rect 673552 285262 673604 285268
rect 673460 243772 673512 243778
rect 673460 243714 673512 243720
rect 42708 238332 42760 238338
rect 42708 238274 42760 238280
rect 42616 231940 42668 231946
rect 42616 231882 42668 231888
rect 42628 231826 42656 231882
rect 42628 231798 42840 231826
rect 42524 228880 42576 228886
rect 42524 228822 42576 228828
rect 42536 226334 42564 228822
rect 42536 226306 42748 226334
rect 42432 195152 42484 195158
rect 42432 195094 42484 195100
rect 41892 188958 42380 188986
rect 41892 188850 41920 188958
rect 41722 188822 41920 188850
rect 41788 188760 41840 188766
rect 41788 188702 41840 188708
rect 41800 188211 41828 188702
rect 41722 188183 41828 188211
rect 41713 187617 42193 187673
rect 41713 186973 42193 187029
rect 41713 186329 42193 186385
rect 41713 185777 42193 185833
rect 41788 185700 41840 185706
rect 41788 185642 41840 185648
rect 41800 185178 41828 185642
rect 41722 185150 41828 185178
rect 42260 184531 42288 188958
rect 41722 184503 42380 184531
rect 42248 184408 42300 184414
rect 42248 184350 42300 184356
rect 41713 183937 42193 183993
rect 41713 183293 42193 183349
rect 41713 182649 42193 182705
rect 41713 182097 42193 182153
rect 39670 80200 39726 80209
rect 39670 80135 39726 80144
rect 39684 78305 39712 80135
rect 39670 78296 39726 78305
rect 39670 78231 39726 78240
rect 42260 45694 42288 184350
rect 42248 45688 42300 45694
rect 42248 45630 42300 45636
rect 42352 45626 42380 184503
rect 42444 106078 42472 195094
rect 42524 188760 42576 188766
rect 42524 188702 42576 188708
rect 42536 121514 42564 188702
rect 42720 185706 42748 226306
rect 42812 188766 42840 231798
rect 673472 199170 673500 243714
rect 673564 240310 673592 285262
rect 673656 277370 673684 322458
rect 673748 289338 673776 328238
rect 674024 322522 674052 365706
rect 675312 364325 675340 372286
rect 675407 371643 675887 371699
rect 675407 371091 675887 371147
rect 675407 370447 675887 370503
rect 675407 369803 675887 369859
rect 675407 368607 675887 368663
rect 675407 366767 675887 366823
rect 675404 365770 675432 366151
rect 675392 365764 675444 365770
rect 675392 365706 675444 365712
rect 675407 364927 675887 364983
rect 675312 364297 675418 364325
rect 675407 335447 675887 335503
rect 675407 334895 675887 334951
rect 675407 334251 675887 334307
rect 675208 334008 675260 334014
rect 675208 333950 675260 333956
rect 675220 328914 675248 333950
rect 675407 333607 675887 333663
rect 675312 333130 675340 333180
rect 675300 333124 675352 333130
rect 675352 333072 675418 333097
rect 675300 333069 675418 333072
rect 675300 333066 675352 333069
rect 675208 328908 675260 328914
rect 675208 328850 675260 328856
rect 675312 328658 675340 333066
rect 675404 331974 675432 332452
rect 675392 331968 675444 331974
rect 675392 331910 675444 331916
rect 675407 331767 675887 331823
rect 675407 331215 675887 331271
rect 675407 330571 675887 330627
rect 675407 329927 675887 329983
rect 675404 328914 675432 329403
rect 675392 328908 675444 328914
rect 675392 328850 675444 328856
rect 675404 328658 675432 328780
rect 675312 328630 675432 328658
rect 675404 328302 675432 328630
rect 675392 328296 675444 328302
rect 675392 328238 675444 328244
rect 675312 328086 675418 328114
rect 674012 322516 674064 322522
rect 674012 322458 674064 322464
rect 675312 320125 675340 328086
rect 675407 327443 675887 327499
rect 675407 326891 675887 326947
rect 675407 326247 675887 326303
rect 675407 325603 675887 325659
rect 675407 324407 675887 324463
rect 675407 322567 675887 322623
rect 675392 322516 675444 322522
rect 675392 322458 675444 322464
rect 675404 321951 675432 322458
rect 675407 320727 675887 320783
rect 675312 320097 675418 320125
rect 675407 291247 675887 291303
rect 675407 290695 675887 290751
rect 675407 290051 675887 290107
rect 675407 289407 675887 289463
rect 673736 289332 673788 289338
rect 673736 289274 673788 289280
rect 675392 289332 675444 289338
rect 675392 289274 675444 289280
rect 675404 288897 675432 289274
rect 675312 288883 675432 288897
rect 675312 288869 675418 288883
rect 675312 285138 675340 288869
rect 675392 288788 675444 288794
rect 675392 288730 675444 288736
rect 675404 288252 675432 288730
rect 675407 287567 675887 287623
rect 675407 287015 675887 287071
rect 675407 286371 675887 286427
rect 675407 285727 675887 285783
rect 675392 285320 675444 285326
rect 675392 285262 675444 285268
rect 675404 285203 675432 285262
rect 675312 285110 675432 285138
rect 675404 284102 675432 285110
rect 673736 284096 673788 284102
rect 673736 284038 673788 284044
rect 675392 284096 675444 284102
rect 675392 284038 675444 284044
rect 673644 277364 673696 277370
rect 673644 277306 673696 277312
rect 673552 240304 673604 240310
rect 673552 240246 673604 240252
rect 673460 199164 673512 199170
rect 673460 199106 673512 199112
rect 42800 188760 42852 188766
rect 42800 188702 42852 188708
rect 42708 185700 42760 185706
rect 42708 185642 42760 185648
rect 42720 184414 42748 185642
rect 42708 184408 42760 184414
rect 42708 184350 42760 184356
rect 673472 155990 673500 199106
rect 673564 197062 673592 240246
rect 673656 233918 673684 277306
rect 673748 244662 673776 284038
rect 675312 283886 675418 283914
rect 675312 275925 675340 283886
rect 675407 283243 675887 283299
rect 675407 282691 675887 282747
rect 675407 282047 675887 282103
rect 675407 281403 675887 281459
rect 675407 280207 675887 280263
rect 675407 278367 675887 278423
rect 675404 277370 675432 277751
rect 675392 277364 675444 277370
rect 675392 277306 675444 277312
rect 675407 276527 675887 276583
rect 675312 275897 675418 275925
rect 675407 246847 675887 246903
rect 675407 246295 675887 246351
rect 675407 245651 675887 245707
rect 675407 245007 675887 245063
rect 673736 244656 673788 244662
rect 673736 244598 673788 244604
rect 675392 244656 675444 244662
rect 675392 244598 675444 244604
rect 675404 243930 675432 244598
rect 675312 243902 675432 243930
rect 675312 240173 675340 243902
rect 675404 243778 675432 243839
rect 675392 243772 675444 243778
rect 675392 243714 675444 243720
rect 675407 243167 675887 243223
rect 675407 242615 675887 242671
rect 675407 241971 675887 242027
rect 675407 241327 675887 241383
rect 675404 240310 675432 240788
rect 675392 240304 675444 240310
rect 675392 240246 675444 240252
rect 675312 240159 675418 240173
rect 675312 240145 675432 240159
rect 675404 239698 675432 240145
rect 673736 239692 673788 239698
rect 673736 239634 673788 239640
rect 675392 239692 675444 239698
rect 675392 239634 675444 239640
rect 673644 233912 673696 233918
rect 673644 233854 673696 233860
rect 673552 197056 673604 197062
rect 673552 196998 673604 197004
rect 673460 155984 673512 155990
rect 673460 155926 673512 155932
rect 673564 152862 673592 196998
rect 673656 189310 673684 233854
rect 673748 200462 673776 239634
rect 675312 239501 675418 239529
rect 675312 231525 675340 239501
rect 675407 238843 675887 238899
rect 675407 238291 675887 238347
rect 675407 237647 675887 237703
rect 675407 237003 675887 237059
rect 675407 235807 675887 235863
rect 675407 233967 675887 234023
rect 675392 233912 675444 233918
rect 675392 233854 675444 233860
rect 675404 233351 675432 233854
rect 675407 232127 675887 232183
rect 675312 231497 675418 231525
rect 675407 202647 675887 202703
rect 675407 202095 675887 202151
rect 675407 201451 675887 201507
rect 675407 200807 675887 200863
rect 673736 200456 673788 200462
rect 673736 200398 673788 200404
rect 675392 200456 675444 200462
rect 675392 200398 675444 200404
rect 675404 199730 675432 200398
rect 675312 199702 675432 199730
rect 675312 195973 675340 199702
rect 675404 199170 675432 199639
rect 675392 199164 675444 199170
rect 675392 199106 675444 199112
rect 675407 198967 675887 199023
rect 675407 198415 675887 198471
rect 675407 197771 675887 197827
rect 675407 197127 675887 197183
rect 675392 197056 675444 197062
rect 675392 196998 675444 197004
rect 675404 196588 675432 196998
rect 675312 195959 675418 195973
rect 675312 195945 675432 195959
rect 675404 195838 675432 195945
rect 673736 195832 673788 195838
rect 673736 195774 673788 195780
rect 675392 195832 675444 195838
rect 675392 195774 675444 195780
rect 673644 189304 673696 189310
rect 673644 189246 673696 189252
rect 673552 152856 673604 152862
rect 673552 152798 673604 152804
rect 42524 121508 42576 121514
rect 42524 121450 42576 121456
rect 44180 121508 44232 121514
rect 44180 121450 44232 121456
rect 44192 110537 44220 121450
rect 673460 111580 673512 111586
rect 673460 111522 673512 111528
rect 44178 110528 44234 110537
rect 44178 110463 44234 110472
rect 44822 110528 44878 110537
rect 44822 110463 44878 110472
rect 44836 110414 44864 110463
rect 44836 110386 44956 110414
rect 42432 106072 42484 106078
rect 42432 106014 42484 106020
rect 44180 106072 44232 106078
rect 44180 106014 44232 106020
rect 44192 80209 44220 106014
rect 44178 80200 44234 80209
rect 44178 80135 44234 80144
rect 44822 80200 44878 80209
rect 44822 80135 44878 80144
rect 44836 46986 44864 80135
rect 44824 46980 44876 46986
rect 44824 46922 44876 46928
rect 42340 45620 42392 45626
rect 42340 45562 42392 45568
rect 44928 45558 44956 110386
rect 143540 46912 143592 46918
rect 200856 46912 200908 46918
rect 143540 46854 143592 46860
rect 151726 46880 151782 46889
rect 140964 45688 141016 45694
rect 140964 45630 141016 45636
rect 44916 45552 44968 45558
rect 44916 45494 44968 45500
rect 93768 41540 93820 41546
rect 93768 41482 93820 41488
rect 93780 40225 93808 41482
rect 135168 40248 135220 40254
rect 93766 40216 93822 40225
rect 93766 40151 93822 40160
rect 135166 40216 135168 40225
rect 135220 40216 135222 40225
rect 140976 40202 141004 45630
rect 143552 40497 143580 46854
rect 151726 46815 151782 46824
rect 188526 46880 188582 46889
rect 200856 46854 200908 46860
rect 256240 46912 256292 46918
rect 256240 46854 256292 46860
rect 297732 46912 297784 46918
rect 297732 46854 297784 46860
rect 309416 46912 309468 46918
rect 309416 46854 309468 46860
rect 352564 46912 352616 46918
rect 352564 46854 352616 46860
rect 364248 46912 364300 46918
rect 364248 46854 364300 46860
rect 407396 46912 407448 46918
rect 407396 46854 407448 46860
rect 419080 46912 419132 46918
rect 419080 46854 419132 46860
rect 462136 46912 462188 46918
rect 462136 46854 462188 46860
rect 473820 46912 473872 46918
rect 473820 46854 473872 46860
rect 516968 46912 517020 46918
rect 516968 46854 517020 46860
rect 527456 46912 527508 46918
rect 527456 46854 527508 46860
rect 188526 46815 188582 46824
rect 143632 45620 143684 45626
rect 143632 45562 143684 45568
rect 143644 44198 143672 45562
rect 143632 44192 143684 44198
rect 143632 44134 143684 44140
rect 145104 44192 145156 44198
rect 145104 44134 145156 44140
rect 143538 40488 143594 40497
rect 143538 40423 143594 40432
rect 143540 40248 143592 40254
rect 143078 40216 143134 40225
rect 140976 40174 141036 40202
rect 135166 40151 135222 40160
rect 141008 40118 141036 40174
rect 143078 40151 143134 40160
rect 143538 40216 143540 40225
rect 143592 40216 143594 40225
rect 145116 40202 145144 44134
rect 146300 41880 146352 41886
rect 146300 41822 146352 41828
rect 143538 40151 143594 40160
rect 145103 40174 145144 40202
rect 143084 40118 143112 40151
rect 140996 40112 141048 40118
rect 140996 40054 141048 40060
rect 143072 40112 143124 40118
rect 143072 40054 143124 40060
rect 144552 40112 144604 40118
rect 144552 40054 144604 40060
rect 141008 39984 141036 40054
rect 143084 39916 143112 40054
rect 144564 39916 144592 40054
rect 145103 40000 145131 40174
rect 146312 40118 146340 41822
rect 151740 40497 151768 46815
rect 186688 45620 186740 45626
rect 186688 45562 186740 45568
rect 186700 41820 186728 45562
rect 188540 44402 188568 46815
rect 194692 45620 194744 45626
rect 194692 45562 194744 45568
rect 188528 44396 188580 44402
rect 188528 44338 188580 44344
rect 192852 44396 192904 44402
rect 192852 44338 192904 44344
rect 187327 41713 187383 42193
rect 188540 41820 188568 44338
rect 189264 41948 189316 41954
rect 189264 41890 189316 41896
rect 191104 41948 191156 41954
rect 191104 41890 191156 41896
rect 192300 41948 192352 41954
rect 192300 41890 192352 41896
rect 189276 41834 189304 41890
rect 191116 41834 191144 41890
rect 192312 41834 192340 41890
rect 189198 41806 189304 41834
rect 191038 41806 191144 41834
rect 192234 41806 192340 41834
rect 192864 41820 192892 44338
rect 193588 41948 193640 41954
rect 193588 41890 193640 41896
rect 193600 41834 193628 41890
rect 193522 41806 193628 41834
rect 194043 41713 194099 42193
rect 194704 41820 194732 45562
rect 195980 45552 196032 45558
rect 195980 45494 196032 45500
rect 195992 44334 196020 45494
rect 195980 44328 196032 44334
rect 195980 44270 196032 44276
rect 195336 44192 195388 44198
rect 195336 44134 195388 44140
rect 195348 41820 195376 44134
rect 195992 41820 196020 44270
rect 199844 44260 199896 44266
rect 199844 44202 199896 44208
rect 199660 44192 199712 44198
rect 199856 44146 199884 44202
rect 199712 44140 199884 44146
rect 199660 44134 199884 44140
rect 199672 44118 199884 44134
rect 196440 41948 196492 41954
rect 196440 41890 196492 41896
rect 198464 41948 198516 41954
rect 198464 41890 198516 41896
rect 196452 41834 196480 41890
rect 198476 41834 198504 41890
rect 196452 41806 198504 41834
rect 198936 41818 199042 41834
rect 199672 41820 199700 44118
rect 200120 41948 200172 41954
rect 200120 41890 200172 41896
rect 200132 41834 200160 41890
rect 200868 41834 200896 46854
rect 201500 44328 201552 44334
rect 201500 44270 201552 44276
rect 200132 41820 200896 41834
rect 201512 41820 201540 44270
rect 198924 41812 199042 41818
rect 198976 41806 199042 41812
rect 200132 41806 200882 41820
rect 198924 41754 198976 41760
rect 151726 40488 151782 40497
rect 151726 40423 151782 40432
rect 146300 40112 146352 40118
rect 146300 40054 146352 40060
rect 145091 39706 145143 40000
rect 256252 39545 256280 46854
rect 297088 44396 297140 44402
rect 297088 44338 297140 44344
rect 295248 44328 295300 44334
rect 295248 44270 295300 44276
rect 295260 41834 295288 44270
rect 297100 41834 297128 44338
rect 297744 41834 297772 46854
rect 299572 44396 299624 44402
rect 299572 44338 299624 44344
rect 305736 44396 305788 44402
rect 305736 44338 305788 44344
rect 297916 41948 297968 41954
rect 297916 41890 297968 41896
rect 297928 41834 297956 41890
rect 295260 41806 295311 41834
rect 297100 41806 297151 41834
rect 297744 41806 297956 41834
rect 299584 41834 299612 44338
rect 303252 44328 303304 44334
rect 303252 44270 303304 44276
rect 300676 41948 300728 41954
rect 300676 41890 300728 41896
rect 302240 41948 302292 41954
rect 302240 41890 302292 41896
rect 300688 41834 300716 41890
rect 302252 41834 302280 41890
rect 299584 41806 299635 41834
rect 300688 41806 302280 41834
rect 302643 41713 302699 42193
rect 303264 41834 303292 44270
rect 303896 44260 303948 44266
rect 303896 44202 303948 44208
rect 303908 41834 303936 44202
rect 304540 44192 304592 44198
rect 304540 44134 304592 44140
rect 304552 41834 304580 44134
rect 305276 41948 305328 41954
rect 305276 41890 305328 41896
rect 305288 41834 305316 41890
rect 303264 41806 303315 41834
rect 303908 41806 303959 41834
rect 304552 41806 304603 41834
rect 305155 41806 305316 41834
rect 305748 41834 305776 44338
rect 308220 44260 308272 44266
rect 308220 44202 308272 44208
rect 306564 41948 306616 41954
rect 306564 41890 306616 41896
rect 306576 41834 306604 41890
rect 305748 41806 305799 41834
rect 306443 41806 306604 41834
rect 306967 41713 307023 42193
rect 308232 41834 308260 44202
rect 308680 41948 308732 41954
rect 308680 41890 308732 41896
rect 308692 41834 308720 41890
rect 309428 41834 309456 46854
rect 349988 44464 350040 44470
rect 349988 44406 350040 44412
rect 350000 44198 350028 44406
rect 351920 44328 351972 44334
rect 351920 44270 351972 44276
rect 349988 44192 350040 44198
rect 349988 44134 350040 44140
rect 350080 44192 350132 44198
rect 350080 44134 350132 44140
rect 307639 41818 307800 41834
rect 307639 41812 307812 41818
rect 307639 41806 307760 41812
rect 308232 41806 308283 41834
rect 308692 41806 309479 41834
rect 307760 41754 307812 41760
rect 310095 41713 310151 42193
rect 350092 41820 350120 44134
rect 351932 41820 351960 44270
rect 352576 41970 352604 46854
rect 359372 44464 359424 44470
rect 359372 44406 359424 44412
rect 354404 44328 354456 44334
rect 354404 44270 354456 44276
rect 352576 41954 352696 41970
rect 352576 41948 352708 41954
rect 352576 41942 352656 41948
rect 352576 41820 352604 41942
rect 352656 41890 352708 41896
rect 354416 41820 354444 44270
rect 358728 44260 358780 44266
rect 358728 44202 358780 44208
rect 358084 44192 358136 44198
rect 358084 44134 358136 44140
rect 355508 41948 355560 41954
rect 355508 41890 355560 41896
rect 356980 41948 357032 41954
rect 356980 41890 357032 41896
rect 355520 41834 355548 41890
rect 356992 41834 357020 41890
rect 355520 41806 357020 41834
rect 357443 41713 357499 42193
rect 358096 41820 358124 44134
rect 358740 41820 358768 44202
rect 359384 41820 359412 44406
rect 360568 44328 360620 44334
rect 360568 44270 360620 44276
rect 363052 44328 363104 44334
rect 363052 44270 363104 44276
rect 360580 44198 360608 44270
rect 360568 44192 360620 44198
rect 360568 44134 360620 44140
rect 359832 41948 359884 41954
rect 359832 41890 359884 41896
rect 359844 41834 359872 41890
rect 359844 41806 359950 41834
rect 360580 41820 360608 44134
rect 361120 41948 361172 41954
rect 361120 41890 361172 41896
rect 361132 41834 361160 41890
rect 361132 41806 361238 41834
rect 361767 41713 361823 42193
rect 362434 41818 362540 41834
rect 363064 41820 363092 44270
rect 363512 41948 363564 41954
rect 363512 41890 363564 41896
rect 363524 41834 363552 41890
rect 364260 41834 364288 46854
rect 404910 44296 404966 44305
rect 404910 44231 404966 44240
rect 406752 44260 406804 44266
rect 363524 41820 364288 41834
rect 362434 41812 362552 41818
rect 362434 41806 362500 41812
rect 363524 41806 364274 41820
rect 362500 41754 362552 41760
rect 364895 41713 364951 42193
rect 404924 41820 404952 44231
rect 406752 44202 406804 44208
rect 405527 41713 405583 42193
rect 406764 41820 406792 44202
rect 407408 41970 407436 46854
rect 414204 44464 414256 44470
rect 411074 44432 411130 44441
rect 414204 44406 414256 44412
rect 411074 44367 411130 44376
rect 407408 41954 407528 41970
rect 407408 41948 407540 41954
rect 407408 41942 407488 41948
rect 407408 41820 407436 41942
rect 407488 41890 407540 41896
rect 410248 41948 410300 41954
rect 410248 41890 410300 41896
rect 410260 41834 410288 41890
rect 409262 41818 409368 41834
rect 409262 41812 409380 41818
rect 409262 41806 409328 41812
rect 410260 41806 410458 41834
rect 411088 41820 411116 44367
rect 413560 44328 413612 44334
rect 412914 44296 412970 44305
rect 413560 44270 413612 44276
rect 412914 44231 412970 44240
rect 411536 41948 411588 41954
rect 411536 41890 411588 41896
rect 411548 41834 411576 41890
rect 412243 41834 412299 42193
rect 411548 41806 411746 41834
rect 412243 41818 412404 41834
rect 412928 41820 412956 44231
rect 413572 41820 413600 44270
rect 414216 44198 414244 44406
rect 417884 44328 417936 44334
rect 417884 44270 417936 44276
rect 414204 44192 414256 44198
rect 414204 44134 414256 44140
rect 414216 41820 414244 44134
rect 414572 41948 414624 41954
rect 414572 41890 414624 41896
rect 415860 41948 415912 41954
rect 415860 41890 415912 41896
rect 414584 41834 414612 41890
rect 415872 41834 415900 41890
rect 412243 41812 412416 41818
rect 412243 41806 412364 41812
rect 409328 41754 409380 41760
rect 412243 41713 412299 41806
rect 414584 41806 414782 41834
rect 415228 41818 415426 41834
rect 415216 41812 415426 41818
rect 412364 41754 412416 41760
rect 415268 41806 415426 41812
rect 415872 41806 416070 41834
rect 415216 41754 415268 41760
rect 416567 41713 416623 42193
rect 417266 41818 417372 41834
rect 417896 41820 417924 44270
rect 418252 41948 418304 41954
rect 418252 41890 418304 41896
rect 418264 41834 418292 41890
rect 419092 41834 419120 46854
rect 419722 44296 419778 44305
rect 419722 44231 419778 44240
rect 459650 44296 459706 44305
rect 459650 44231 459706 44240
rect 461492 44260 461544 44266
rect 419736 42193 419764 44231
rect 418264 41820 419120 41834
rect 419695 41820 419764 42193
rect 459664 41834 459692 44231
rect 461492 44202 461544 44208
rect 417266 41812 417384 41818
rect 417266 41806 417332 41812
rect 418264 41806 419106 41820
rect 417332 41754 417384 41760
rect 419695 41713 419751 41820
rect 459664 41806 459711 41834
rect 460327 41713 460383 42193
rect 461504 41834 461532 44202
rect 462148 41834 462176 46854
rect 465814 44432 465870 44441
rect 465814 44367 465870 44376
rect 468944 44396 468996 44402
rect 462320 41948 462372 41954
rect 462320 41890 462372 41896
rect 465080 41948 465132 41954
rect 465080 41890 465132 41896
rect 462332 41834 462360 41890
rect 465092 41834 465120 41890
rect 465828 41834 465856 44367
rect 468944 44338 468996 44344
rect 468300 44328 468352 44334
rect 467654 44296 467710 44305
rect 468300 44270 468352 44276
rect 467654 44231 467710 44240
rect 466368 41948 466420 41954
rect 466368 41890 466420 41896
rect 466380 41834 466408 41890
rect 467043 41834 467099 42193
rect 467668 41834 467696 44231
rect 468312 41834 468340 44270
rect 468956 44198 468984 44338
rect 472624 44328 472676 44334
rect 472624 44270 472676 44276
rect 468944 44192 468996 44198
rect 468944 44134 468996 44140
rect 468956 41834 468984 44134
rect 469404 41948 469456 41954
rect 469404 41890 469456 41896
rect 470692 41948 470744 41954
rect 470692 41890 470744 41896
rect 469416 41834 469444 41890
rect 470704 41834 470732 41890
rect 461504 41806 461551 41834
rect 462148 41806 462360 41834
rect 464035 41818 464200 41834
rect 464035 41812 464212 41818
rect 464035 41806 464160 41812
rect 465092 41806 465231 41834
rect 465828 41806 465875 41834
rect 466380 41806 466519 41834
rect 467043 41818 467236 41834
rect 467043 41812 467248 41818
rect 467043 41806 467196 41812
rect 464160 41754 464212 41760
rect 467043 41713 467099 41806
rect 467668 41806 467715 41834
rect 468312 41806 468359 41834
rect 468956 41806 469003 41834
rect 469416 41806 469555 41834
rect 470060 41818 470199 41834
rect 470048 41812 470199 41818
rect 467196 41754 467248 41760
rect 470100 41806 470199 41812
rect 470704 41806 470843 41834
rect 470048 41754 470100 41760
rect 471367 41713 471423 42193
rect 472636 41834 472664 44270
rect 473084 41948 473136 41954
rect 473084 41890 473136 41896
rect 473096 41834 473124 41890
rect 473832 41834 473860 46854
rect 474462 44432 474518 44441
rect 474462 44367 474518 44376
rect 474476 42193 474504 44367
rect 514482 44296 514538 44305
rect 514482 44231 514538 44240
rect 516324 44260 516376 44266
rect 472039 41818 472204 41834
rect 472039 41812 472216 41818
rect 472039 41806 472164 41812
rect 472636 41806 472683 41834
rect 473096 41806 473879 41834
rect 474476 41806 474551 42193
rect 514496 41820 514524 44231
rect 516324 44202 516376 44208
rect 472164 41754 472216 41760
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 516336 41820 516364 44202
rect 516980 41970 517008 46854
rect 523776 45620 523828 45626
rect 523776 45562 523828 45568
rect 518716 45552 518768 45558
rect 518716 45494 518768 45500
rect 518728 44266 518756 45494
rect 522486 44432 522542 44441
rect 523788 44402 523816 45562
rect 522486 44367 522542 44376
rect 523776 44396 523828 44402
rect 518806 44296 518862 44305
rect 518716 44260 518768 44266
rect 518806 44231 518862 44240
rect 518716 44202 518768 44208
rect 516980 41954 517100 41970
rect 516980 41948 517112 41954
rect 516980 41942 517060 41948
rect 516980 41820 517008 41942
rect 517060 41890 517112 41896
rect 518820 41820 518848 44231
rect 519912 41948 519964 41954
rect 519912 41890 519964 41896
rect 519924 41834 519952 41890
rect 519924 41806 520030 41834
rect 520647 41713 520703 42193
rect 521200 41948 521252 41954
rect 521200 41890 521252 41896
rect 521212 41834 521240 41890
rect 521212 41806 521318 41834
rect 521843 41713 521899 42193
rect 522500 41820 522528 44367
rect 523776 44338 523828 44344
rect 523132 44192 523184 44198
rect 523132 44134 523184 44140
rect 523144 41820 523172 44134
rect 523788 41820 523816 44338
rect 524970 44296 525026 44305
rect 524970 44231 525026 44240
rect 524984 42193 525012 44231
rect 527468 44198 527496 46854
rect 527456 44192 527508 44198
rect 527456 44134 527508 44140
rect 524236 41948 524288 41954
rect 524236 41890 524288 41896
rect 524248 41834 524276 41890
rect 524248 41806 524354 41834
rect 524971 41713 525027 42193
rect 525524 41948 525576 41954
rect 525524 41890 525576 41896
rect 525536 41834 525564 41890
rect 525536 41806 525642 41834
rect 526167 41713 526223 42193
rect 526732 41818 526838 41834
rect 527468 41820 527496 44134
rect 673472 42770 673500 111522
rect 673564 108458 673592 152798
rect 673656 149054 673684 189246
rect 673748 156330 673776 195774
rect 675312 195301 675418 195329
rect 675312 187325 675340 195301
rect 675407 194643 675887 194699
rect 675407 194091 675887 194147
rect 675407 193447 675887 193503
rect 675407 192803 675887 192859
rect 675407 191607 675887 191663
rect 675407 189767 675887 189823
rect 675392 189304 675444 189310
rect 675392 189246 675444 189252
rect 675404 189151 675432 189246
rect 675407 187927 675887 187983
rect 675312 187297 675418 187325
rect 675407 158447 675887 158503
rect 675407 157895 675887 157951
rect 675407 157251 675887 157307
rect 675407 156607 675887 156663
rect 673736 156324 673788 156330
rect 673736 156266 673788 156272
rect 675392 156324 675444 156330
rect 675392 156266 675444 156272
rect 675404 156210 675432 156266
rect 675312 156182 675432 156210
rect 673920 155984 673972 155990
rect 673920 155926 673972 155932
rect 673828 151768 673880 151774
rect 673828 151710 673880 151716
rect 673656 149026 673776 149054
rect 673748 144566 673776 149026
rect 673736 144560 673788 144566
rect 673736 144502 673788 144508
rect 673552 108452 673604 108458
rect 673552 108394 673604 108400
rect 673564 45626 673592 108394
rect 673644 107364 673696 107370
rect 673644 107306 673696 107312
rect 673656 46986 673684 107306
rect 673748 100609 673776 144502
rect 673840 111858 673868 151710
rect 673828 111852 673880 111858
rect 673828 111794 673880 111800
rect 673932 111586 673960 155926
rect 675312 151774 675340 156182
rect 675404 156060 675432 156182
rect 675392 155984 675444 155990
rect 675392 155926 675444 155932
rect 675404 155439 675432 155926
rect 675407 154767 675887 154823
rect 675407 154215 675887 154271
rect 675407 153571 675887 153627
rect 675407 152927 675887 152983
rect 675392 152856 675444 152862
rect 675392 152798 675444 152804
rect 675404 152388 675432 152798
rect 675300 151773 675352 151774
rect 675300 151768 675418 151773
rect 675352 151745 675418 151768
rect 675300 151710 675352 151716
rect 675312 151662 675340 151710
rect 675312 151101 675418 151129
rect 675312 143125 675340 151101
rect 675407 150443 675887 150499
rect 675407 149891 675887 149947
rect 675407 149247 675887 149303
rect 675407 148603 675887 148659
rect 675407 147407 675887 147463
rect 675407 145567 675887 145623
rect 675404 144566 675432 144951
rect 675392 144560 675444 144566
rect 675392 144502 675444 144508
rect 675407 143727 675887 143783
rect 675312 143097 675418 143125
rect 675407 114047 675887 114103
rect 675407 113495 675887 113551
rect 675407 112851 675887 112907
rect 675407 112207 675887 112263
rect 675392 111852 675444 111858
rect 675392 111794 675444 111800
rect 675404 111697 675432 111794
rect 675312 111683 675432 111697
rect 675312 111669 675418 111683
rect 673920 111580 673972 111586
rect 673920 111522 673972 111528
rect 675312 107386 675340 111669
rect 675392 111580 675444 111586
rect 675392 111522 675444 111528
rect 675404 111044 675432 111522
rect 675407 110367 675887 110423
rect 675407 109815 675887 109871
rect 675407 109171 675887 109227
rect 675407 108527 675887 108583
rect 675392 108452 675444 108458
rect 675392 108394 675444 108400
rect 675404 108003 675432 108394
rect 675312 107370 675418 107386
rect 675300 107364 675418 107370
rect 675352 107358 675418 107364
rect 675300 107306 675352 107312
rect 675312 107275 675340 107306
rect 675312 106814 675432 106842
rect 673734 100600 673790 100609
rect 673734 100535 673790 100544
rect 673644 46980 673696 46986
rect 673644 46922 673696 46928
rect 673552 45620 673604 45626
rect 673552 45562 673604 45568
rect 673748 45558 673776 100535
rect 675312 98725 675340 106814
rect 675404 106692 675432 106814
rect 675407 106043 675887 106099
rect 675407 105491 675887 105547
rect 675407 104847 675887 104903
rect 675407 104203 675887 104259
rect 675407 103007 675887 103063
rect 675407 101167 675887 101223
rect 675390 100600 675446 100609
rect 675390 100535 675446 100544
rect 675407 99327 675887 99383
rect 675312 98697 675418 98725
rect 673736 45552 673788 45558
rect 673736 45494 673788 45500
rect 579896 42764 579948 42770
rect 579896 42706 579948 42712
rect 673460 42764 673512 42770
rect 673460 42706 673512 42712
rect 527916 41948 527968 41954
rect 527916 41890 527968 41896
rect 527928 41834 527956 41890
rect 526720 41812 526838 41818
rect 526772 41806 526838 41812
rect 527928 41806 528678 41834
rect 526720 41754 526772 41760
rect 529295 41713 529351 42193
rect 579908 41886 579936 42706
rect 568856 41880 568908 41886
rect 568856 41822 568908 41828
rect 579896 41880 579948 41886
rect 579896 41822 579948 41828
rect 568868 39681 568896 41822
rect 568854 39672 568910 39681
rect 568854 39607 568910 39616
rect 256238 39536 256294 39545
rect 256238 39471 256294 39480
<< via2 >>
rect 585782 997464 585838 997520
rect 339498 997056 339554 997112
rect 44178 885808 44234 885864
rect 44822 885808 44878 885864
rect 44178 870984 44234 871040
rect 677598 803820 677654 803856
rect 677598 803800 677600 803820
rect 677600 803800 677652 803820
rect 677652 803800 677654 803820
rect 677966 494844 677968 494864
rect 677968 494844 678020 494864
rect 678020 494844 678022 494864
rect 677966 494808 678022 494844
rect 674010 419872 674066 419928
rect 674010 419212 674066 419248
rect 674010 419192 674012 419212
rect 674012 419192 674064 419212
rect 674064 419192 674066 419212
rect 677506 418376 677562 418432
rect 39670 80144 39726 80200
rect 39670 78240 39726 78296
rect 44178 110472 44234 110528
rect 44822 110472 44878 110528
rect 44178 80144 44234 80200
rect 44822 80144 44878 80200
rect 93766 40160 93822 40216
rect 135166 40196 135168 40216
rect 135168 40196 135220 40216
rect 135220 40196 135222 40216
rect 135166 40160 135222 40196
rect 151726 46824 151782 46880
rect 188526 46824 188582 46880
rect 143538 40432 143594 40488
rect 143078 40160 143134 40216
rect 143538 40196 143540 40216
rect 143540 40196 143592 40216
rect 143592 40196 143594 40216
rect 143538 40160 143594 40196
rect 151726 40432 151782 40488
rect 404910 44240 404966 44296
rect 411074 44376 411130 44432
rect 412914 44240 412970 44296
rect 419722 44240 419778 44296
rect 459650 44240 459706 44296
rect 465814 44376 465870 44432
rect 467654 44240 467710 44296
rect 474462 44376 474518 44432
rect 514482 44240 514538 44296
rect 522486 44376 522542 44432
rect 518806 44240 518862 44296
rect 524970 44240 525026 44296
rect 673734 100544 673790 100600
rect 675390 100544 675446 100600
rect 568854 39616 568910 39672
rect 256238 39480 256294 39536
<< metal3 >>
rect 79944 997600 84944 1014070
rect 127944 997600 132944 1014070
rect 175944 997600 180944 1014070
rect 239478 997600 253800 1000736
rect 290878 997600 305200 1000736
rect 339542 997117 339602 997628
rect 429744 997600 434744 1014070
rect 479144 997600 484144 1014070
rect 530744 997600 535744 1014070
rect 585734 997525 585794 997628
rect 631944 997600 636944 1014070
rect 585734 997520 585843 997525
rect 585734 997464 585782 997520
rect 585838 997464 585843 997520
rect 585734 997462 585843 997464
rect 585777 997459 585843 997462
rect 339493 997112 339602 997117
rect 339493 997056 339498 997112
rect 339554 997056 339602 997112
rect 339493 997054 339602 997056
rect 339493 997051 339559 997054
rect 23530 960144 40000 965144
rect 677600 934600 680736 948922
rect 44173 885866 44239 885869
rect 44817 885866 44883 885869
rect 44173 885864 44883 885866
rect 44173 885808 44178 885864
rect 44234 885808 44822 885864
rect 44878 885808 44883 885864
rect 44173 885806 44883 885808
rect 44173 885803 44239 885806
rect 44817 885803 44883 885806
rect 44173 871042 44239 871045
rect 39652 871040 44239 871042
rect 39652 870984 44178 871040
rect 44234 870984 44239 871040
rect 39652 870982 44239 870984
rect 44173 870979 44239 870982
rect 677593 803858 677659 803861
rect 677734 803858 677794 803964
rect 677593 803856 677794 803858
rect 677593 803800 677598 803856
rect 677654 803800 677794 803856
rect 677593 803798 677794 803800
rect 677593 803795 677659 803798
rect 677764 495214 677978 495274
rect 677918 494869 677978 495214
rect 677918 494864 678027 494869
rect 677918 494808 677966 494864
rect 678022 494808 678027 494864
rect 677918 494806 678027 494808
rect 677961 494803 678027 494806
rect 678000 461700 685920 466500
rect 31680 441300 39600 446100
rect 673862 419868 673868 419932
rect 673932 419930 673938 419932
rect 674005 419930 674071 419933
rect 673932 419928 674071 419930
rect 673932 419872 674010 419928
rect 674066 419872 674071 419928
rect 673932 419870 674071 419872
rect 673932 419868 673938 419870
rect 674005 419867 674071 419870
rect 673862 419188 673868 419252
rect 673932 419250 673938 419252
rect 674005 419250 674071 419253
rect 673932 419248 674071 419250
rect 673932 419192 674010 419248
rect 674066 419192 674071 419248
rect 673932 419190 674071 419192
rect 673932 419188 673938 419190
rect 674005 419187 674071 419190
rect 677501 418434 677567 418437
rect 677734 418434 677794 418540
rect 677501 418432 677794 418434
rect 677501 418376 677506 418432
rect 677562 418376 677794 418432
rect 677501 418374 677794 418376
rect 677501 418371 677567 418374
rect 44173 110530 44239 110533
rect 44817 110530 44883 110533
rect 39652 110528 44883 110530
rect 39652 110472 44178 110528
rect 44234 110472 44822 110528
rect 44878 110472 44883 110528
rect 39652 110470 44883 110472
rect 44173 110467 44239 110470
rect 44817 110467 44883 110470
rect 673729 100602 673795 100605
rect 675385 100602 675451 100605
rect 673729 100600 675451 100602
rect 673729 100544 673734 100600
rect 673790 100544 675390 100600
rect 675446 100544 675451 100600
rect 673729 100542 675451 100544
rect 673729 100539 673795 100542
rect 675385 100539 675451 100542
rect 39665 80202 39731 80205
rect 44173 80202 44239 80205
rect 44817 80202 44883 80205
rect 39665 80200 44883 80202
rect 39665 80144 39670 80200
rect 39726 80144 44178 80200
rect 44234 80144 44822 80200
rect 44878 80144 44883 80200
rect 39665 80142 44883 80144
rect 39665 80139 39731 80142
rect 44173 80139 44239 80142
rect 44817 80139 44883 80142
rect 39665 78298 39731 78301
rect 39468 78296 39731 78298
rect 39468 78240 39670 78296
rect 39726 78240 39731 78296
rect 39468 78238 39731 78240
rect 39665 78235 39731 78238
rect 151721 46882 151787 46885
rect 188521 46882 188587 46885
rect 151721 46880 188587 46882
rect 151721 46824 151726 46880
rect 151782 46824 188526 46880
rect 188582 46824 188587 46880
rect 151721 46822 188587 46824
rect 151721 46819 151787 46822
rect 188521 46819 188587 46822
rect 411069 44434 411135 44437
rect 465809 44434 465875 44437
rect 474457 44434 474523 44437
rect 522481 44434 522547 44437
rect 411069 44432 419550 44434
rect 411069 44376 411074 44432
rect 411130 44376 419550 44432
rect 411069 44374 419550 44376
rect 411069 44371 411135 44374
rect 404905 44298 404971 44301
rect 412909 44298 412975 44301
rect 404905 44296 412975 44298
rect 404905 44240 404910 44296
rect 404966 44240 412914 44296
rect 412970 44240 412975 44296
rect 404905 44238 412975 44240
rect 419490 44298 419550 44374
rect 465809 44432 474523 44434
rect 465809 44376 465814 44432
rect 465870 44376 474462 44432
rect 474518 44376 474523 44432
rect 465809 44374 474523 44376
rect 465809 44371 465875 44374
rect 474457 44371 474523 44374
rect 516090 44432 522547 44434
rect 516090 44376 522486 44432
rect 522542 44376 522547 44432
rect 516090 44374 522547 44376
rect 419717 44298 419783 44301
rect 419490 44296 419783 44298
rect 419490 44240 419722 44296
rect 419778 44240 419783 44296
rect 419490 44238 419783 44240
rect 404905 44235 404971 44238
rect 412909 44235 412975 44238
rect 419717 44235 419783 44238
rect 459645 44298 459711 44301
rect 467649 44298 467715 44301
rect 459645 44296 467715 44298
rect 459645 44240 459650 44296
rect 459706 44240 467654 44296
rect 467710 44240 467715 44296
rect 459645 44238 467715 44240
rect 459645 44235 459711 44238
rect 467649 44235 467715 44238
rect 514477 44298 514543 44301
rect 516090 44298 516150 44374
rect 522481 44371 522547 44374
rect 514477 44296 516150 44298
rect 514477 44240 514482 44296
rect 514538 44240 516150 44296
rect 514477 44238 516150 44240
rect 518801 44298 518867 44301
rect 524965 44298 525031 44301
rect 518801 44296 525031 44298
rect 518801 44240 518806 44296
rect 518862 44240 524970 44296
rect 525026 44240 525031 44296
rect 518801 44238 525031 44240
rect 514477 44235 514543 44238
rect 518801 44235 518867 44238
rect 524965 44235 525031 44238
rect 143533 40490 143599 40493
rect 151721 40490 151787 40493
rect 143533 40488 151787 40490
rect 143533 40432 143538 40488
rect 143594 40432 151726 40488
rect 151782 40432 151787 40488
rect 143533 40430 151787 40432
rect 143533 40427 143599 40430
rect 145790 40354 145850 40430
rect 151721 40427 151787 40430
rect 145790 40294 145898 40354
rect 93761 40218 93827 40221
rect 135161 40218 135227 40221
rect 91142 40216 93827 40218
rect 91142 40160 93766 40216
rect 93822 40160 93827 40216
rect 91142 40158 93827 40160
rect 91142 39644 91202 40158
rect 93761 40155 93827 40158
rect 133094 40216 135227 40218
rect 133094 40160 135166 40216
rect 135222 40160 135227 40216
rect 133094 40158 135227 40160
rect 133094 39984 133154 40158
rect 135161 40155 135227 40158
rect 143073 40218 143139 40221
rect 143533 40218 143599 40221
rect 143073 40216 143458 40218
rect 143073 40160 143078 40216
rect 143134 40160 143458 40216
rect 143073 40158 143458 40160
rect 143073 40155 143139 40158
rect 141667 38031 141813 39999
rect 143398 39984 143458 40158
rect 143533 40216 144010 40218
rect 143533 40160 143538 40216
rect 143594 40160 144010 40216
rect 143533 40158 144010 40160
rect 143533 40155 143599 40158
rect 143950 39984 144010 40158
rect 145838 40014 145898 40294
rect 145820 39954 145898 40014
rect 568849 39674 568915 39677
rect 568849 39672 569204 39674
rect 568849 39616 568854 39672
rect 568910 39616 569204 39672
rect 568849 39614 569204 39616
rect 568849 39611 568915 39614
rect 256233 39538 256299 39541
rect 251406 39536 256299 39538
rect 251406 39480 256238 39536
rect 256294 39480 256299 39536
rect 251406 39478 256299 39480
rect 251406 39372 251466 39478
rect 256233 39475 256299 39478
<< via3 >>
rect 673868 419868 673932 419932
rect 673868 419188 673932 419252
<< metal4 >>
rect 7 456045 4843 456493
rect 28653 441200 28719 456200
rect 32933 455946 33623 456200
rect 36323 456007 37013 456199
rect 37293 455946 38223 456200
rect 38503 455946 39593 456200
rect 679377 451600 680307 451854
rect 680587 451600 681277 451792
rect 688881 451600 688947 466600
rect 673867 419932 673933 419933
rect 673867 419868 673868 419932
rect 673932 419930 673933 419932
rect 673932 419870 674114 419930
rect 673932 419868 673933 419870
rect 673867 419867 673933 419868
rect 673867 419252 673933 419253
rect 673867 419188 673868 419252
rect 673932 419250 673933 419252
rect 674054 419250 674114 419870
rect 673932 419190 674114 419250
rect 673932 419188 673933 419190
rect 673867 419187 673933 419188
rect 132600 36323 132792 37013
rect 132600 30762 132868 31674
rect 132600 28653 147600 28719
<< metal5 >>
rect 76410 1018624 88578 1030788
rect 124410 1018624 136578 1030788
rect 172410 1018624 184578 1030788
rect 230810 1018624 242978 1030788
rect 282210 1018624 294378 1030788
rect 340810 1018624 352978 1030788
rect 426210 1018624 438378 1030788
rect 475610 1018624 487778 1030788
rect 527210 1018624 539378 1030788
rect 577010 1018624 589178 1030788
rect 628410 1018624 640578 1030788
rect 6811 956610 18975 968778
rect 698624 945422 710788 957590
rect 6167 915054 19619 925934
rect 697980 893466 711432 904346
rect 6811 872210 18975 884378
rect 698512 848240 711002 860780
rect 6811 829810 18975 841978
rect 698624 805222 710788 817390
rect 6598 787420 19088 799960
rect 698512 760840 711002 773380
rect 6598 744220 19088 756760
rect 698512 716440 711002 728980
rect 6598 701020 19088 713560
rect 698512 672240 711002 684780
rect 6598 657620 19088 670160
rect 698512 628040 711002 640580
rect 6598 614420 19088 626960
rect 6598 571220 19088 583760
rect 698512 583640 711002 596180
rect 6598 528020 19088 540560
rect 698512 539440 711002 551980
rect 6811 484810 18975 496978
rect 698624 496422 710788 508590
rect 6167 443254 19619 454134
rect 697980 453666 711432 464546
rect 6598 400220 19088 412760
rect 698624 409822 710788 421990
rect 6598 357020 19088 369560
rect 698512 365240 711002 377780
rect 6598 313620 19088 326160
rect 698512 321040 711002 333580
rect 6598 270420 19088 282960
rect 698512 276840 711002 289380
rect 6598 227220 19088 239760
rect 698512 232440 711002 244980
rect 6598 184020 19088 196560
rect 698512 188240 711002 200780
rect 698512 144040 711002 156580
rect 6811 111610 18975 123778
rect 698512 99640 711002 112180
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200180 19088
rect 243266 6167 254146 19619
rect 296240 6598 308780 19088
rect 351040 6598 363580 19088
rect 405840 6598 418380 19088
rect 460640 6598 473180 19088
rect 515440 6598 527980 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use sky130_ef_io__corner_pad  mgmt_corner\[0\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_153 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_357
timestamp 1624635410
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1624635410
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1
timestamp 1624635410
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_157 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_156
timestamp 1624635410
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_155 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_154 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_164
timestamp 1624635410
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1624635410
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1624635410
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1624635410
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_168
timestamp 1624635410
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_167
timestamp 1624635410
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_166
timestamp 1624635410
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_165
timestamp 1624635410
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  mgmt_vssa_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 93800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_170
timestamp 1624635410
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_172
timestamp 1624635410
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_171
timestamp 1624635410
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1624635410
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_174
timestamp 1624635410
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_173
timestamp 1624635410
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1624635410
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1624635410
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1624635410
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1624635410
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1624635410
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_181
timestamp 1624635410
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_185
timestamp 1624635410
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_184
timestamp 1624635410
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_183
timestamp 1624635410
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_182
timestamp 1624635410
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_fd_io__top_xres4v2  resetb_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 147600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1624635410
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_191
timestamp 1624635410
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_190
timestamp 1624635410
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_189
timestamp 1624635410
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_188
timestamp 1624635410
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_187
timestamp 1624635410
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1624635410
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1624635410
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1624635410
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_200
timestamp 1624635410
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_199
timestamp 1624635410
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_198
timestamp 1624635410
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1624635410
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1624635410
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_202
timestamp 1624635410
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_201
timestamp 1624635410
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 202400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1624635410
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_208
timestamp 1624635410
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_207
timestamp 1624635410
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_206
timestamp 1624635410
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_205
timestamp 1624635410
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_204
timestamp 1624635410
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1624635410
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1624635410
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1624635410
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1624635410
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_219
timestamp 1624635410
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_218
timestamp 1624635410
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_217
timestamp 1624635410
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_216
timestamp 1624635410
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_215
timestamp 1624635410
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1624635410
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_clamped_pad  mgmt_vssd_lvclmap_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 256200 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1624635410
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1624635410
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_225
timestamp 1624635410
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_224
timestamp 1624635410
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_223
timestamp 1624635410
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_222
timestamp 1624635410
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_221
timestamp 1624635410
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1624635410
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1624635410
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1624635410
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1624635410
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_236
timestamp 1624635410
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_235
timestamp 1624635410
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_234
timestamp 1624635410
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_233
timestamp 1624635410
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_232
timestamp 1624635410
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1624635410
transform -1 0 311000 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_238
timestamp 1624635410
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_239
timestamp 1624635410
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1624635410
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_242
timestamp 1624635410
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_241
timestamp 1624635410
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_240
timestamp 1624635410
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1624635410
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1624635410
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1624635410
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1624635410
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_253
timestamp 1624635410
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_252
timestamp 1624635410
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_251
timestamp 1624635410
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_250
timestamp 1624635410
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_249
timestamp 1624635410
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1624635410
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1624635410
transform -1 0 365800 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_256
timestamp 1624635410
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_255
timestamp 1624635410
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1624635410
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1624635410
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_259
timestamp 1624635410
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_258
timestamp 1624635410
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_257
timestamp 1624635410
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1624635410
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1624635410
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1624635410
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1624635410
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_270
timestamp 1624635410
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_269
timestamp 1624635410
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_268
timestamp 1624635410
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_267
timestamp 1624635410
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_266
timestamp 1624635410
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1624635410
transform -1 0 420600 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_272
timestamp 1624635410
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1624635410
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1624635410
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1624635410
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_276
timestamp 1624635410
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_275
timestamp 1624635410
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_274
timestamp 1624635410
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_273
timestamp 1624635410
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_283
timestamp 1624635410
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1624635410
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1624635410
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1624635410
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_287
timestamp 1624635410
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_286
timestamp 1624635410
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_285
timestamp 1624635410
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_284
timestamp 1624635410
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1624635410
transform -1 0 475400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_289
timestamp 1624635410
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_290
timestamp 1624635410
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1624635410
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_293
timestamp 1624635410
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_292
timestamp 1624635410
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_291
timestamp 1624635410
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1624635410
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1624635410
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1624635410
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1624635410
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1624635410
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_304
timestamp 1624635410
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_303
timestamp 1624635410
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_302
timestamp 1624635410
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_301
timestamp 1624635410
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_300
timestamp 1624635410
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1624635410
transform -1 0 530200 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1624635410
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_310
timestamp 1624635410
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_309
timestamp 1624635410
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_308
timestamp 1624635410
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_307
timestamp 1624635410
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_306
timestamp 1624635410
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1624635410
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1624635410
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_317
timestamp 1624635410
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1624635410
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1624635410
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1624635410
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_321
timestamp 1624635410
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_320
timestamp 1624635410
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_319
timestamp 1624635410
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_318
timestamp 1624635410
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 584000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_325
timestamp 1624635410
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_324
timestamp 1624635410
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_323
timestamp 1624635410
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1624635410
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1624635410
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1624635410
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1624635410
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_327
timestamp 1624635410
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_326
timestamp 1624635410
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_335
timestamp 1624635410
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_334
timestamp 1624635410
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1624635410
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1624635410
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_338
timestamp 1624635410
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_337
timestamp 1624635410
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_336
timestamp 1624635410
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  mgmt_vdda_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_340
timestamp 1624635410
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_343
timestamp 1624635410
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_342
timestamp 1624635410
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_341
timestamp 1624635410
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1624635410
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_344
timestamp 1624635410
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1624635410
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1624635410
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1624635410
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1624635410
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1624635410
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_351
timestamp 1624635410
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_352
timestamp 1624635410
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1624635410
transform 0 1 676800 -1 0 40000
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_5um  FILLER_353
timestamp 1624635410
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_354
timestamp 1624635410
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_355
timestamp 1624635410
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_356
timestamp 1624635410
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_593
timestamp 1624635410
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_361
timestamp 1624635410
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_360
timestamp 1624635410
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_359
timestamp 1624635410
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_358
timestamp 1624635410
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_365
timestamp 1624635410
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_364
timestamp 1624635410
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_363
timestamp 1624635410
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_362
timestamp 1624635410
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_clamped_pad  mgmt_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 -1 39593 1 0 68000
box 0 -2107 17239 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_367
timestamp 1624635410
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_594
timestamp 1624635410
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1624635410
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1624635410
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_597
timestamp 1624635410
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_598
timestamp 1624635410
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_599
timestamp 1624635410
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_603
timestamp 1624635410
transform 0 1 678007 -1 0 74200
box 0 0 4000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_1 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 1 678007 -1 0 70200
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 1 678007 -1 0 69200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_600
timestamp 1624635410
transform 0 1 678007 -1 0 68200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_604
timestamp 1624635410
transform 0 1 678007 -1 0 78200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1624635410
transform 0 1 678007 -1 0 82200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_606
timestamp 1624635410
transform 0 1 678007 -1 0 86200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_371
timestamp 1624635410
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_370
timestamp 1624635410
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_369
timestamp 1624635410
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_368
timestamp 1624635410
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_375
timestamp 1624635410
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_374
timestamp 1624635410
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_373
timestamp 1624635410
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_372
timestamp 1624635410
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_377
timestamp 1624635410
transform 0 -1 39593 1 0 125200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[0\]
timestamp 1624635410
transform 0 1 675407 -1 0 114400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_607
timestamp 1624635410
transform 0 1 678007 -1 0 90200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_608
timestamp 1624635410
transform 0 1 678007 -1 0 94200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_609
timestamp 1624635410
transform 0 1 678007 -1 0 98200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_610
timestamp 1624635410
transform 0 1 678007 -1 0 98400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_612
timestamp 1624635410
transform 0 1 678007 -1 0 118400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_613
timestamp 1624635410
transform 0 1 678007 -1 0 122400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_614
timestamp 1624635410
transform 0 1 678007 -1 0 126400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1624635410
transform 0 1 678007 -1 0 130400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_378
timestamp 1624635410
transform 0 -1 39593 1 0 129200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_379
timestamp 1624635410
transform 0 -1 39593 1 0 133200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_380
timestamp 1624635410
transform 0 -1 39593 1 0 137200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_381
timestamp 1624635410
transform 0 -1 39593 1 0 141200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_382
timestamp 1624635410
transform 0 -1 39593 1 0 145200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_383
timestamp 1624635410
transform 0 -1 39593 1 0 149200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_388
timestamp 1624635410
transform 0 -1 39593 1 0 154400
box 0 0 4000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_2
timestamp 1624635410
transform 0 -1 39593 1 0 153400
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1624635410
transform 0 -1 39593 1 0 152400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_385
timestamp 1624635410
transform 0 -1 39593 1 0 152200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_384
timestamp 1624635410
transform 0 -1 39593 1 0 151200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_389
timestamp 1624635410
transform 0 -1 39593 1 0 158400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_390
timestamp 1624635410
transform 0 -1 39593 1 0 162400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_391
timestamp 1624635410
transform 0 -1 39593 1 0 166400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[1\]
timestamp 1624635410
transform 0 1 675407 -1 0 158800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_616
timestamp 1624635410
transform 0 1 678007 -1 0 134400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_617
timestamp 1624635410
transform 0 1 678007 -1 0 138400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1624635410
transform 0 1 678007 -1 0 142400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_619
timestamp 1624635410
transform 0 1 678007 -1 0 142600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_620
timestamp 1624635410
transform 0 1 678007 -1 0 142800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_622
timestamp 1624635410
transform 0 1 678007 -1 0 162800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_623
timestamp 1624635410
transform 0 1 678007 -1 0 166800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1624635410
transform 0 1 678007 -1 0 170800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_397
timestamp 1624635410
transform 0 -1 39593 1 0 181600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_396
timestamp 1624635410
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_395
timestamp 1624635410
transform 0 -1 39593 1 0 180400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_394
timestamp 1624635410
transform 0 -1 39593 1 0 178400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_393
timestamp 1624635410
transform 0 -1 39593 1 0 174400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_392
timestamp 1624635410
transform 0 -1 39593 1 0 170400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[12\]
timestamp 1624635410
transform 0 -1 42193 1 0 181800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_399
timestamp 1624635410
transform 0 -1 39593 1 0 197800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_402
timestamp 1624635410
transform 0 -1 39593 1 0 209800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_401
timestamp 1624635410
transform 0 -1 39593 1 0 205800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_400
timestamp 1624635410
transform 0 -1 39593 1 0 201800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[2\]
timestamp 1624635410
transform 0 1 675407 -1 0 203000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_625
timestamp 1624635410
transform 0 1 678007 -1 0 174800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_626
timestamp 1624635410
transform 0 1 678007 -1 0 178800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_627
timestamp 1624635410
transform 0 1 678007 -1 0 182800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1624635410
transform 0 1 678007 -1 0 186800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_629
timestamp 1624635410
transform 0 1 678007 -1 0 187000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_631
timestamp 1624635410
transform 0 1 678007 -1 0 207000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_632
timestamp 1624635410
transform 0 1 678007 -1 0 211000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_407
timestamp 1624635410
transform 0 -1 39593 1 0 224800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_406
timestamp 1624635410
transform 0 -1 39593 1 0 223800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_405
timestamp 1624635410
transform 0 -1 39593 1 0 221800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_404
timestamp 1624635410
transform 0 -1 39593 1 0 217800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_403
timestamp 1624635410
transform 0 -1 39593 1 0 213800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[11\]
timestamp 1624635410
transform 0 -1 42193 1 0 225000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_409
timestamp 1624635410
transform 0 -1 39593 1 0 241000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_412
timestamp 1624635410
transform 0 -1 39593 1 0 253000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_411
timestamp 1624635410
transform 0 -1 39593 1 0 249000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_410
timestamp 1624635410
transform 0 -1 39593 1 0 245000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[3\]
timestamp 1624635410
transform 0 1 675407 -1 0 247200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_633
timestamp 1624635410
transform 0 1 678007 -1 0 215000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1624635410
transform 0 1 678007 -1 0 219000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_635
timestamp 1624635410
transform 0 1 678007 -1 0 223000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_636
timestamp 1624635410
transform 0 1 678007 -1 0 227000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1624635410
transform 0 1 678007 -1 0 231000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_638
timestamp 1624635410
transform 0 1 678007 -1 0 231200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_640
timestamp 1624635410
transform 0 1 678007 -1 0 251200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_641
timestamp 1624635410
transform 0 1 678007 -1 0 255200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[10\]
timestamp 1624635410
transform 0 -1 42193 1 0 268200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_413
timestamp 1624635410
transform 0 -1 39593 1 0 257000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_414
timestamp 1624635410
transform 0 -1 39593 1 0 261000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_415
timestamp 1624635410
transform 0 -1 39593 1 0 265000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_416
timestamp 1624635410
transform 0 -1 39593 1 0 267000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_417
timestamp 1624635410
transform 0 -1 39593 1 0 268000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_419
timestamp 1624635410
transform 0 -1 39593 1 0 284200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_420
timestamp 1624635410
transform 0 -1 39593 1 0 288200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_421
timestamp 1624635410
transform 0 -1 39593 1 0 292200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[4\]
timestamp 1624635410
transform 0 1 675407 -1 0 291600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_642
timestamp 1624635410
transform 0 1 678007 -1 0 259200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1624635410
transform 0 1 678007 -1 0 263200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_644
timestamp 1624635410
transform 0 1 678007 -1 0 267200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_645
timestamp 1624635410
transform 0 1 678007 -1 0 271200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1624635410
transform 0 1 678007 -1 0 275200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_647
timestamp 1624635410
transform 0 1 678007 -1 0 275400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_648
timestamp 1624635410
transform 0 1 678007 -1 0 275600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_650
timestamp 1624635410
transform 0 1 678007 -1 0 295600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_427
timestamp 1624635410
transform 0 -1 39593 1 0 311200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_426
timestamp 1624635410
transform 0 -1 39593 1 0 310200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_425
timestamp 1624635410
transform 0 -1 39593 1 0 308200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_424
timestamp 1624635410
transform 0 -1 39593 1 0 304200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_423
timestamp 1624635410
transform 0 -1 39593 1 0 300200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_422
timestamp 1624635410
transform 0 -1 39593 1 0 296200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[9\]
timestamp 1624635410
transform 0 -1 42193 1 0 311400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_429
timestamp 1624635410
transform 0 -1 39593 1 0 327400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_431
timestamp 1624635410
transform 0 -1 39593 1 0 335400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_430
timestamp 1624635410
transform 0 -1 39593 1 0 331400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[5\]
timestamp 1624635410
transform 0 1 675407 -1 0 335800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_651
timestamp 1624635410
transform 0 1 678007 -1 0 299600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_652
timestamp 1624635410
transform 0 1 678007 -1 0 303600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_653
timestamp 1624635410
transform 0 1 678007 -1 0 307600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_654
timestamp 1624635410
transform 0 1 678007 -1 0 311600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_655
timestamp 1624635410
transform 0 1 678007 -1 0 315600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1624635410
transform 0 1 678007 -1 0 319600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_657
timestamp 1624635410
transform 0 1 678007 -1 0 319800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_659
timestamp 1624635410
transform 0 1 678007 -1 0 339800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_436
timestamp 1624635410
transform 0 -1 39593 1 0 353400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_435
timestamp 1624635410
transform 0 -1 39593 1 0 351400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_434
timestamp 1624635410
transform 0 -1 39593 1 0 347400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_433
timestamp 1624635410
transform 0 -1 39593 1 0 343400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_432
timestamp 1624635410
transform 0 -1 39593 1 0 339400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_438
timestamp 1624635410
transform 0 -1 39593 1 0 354600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_437
timestamp 1624635410
transform 0 -1 39593 1 0 354400
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[8\]
timestamp 1624635410
transform 0 -1 42193 1 0 354800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_442
timestamp 1624635410
transform 0 -1 39593 1 0 378800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_441
timestamp 1624635410
transform 0 -1 39593 1 0 374800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_440
timestamp 1624635410
transform 0 -1 39593 1 0 370800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[6\]
timestamp 1624635410
transform 0 1 675407 -1 0 380000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_660
timestamp 1624635410
transform 0 1 678007 -1 0 343800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_661
timestamp 1624635410
transform 0 1 678007 -1 0 347800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1624635410
transform 0 1 678007 -1 0 351800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_663
timestamp 1624635410
transform 0 1 678007 -1 0 355800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_664
timestamp 1624635410
transform 0 1 678007 -1 0 359800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1624635410
transform 0 1 678007 -1 0 363800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_666
timestamp 1624635410
transform 0 1 678007 -1 0 364000
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[7\]
timestamp 1624635410
transform 0 -1 42193 1 0 398000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_443
timestamp 1624635410
transform 0 -1 39593 1 0 382800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_444
timestamp 1624635410
transform 0 -1 39593 1 0 386800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1624635410
transform 0 -1 39593 1 0 390800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_446
timestamp 1624635410
transform 0 -1 39593 1 0 394800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_447
timestamp 1624635410
transform 0 -1 39593 1 0 396800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_448
timestamp 1624635410
transform 0 -1 39593 1 0 397800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_450
timestamp 1624635410
transform 0 -1 39593 1 0 414000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_451
timestamp 1624635410
transform 0 -1 39593 1 0 418000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1624635410
transform 0 1 678007 -1 0 396000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_670
timestamp 1624635410
transform 0 1 678007 -1 0 392000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_669
timestamp 1624635410
transform 0 1 678007 -1 0 388000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_668
timestamp 1624635410
transform 0 1 678007 -1 0 384000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_676
timestamp 1624635410
transform 0 1 678007 -1 0 408400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_675
timestamp 1624635410
transform 0 1 678007 -1 0 408200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_674
timestamp 1624635410
transform 0 1 678007 -1 0 408000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_673
timestamp 1624635410
transform 0 1 678007 -1 0 404000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_672
timestamp 1624635410
transform 0 1 678007 -1 0 400000
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1624635410
transform 0 1 678007 -1 0 423400
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_458
timestamp 1624635410
transform 0 -1 39593 1 0 441000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_457
timestamp 1624635410
transform 0 -1 39593 1 0 440000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_456
timestamp 1624635410
transform 0 -1 39593 1 0 438000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1624635410
transform 0 -1 39593 1 0 434000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_454
timestamp 1624635410
transform 0 -1 39593 1 0 430000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_453
timestamp 1624635410
transform 0 -1 39593 1 0 426000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_452
timestamp 1624635410
transform 0 -1 39593 1 0 422000
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_clamped2_pad  user2_vssd_lvclmap_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 -1 39593 1 0 441200
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_461
timestamp 1624635410
transform 0 -1 39593 1 0 460200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_460
timestamp 1624635410
transform 0 -1 39593 1 0 456200
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_clamped2_pad  user1_vssd_lvclmap_pad
timestamp 1624635410
transform 0 1 678007 -1 0 466600
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_678
timestamp 1624635410
transform 0 1 678007 -1 0 427400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_679
timestamp 1624635410
transform 0 1 678007 -1 0 431400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_680
timestamp 1624635410
transform 0 1 678007 -1 0 435400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1624635410
transform 0 1 678007 -1 0 439400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_682
timestamp 1624635410
transform 0 1 678007 -1 0 443400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_683
timestamp 1624635410
transform 0 1 678007 -1 0 447400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1624635410
transform 0 1 678007 -1 0 451400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_685
timestamp 1624635410
transform 0 1 678007 -1 0 451600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1624635410
transform 0 -1 39593 1 0 476200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_464
timestamp 1624635410
transform 0 -1 39593 1 0 472200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_463
timestamp 1624635410
transform 0 -1 39593 1 0 468200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_462
timestamp 1624635410
transform 0 -1 39593 1 0 464200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_468
timestamp 1624635410
transform 0 -1 39593 1 0 483200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_467
timestamp 1624635410
transform 0 -1 39593 1 0 482200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_466
timestamp 1624635410
transform 0 -1 39593 1 0 480200
box 0 0 2000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user2_vdda_hvclamp_pad
timestamp 1624635410
transform 0 -1 39593 1 0 483400
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_471
timestamp 1624635410
transform 0 -1 39593 1 0 502400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_470
timestamp 1624635410
transform 0 -1 39593 1 0 498400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1624635410
transform 0 1 678007 -1 0 482600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_689
timestamp 1624635410
transform 0 1 678007 -1 0 478600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_688
timestamp 1624635410
transform 0 1 678007 -1 0 474600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_687
timestamp 1624635410
transform 0 1 678007 -1 0 470600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1624635410
transform 0 1 678007 -1 0 494600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_692
timestamp 1624635410
transform 0 1 678007 -1 0 490600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_691
timestamp 1624635410
transform 0 1 678007 -1 0 486600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_695
timestamp 1624635410
transform 0 1 678007 -1 0 495000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_694
timestamp 1624635410
transform 0 1 678007 -1 0 494800
box 0 0 200 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1624635410
transform 0 1 678007 -1 0 510000
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_476
timestamp 1624635410
transform 0 -1 39593 1 0 522400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1624635410
transform 0 -1 39593 1 0 518400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_474
timestamp 1624635410
transform 0 -1 39593 1 0 514400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_473
timestamp 1624635410
transform 0 -1 39593 1 0 510400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_472
timestamp 1624635410
transform 0 -1 39593 1 0 506400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_479
timestamp 1624635410
transform 0 -1 39593 1 0 525600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_478
timestamp 1624635410
transform 0 -1 39593 1 0 525400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_477
timestamp 1624635410
transform 0 -1 39593 1 0 524400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[6\]
timestamp 1624635410
transform 0 -1 42193 1 0 525800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_482
timestamp 1624635410
transform 0 -1 39593 1 0 545800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_481
timestamp 1624635410
transform 0 -1 39593 1 0 541800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[7\]
timestamp 1624635410
transform 0 1 675407 -1 0 554200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_697
timestamp 1624635410
transform 0 1 678007 -1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_698
timestamp 1624635410
transform 0 1 678007 -1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_699
timestamp 1624635410
transform 0 1 678007 -1 0 522000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_700
timestamp 1624635410
transform 0 1 678007 -1 0 526000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_701
timestamp 1624635410
transform 0 1 678007 -1 0 530000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_702
timestamp 1624635410
transform 0 1 678007 -1 0 534000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1624635410
transform 0 1 678007 -1 0 538000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_704
timestamp 1624635410
transform 0 1 678007 -1 0 538200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1624635410
transform 0 -1 39593 1 0 561800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1624635410
transform 0 -1 39593 1 0 557800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_484
timestamp 1624635410
transform 0 -1 39593 1 0 553800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_483
timestamp 1624635410
transform 0 -1 39593 1 0 549800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_489
timestamp 1624635410
transform 0 -1 39593 1 0 568800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_488
timestamp 1624635410
transform 0 -1 39593 1 0 567800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_487
timestamp 1624635410
transform 0 -1 39593 1 0 565800
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[5\]
timestamp 1624635410
transform 0 -1 42193 1 0 569000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_492
timestamp 1624635410
transform 0 -1 39593 1 0 589000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_491
timestamp 1624635410
transform 0 -1 39593 1 0 585000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[8\]
timestamp 1624635410
transform 0 1 675407 -1 0 598400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_706
timestamp 1624635410
transform 0 1 678007 -1 0 558200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_707
timestamp 1624635410
transform 0 1 678007 -1 0 562200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_708
timestamp 1624635410
transform 0 1 678007 -1 0 566200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1624635410
transform 0 1 678007 -1 0 570200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_710
timestamp 1624635410
transform 0 1 678007 -1 0 574200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_711
timestamp 1624635410
transform 0 1 678007 -1 0 578200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1624635410
transform 0 1 678007 -1 0 582200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_713
timestamp 1624635410
transform 0 1 678007 -1 0 582400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1624635410
transform 0 -1 39593 1 0 605000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1624635410
transform 0 -1 39593 1 0 601000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_494
timestamp 1624635410
transform 0 -1 39593 1 0 597000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_493
timestamp 1624635410
transform 0 -1 39593 1 0 593000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_499
timestamp 1624635410
transform 0 -1 39593 1 0 612000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_498
timestamp 1624635410
transform 0 -1 39593 1 0 611000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_497
timestamp 1624635410
transform 0 -1 39593 1 0 609000
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[4\]
timestamp 1624635410
transform 0 -1 42193 1 0 612200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_502
timestamp 1624635410
transform 0 -1 39593 1 0 632200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_501
timestamp 1624635410
transform 0 -1 39593 1 0 628200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_717
timestamp 1624635410
transform 0 1 678007 -1 0 610400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_716
timestamp 1624635410
transform 0 1 678007 -1 0 606400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_715
timestamp 1624635410
transform 0 1 678007 -1 0 602400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_721
timestamp 1624635410
transform 0 1 678007 -1 0 626400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_720
timestamp 1624635410
transform 0 1 678007 -1 0 622400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_719
timestamp 1624635410
transform 0 1 678007 -1 0 618400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1624635410
transform 0 1 678007 -1 0 614400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_723
timestamp 1624635410
transform 0 1 678007 -1 0 626800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_722
timestamp 1624635410
transform 0 1 678007 -1 0 626600
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[9\]
timestamp 1624635410
transform 0 1 675407 -1 0 642800
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[3\]
timestamp 1624635410
transform 0 -1 42193 1 0 655400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_503
timestamp 1624635410
transform 0 -1 39593 1 0 636200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_504
timestamp 1624635410
transform 0 -1 39593 1 0 640200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1624635410
transform 0 -1 39593 1 0 644200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1624635410
transform 0 -1 39593 1 0 648200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_507
timestamp 1624635410
transform 0 -1 39593 1 0 652200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_508
timestamp 1624635410
transform 0 -1 39593 1 0 654200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_509
timestamp 1624635410
transform 0 -1 39593 1 0 655200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_511
timestamp 1624635410
transform 0 -1 39593 1 0 671400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[10\]
timestamp 1624635410
transform 0 1 675407 -1 0 687000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_725
timestamp 1624635410
transform 0 1 678007 -1 0 646800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_726
timestamp 1624635410
transform 0 1 678007 -1 0 650800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_727
timestamp 1624635410
transform 0 1 678007 -1 0 654800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1624635410
transform 0 1 678007 -1 0 658800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_729
timestamp 1624635410
transform 0 1 678007 -1 0 662800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_730
timestamp 1624635410
transform 0 1 678007 -1 0 666800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1624635410
transform 0 1 678007 -1 0 670800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_732
timestamp 1624635410
transform 0 1 678007 -1 0 671000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1624635410
transform 0 -1 39593 1 0 687400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_514
timestamp 1624635410
transform 0 -1 39593 1 0 683400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_513
timestamp 1624635410
transform 0 -1 39593 1 0 679400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_512
timestamp 1624635410
transform 0 -1 39593 1 0 675400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_520
timestamp 1624635410
transform 0 -1 39593 1 0 698600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_519
timestamp 1624635410
transform 0 -1 39593 1 0 698400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_518
timestamp 1624635410
transform 0 -1 39593 1 0 697400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_517
timestamp 1624635410
transform 0 -1 39593 1 0 695400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1624635410
transform 0 -1 39593 1 0 691400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[2\]
timestamp 1624635410
transform 0 -1 42193 1 0 698800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_522
timestamp 1624635410
transform 0 -1 39593 1 0 714800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[11\]
timestamp 1624635410
transform 0 1 675407 -1 0 731200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_734
timestamp 1624635410
transform 0 1 678007 -1 0 691000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_735
timestamp 1624635410
transform 0 1 678007 -1 0 695000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_736
timestamp 1624635410
transform 0 1 678007 -1 0 699000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1624635410
transform 0 1 678007 -1 0 703000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_738
timestamp 1624635410
transform 0 1 678007 -1 0 707000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_739
timestamp 1624635410
transform 0 1 678007 -1 0 711000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1624635410
transform 0 1 678007 -1 0 715000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_741
timestamp 1624635410
transform 0 1 678007 -1 0 715200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1624635410
transform 0 -1 39593 1 0 730800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1624635410
transform 0 -1 39593 1 0 726800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_524
timestamp 1624635410
transform 0 -1 39593 1 0 722800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_523
timestamp 1624635410
transform 0 -1 39593 1 0 718800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_530
timestamp 1624635410
transform 0 -1 39593 1 0 741800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_529
timestamp 1624635410
transform 0 -1 39593 1 0 740800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_528
timestamp 1624635410
transform 0 -1 39593 1 0 738800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_527
timestamp 1624635410
transform 0 -1 39593 1 0 734800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[1\]
timestamp 1624635410
transform 0 -1 42193 1 0 742000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_532
timestamp 1624635410
transform 0 -1 39593 1 0 758000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_743
timestamp 1624635410
transform 0 1 678007 -1 0 735200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_747
timestamp 1624635410
transform 0 1 678007 -1 0 751200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_746
timestamp 1624635410
transform 0 1 678007 -1 0 747200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_745
timestamp 1624635410
transform 0 1 678007 -1 0 743200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_744
timestamp 1624635410
transform 0 1 678007 -1 0 739200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_751
timestamp 1624635410
transform 0 1 678007 -1 0 759600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_750
timestamp 1624635410
transform 0 1 678007 -1 0 759400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_749
timestamp 1624635410
transform 0 1 678007 -1 0 759200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_748
timestamp 1624635410
transform 0 1 678007 -1 0 755200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[12\]
timestamp 1624635410
transform 0 1 675407 -1 0 775600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1624635410
transform 0 -1 39593 1 0 774000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1624635410
transform 0 -1 39593 1 0 770000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_534
timestamp 1624635410
transform 0 -1 39593 1 0 766000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_533
timestamp 1624635410
transform 0 -1 39593 1 0 762000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_540
timestamp 1624635410
transform 0 -1 39593 1 0 785000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_539
timestamp 1624635410
transform 0 -1 39593 1 0 784000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_538
timestamp 1624635410
transform 0 -1 39593 1 0 782000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_537
timestamp 1624635410
transform 0 -1 39593 1 0 778000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[0\]
timestamp 1624635410
transform 0 -1 42193 1 0 785200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_542
timestamp 1624635410
transform 0 -1 39593 1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_753
timestamp 1624635410
transform 0 1 678007 -1 0 779600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_754
timestamp 1624635410
transform 0 1 678007 -1 0 783600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_755
timestamp 1624635410
transform 0 1 678007 -1 0 787600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1624635410
transform 0 1 678007 -1 0 791600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_757
timestamp 1624635410
transform 0 1 678007 -1 0 795600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_758
timestamp 1624635410
transform 0 1 678007 -1 0 799600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1624635410
transform 0 1 678007 -1 0 803600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1624635410
transform 0 -1 39593 1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_544
timestamp 1624635410
transform 0 -1 39593 1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_543
timestamp 1624635410
transform 0 -1 39593 1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_550
timestamp 1624635410
transform 0 -1 39593 1 0 828200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_549
timestamp 1624635410
transform 0 -1 39593 1 0 827200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_548
timestamp 1624635410
transform 0 -1 39593 1 0 825200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_547
timestamp 1624635410
transform 0 -1 39593 1 0 821200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1624635410
transform 0 -1 39593 1 0 817200
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user2_vssa_hvclamp_pad
timestamp 1624635410
transform 0 -1 39593 1 0 828400
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_552
timestamp 1624635410
transform 0 -1 39593 1 0 843400
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1624635410
transform 0 1 678007 -1 0 818800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_760
timestamp 1624635410
transform 0 1 678007 -1 0 803800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_762
timestamp 1624635410
transform 0 1 678007 -1 0 822800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_763
timestamp 1624635410
transform 0 1 678007 -1 0 826800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_764
timestamp 1624635410
transform 0 1 678007 -1 0 830800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1624635410
transform 0 1 678007 -1 0 834800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_766
timestamp 1624635410
transform 0 1 678007 -1 0 838800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_767
timestamp 1624635410
transform 0 1 678007 -1 0 842800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_768
timestamp 1624635410
transform 0 1 678007 -1 0 846800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1624635410
transform 0 -1 39593 1 0 855400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_554
timestamp 1624635410
transform 0 -1 39593 1 0 851400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_553
timestamp 1624635410
transform 0 -1 39593 1 0 847400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_561
timestamp 1624635410
transform 0 -1 39593 1 0 870600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_560
timestamp 1624635410
transform 0 -1 39593 1 0 870400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_559
timestamp 1624635410
transform 0 -1 39593 1 0 869400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_558
timestamp 1624635410
transform 0 -1 39593 1 0 867400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_557
timestamp 1624635410
transform 0 -1 39593 1 0 863400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1624635410
transform 0 -1 39593 1 0 859400
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1624635410
transform 0 -1 39593 1 0 870800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_563
timestamp 1624635410
transform 0 -1 39593 1 0 885800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[13\]
timestamp 1624635410
transform 0 1 675407 -1 0 863000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_769
timestamp 1624635410
transform 0 1 678007 -1 0 847000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_771
timestamp 1624635410
transform 0 1 678007 -1 0 867000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_772
timestamp 1624635410
transform 0 1 678007 -1 0 871000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_773
timestamp 1624635410
transform 0 1 678007 -1 0 875000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_774
timestamp 1624635410
transform 0 1 678007 -1 0 879000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1624635410
transform 0 1 678007 -1 0 883000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_776
timestamp 1624635410
transform 0 1 678007 -1 0 887000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1624635410
transform 0 -1 39593 1 0 901800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1624635410
transform 0 -1 39593 1 0 897800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1624635410
transform 0 -1 39593 1 0 893800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_564
timestamp 1624635410
transform 0 -1 39593 1 0 889800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_571
timestamp 1624635410
transform 0 -1 39593 1 0 912800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_570
timestamp 1624635410
transform 0 -1 39593 1 0 911800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_569
timestamp 1624635410
transform 0 -1 39593 1 0 909800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_568
timestamp 1624635410
transform 0 -1 39593 1 0 905800
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_clamped2_pad  user2_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 -1 39593 1 0 913000
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_573
timestamp 1624635410
transform 0 -1 39593 1 0 928000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_779
timestamp 1624635410
transform 0 1 678007 -1 0 891400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_778
timestamp 1624635410
transform 0 1 678007 -1 0 891200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_777
timestamp 1624635410
transform 0 1 678007 -1 0 891000
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_clamped2_pad  user1_vccd_lvclamp_pad
timestamp 1624635410
transform 0 1 678007 -1 0 906400
box -2195 -2184 17228 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1624635410
transform 0 1 678007 -1 0 926400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1624635410
transform 0 1 678007 -1 0 922400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_783
timestamp 1624635410
transform 0 1 678007 -1 0 918400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_782
timestamp 1624635410
transform 0 1 678007 -1 0 914400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_781
timestamp 1624635410
transform 0 1 678007 -1 0 910400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_786
timestamp 1624635410
transform 0 1 678007 -1 0 930400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_576
timestamp 1624635410
transform 0 -1 39593 1 0 940000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1624635410
transform 0 -1 39593 1 0 936000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_574
timestamp 1624635410
transform 0 -1 39593 1 0 932000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_581
timestamp 1624635410
transform 0 -1 39593 1 0 955000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_580
timestamp 1624635410
transform 0 -1 39593 1 0 954000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_579
timestamp 1624635410
transform 0 -1 39593 1 0 952000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_578
timestamp 1624635410
transform 0 -1 39593 1 0 948000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_577
timestamp 1624635410
transform 0 -1 39593 1 0 944000
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[3\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 -1 40000 1 0 955200
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_583
timestamp 1624635410
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__top_power_hvc  user1_analog_pad_with_clamp $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1624635410
transform 0 1 678007 -1 0 968400
box 0 -407 33800 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_787
timestamp 1624635410
transform 0 1 678007 -1 0 934400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_788
timestamp 1624635410
transform 0 1 678007 -1 0 934600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_790
timestamp 1624635410
transform 0 1 678007 -1 0 972400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_588
timestamp 1624635410
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_587
timestamp 1624635410
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1624635410
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1624635410
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_584
timestamp 1624635410
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_592
timestamp 1624635410
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_591
timestamp 1624635410
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_590
timestamp 1624635410
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_589
timestamp 1624635410
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_5
timestamp 1624635410
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1624635410
transform 0 -1 40800 1 0 997600
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1624635410
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1624635410
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1624635410
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1624635410
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1624635410
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1624635410
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1624635410
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_14
timestamp 1624635410
transform 1 0 74800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_13
timestamp 1624635410
transform 1 0 72800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[2\]
timestamp 1624635410
transform 1 0 75000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1624635410
transform 1 0 98000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_17
timestamp 1624635410
transform 1 0 94000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_16
timestamp 1624635410
transform 1 0 90000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1624635410
transform 1 0 114000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1624635410
transform 1 0 110000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1624635410
transform 1 0 106000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1624635410
transform 1 0 102000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_24
timestamp 1624635410
transform 1 0 122000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1624635410
transform 1 0 118000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[1\]
timestamp 1624635410
transform 1 0 123000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_26
timestamp 1624635410
transform 1 0 138000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_27
timestamp 1624635410
transform 1 0 142000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_28
timestamp 1624635410
transform 1 0 146000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_29
timestamp 1624635410
transform 1 0 150000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_30
timestamp 1624635410
transform 1 0 154000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1624635410
transform 1 0 158000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1624635410
transform 1 0 162000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1624635410
transform 1 0 166000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[0\]
timestamp 1624635410
transform 1 0 171000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_5um  FILLER_34
timestamp 1624635410
transform 1 0 170000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1624635410
transform 1 0 186000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1624635410
transform 1 0 190000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_38
timestamp 1624635410
transform 1 0 194000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_39
timestamp 1624635410
transform 1 0 198000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_40
timestamp 1624635410
transform 1 0 202000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_41
timestamp 1624635410
transform 1 0 206000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_42
timestamp 1624635410
transform 1 0 210000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__top_power_hvc  user2_analog_pad_with_clamp\[1\]
timestamp 1624635410
transform 1 0 220000 0 1 998007
box 0 -407 33800 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_43
timestamp 1624635410
transform 1 0 214000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_44
timestamp 1624635410
transform 1 0 218000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__top_power_hvc  user2_analog_pad_with_clamp\[0\]
timestamp 1624635410
transform 1 0 271400 0 1 998007
box 0 -407 33800 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1624635410
transform 1 0 253800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_47
timestamp 1624635410
transform 1 0 257800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_48
timestamp 1624635410
transform 1 0 261800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1624635410
transform 1 0 265800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_50
timestamp 1624635410
transform 1 0 269800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_51
timestamp 1624635410
transform 1 0 270800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_52
timestamp 1624635410
transform 1 0 271000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_53
timestamp 1624635410
transform 1 0 271200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_55
timestamp 1624635410
transform 1 0 305200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_56
timestamp 1624635410
transform 1 0 309200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_57
timestamp 1624635410
transform 1 0 313200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_58
timestamp 1624635410
transform 1 0 317200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_59
timestamp 1624635410
transform 1 0 321200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1624635410
transform 1 0 325200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1624635410
transform 1 0 329200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1624635410
transform 1 0 333200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_63
timestamp 1624635410
transform 1 0 337200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[1\]
timestamp 1624635410
transform 1 0 339400 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_64
timestamp 1624635410
transform 1 0 339200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_66
timestamp 1624635410
transform 1 0 354400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_67
timestamp 1624635410
transform 1 0 358400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_68
timestamp 1624635410
transform 1 0 362400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_69
timestamp 1624635410
transform 1 0 366400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_70
timestamp 1624635410
transform 1 0 370400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1624635410
transform 1 0 374400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1624635410
transform 1 0 378400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1624635410
transform 1 0 382400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_74
timestamp 1624635410
transform 1 0 386400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1624635410
transform 1 0 390600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_0
timestamp 1624635410
transform 1 0 389600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0
timestamp 1624635410
transform 1 0 388600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_75
timestamp 1624635410
transform 1 0 388400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_79
timestamp 1624635410
transform 1 0 394600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_80
timestamp 1624635410
transform 1 0 398600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_81
timestamp 1624635410
transform 1 0 402600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_82
timestamp 1624635410
transform 1 0 406600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_83
timestamp 1624635410
transform 1 0 410600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_84
timestamp 1624635410
transform 1 0 414600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_85
timestamp 1624635410
transform 1 0 418600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_87
timestamp 1624635410
transform 1 0 424600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_86
timestamp 1624635410
transform 1 0 422600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[3\]
timestamp 1624635410
transform 1 0 424800 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_92
timestamp 1624635410
transform 1 0 451800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1624635410
transform 1 0 447800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1624635410
transform 1 0 443800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1624635410
transform 1 0 439800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_95
timestamp 1624635410
transform 1 0 463800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_94
timestamp 1624635410
transform 1 0 459800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_93
timestamp 1624635410
transform 1 0 455800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_99
timestamp 1624635410
transform 1 0 474000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_98
timestamp 1624635410
transform 1 0 473800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_97
timestamp 1624635410
transform 1 0 471800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_96
timestamp 1624635410
transform 1 0 467800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[2\]
timestamp 1624635410
transform 1 0 474200 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1624635410
transform 1 0 493200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1624635410
transform 1 0 489200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_105
timestamp 1624635410
transform 1 0 505200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1624635410
transform 1 0 501200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1624635410
transform 1 0 497200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_109
timestamp 1624635410
transform 1 0 521200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_108
timestamp 1624635410
transform 1 0 517200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_107
timestamp 1624635410
transform 1 0 513200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_106
timestamp 1624635410
transform 1 0 509200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_112
timestamp 1624635410
transform 1 0 525600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_111
timestamp 1624635410
transform 1 0 525400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_110
timestamp 1624635410
transform 1 0 525200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[1\]
timestamp 1624635410
transform 1 0 525800 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1624635410
transform 1 0 544800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1624635410
transform 1 0 540800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_119
timestamp 1624635410
transform 1 0 560800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_118
timestamp 1624635410
transform 1 0 556800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_117
timestamp 1624635410
transform 1 0 552800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_116
timestamp 1624635410
transform 1 0 548800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_126
timestamp 1624635410
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_125
timestamp 1624635410
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_124
timestamp 1624635410
transform 1 0 575000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_123
timestamp 1624635410
transform 1 0 574800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_122
timestamp 1624635410
transform 1 0 572800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_121
timestamp 1624635410
transform 1 0 568800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_120
timestamp 1624635410
transform 1 0 564800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1624635410
transform 1 0 575600 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_128
timestamp 1624635410
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1624635410
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_130
timestamp 1624635410
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_129
timestamp 1624635410
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_135
timestamp 1624635410
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_134
timestamp 1624635410
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_133
timestamp 1624635410
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_132
timestamp 1624635410
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_138
timestamp 1624635410
transform 1 0 626800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_137
timestamp 1624635410
transform 1 0 626600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_136
timestamp 1624635410
transform 1 0 622600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[0\]
timestamp 1624635410
transform 1 0 627000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_140
timestamp 1624635410
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_141
timestamp 1624635410
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_142
timestamp 1624635410
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_143
timestamp 1624635410
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_144
timestamp 1624635410
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_145
timestamp 1624635410
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_146
timestamp 1624635410
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_147
timestamp 1624635410
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_148
timestamp 1624635410
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_795
timestamp 1624635410
transform 0 1 678007 -1 0 992400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_794
timestamp 1624635410
transform 0 1 678007 -1 0 988400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_793
timestamp 1624635410
transform 0 1 678007 -1 0 984400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_792
timestamp 1624635410
transform 0 1 678007 -1 0 980400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_791
timestamp 1624635410
transform 0 1 678007 -1 0 976400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_798
timestamp 1624635410
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_797
timestamp 1624635410
transform 0 1 678007 -1 0 996600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_796
timestamp 1624635410
transform 0 1 678007 -1 0 996400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_152
timestamp 1624635410
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_151
timestamp 1624635410
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_150
timestamp 1624635410
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_149
timestamp 1624635410
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__corner_pad  user1_corner
timestamp 1624635410
transform 1 0 677600 0 1 996800
box 0 0 40000 40800
<< labels >>
rlabel metal5 s 187640 6598 200180 19088 6 clock
port 0 nsew signal input
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 1 nsew signal tristate
rlabel metal2 s 194043 41713 194099 42193 6 por
port 2 nsew signal input
rlabel metal5 s 351040 6598 363580 19088 6 flash_clk
port 3 nsew signal tristate
rlabel metal2 s 361767 41713 361823 42193 6 flash_clk_core
port 4 nsew signal input
rlabel metal2 s 357443 41713 357499 42193 6 flash_clk_ieb_core
port 5 nsew signal input
rlabel metal2 s 364895 41713 364951 42193 6 flash_clk_oeb_core
port 6 nsew signal input
rlabel metal5 s 296240 6598 308780 19088 6 flash_csb
port 7 nsew signal tristate
rlabel metal2 s 306967 41713 307023 42193 6 flash_csb_core
port 8 nsew signal input
rlabel metal2 s 302643 41713 302699 42193 6 flash_csb_ieb_core
port 9 nsew signal input
rlabel metal2 s 310095 41713 310151 42193 6 flash_csb_oeb_core
port 10 nsew signal input
rlabel metal5 s 405840 6598 418380 19088 6 flash_io0
port 11 nsew signal bidirectional
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 12 nsew signal tristate
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 13 nsew signal input
rlabel metal2 s 412243 41713 412299 42193 6 flash_io0_ieb_core
port 14 nsew signal input
rlabel metal2 s 419695 41713 419751 42193 6 flash_io0_oeb_core
port 15 nsew signal input
rlabel metal5 s 460640 6598 473180 19088 6 flash_io1
port 16 nsew signal bidirectional
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 17 nsew signal tristate
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 18 nsew signal input
rlabel metal2 s 467043 41713 467099 42193 6 flash_io1_ieb_core
port 19 nsew signal input
rlabel metal2 s 474495 41713 474551 42193 6 flash_io1_oeb_core
port 20 nsew signal input
rlabel metal5 s 515440 6598 527980 19088 6 gpio
port 21 nsew signal bidirectional
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 22 nsew signal tristate
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 23 nsew signal input
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 24 nsew signal input
rlabel metal2 s 524971 41713 525027 42193 6 gpio_mode1_core
port 25 nsew signal input
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 26 nsew signal input
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 27 nsew signal input
rlabel metal5 s 6167 70054 19619 80934 6 vccd_pad
port 28 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18975 6 vdda_pad
port 29 nsew signal bidirectional
rlabel metal5 s 6811 111610 18975 123778 6 vddio_pad
port 30 nsew signal bidirectional
rlabel metal5 s 6811 872210 18975 884378 6 vddio_pad2
port 31 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18975 6 vssa_pad
port 32 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19619 6 vssd_pad
port 33 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18975 6 vssio_pad
port 34 nsew signal bidirectional
rlabel metal5 s 340810 1018624 352978 1030788 6 vssio_pad2
port 35 nsew signal bidirectional
rlabel metal5 s 698512 99640 711002 112180 6 mprj_io[0]
port 36 nsew signal bidirectional
rlabel metal2 s 675407 104203 675887 104259 6 mprj_io_analog_en[0]
port 37 nsew signal input
rlabel metal2 s 675407 105491 675887 105547 6 mprj_io_analog_pol[0]
port 38 nsew signal input
rlabel metal2 s 675407 108527 675887 108583 6 mprj_io_analog_sel[0]
port 39 nsew signal input
rlabel metal2 s 675407 104847 675887 104903 6 mprj_io_dm[0]
port 40 nsew signal input
rlabel metal2 s 675407 103007 675887 103063 6 mprj_io_dm[1]
port 41 nsew signal input
rlabel metal2 s 675407 109171 675887 109227 6 mprj_io_dm[2]
port 42 nsew signal input
rlabel metal2 s 675407 109815 675887 109871 6 mprj_io_holdover[0]
port 43 nsew signal input
rlabel metal2 s 675407 112851 675887 112907 6 mprj_io_ib_mode_sel[0]
port 44 nsew signal input
rlabel metal2 s 675407 106043 675887 106099 6 mprj_io_inp_dis[0]
port 45 nsew signal input
rlabel metal2 s 675407 113495 675887 113551 6 mprj_io_oeb[0]
port 46 nsew signal input
rlabel metal2 s 675407 110367 675887 110423 6 mprj_io_out[0]
port 47 nsew signal input
rlabel metal2 s 675407 101167 675887 101223 6 mprj_io_slow_sel[0]
port 48 nsew signal input
rlabel metal2 s 675407 112207 675887 112263 6 mprj_io_vtrip_sel[0]
port 49 nsew signal input
rlabel metal2 s 675407 99327 675887 99383 6 mprj_io_in[0]
port 50 nsew signal tristate
rlabel metal2 s 675407 114047 675887 114103 6 mprj_io_in_3v3[0]
port 51 nsew signal tristate
rlabel metal2 s 675407 674411 675887 674467 6 mprj_gpio_analog[3]
port 52 nsew signal bidirectional
rlabel metal2 s 675407 676251 675887 676307 6 mprj_gpio_noesd[3]
port 53 nsew signal bidirectional
rlabel metal5 s 698512 672240 711002 684780 6 mprj_io[10]
port 54 nsew signal bidirectional
rlabel metal2 s 675407 676803 675887 676859 6 mprj_io_analog_en[10]
port 55 nsew signal input
rlabel metal2 s 675407 678091 675887 678147 6 mprj_io_analog_pol[10]
port 56 nsew signal input
rlabel metal2 s 675407 681127 675887 681183 6 mprj_io_analog_sel[10]
port 57 nsew signal input
rlabel metal2 s 675407 677447 675887 677503 6 mprj_io_dm[30]
port 58 nsew signal input
rlabel metal2 s 675407 675607 675887 675663 6 mprj_io_dm[31]
port 59 nsew signal input
rlabel metal2 s 675407 681771 675887 681827 6 mprj_io_dm[32]
port 60 nsew signal input
rlabel metal2 s 675407 682415 675887 682471 6 mprj_io_holdover[10]
port 61 nsew signal input
rlabel metal2 s 675407 685451 675887 685507 6 mprj_io_ib_mode_sel[10]
port 62 nsew signal input
rlabel metal2 s 675407 678643 675887 678699 6 mprj_io_inp_dis[10]
port 63 nsew signal input
rlabel metal2 s 675407 686095 675887 686151 6 mprj_io_oeb[10]
port 64 nsew signal input
rlabel metal2 s 675407 682967 675887 683023 6 mprj_io_out[10]
port 65 nsew signal input
rlabel metal2 s 675407 673767 675887 673823 6 mprj_io_slow_sel[10]
port 66 nsew signal input
rlabel metal2 s 675407 684807 675887 684863 6 mprj_io_vtrip_sel[10]
port 67 nsew signal input
rlabel metal2 s 675407 671927 675887 671983 6 mprj_io_in[10]
port 68 nsew signal tristate
rlabel metal2 s 675407 686647 675887 686703 6 mprj_io_in_3v3[10]
port 69 nsew signal tristate
rlabel metal2 s 675407 718611 675887 718667 6 mprj_gpio_analog[4]
port 70 nsew signal bidirectional
rlabel metal2 s 675407 720451 675887 720507 6 mprj_gpio_noesd[4]
port 71 nsew signal bidirectional
rlabel metal5 s 698512 716440 711002 728980 6 mprj_io[11]
port 72 nsew signal bidirectional
rlabel metal2 s 675407 721003 675887 721059 6 mprj_io_analog_en[11]
port 73 nsew signal input
rlabel metal2 s 675407 722291 675887 722347 6 mprj_io_analog_pol[11]
port 74 nsew signal input
rlabel metal2 s 675407 725327 675887 725383 6 mprj_io_analog_sel[11]
port 75 nsew signal input
rlabel metal2 s 675407 721647 675887 721703 6 mprj_io_dm[33]
port 76 nsew signal input
rlabel metal2 s 675407 719807 675887 719863 6 mprj_io_dm[34]
port 77 nsew signal input
rlabel metal2 s 675407 725971 675887 726027 6 mprj_io_dm[35]
port 78 nsew signal input
rlabel metal2 s 675407 726615 675887 726671 6 mprj_io_holdover[11]
port 79 nsew signal input
rlabel metal2 s 675407 729651 675887 729707 6 mprj_io_ib_mode_sel[11]
port 80 nsew signal input
rlabel metal2 s 675407 722843 675887 722899 6 mprj_io_inp_dis[11]
port 81 nsew signal input
rlabel metal2 s 675407 730295 675887 730351 6 mprj_io_oeb[11]
port 82 nsew signal input
rlabel metal2 s 675407 727167 675887 727223 6 mprj_io_out[11]
port 83 nsew signal input
rlabel metal2 s 675407 717967 675887 718023 6 mprj_io_slow_sel[11]
port 84 nsew signal input
rlabel metal2 s 675407 729007 675887 729063 6 mprj_io_vtrip_sel[11]
port 85 nsew signal input
rlabel metal2 s 675407 716127 675887 716183 6 mprj_io_in[11]
port 86 nsew signal tristate
rlabel metal2 s 675407 730847 675887 730903 6 mprj_io_in_3v3[11]
port 87 nsew signal tristate
rlabel metal2 s 675407 763011 675887 763067 6 mprj_gpio_analog[5]
port 88 nsew signal bidirectional
rlabel metal2 s 675407 764851 675887 764907 6 mprj_gpio_noesd[5]
port 89 nsew signal bidirectional
rlabel metal5 s 698512 760840 711002 773380 6 mprj_io[12]
port 90 nsew signal bidirectional
rlabel metal2 s 675407 765403 675887 765459 6 mprj_io_analog_en[12]
port 91 nsew signal input
rlabel metal2 s 675407 766691 675887 766747 6 mprj_io_analog_pol[12]
port 92 nsew signal input
rlabel metal2 s 675407 769727 675887 769783 6 mprj_io_analog_sel[12]
port 93 nsew signal input
rlabel metal2 s 675407 766047 675887 766103 6 mprj_io_dm[36]
port 94 nsew signal input
rlabel metal2 s 675407 764207 675887 764263 6 mprj_io_dm[37]
port 95 nsew signal input
rlabel metal2 s 675407 770371 675887 770427 6 mprj_io_dm[38]
port 96 nsew signal input
rlabel metal2 s 675407 771015 675887 771071 6 mprj_io_holdover[12]
port 97 nsew signal input
rlabel metal2 s 675407 774051 675887 774107 6 mprj_io_ib_mode_sel[12]
port 98 nsew signal input
rlabel metal2 s 675407 767243 675887 767299 6 mprj_io_inp_dis[12]
port 99 nsew signal input
rlabel metal2 s 675407 774695 675887 774751 6 mprj_io_oeb[12]
port 100 nsew signal input
rlabel metal2 s 675407 771567 675887 771623 6 mprj_io_out[12]
port 101 nsew signal input
rlabel metal2 s 675407 762367 675887 762423 6 mprj_io_slow_sel[12]
port 102 nsew signal input
rlabel metal2 s 675407 773407 675887 773463 6 mprj_io_vtrip_sel[12]
port 103 nsew signal input
rlabel metal2 s 675407 760527 675887 760583 6 mprj_io_in[12]
port 104 nsew signal tristate
rlabel metal2 s 675407 775247 675887 775303 6 mprj_io_in_3v3[12]
port 105 nsew signal tristate
rlabel metal2 s 675407 850411 675887 850467 6 mprj_gpio_analog[6]
port 106 nsew signal bidirectional
rlabel metal2 s 675407 852251 675887 852307 6 mprj_gpio_noesd[6]
port 107 nsew signal bidirectional
rlabel metal5 s 698512 848240 711002 860780 6 mprj_io[13]
port 108 nsew signal bidirectional
rlabel metal2 s 675407 852803 675887 852859 6 mprj_io_analog_en[13]
port 109 nsew signal input
rlabel metal2 s 675407 854091 675887 854147 6 mprj_io_analog_pol[13]
port 110 nsew signal input
rlabel metal2 s 675407 857127 675887 857183 6 mprj_io_analog_sel[13]
port 111 nsew signal input
rlabel metal2 s 675407 853447 675887 853503 6 mprj_io_dm[39]
port 112 nsew signal input
rlabel metal2 s 675407 851607 675887 851663 6 mprj_io_dm[40]
port 113 nsew signal input
rlabel metal2 s 675407 857771 675887 857827 6 mprj_io_dm[41]
port 114 nsew signal input
rlabel metal2 s 675407 858415 675887 858471 6 mprj_io_holdover[13]
port 115 nsew signal input
rlabel metal2 s 675407 861451 675887 861507 6 mprj_io_ib_mode_sel[13]
port 116 nsew signal input
rlabel metal2 s 675407 854643 675887 854699 6 mprj_io_inp_dis[13]
port 117 nsew signal input
rlabel metal2 s 675407 862095 675887 862151 6 mprj_io_oeb[13]
port 118 nsew signal input
rlabel metal2 s 675407 858967 675887 859023 6 mprj_io_out[13]
port 119 nsew signal input
rlabel metal2 s 675407 849767 675887 849823 6 mprj_io_slow_sel[13]
port 120 nsew signal input
rlabel metal2 s 675407 860807 675887 860863 6 mprj_io_vtrip_sel[13]
port 121 nsew signal input
rlabel metal2 s 675407 847927 675887 847983 6 mprj_io_in[13]
port 122 nsew signal tristate
rlabel metal2 s 675407 862647 675887 862703 6 mprj_io_in_3v3[13]
port 123 nsew signal tristate
rlabel metal5 s 698512 144040 711002 156580 6 mprj_io[1]
port 124 nsew signal bidirectional
rlabel metal2 s 675407 148603 675887 148659 6 mprj_io_analog_en[1]
port 125 nsew signal input
rlabel metal2 s 675407 149891 675887 149947 6 mprj_io_analog_pol[1]
port 126 nsew signal input
rlabel metal2 s 675407 152927 675887 152983 6 mprj_io_analog_sel[1]
port 127 nsew signal input
rlabel metal2 s 675407 149247 675887 149303 6 mprj_io_dm[3]
port 128 nsew signal input
rlabel metal2 s 675407 147407 675887 147463 6 mprj_io_dm[4]
port 129 nsew signal input
rlabel metal2 s 675407 153571 675887 153627 6 mprj_io_dm[5]
port 130 nsew signal input
rlabel metal2 s 675407 154215 675887 154271 6 mprj_io_holdover[1]
port 131 nsew signal input
rlabel metal2 s 675407 157251 675887 157307 6 mprj_io_ib_mode_sel[1]
port 132 nsew signal input
rlabel metal2 s 675407 150443 675887 150499 6 mprj_io_inp_dis[1]
port 133 nsew signal input
rlabel metal2 s 675407 157895 675887 157951 6 mprj_io_oeb[1]
port 134 nsew signal input
rlabel metal2 s 675407 154767 675887 154823 6 mprj_io_out[1]
port 135 nsew signal input
rlabel metal2 s 675407 145567 675887 145623 6 mprj_io_slow_sel[1]
port 136 nsew signal input
rlabel metal2 s 675407 156607 675887 156663 6 mprj_io_vtrip_sel[1]
port 137 nsew signal input
rlabel metal2 s 675407 143727 675887 143783 6 mprj_io_in[1]
port 138 nsew signal tristate
rlabel metal2 s 675407 158447 675887 158503 6 mprj_io_in_3v3[1]
port 139 nsew signal tristate
rlabel metal5 s 698512 188240 711002 200780 6 mprj_io[2]
port 140 nsew signal bidirectional
rlabel metal2 s 675407 192803 675887 192859 6 mprj_io_analog_en[2]
port 141 nsew signal input
rlabel metal2 s 675407 194091 675887 194147 6 mprj_io_analog_pol[2]
port 142 nsew signal input
rlabel metal2 s 675407 197127 675887 197183 6 mprj_io_analog_sel[2]
port 143 nsew signal input
rlabel metal2 s 675407 193447 675887 193503 6 mprj_io_dm[6]
port 144 nsew signal input
rlabel metal2 s 675407 191607 675887 191663 6 mprj_io_dm[7]
port 145 nsew signal input
rlabel metal2 s 675407 197771 675887 197827 6 mprj_io_dm[8]
port 146 nsew signal input
rlabel metal2 s 675407 198415 675887 198471 6 mprj_io_holdover[2]
port 147 nsew signal input
rlabel metal2 s 675407 201451 675887 201507 6 mprj_io_ib_mode_sel[2]
port 148 nsew signal input
rlabel metal2 s 675407 194643 675887 194699 6 mprj_io_inp_dis[2]
port 149 nsew signal input
rlabel metal2 s 675407 202095 675887 202151 6 mprj_io_oeb[2]
port 150 nsew signal input
rlabel metal2 s 675407 198967 675887 199023 6 mprj_io_out[2]
port 151 nsew signal input
rlabel metal2 s 675407 189767 675887 189823 6 mprj_io_slow_sel[2]
port 152 nsew signal input
rlabel metal2 s 675407 200807 675887 200863 6 mprj_io_vtrip_sel[2]
port 153 nsew signal input
rlabel metal2 s 675407 187927 675887 187983 6 mprj_io_in[2]
port 154 nsew signal tristate
rlabel metal2 s 675407 202647 675887 202703 6 mprj_io_in_3v3[2]
port 155 nsew signal tristate
rlabel metal5 s 698512 232440 711002 244980 6 mprj_io[3]
port 156 nsew signal bidirectional
rlabel metal2 s 675407 237003 675887 237059 6 mprj_io_analog_en[3]
port 157 nsew signal input
rlabel metal2 s 675407 238291 675887 238347 6 mprj_io_analog_pol[3]
port 158 nsew signal input
rlabel metal2 s 675407 241327 675887 241383 6 mprj_io_analog_sel[3]
port 159 nsew signal input
rlabel metal2 s 675407 235807 675887 235863 6 mprj_io_dm[10]
port 160 nsew signal input
rlabel metal2 s 675407 241971 675887 242027 6 mprj_io_dm[11]
port 161 nsew signal input
rlabel metal2 s 675407 237647 675887 237703 6 mprj_io_dm[9]
port 162 nsew signal input
rlabel metal2 s 675407 242615 675887 242671 6 mprj_io_holdover[3]
port 163 nsew signal input
rlabel metal2 s 675407 245651 675887 245707 6 mprj_io_ib_mode_sel[3]
port 164 nsew signal input
rlabel metal2 s 675407 238843 675887 238899 6 mprj_io_inp_dis[3]
port 165 nsew signal input
rlabel metal2 s 675407 246295 675887 246351 6 mprj_io_oeb[3]
port 166 nsew signal input
rlabel metal2 s 675407 243167 675887 243223 6 mprj_io_out[3]
port 167 nsew signal input
rlabel metal2 s 675407 233967 675887 234023 6 mprj_io_slow_sel[3]
port 168 nsew signal input
rlabel metal2 s 675407 245007 675887 245063 6 mprj_io_vtrip_sel[3]
port 169 nsew signal input
rlabel metal2 s 675407 232127 675887 232183 6 mprj_io_in[3]
port 170 nsew signal tristate
rlabel metal2 s 675407 246847 675887 246903 6 mprj_io_in_3v3[3]
port 171 nsew signal tristate
rlabel metal5 s 698512 276840 711002 289380 6 mprj_io[4]
port 172 nsew signal bidirectional
rlabel metal2 s 675407 281403 675887 281459 6 mprj_io_analog_en[4]
port 173 nsew signal input
rlabel metal2 s 675407 282691 675887 282747 6 mprj_io_analog_pol[4]
port 174 nsew signal input
rlabel metal2 s 675407 285727 675887 285783 6 mprj_io_analog_sel[4]
port 175 nsew signal input
rlabel metal2 s 675407 282047 675887 282103 6 mprj_io_dm[12]
port 176 nsew signal input
rlabel metal2 s 675407 280207 675887 280263 6 mprj_io_dm[13]
port 177 nsew signal input
rlabel metal2 s 675407 286371 675887 286427 6 mprj_io_dm[14]
port 178 nsew signal input
rlabel metal2 s 675407 287015 675887 287071 6 mprj_io_holdover[4]
port 179 nsew signal input
rlabel metal2 s 675407 290051 675887 290107 6 mprj_io_ib_mode_sel[4]
port 180 nsew signal input
rlabel metal2 s 675407 283243 675887 283299 6 mprj_io_inp_dis[4]
port 181 nsew signal input
rlabel metal2 s 675407 290695 675887 290751 6 mprj_io_oeb[4]
port 182 nsew signal input
rlabel metal2 s 675407 287567 675887 287623 6 mprj_io_out[4]
port 183 nsew signal input
rlabel metal2 s 675407 278367 675887 278423 6 mprj_io_slow_sel[4]
port 184 nsew signal input
rlabel metal2 s 675407 289407 675887 289463 6 mprj_io_vtrip_sel[4]
port 185 nsew signal input
rlabel metal2 s 675407 276527 675887 276583 6 mprj_io_in[4]
port 186 nsew signal tristate
rlabel metal2 s 675407 291247 675887 291303 6 mprj_io_in_3v3[4]
port 187 nsew signal tristate
rlabel metal5 s 698512 321040 711002 333580 6 mprj_io[5]
port 188 nsew signal bidirectional
rlabel metal2 s 675407 325603 675887 325659 6 mprj_io_analog_en[5]
port 189 nsew signal input
rlabel metal2 s 675407 326891 675887 326947 6 mprj_io_analog_pol[5]
port 190 nsew signal input
rlabel metal2 s 675407 329927 675887 329983 6 mprj_io_analog_sel[5]
port 191 nsew signal input
rlabel metal2 s 675407 326247 675887 326303 6 mprj_io_dm[15]
port 192 nsew signal input
rlabel metal2 s 675407 324407 675887 324463 6 mprj_io_dm[16]
port 193 nsew signal input
rlabel metal2 s 675407 330571 675887 330627 6 mprj_io_dm[17]
port 194 nsew signal input
rlabel metal2 s 675407 331215 675887 331271 6 mprj_io_holdover[5]
port 195 nsew signal input
rlabel metal2 s 675407 334251 675887 334307 6 mprj_io_ib_mode_sel[5]
port 196 nsew signal input
rlabel metal2 s 675407 327443 675887 327499 6 mprj_io_inp_dis[5]
port 197 nsew signal input
rlabel metal2 s 675407 334895 675887 334951 6 mprj_io_oeb[5]
port 198 nsew signal input
rlabel metal2 s 675407 331767 675887 331823 6 mprj_io_out[5]
port 199 nsew signal input
rlabel metal2 s 675407 322567 675887 322623 6 mprj_io_slow_sel[5]
port 200 nsew signal input
rlabel metal2 s 675407 333607 675887 333663 6 mprj_io_vtrip_sel[5]
port 201 nsew signal input
rlabel metal2 s 675407 320727 675887 320783 6 mprj_io_in[5]
port 202 nsew signal tristate
rlabel metal2 s 675407 335447 675887 335503 6 mprj_io_in_3v3[5]
port 203 nsew signal tristate
rlabel metal5 s 698512 365240 711002 377780 6 mprj_io[6]
port 204 nsew signal bidirectional
rlabel metal2 s 675407 369803 675887 369859 6 mprj_io_analog_en[6]
port 205 nsew signal input
rlabel metal2 s 675407 371091 675887 371147 6 mprj_io_analog_pol[6]
port 206 nsew signal input
rlabel metal2 s 675407 374127 675887 374183 6 mprj_io_analog_sel[6]
port 207 nsew signal input
rlabel metal2 s 675407 370447 675887 370503 6 mprj_io_dm[18]
port 208 nsew signal input
rlabel metal2 s 675407 368607 675887 368663 6 mprj_io_dm[19]
port 209 nsew signal input
rlabel metal2 s 675407 374771 675887 374827 6 mprj_io_dm[20]
port 210 nsew signal input
rlabel metal2 s 675407 375415 675887 375471 6 mprj_io_holdover[6]
port 211 nsew signal input
rlabel metal2 s 675407 378451 675887 378507 6 mprj_io_ib_mode_sel[6]
port 212 nsew signal input
rlabel metal2 s 675407 371643 675887 371699 6 mprj_io_inp_dis[6]
port 213 nsew signal input
rlabel metal2 s 675407 379095 675887 379151 6 mprj_io_oeb[6]
port 214 nsew signal input
rlabel metal2 s 675407 375967 675887 376023 6 mprj_io_out[6]
port 215 nsew signal input
rlabel metal2 s 675407 366767 675887 366823 6 mprj_io_slow_sel[6]
port 216 nsew signal input
rlabel metal2 s 675407 377807 675887 377863 6 mprj_io_vtrip_sel[6]
port 217 nsew signal input
rlabel metal2 s 675407 364927 675887 364983 6 mprj_io_in[6]
port 218 nsew signal tristate
rlabel metal2 s 675407 379647 675887 379703 6 mprj_io_in_3v3[6]
port 219 nsew signal tristate
rlabel metal2 s 675407 541611 675887 541667 6 mprj_gpio_analog[0]
port 220 nsew signal bidirectional
rlabel metal2 s 675407 543451 675887 543507 6 mprj_gpio_noesd[0]
port 221 nsew signal bidirectional
rlabel metal5 s 698512 539440 711002 551980 6 mprj_io[7]
port 222 nsew signal bidirectional
rlabel metal2 s 675407 544003 675887 544059 6 mprj_io_analog_en[7]
port 223 nsew signal input
rlabel metal2 s 675407 545291 675887 545347 6 mprj_io_analog_pol[7]
port 224 nsew signal input
rlabel metal2 s 675407 548327 675887 548383 6 mprj_io_analog_sel[7]
port 225 nsew signal input
rlabel metal2 s 675407 544647 675887 544703 6 mprj_io_dm[21]
port 226 nsew signal input
rlabel metal2 s 675407 542807 675887 542863 6 mprj_io_dm[22]
port 227 nsew signal input
rlabel metal2 s 675407 548971 675887 549027 6 mprj_io_dm[23]
port 228 nsew signal input
rlabel metal2 s 675407 549615 675887 549671 6 mprj_io_holdover[7]
port 229 nsew signal input
rlabel metal2 s 675407 552651 675887 552707 6 mprj_io_ib_mode_sel[7]
port 230 nsew signal input
rlabel metal2 s 675407 545843 675887 545899 6 mprj_io_inp_dis[7]
port 231 nsew signal input
rlabel metal2 s 675407 553295 675887 553351 6 mprj_io_oeb[7]
port 232 nsew signal input
rlabel metal2 s 675407 550167 675887 550223 6 mprj_io_out[7]
port 233 nsew signal input
rlabel metal2 s 675407 540967 675887 541023 6 mprj_io_slow_sel[7]
port 234 nsew signal input
rlabel metal2 s 675407 552007 675887 552063 6 mprj_io_vtrip_sel[7]
port 235 nsew signal input
rlabel metal2 s 675407 539127 675887 539183 6 mprj_io_in[7]
port 236 nsew signal tristate
rlabel metal2 s 675407 553847 675887 553903 6 mprj_io_in_3v3[7]
port 237 nsew signal tristate
rlabel metal2 s 675407 585811 675887 585867 6 mprj_gpio_analog[1]
port 238 nsew signal bidirectional
rlabel metal2 s 675407 587651 675887 587707 6 mprj_gpio_noesd[1]
port 239 nsew signal bidirectional
rlabel metal5 s 698512 583640 711002 596180 6 mprj_io[8]
port 240 nsew signal bidirectional
rlabel metal2 s 675407 588203 675887 588259 6 mprj_io_analog_en[8]
port 241 nsew signal input
rlabel metal2 s 675407 589491 675887 589547 6 mprj_io_analog_pol[8]
port 242 nsew signal input
rlabel metal2 s 675407 592527 675887 592583 6 mprj_io_analog_sel[8]
port 243 nsew signal input
rlabel metal2 s 675407 588847 675887 588903 6 mprj_io_dm[24]
port 244 nsew signal input
rlabel metal2 s 675407 587007 675887 587063 6 mprj_io_dm[25]
port 245 nsew signal input
rlabel metal2 s 675407 593171 675887 593227 6 mprj_io_dm[26]
port 246 nsew signal input
rlabel metal2 s 675407 593815 675887 593871 6 mprj_io_holdover[8]
port 247 nsew signal input
rlabel metal2 s 675407 596851 675887 596907 6 mprj_io_ib_mode_sel[8]
port 248 nsew signal input
rlabel metal2 s 675407 590043 675887 590099 6 mprj_io_inp_dis[8]
port 249 nsew signal input
rlabel metal2 s 675407 597495 675887 597551 6 mprj_io_oeb[8]
port 250 nsew signal input
rlabel metal2 s 675407 594367 675887 594423 6 mprj_io_out[8]
port 251 nsew signal input
rlabel metal2 s 675407 585167 675887 585223 6 mprj_io_slow_sel[8]
port 252 nsew signal input
rlabel metal2 s 675407 596207 675887 596263 6 mprj_io_vtrip_sel[8]
port 253 nsew signal input
rlabel metal2 s 675407 583327 675887 583383 6 mprj_io_in[8]
port 254 nsew signal tristate
rlabel metal2 s 675407 598047 675887 598103 6 mprj_io_in_3v3[8]
port 255 nsew signal tristate
rlabel metal2 s 675407 630211 675887 630267 6 mprj_gpio_analog[2]
port 256 nsew signal bidirectional
rlabel metal2 s 675407 632051 675887 632107 6 mprj_gpio_noesd[2]
port 257 nsew signal bidirectional
rlabel metal5 s 698512 628040 711002 640580 6 mprj_io[9]
port 258 nsew signal bidirectional
rlabel metal2 s 675407 632603 675887 632659 6 mprj_io_analog_en[9]
port 259 nsew signal input
rlabel metal2 s 675407 633891 675887 633947 6 mprj_io_analog_pol[9]
port 260 nsew signal input
rlabel metal2 s 675407 636927 675887 636983 6 mprj_io_analog_sel[9]
port 261 nsew signal input
rlabel metal2 s 675407 633247 675887 633303 6 mprj_io_dm[27]
port 262 nsew signal input
rlabel metal2 s 675407 631407 675887 631463 6 mprj_io_dm[28]
port 263 nsew signal input
rlabel metal2 s 675407 637571 675887 637627 6 mprj_io_dm[29]
port 264 nsew signal input
rlabel metal2 s 675407 638215 675887 638271 6 mprj_io_holdover[9]
port 265 nsew signal input
rlabel metal2 s 675407 641251 675887 641307 6 mprj_io_ib_mode_sel[9]
port 266 nsew signal input
rlabel metal2 s 675407 634443 675887 634499 6 mprj_io_inp_dis[9]
port 267 nsew signal input
rlabel metal2 s 675407 641895 675887 641951 6 mprj_io_oeb[9]
port 268 nsew signal input
rlabel metal2 s 675407 638767 675887 638823 6 mprj_io_out[9]
port 269 nsew signal input
rlabel metal2 s 675407 629567 675887 629623 6 mprj_io_slow_sel[9]
port 270 nsew signal input
rlabel metal2 s 675407 640607 675887 640663 6 mprj_io_vtrip_sel[9]
port 271 nsew signal input
rlabel metal2 s 675407 627727 675887 627783 6 mprj_io_in[9]
port 272 nsew signal tristate
rlabel metal2 s 675407 642447 675887 642503 6 mprj_io_in_3v3[9]
port 273 nsew signal tristate
rlabel metal2 s 41713 797733 42193 797789 6 mprj_gpio_analog[7]
port 274 nsew signal bidirectional
rlabel metal2 s 41713 795893 42193 795949 6 mprj_gpio_noesd[7]
port 275 nsew signal bidirectional
rlabel metal5 s 6598 787420 19088 799960 6 mprj_io[25]
port 276 nsew signal bidirectional
rlabel metal2 s 41713 795341 42193 795397 6 mprj_io_analog_en[14]
port 277 nsew signal input
rlabel metal2 s 41713 794053 42193 794109 6 mprj_io_analog_pol[14]
port 278 nsew signal input
rlabel metal2 s 41713 791017 42193 791073 6 mprj_io_analog_sel[14]
port 279 nsew signal input
rlabel metal2 s 41713 794697 42193 794753 6 mprj_io_dm[42]
port 280 nsew signal input
rlabel metal2 s 41713 796537 42193 796593 6 mprj_io_dm[43]
port 281 nsew signal input
rlabel metal2 s 41713 790373 42193 790429 6 mprj_io_dm[44]
port 282 nsew signal input
rlabel metal2 s 41713 789729 42193 789785 6 mprj_io_holdover[14]
port 283 nsew signal input
rlabel metal2 s 41713 786693 42193 786749 6 mprj_io_ib_mode_sel[14]
port 284 nsew signal input
rlabel metal2 s 41713 793501 42193 793557 6 mprj_io_inp_dis[14]
port 285 nsew signal input
rlabel metal2 s 41713 786049 42193 786105 6 mprj_io_oeb[14]
port 286 nsew signal input
rlabel metal2 s 41713 789177 42193 789233 6 mprj_io_out[14]
port 287 nsew signal input
rlabel metal2 s 41713 798377 42193 798433 6 mprj_io_slow_sel[14]
port 288 nsew signal input
rlabel metal2 s 41713 787337 42193 787393 6 mprj_io_vtrip_sel[14]
port 289 nsew signal input
rlabel metal2 s 41713 800217 42193 800273 6 mprj_io_in[14]
port 290 nsew signal tristate
rlabel metal2 s 41713 785497 42193 785553 6 mprj_io_in_3v3[14]
port 291 nsew signal tristate
rlabel metal2 s 41713 280733 42193 280789 6 mprj_gpio_analog[17]
port 292 nsew signal bidirectional
rlabel metal2 s 41713 278893 42193 278949 6 mprj_gpio_noesd[17]
port 293 nsew signal bidirectional
rlabel metal5 s 6598 270420 19088 282960 6 mprj_io[35]
port 294 nsew signal bidirectional
rlabel metal2 s 41713 278341 42193 278397 6 mprj_io_analog_en[24]
port 295 nsew signal input
rlabel metal2 s 41713 277053 42193 277109 6 mprj_io_analog_pol[24]
port 296 nsew signal input
rlabel metal2 s 41713 274017 42193 274073 6 mprj_io_analog_sel[24]
port 297 nsew signal input
rlabel metal2 s 41713 277697 42193 277753 6 mprj_io_dm[72]
port 298 nsew signal input
rlabel metal2 s 41713 279537 42193 279593 6 mprj_io_dm[73]
port 299 nsew signal input
rlabel metal2 s 41713 273373 42193 273429 6 mprj_io_dm[74]
port 300 nsew signal input
rlabel metal2 s 41713 272729 42193 272785 6 mprj_io_holdover[24]
port 301 nsew signal input
rlabel metal2 s 41713 269693 42193 269749 6 mprj_io_ib_mode_sel[24]
port 302 nsew signal input
rlabel metal2 s 41713 276501 42193 276557 6 mprj_io_inp_dis[24]
port 303 nsew signal input
rlabel metal2 s 41713 269049 42193 269105 6 mprj_io_oeb[24]
port 304 nsew signal input
rlabel metal2 s 41713 272177 42193 272233 6 mprj_io_out[24]
port 305 nsew signal input
rlabel metal2 s 41713 281377 42193 281433 6 mprj_io_slow_sel[24]
port 306 nsew signal input
rlabel metal2 s 41713 270337 42193 270393 6 mprj_io_vtrip_sel[24]
port 307 nsew signal input
rlabel metal2 s 41713 283217 42193 283273 6 mprj_io_in[24]
port 308 nsew signal tristate
rlabel metal2 s 41713 268497 42193 268553 6 mprj_io_in_3v3[24]
port 309 nsew signal tristate
rlabel metal5 s 6598 227220 19088 239760 6 mprj_io[36]
port 310 nsew signal bidirectional
rlabel metal2 s 41713 235141 42193 235197 6 mprj_io_analog_en[25]
port 311 nsew signal input
rlabel metal2 s 41713 233853 42193 233909 6 mprj_io_analog_pol[25]
port 312 nsew signal input
rlabel metal2 s 41713 230817 42193 230873 6 mprj_io_analog_sel[25]
port 313 nsew signal input
rlabel metal2 s 41713 234497 42193 234553 6 mprj_io_dm[75]
port 314 nsew signal input
rlabel metal2 s 41713 236337 42193 236393 6 mprj_io_dm[76]
port 315 nsew signal input
rlabel metal2 s 41713 230173 42193 230229 6 mprj_io_dm[77]
port 316 nsew signal input
rlabel metal2 s 41713 229529 42193 229585 6 mprj_io_holdover[25]
port 317 nsew signal input
rlabel metal2 s 41713 226493 42193 226549 6 mprj_io_ib_mode_sel[25]
port 318 nsew signal input
rlabel metal2 s 41713 233301 42193 233357 6 mprj_io_inp_dis[25]
port 319 nsew signal input
rlabel metal2 s 41713 225849 42193 225905 6 mprj_io_oeb[25]
port 320 nsew signal input
rlabel metal2 s 41713 228977 42193 229033 6 mprj_io_out[25]
port 321 nsew signal input
rlabel metal2 s 41713 238177 42193 238233 6 mprj_io_slow_sel[25]
port 322 nsew signal input
rlabel metal2 s 41713 227137 42193 227193 6 mprj_io_vtrip_sel[25]
port 323 nsew signal input
rlabel metal2 s 41713 240017 42193 240073 6 mprj_io_in[25]
port 324 nsew signal tristate
rlabel metal2 s 41713 225297 42193 225353 6 mprj_io_in_3v3[25]
port 325 nsew signal tristate
rlabel metal5 s 6598 184020 19088 196560 6 mprj_io[37]
port 326 nsew signal bidirectional
rlabel metal2 s 41713 191941 42193 191997 6 mprj_io_analog_en[26]
port 327 nsew signal input
rlabel metal2 s 41713 190653 42193 190709 6 mprj_io_analog_pol[26]
port 328 nsew signal input
rlabel metal2 s 41713 187617 42193 187673 6 mprj_io_analog_sel[26]
port 329 nsew signal input
rlabel metal2 s 41713 191297 42193 191353 6 mprj_io_dm[78]
port 330 nsew signal input
rlabel metal2 s 41713 193137 42193 193193 6 mprj_io_dm[79]
port 331 nsew signal input
rlabel metal2 s 41713 186973 42193 187029 6 mprj_io_dm[80]
port 332 nsew signal input
rlabel metal2 s 41713 186329 42193 186385 6 mprj_io_holdover[26]
port 333 nsew signal input
rlabel metal2 s 41713 183293 42193 183349 6 mprj_io_ib_mode_sel[26]
port 334 nsew signal input
rlabel metal2 s 41713 190101 42193 190157 6 mprj_io_inp_dis[26]
port 335 nsew signal input
rlabel metal2 s 41713 182649 42193 182705 6 mprj_io_oeb[26]
port 336 nsew signal input
rlabel metal2 s 41713 185777 42193 185833 6 mprj_io_out[26]
port 337 nsew signal input
rlabel metal2 s 41713 194977 42193 195033 6 mprj_io_slow_sel[26]
port 338 nsew signal input
rlabel metal2 s 41713 183937 42193 183993 6 mprj_io_vtrip_sel[26]
port 339 nsew signal input
rlabel metal2 s 41713 196817 42193 196873 6 mprj_io_in[26]
port 340 nsew signal tristate
rlabel metal2 s 41713 182097 42193 182153 6 mprj_io_in_3v3[26]
port 341 nsew signal tristate
rlabel metal2 s 41713 754533 42193 754589 6 mprj_gpio_analog[8]
port 342 nsew signal bidirectional
rlabel metal2 s 41713 752693 42193 752749 6 mprj_gpio_noesd[8]
port 343 nsew signal bidirectional
rlabel metal5 s 6598 744220 19088 756760 6 mprj_io[26]
port 344 nsew signal bidirectional
rlabel metal2 s 41713 752141 42193 752197 6 mprj_io_analog_en[15]
port 345 nsew signal input
rlabel metal2 s 41713 750853 42193 750909 6 mprj_io_analog_pol[15]
port 346 nsew signal input
rlabel metal2 s 41713 747817 42193 747873 6 mprj_io_analog_sel[15]
port 347 nsew signal input
rlabel metal2 s 41713 751497 42193 751553 6 mprj_io_dm[45]
port 348 nsew signal input
rlabel metal2 s 41713 753337 42193 753393 6 mprj_io_dm[46]
port 349 nsew signal input
rlabel metal2 s 41713 747173 42193 747229 6 mprj_io_dm[47]
port 350 nsew signal input
rlabel metal2 s 41713 746529 42193 746585 6 mprj_io_holdover[15]
port 351 nsew signal input
rlabel metal2 s 41713 743493 42193 743549 6 mprj_io_ib_mode_sel[15]
port 352 nsew signal input
rlabel metal2 s 41713 750301 42193 750357 6 mprj_io_inp_dis[15]
port 353 nsew signal input
rlabel metal2 s 41713 742849 42193 742905 6 mprj_io_oeb[15]
port 354 nsew signal input
rlabel metal2 s 41713 745977 42193 746033 6 mprj_io_out[15]
port 355 nsew signal input
rlabel metal2 s 41713 755177 42193 755233 6 mprj_io_slow_sel[15]
port 356 nsew signal input
rlabel metal2 s 41713 744137 42193 744193 6 mprj_io_vtrip_sel[15]
port 357 nsew signal input
rlabel metal2 s 41713 757017 42193 757073 6 mprj_io_in[15]
port 358 nsew signal tristate
rlabel metal2 s 41713 742297 42193 742353 6 mprj_io_in_3v3[15]
port 359 nsew signal tristate
rlabel metal2 s 41713 711333 42193 711389 6 mprj_gpio_analog[9]
port 360 nsew signal bidirectional
rlabel metal2 s 41713 709493 42193 709549 6 mprj_gpio_noesd[9]
port 361 nsew signal bidirectional
rlabel metal5 s 6598 701020 19088 713560 6 mprj_io[27]
port 362 nsew signal bidirectional
rlabel metal2 s 41713 708941 42193 708997 6 mprj_io_analog_en[16]
port 363 nsew signal input
rlabel metal2 s 41713 707653 42193 707709 6 mprj_io_analog_pol[16]
port 364 nsew signal input
rlabel metal2 s 41713 704617 42193 704673 6 mprj_io_analog_sel[16]
port 365 nsew signal input
rlabel metal2 s 41713 708297 42193 708353 6 mprj_io_dm[48]
port 366 nsew signal input
rlabel metal2 s 41713 710137 42193 710193 6 mprj_io_dm[49]
port 367 nsew signal input
rlabel metal2 s 41713 703973 42193 704029 6 mprj_io_dm[50]
port 368 nsew signal input
rlabel metal2 s 41713 703329 42193 703385 6 mprj_io_holdover[16]
port 369 nsew signal input
rlabel metal2 s 41713 700293 42193 700349 6 mprj_io_ib_mode_sel[16]
port 370 nsew signal input
rlabel metal2 s 41713 707101 42193 707157 6 mprj_io_inp_dis[16]
port 371 nsew signal input
rlabel metal2 s 41713 699649 42193 699705 6 mprj_io_oeb[16]
port 372 nsew signal input
rlabel metal2 s 41713 702777 42193 702833 6 mprj_io_out[16]
port 373 nsew signal input
rlabel metal2 s 41713 711977 42193 712033 6 mprj_io_slow_sel[16]
port 374 nsew signal input
rlabel metal2 s 41713 700937 42193 700993 6 mprj_io_vtrip_sel[16]
port 375 nsew signal input
rlabel metal2 s 41713 713817 42193 713873 6 mprj_io_in[16]
port 376 nsew signal tristate
rlabel metal2 s 41713 699097 42193 699153 6 mprj_io_in_3v3[16]
port 377 nsew signal tristate
rlabel metal2 s 41713 667933 42193 667989 6 mprj_gpio_analog[10]
port 378 nsew signal bidirectional
rlabel metal2 s 41713 666093 42193 666149 6 mprj_gpio_noesd[10]
port 379 nsew signal bidirectional
rlabel metal5 s 6598 657620 19088 670160 6 mprj_io[28]
port 380 nsew signal bidirectional
rlabel metal2 s 41713 665541 42193 665597 6 mprj_io_analog_en[17]
port 381 nsew signal input
rlabel metal2 s 41713 664253 42193 664309 6 mprj_io_analog_pol[17]
port 382 nsew signal input
rlabel metal2 s 41713 661217 42193 661273 6 mprj_io_analog_sel[17]
port 383 nsew signal input
rlabel metal2 s 41713 664897 42193 664953 6 mprj_io_dm[51]
port 384 nsew signal input
rlabel metal2 s 41713 666737 42193 666793 6 mprj_io_dm[52]
port 385 nsew signal input
rlabel metal2 s 41713 660573 42193 660629 6 mprj_io_dm[53]
port 386 nsew signal input
rlabel metal2 s 41713 659929 42193 659985 6 mprj_io_holdover[17]
port 387 nsew signal input
rlabel metal2 s 41713 656893 42193 656949 6 mprj_io_ib_mode_sel[17]
port 388 nsew signal input
rlabel metal2 s 41713 663701 42193 663757 6 mprj_io_inp_dis[17]
port 389 nsew signal input
rlabel metal2 s 41713 656249 42193 656305 6 mprj_io_oeb[17]
port 390 nsew signal input
rlabel metal2 s 41713 659377 42193 659433 6 mprj_io_out[17]
port 391 nsew signal input
rlabel metal2 s 41713 668577 42193 668633 6 mprj_io_slow_sel[17]
port 392 nsew signal input
rlabel metal2 s 41713 657537 42193 657593 6 mprj_io_vtrip_sel[17]
port 393 nsew signal input
rlabel metal2 s 41713 670417 42193 670473 6 mprj_io_in[17]
port 394 nsew signal tristate
rlabel metal2 s 41713 655697 42193 655753 6 mprj_io_in_3v3[17]
port 395 nsew signal tristate
rlabel metal2 s 41713 624733 42193 624789 6 mprj_gpio_analog[11]
port 396 nsew signal bidirectional
rlabel metal2 s 41713 622893 42193 622949 6 mprj_gpio_noesd[11]
port 397 nsew signal bidirectional
rlabel metal5 s 6598 614420 19088 626960 6 mprj_io[29]
port 398 nsew signal bidirectional
rlabel metal2 s 41713 622341 42193 622397 6 mprj_io_analog_en[18]
port 399 nsew signal input
rlabel metal2 s 41713 621053 42193 621109 6 mprj_io_analog_pol[18]
port 400 nsew signal input
rlabel metal2 s 41713 618017 42193 618073 6 mprj_io_analog_sel[18]
port 401 nsew signal input
rlabel metal2 s 41713 621697 42193 621753 6 mprj_io_dm[54]
port 402 nsew signal input
rlabel metal2 s 41713 623537 42193 623593 6 mprj_io_dm[55]
port 403 nsew signal input
rlabel metal2 s 41713 617373 42193 617429 6 mprj_io_dm[56]
port 404 nsew signal input
rlabel metal2 s 41713 616729 42193 616785 6 mprj_io_holdover[18]
port 405 nsew signal input
rlabel metal2 s 41713 613693 42193 613749 6 mprj_io_ib_mode_sel[18]
port 406 nsew signal input
rlabel metal2 s 41713 620501 42193 620557 6 mprj_io_inp_dis[18]
port 407 nsew signal input
rlabel metal2 s 41713 613049 42193 613105 6 mprj_io_oeb[18]
port 408 nsew signal input
rlabel metal2 s 41713 616177 42193 616233 6 mprj_io_out[18]
port 409 nsew signal input
rlabel metal2 s 41713 625377 42193 625433 6 mprj_io_slow_sel[18]
port 410 nsew signal input
rlabel metal2 s 41713 614337 42193 614393 6 mprj_io_vtrip_sel[18]
port 411 nsew signal input
rlabel metal2 s 41713 627217 42193 627273 6 mprj_io_in[18]
port 412 nsew signal tristate
rlabel metal2 s 41713 612497 42193 612553 6 mprj_io_in_3v3[18]
port 413 nsew signal tristate
rlabel metal2 s 41713 581533 42193 581589 6 mprj_gpio_analog[12]
port 414 nsew signal bidirectional
rlabel metal2 s 41713 579693 42193 579749 6 mprj_gpio_noesd[12]
port 415 nsew signal bidirectional
rlabel metal5 s 6598 571220 19088 583760 6 mprj_io[30]
port 416 nsew signal bidirectional
rlabel metal2 s 41713 579141 42193 579197 6 mprj_io_analog_en[19]
port 417 nsew signal input
rlabel metal2 s 41713 577853 42193 577909 6 mprj_io_analog_pol[19]
port 418 nsew signal input
rlabel metal2 s 41713 574817 42193 574873 6 mprj_io_analog_sel[19]
port 419 nsew signal input
rlabel metal2 s 41713 578497 42193 578553 6 mprj_io_dm[57]
port 420 nsew signal input
rlabel metal2 s 41713 580337 42193 580393 6 mprj_io_dm[58]
port 421 nsew signal input
rlabel metal2 s 41713 574173 42193 574229 6 mprj_io_dm[59]
port 422 nsew signal input
rlabel metal2 s 41713 573529 42193 573585 6 mprj_io_holdover[19]
port 423 nsew signal input
rlabel metal2 s 41713 570493 42193 570549 6 mprj_io_ib_mode_sel[19]
port 424 nsew signal input
rlabel metal2 s 41713 577301 42193 577357 6 mprj_io_inp_dis[19]
port 425 nsew signal input
rlabel metal2 s 41713 569849 42193 569905 6 mprj_io_oeb[19]
port 426 nsew signal input
rlabel metal2 s 41713 572977 42193 573033 6 mprj_io_out[19]
port 427 nsew signal input
rlabel metal2 s 41713 582177 42193 582233 6 mprj_io_slow_sel[19]
port 428 nsew signal input
rlabel metal2 s 41713 571137 42193 571193 6 mprj_io_vtrip_sel[19]
port 429 nsew signal input
rlabel metal2 s 41713 584017 42193 584073 6 mprj_io_in[19]
port 430 nsew signal tristate
rlabel metal2 s 41713 569297 42193 569353 6 mprj_io_in_3v3[19]
port 431 nsew signal tristate
rlabel metal2 s 41713 538333 42193 538389 6 mprj_gpio_analog[13]
port 432 nsew signal bidirectional
rlabel metal2 s 41713 536493 42193 536549 6 mprj_gpio_noesd[13]
port 433 nsew signal bidirectional
rlabel metal5 s 6598 528020 19088 540560 6 mprj_io[31]
port 434 nsew signal bidirectional
rlabel metal2 s 41713 535941 42193 535997 6 mprj_io_analog_en[20]
port 435 nsew signal input
rlabel metal2 s 41713 534653 42193 534709 6 mprj_io_analog_pol[20]
port 436 nsew signal input
rlabel metal2 s 41713 531617 42193 531673 6 mprj_io_analog_sel[20]
port 437 nsew signal input
rlabel metal2 s 41713 535297 42193 535353 6 mprj_io_dm[60]
port 438 nsew signal input
rlabel metal2 s 41713 537137 42193 537193 6 mprj_io_dm[61]
port 439 nsew signal input
rlabel metal2 s 41713 530973 42193 531029 6 mprj_io_dm[62]
port 440 nsew signal input
rlabel metal2 s 41713 530329 42193 530385 6 mprj_io_holdover[20]
port 441 nsew signal input
rlabel metal2 s 41713 527293 42193 527349 6 mprj_io_ib_mode_sel[20]
port 442 nsew signal input
rlabel metal2 s 41713 534101 42193 534157 6 mprj_io_inp_dis[20]
port 443 nsew signal input
rlabel metal2 s 41713 526649 42193 526705 6 mprj_io_oeb[20]
port 444 nsew signal input
rlabel metal2 s 41713 529777 42193 529833 6 mprj_io_out[20]
port 445 nsew signal input
rlabel metal2 s 41713 538977 42193 539033 6 mprj_io_slow_sel[20]
port 446 nsew signal input
rlabel metal2 s 41713 527937 42193 527993 6 mprj_io_vtrip_sel[20]
port 447 nsew signal input
rlabel metal2 s 41713 540817 42193 540873 6 mprj_io_in[20]
port 448 nsew signal tristate
rlabel metal2 s 41713 526097 42193 526153 6 mprj_io_in_3v3[20]
port 449 nsew signal tristate
rlabel metal2 s 41713 410533 42193 410589 6 mprj_gpio_analog[14]
port 450 nsew signal bidirectional
rlabel metal2 s 41713 408693 42193 408749 6 mprj_gpio_noesd[14]
port 451 nsew signal bidirectional
rlabel metal5 s 6598 400220 19088 412760 6 mprj_io[32]
port 452 nsew signal bidirectional
rlabel metal2 s 41713 408141 42193 408197 6 mprj_io_analog_en[21]
port 453 nsew signal input
rlabel metal2 s 41713 406853 42193 406909 6 mprj_io_analog_pol[21]
port 454 nsew signal input
rlabel metal2 s 41713 403817 42193 403873 6 mprj_io_analog_sel[21]
port 455 nsew signal input
rlabel metal2 s 41713 407497 42193 407553 6 mprj_io_dm[63]
port 456 nsew signal input
rlabel metal2 s 41713 409337 42193 409393 6 mprj_io_dm[64]
port 457 nsew signal input
rlabel metal2 s 41713 403173 42193 403229 6 mprj_io_dm[65]
port 458 nsew signal input
rlabel metal2 s 41713 402529 42193 402585 6 mprj_io_holdover[21]
port 459 nsew signal input
rlabel metal2 s 41713 399493 42193 399549 6 mprj_io_ib_mode_sel[21]
port 460 nsew signal input
rlabel metal2 s 41713 406301 42193 406357 6 mprj_io_inp_dis[21]
port 461 nsew signal input
rlabel metal2 s 41713 398849 42193 398905 6 mprj_io_oeb[21]
port 462 nsew signal input
rlabel metal2 s 41713 401977 42193 402033 6 mprj_io_out[21]
port 463 nsew signal input
rlabel metal2 s 41713 411177 42193 411233 6 mprj_io_slow_sel[21]
port 464 nsew signal input
rlabel metal2 s 41713 400137 42193 400193 6 mprj_io_vtrip_sel[21]
port 465 nsew signal input
rlabel metal2 s 41713 413017 42193 413073 6 mprj_io_in[21]
port 466 nsew signal tristate
rlabel metal2 s 41713 398297 42193 398353 6 mprj_io_in_3v3[21]
port 467 nsew signal tristate
rlabel metal2 s 41713 367333 42193 367389 6 mprj_gpio_analog[15]
port 468 nsew signal bidirectional
rlabel metal2 s 41713 365493 42193 365549 6 mprj_gpio_noesd[15]
port 469 nsew signal bidirectional
rlabel metal5 s 6598 357020 19088 369560 6 mprj_io[33]
port 470 nsew signal bidirectional
rlabel metal2 s 41713 364941 42193 364997 6 mprj_io_analog_en[22]
port 471 nsew signal input
rlabel metal2 s 41713 363653 42193 363709 6 mprj_io_analog_pol[22]
port 472 nsew signal input
rlabel metal2 s 41713 360617 42193 360673 6 mprj_io_analog_sel[22]
port 473 nsew signal input
rlabel metal2 s 41713 364297 42193 364353 6 mprj_io_dm[66]
port 474 nsew signal input
rlabel metal2 s 41713 366137 42193 366193 6 mprj_io_dm[67]
port 475 nsew signal input
rlabel metal2 s 41713 359973 42193 360029 6 mprj_io_dm[68]
port 476 nsew signal input
rlabel metal2 s 41713 359329 42193 359385 6 mprj_io_holdover[22]
port 477 nsew signal input
rlabel metal2 s 41713 356293 42193 356349 6 mprj_io_ib_mode_sel[22]
port 478 nsew signal input
rlabel metal2 s 41713 363101 42193 363157 6 mprj_io_inp_dis[22]
port 479 nsew signal input
rlabel metal2 s 41713 355649 42193 355705 6 mprj_io_oeb[22]
port 480 nsew signal input
rlabel metal2 s 41713 358777 42193 358833 6 mprj_io_out[22]
port 481 nsew signal input
rlabel metal2 s 41713 367977 42193 368033 6 mprj_io_slow_sel[22]
port 482 nsew signal input
rlabel metal2 s 41713 356937 42193 356993 6 mprj_io_vtrip_sel[22]
port 483 nsew signal input
rlabel metal2 s 41713 369817 42193 369873 6 mprj_io_in[22]
port 484 nsew signal tristate
rlabel metal2 s 41713 355097 42193 355153 6 mprj_io_in_3v3[22]
port 485 nsew signal tristate
rlabel metal2 s 41713 323933 42193 323989 6 mprj_gpio_analog[16]
port 486 nsew signal bidirectional
rlabel metal2 s 41713 322093 42193 322149 6 mprj_gpio_noesd[16]
port 487 nsew signal bidirectional
rlabel metal5 s 6598 313620 19088 326160 6 mprj_io[34]
port 488 nsew signal bidirectional
rlabel metal2 s 41713 321541 42193 321597 6 mprj_io_analog_en[23]
port 489 nsew signal input
rlabel metal2 s 41713 320253 42193 320309 6 mprj_io_analog_pol[23]
port 490 nsew signal input
rlabel metal2 s 41713 317217 42193 317273 6 mprj_io_analog_sel[23]
port 491 nsew signal input
rlabel metal2 s 41713 320897 42193 320953 6 mprj_io_dm[69]
port 492 nsew signal input
rlabel metal2 s 41713 322737 42193 322793 6 mprj_io_dm[70]
port 493 nsew signal input
rlabel metal2 s 41713 316573 42193 316629 6 mprj_io_dm[71]
port 494 nsew signal input
rlabel metal2 s 41713 315929 42193 315985 6 mprj_io_holdover[23]
port 495 nsew signal input
rlabel metal2 s 41713 312893 42193 312949 6 mprj_io_ib_mode_sel[23]
port 496 nsew signal input
rlabel metal2 s 41713 319701 42193 319757 6 mprj_io_inp_dis[23]
port 497 nsew signal input
rlabel metal2 s 41713 312249 42193 312305 6 mprj_io_oeb[23]
port 498 nsew signal input
rlabel metal2 s 41713 315377 42193 315433 6 mprj_io_out[23]
port 499 nsew signal input
rlabel metal2 s 41713 324577 42193 324633 6 mprj_io_slow_sel[23]
port 500 nsew signal input
rlabel metal2 s 41713 313537 42193 313593 6 mprj_io_vtrip_sel[23]
port 501 nsew signal input
rlabel metal2 s 41713 326417 42193 326473 6 mprj_io_in[23]
port 502 nsew signal tristate
rlabel metal2 s 41713 311697 42193 311753 6 mprj_io_in_3v3[23]
port 503 nsew signal tristate
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 504 nsew signal input
rlabel metal5 s 136713 7143 144149 18309 6 resetb
port 505 nsew signal input
rlabel metal3 s 141667 38031 141813 39999 6 resetb_core_h
port 506 nsew signal tristate
rlabel metal4 s 132600 36323 132792 37013 6 vdda
port 507 nsew signal bidirectional
rlabel metal4 s 132600 28653 147600 28719 6 vssa
port 508 nsew signal bidirectional
rlabel metal4 s 132600 30762 132868 31674 6 vssd
port 509 nsew signal bidirectional
rlabel metal3 s 631944 997600 636944 1014070 6 mprj_analog[1]
port 510 nsew signal bidirectional
rlabel metal5 s 628410 1018624 640578 1030788 6 mprj_io[15]
port 511 nsew signal bidirectional
rlabel metal3 s 530744 997600 535744 1014070 6 mprj_analog[2]
port 512 nsew signal bidirectional
rlabel metal5 s 527210 1018624 539378 1030788 6 mprj_io[16]
port 513 nsew signal bidirectional
rlabel metal3 s 479144 997600 484144 1014070 6 mprj_analog[3]
port 514 nsew signal bidirectional
rlabel metal5 s 475610 1018624 487778 1030788 6 mprj_io[17]
port 515 nsew signal bidirectional
rlabel metal3 s 429744 997600 434744 1014070 6 mprj_analog[4]
port 516 nsew signal bidirectional
rlabel metal5 s 426210 1018624 438378 1030788 6 mprj_io[18]
port 517 nsew signal bidirectional
rlabel metal3 s 677600 934600 680736 948922 6 mprj_analog[0]
port 518 nsew signal bidirectional
rlabel metal2 s 677600 944142 682732 948922 6 mprj_clamp_high[0]
port 519 nsew signal input
rlabel metal2 s 677600 954121 678010 958901 6 mprj_clamp_low[0]
port 520 nsew signal input
rlabel metal5 s 698624 945422 710788 957590 6 mprj_io[14]
port 521 nsew signal bidirectional
rlabel metal5 s 697980 893466 711432 904346 6 vccd1_pad
port 522 nsew signal bidirectional
rlabel metal5 s 698624 805222 710788 817390 6 vdda1_pad
port 523 nsew signal bidirectional
rlabel metal5 s 698624 496422 710788 508590 6 vdda1_pad2
port 524 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030788 6 vssa1_pad
port 525 nsew signal bidirectional
rlabel metal5 s 698624 409822 710788 421990 6 vssa1_pad2
port 526 nsew signal bidirectional
rlabel metal4 s 679377 451600 680307 451854 6 vccd1
port 527 nsew signal bidirectional
rlabel metal4 s 680587 451600 681277 451792 6 vdda1
port 528 nsew signal bidirectional
rlabel metal4 s 688881 451600 688947 466600 6 vssa1
port 529 nsew signal bidirectional
rlabel metal3 s 678000 461700 685920 466500 6 vssd1
port 530 nsew signal bidirectional
rlabel metal5 s 697980 453666 711432 464546 6 vssd1_pad
port 531 nsew signal bidirectional
rlabel metal3 s 175944 997600 180944 1014070 6 mprj_analog[7]
port 532 nsew signal bidirectional
rlabel metal5 s 172410 1018624 184578 1030788 6 mprj_io[21]
port 533 nsew signal bidirectional
rlabel metal3 s 127944 997600 132944 1014070 6 mprj_analog[8]
port 534 nsew signal bidirectional
rlabel metal5 s 124410 1018624 136578 1030788 6 mprj_io[22]
port 535 nsew signal bidirectional
rlabel metal3 s 79944 997600 84944 1014070 6 mprj_analog[9]
port 536 nsew signal bidirectional
rlabel metal5 s 76410 1018624 88578 1030788 6 mprj_io[23]
port 537 nsew signal bidirectional
rlabel metal3 s 23530 960144 40000 965144 6 mprj_analog[10]
port 538 nsew signal bidirectional
rlabel metal5 s 6811 956610 18975 968778 6 mprj_io[24]
port 539 nsew signal bidirectional
rlabel metal3 s 290878 997600 305200 1000736 6 mprj_analog[5]
port 540 nsew signal bidirectional
rlabel metal2 s 290878 997600 295658 1002732 6 mprj_clamp_high[1]
port 541 nsew signal input
rlabel metal2 s 280899 997600 285679 998010 6 mprj_clamp_low[1]
port 542 nsew signal input
rlabel metal5 s 282210 1018624 294378 1030788 6 mprj_io[19]
port 543 nsew signal bidirectional
rlabel metal3 s 239478 997600 253800 1000736 6 mprj_analog[6]
port 544 nsew signal bidirectional
rlabel metal2 s 239478 997600 244258 1002732 6 mprj_clamp_high[2]
port 545 nsew signal input
rlabel metal2 s 229499 997600 234279 998010 6 mprj_clamp_low[2]
port 546 nsew signal input
rlabel metal5 s 230810 1018624 242978 1030788 6 mprj_io[20]
port 547 nsew signal bidirectional
rlabel metal5 s 6167 915054 19619 925934 6 vccd2_pad
port 548 nsew signal bidirectional
rlabel metal5 s 6811 484810 18975 496978 6 vdda2_pad
port 549 nsew signal bidirectional
rlabel metal5 s 6811 829810 18975 841978 6 vssa2_pad
port 550 nsew signal bidirectional
rlabel metal4 s 38503 455946 39593 456200 6 vccd
port 551 nsew signal bidirectional
rlabel metal4 s 37293 455946 38223 456200 6 vccd2
port 552 nsew signal bidirectional
rlabel metal4 s 36323 456007 37013 456199 6 vdda2
port 553 nsew signal bidirectional
rlabel metal4 s 32933 455946 33623 456200 6 vddio
port 554 nsew signal bidirectional
rlabel metal4 s 28653 441200 28719 456200 6 vssa2
port 555 nsew signal bidirectional
rlabel metal3 s 31680 441300 39600 446100 6 vssd2
port 556 nsew signal bidirectional
rlabel metal5 s 6167 443254 19619 454134 6 vssd2_pad
port 557 nsew signal bidirectional
rlabel metal4 s 7 456045 4843 456493 6 vssio
port 558 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
