VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 28.980000 2924.800000 30.180000 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2374.980000 2924.800000 2376.180000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2609.580000 2924.800000 2610.780000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2844.180000 2924.800000 2845.380000 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3078.780000 2924.800000 3079.980000 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3313.380000 2924.800000 3314.580000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090000 3520.400000 2879.650000 3524.800000 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790000 3520.400000 2555.350000 3524.800000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490000 3520.400000 2231.050000 3524.800000 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730000 3520.400000 1906.290000 3524.800000 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430000 3520.400000 1581.990000 3524.800000 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 263.580000 2924.800000 264.780000 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130000 3520.400000 1257.690000 3524.800000 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370000 3520.400000 932.930000 3524.800000 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070000 3520.400000 608.630000 3524.800000 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770000 3520.400000 284.330000 3524.800000 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3482.700000 -0.400000 3483.900000 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3195.060000 -0.400000 3196.260000 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2908.100000 -0.400000 2909.300000 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2620.460000 -0.400000 2621.660000 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2333.500000 -0.400000 2334.700000 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2045.860000 -0.400000 2047.060000 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 498.180000 2924.800000 499.380000 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1758.900000 -0.400000 1760.100000 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 732.780000 2924.800000 733.980000 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 967.380000 2924.800000 968.580000 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1201.980000 2924.800000 1203.180000 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1436.580000 2924.800000 1437.780000 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1671.180000 2924.800000 1672.380000 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1905.780000 2924.800000 1906.980000 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2140.380000 2924.800000 2141.580000 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 87.460000 2924.800000 88.660000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2433.460000 2924.800000 2434.660000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2668.740000 2924.800000 2669.940000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2903.340000 2924.800000 2904.540000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3137.940000 2924.800000 3139.140000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3372.540000 2924.800000 3373.740000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2798.130000 3520.400000 2798.690000 3524.800000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.830000 3520.400000 2474.390000 3524.800000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.070000 3520.400000 2149.630000 3524.800000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1824.770000 3520.400000 1825.330000 3524.800000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1500.470000 3520.400000 1501.030000 3524.800000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 322.060000 2924.800000 323.260000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.710000 3520.400000 1176.270000 3524.800000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.410000 3520.400000 851.970000 3524.800000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.110000 3520.400000 527.670000 3524.800000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.350000 3520.400000 202.910000 3524.800000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3410.620000 -0.400000 3411.820000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3123.660000 -0.400000 3124.860000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2836.020000 -0.400000 2837.220000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2549.060000 -0.400000 2550.260000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2261.420000 -0.400000 2262.620000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1974.460000 -0.400000 1975.660000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 556.660000 2924.800000 557.860000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1686.820000 -0.400000 1688.020000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1471.260000 -0.400000 1472.460000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1255.700000 -0.400000 1256.900000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1040.140000 -0.400000 1041.340000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 824.580000 -0.400000 825.780000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 609.700000 -0.400000 610.900000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 394.140000 -0.400000 395.340000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800000 178.580000 -0.400000 179.780000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 791.260000 2924.800000 792.460000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1025.860000 2924.800000 1027.060000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1260.460000 2924.800000 1261.660000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1495.060000 2924.800000 1496.260000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1729.660000 2924.800000 1730.860000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1964.260000 2924.800000 1965.460000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2198.860000 2924.800000 2200.060000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 204.420000 2924.800000 205.620000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2551.100000 2924.800000 2552.300000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2785.700000 2924.800000 2786.900000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3020.300000 2924.800000 3021.500000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3254.900000 2924.800000 3256.100000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3489.500000 2924.800000 3490.700000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750000 3520.400000 2636.310000 3524.800000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450000 3520.400000 2312.010000 3524.800000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150000 3520.400000 1987.710000 3524.800000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390000 3520.400000 1662.950000 3524.800000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090000 3520.400000 1338.650000 3524.800000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 439.020000 2924.800000 440.220000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790000 3520.400000 1014.350000 3524.800000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030000 3520.400000 689.590000 3524.800000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730000 3520.400000 365.290000 3524.800000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430000 3520.400000 40.990000 3524.800000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3267.140000 -0.400000 3268.340000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2979.500000 -0.400000 2980.700000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2692.540000 -0.400000 2693.740000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2404.900000 -0.400000 2406.100000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2117.940000 -0.400000 2119.140000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1830.300000 -0.400000 1831.500000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 673.620000 2924.800000 674.820000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1543.340000 -0.400000 1544.540000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1327.780000 -0.400000 1328.980000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1112.220000 -0.400000 1113.420000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 896.660000 -0.400000 897.860000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 681.100000 -0.400000 682.300000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 465.540000 -0.400000 466.740000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 249.980000 -0.400000 251.180000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 35.100000 -0.400000 36.300000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 908.900000 2924.800000 910.100000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1143.500000 2924.800000 1144.700000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1378.100000 2924.800000 1379.300000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1612.700000 2924.800000 1613.900000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1847.300000 2924.800000 1848.500000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2081.900000 2924.800000 2083.100000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2316.500000 2924.800000 2317.700000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 145.940000 2924.800000 147.140000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2492.620000 2924.800000 2493.820000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2727.220000 2924.800000 2728.420000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2961.820000 2924.800000 2963.020000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3196.420000 2924.800000 3197.620000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 3431.020000 2924.800000 3432.220000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170000 3520.400000 2717.730000 3524.800000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410000 3520.400000 2392.970000 3524.800000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110000 3520.400000 2068.670000 3524.800000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810000 3520.400000 1744.370000 3524.800000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050000 3520.400000 1419.610000 3524.800000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 380.540000 2924.800000 381.740000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.750000 3520.400000 1095.310000 3524.800000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.450000 3520.400000 771.010000 3524.800000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690000 3520.400000 446.250000 3524.800000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390000 3520.400000 121.950000 3524.800000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3339.220000 -0.400000 3340.420000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 3051.580000 -0.400000 3052.780000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2764.620000 -0.400000 2765.820000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2476.980000 -0.400000 2478.180000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 2189.340000 -0.400000 2190.540000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1902.380000 -0.400000 1903.580000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 615.140000 2924.800000 616.340000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1614.740000 -0.400000 1615.940000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1399.860000 -0.400000 1401.060000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 1184.300000 -0.400000 1185.500000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 968.740000 -0.400000 969.940000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 753.180000 -0.400000 754.380000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 537.620000 -0.400000 538.820000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 322.060000 -0.400000 323.260000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800000 106.500000 -0.400000 107.700000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 849.740000 2924.800000 850.940000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1084.340000 2924.800000 1085.540000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1318.940000 2924.800000 1320.140000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1553.540000 2924.800000 1554.740000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 1788.820000 2924.800000 1790.020000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2023.420000 2924.800000 2024.620000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2920.400000 2258.020000 2924.800000 2259.220000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.910000 -4.800000 633.470000 -0.400000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250000 -4.800000 2417.810000 -0.400000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730000 -4.800000 2435.290000 -0.400000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670000 -4.800000 2453.230000 -0.400000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610000 -4.800000 2471.170000 -0.400000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550000 -4.800000 2489.110000 -0.400000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030000 -4.800000 2506.590000 -0.400000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970000 -4.800000 2524.530000 -0.400000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910000 -4.800000 2542.470000 -0.400000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850000 -4.800000 2560.410000 -0.400000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790000 -4.800000 2578.350000 -0.400000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390000 -4.800000 811.950000 -0.400000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270000 -4.800000 2595.830000 -0.400000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210000 -4.800000 2613.770000 -0.400000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150000 -4.800000 2631.710000 -0.400000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090000 -4.800000 2649.650000 -0.400000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030000 -4.800000 2667.590000 -0.400000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510000 -4.800000 2685.070000 -0.400000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450000 -4.800000 2703.010000 -0.400000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390000 -4.800000 2720.950000 -0.400000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330000 -4.800000 2738.890000 -0.400000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810000 -4.800000 2756.370000 -0.400000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330000 -4.800000 829.890000 -0.400000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750000 -4.800000 2774.310000 -0.400000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690000 -4.800000 2792.250000 -0.400000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630000 -4.800000 2810.190000 -0.400000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570000 -4.800000 2828.130000 -0.400000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050000 -4.800000 2845.610000 -0.400000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990000 -4.800000 2863.550000 -0.400000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930000 -4.800000 2881.490000 -0.400000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870000 -4.800000 2899.430000 -0.400000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810000 -4.800000 847.370000 -0.400000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750000 -4.800000 865.310000 -0.400000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690000 -4.800000 883.250000 -0.400000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630000 -4.800000 901.190000 -0.400000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570000 -4.800000 919.130000 -0.400000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050000 -4.800000 936.610000 -0.400000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990000 -4.800000 954.550000 -0.400000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930000 -4.800000 972.490000 -0.400000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.850000 -4.800000 651.410000 -0.400000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870000 -4.800000 990.430000 -0.400000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350000 -4.800000 1007.910000 -0.400000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290000 -4.800000 1025.850000 -0.400000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230000 -4.800000 1043.790000 -0.400000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170000 -4.800000 1061.730000 -0.400000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110000 -4.800000 1079.670000 -0.400000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590000 -4.800000 1097.150000 -0.400000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530000 -4.800000 1115.090000 -0.400000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470000 -4.800000 1133.030000 -0.400000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410000 -4.800000 1150.970000 -0.400000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790000 -4.800000 669.350000 -0.400000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350000 -4.800000 1168.910000 -0.400000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830000 -4.800000 1186.390000 -0.400000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770000 -4.800000 1204.330000 -0.400000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710000 -4.800000 1222.270000 -0.400000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650000 -4.800000 1240.210000 -0.400000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130000 -4.800000 1257.690000 -0.400000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070000 -4.800000 1275.630000 -0.400000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010000 -4.800000 1293.570000 -0.400000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950000 -4.800000 1311.510000 -0.400000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890000 -4.800000 1329.450000 -0.400000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270000 -4.800000 686.830000 -0.400000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370000 -4.800000 1346.930000 -0.400000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310000 -4.800000 1364.870000 -0.400000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250000 -4.800000 1382.810000 -0.400000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190000 -4.800000 1400.750000 -0.400000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130000 -4.800000 1418.690000 -0.400000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610000 -4.800000 1436.170000 -0.400000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550000 -4.800000 1454.110000 -0.400000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490000 -4.800000 1472.050000 -0.400000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430000 -4.800000 1489.990000 -0.400000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910000 -4.800000 1507.470000 -0.400000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210000 -4.800000 704.770000 -0.400000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850000 -4.800000 1525.410000 -0.400000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790000 -4.800000 1543.350000 -0.400000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730000 -4.800000 1561.290000 -0.400000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670000 -4.800000 1579.230000 -0.400000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150000 -4.800000 1596.710000 -0.400000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090000 -4.800000 1614.650000 -0.400000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030000 -4.800000 1632.590000 -0.400000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970000 -4.800000 1650.530000 -0.400000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910000 -4.800000 1668.470000 -0.400000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390000 -4.800000 1685.950000 -0.400000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150000 -4.800000 722.710000 -0.400000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330000 -4.800000 1703.890000 -0.400000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270000 -4.800000 1721.830000 -0.400000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210000 -4.800000 1739.770000 -0.400000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690000 -4.800000 1757.250000 -0.400000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630000 -4.800000 1775.190000 -0.400000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570000 -4.800000 1793.130000 -0.400000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510000 -4.800000 1811.070000 -0.400000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450000 -4.800000 1829.010000 -0.400000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930000 -4.800000 1846.490000 -0.400000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870000 -4.800000 1864.430000 -0.400000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090000 -4.800000 740.650000 -0.400000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810000 -4.800000 1882.370000 -0.400000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750000 -4.800000 1900.310000 -0.400000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690000 -4.800000 1918.250000 -0.400000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170000 -4.800000 1935.730000 -0.400000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110000 -4.800000 1953.670000 -0.400000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050000 -4.800000 1971.610000 -0.400000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990000 -4.800000 1989.550000 -0.400000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470000 -4.800000 2007.030000 -0.400000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410000 -4.800000 2024.970000 -0.400000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350000 -4.800000 2042.910000 -0.400000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570000 -4.800000 758.130000 -0.400000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290000 -4.800000 2060.850000 -0.400000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230000 -4.800000 2078.790000 -0.400000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710000 -4.800000 2096.270000 -0.400000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650000 -4.800000 2114.210000 -0.400000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590000 -4.800000 2132.150000 -0.400000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530000 -4.800000 2150.090000 -0.400000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470000 -4.800000 2168.030000 -0.400000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950000 -4.800000 2185.510000 -0.400000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890000 -4.800000 2203.450000 -0.400000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830000 -4.800000 2221.390000 -0.400000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510000 -4.800000 776.070000 -0.400000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770000 -4.800000 2239.330000 -0.400000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250000 -4.800000 2256.810000 -0.400000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190000 -4.800000 2274.750000 -0.400000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130000 -4.800000 2292.690000 -0.400000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070000 -4.800000 2310.630000 -0.400000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010000 -4.800000 2328.570000 -0.400000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490000 -4.800000 2346.050000 -0.400000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430000 -4.800000 2363.990000 -0.400000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370000 -4.800000 2381.930000 -0.400000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310000 -4.800000 2399.870000 -0.400000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450000 -4.800000 794.010000 -0.400000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.890000 -4.800000 639.450000 -0.400000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770000 -4.800000 2423.330000 -0.400000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710000 -4.800000 2441.270000 -0.400000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650000 -4.800000 2459.210000 -0.400000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590000 -4.800000 2477.150000 -0.400000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530000 -4.800000 2495.090000 -0.400000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010000 -4.800000 2512.570000 -0.400000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950000 -4.800000 2530.510000 -0.400000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890000 -4.800000 2548.450000 -0.400000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830000 -4.800000 2566.390000 -0.400000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770000 -4.800000 2584.330000 -0.400000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370000 -4.800000 817.930000 -0.400000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250000 -4.800000 2601.810000 -0.400000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190000 -4.800000 2619.750000 -0.400000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130000 -4.800000 2637.690000 -0.400000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070000 -4.800000 2655.630000 -0.400000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550000 -4.800000 2673.110000 -0.400000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490000 -4.800000 2691.050000 -0.400000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430000 -4.800000 2708.990000 -0.400000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370000 -4.800000 2726.930000 -0.400000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310000 -4.800000 2744.870000 -0.400000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790000 -4.800000 2762.350000 -0.400000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310000 -4.800000 835.870000 -0.400000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730000 -4.800000 2780.290000 -0.400000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670000 -4.800000 2798.230000 -0.400000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610000 -4.800000 2816.170000 -0.400000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550000 -4.800000 2834.110000 -0.400000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030000 -4.800000 2851.590000 -0.400000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970000 -4.800000 2869.530000 -0.400000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910000 -4.800000 2887.470000 -0.400000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850000 -4.800000 2905.410000 -0.400000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790000 -4.800000 853.350000 -0.400000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730000 -4.800000 871.290000 -0.400000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670000 -4.800000 889.230000 -0.400000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610000 -4.800000 907.170000 -0.400000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090000 -4.800000 924.650000 -0.400000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030000 -4.800000 942.590000 -0.400000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970000 -4.800000 960.530000 -0.400000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910000 -4.800000 978.470000 -0.400000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 656.830000 -4.800000 657.390000 -0.400000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850000 -4.800000 996.410000 -0.400000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330000 -4.800000 1013.890000 -0.400000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270000 -4.800000 1031.830000 -0.400000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210000 -4.800000 1049.770000 -0.400000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150000 -4.800000 1067.710000 -0.400000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090000 -4.800000 1085.650000 -0.400000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570000 -4.800000 1103.130000 -0.400000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510000 -4.800000 1121.070000 -0.400000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450000 -4.800000 1139.010000 -0.400000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390000 -4.800000 1156.950000 -0.400000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 674.310000 -4.800000 674.870000 -0.400000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870000 -4.800000 1174.430000 -0.400000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810000 -4.800000 1192.370000 -0.400000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750000 -4.800000 1210.310000 -0.400000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690000 -4.800000 1228.250000 -0.400000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630000 -4.800000 1246.190000 -0.400000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110000 -4.800000 1263.670000 -0.400000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050000 -4.800000 1281.610000 -0.400000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990000 -4.800000 1299.550000 -0.400000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930000 -4.800000 1317.490000 -0.400000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870000 -4.800000 1335.430000 -0.400000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250000 -4.800000 692.810000 -0.400000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350000 -4.800000 1352.910000 -0.400000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290000 -4.800000 1370.850000 -0.400000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230000 -4.800000 1388.790000 -0.400000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170000 -4.800000 1406.730000 -0.400000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650000 -4.800000 1424.210000 -0.400000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590000 -4.800000 1442.150000 -0.400000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530000 -4.800000 1460.090000 -0.400000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470000 -4.800000 1478.030000 -0.400000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410000 -4.800000 1495.970000 -0.400000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890000 -4.800000 1513.450000 -0.400000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190000 -4.800000 710.750000 -0.400000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830000 -4.800000 1531.390000 -0.400000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770000 -4.800000 1549.330000 -0.400000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710000 -4.800000 1567.270000 -0.400000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650000 -4.800000 1585.210000 -0.400000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130000 -4.800000 1602.690000 -0.400000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070000 -4.800000 1620.630000 -0.400000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010000 -4.800000 1638.570000 -0.400000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950000 -4.800000 1656.510000 -0.400000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430000 -4.800000 1673.990000 -0.400000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370000 -4.800000 1691.930000 -0.400000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130000 -4.800000 728.690000 -0.400000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310000 -4.800000 1709.870000 -0.400000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250000 -4.800000 1727.810000 -0.400000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190000 -4.800000 1745.750000 -0.400000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670000 -4.800000 1763.230000 -0.400000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610000 -4.800000 1781.170000 -0.400000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550000 -4.800000 1799.110000 -0.400000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490000 -4.800000 1817.050000 -0.400000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430000 -4.800000 1834.990000 -0.400000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910000 -4.800000 1852.470000 -0.400000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850000 -4.800000 1870.410000 -0.400000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070000 -4.800000 746.630000 -0.400000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790000 -4.800000 1888.350000 -0.400000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730000 -4.800000 1906.290000 -0.400000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210000 -4.800000 1923.770000 -0.400000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150000 -4.800000 1941.710000 -0.400000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090000 -4.800000 1959.650000 -0.400000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030000 -4.800000 1977.590000 -0.400000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970000 -4.800000 1995.530000 -0.400000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450000 -4.800000 2013.010000 -0.400000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390000 -4.800000 2030.950000 -0.400000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330000 -4.800000 2048.890000 -0.400000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550000 -4.800000 764.110000 -0.400000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270000 -4.800000 2066.830000 -0.400000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210000 -4.800000 2084.770000 -0.400000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690000 -4.800000 2102.250000 -0.400000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630000 -4.800000 2120.190000 -0.400000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570000 -4.800000 2138.130000 -0.400000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510000 -4.800000 2156.070000 -0.400000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990000 -4.800000 2173.550000 -0.400000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930000 -4.800000 2191.490000 -0.400000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870000 -4.800000 2209.430000 -0.400000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810000 -4.800000 2227.370000 -0.400000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490000 -4.800000 782.050000 -0.400000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750000 -4.800000 2245.310000 -0.400000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230000 -4.800000 2262.790000 -0.400000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170000 -4.800000 2280.730000 -0.400000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110000 -4.800000 2298.670000 -0.400000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050000 -4.800000 2316.610000 -0.400000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990000 -4.800000 2334.550000 -0.400000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470000 -4.800000 2352.030000 -0.400000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410000 -4.800000 2369.970000 -0.400000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350000 -4.800000 2387.910000 -0.400000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290000 -4.800000 2405.850000 -0.400000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430000 -4.800000 799.990000 -0.400000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.870000 -4.800000 645.430000 -0.400000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750000 -4.800000 2429.310000 -0.400000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690000 -4.800000 2447.250000 -0.400000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630000 -4.800000 2465.190000 -0.400000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570000 -4.800000 2483.130000 -0.400000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510000 -4.800000 2501.070000 -0.400000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990000 -4.800000 2518.550000 -0.400000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930000 -4.800000 2536.490000 -0.400000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870000 -4.800000 2554.430000 -0.400000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810000 -4.800000 2572.370000 -0.400000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290000 -4.800000 2589.850000 -0.400000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350000 -4.800000 823.910000 -0.400000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230000 -4.800000 2607.790000 -0.400000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170000 -4.800000 2625.730000 -0.400000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110000 -4.800000 2643.670000 -0.400000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050000 -4.800000 2661.610000 -0.400000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530000 -4.800000 2679.090000 -0.400000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470000 -4.800000 2697.030000 -0.400000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410000 -4.800000 2714.970000 -0.400000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350000 -4.800000 2732.910000 -0.400000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290000 -4.800000 2750.850000 -0.400000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770000 -4.800000 2768.330000 -0.400000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830000 -4.800000 841.390000 -0.400000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710000 -4.800000 2786.270000 -0.400000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650000 -4.800000 2804.210000 -0.400000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590000 -4.800000 2822.150000 -0.400000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070000 -4.800000 2839.630000 -0.400000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010000 -4.800000 2857.570000 -0.400000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950000 -4.800000 2875.510000 -0.400000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890000 -4.800000 2893.450000 -0.400000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830000 -4.800000 2911.390000 -0.400000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770000 -4.800000 859.330000 -0.400000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710000 -4.800000 877.270000 -0.400000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650000 -4.800000 895.210000 -0.400000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590000 -4.800000 913.150000 -0.400000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070000 -4.800000 930.630000 -0.400000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010000 -4.800000 948.570000 -0.400000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950000 -4.800000 966.510000 -0.400000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890000 -4.800000 984.450000 -0.400000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.810000 -4.800000 663.370000 -0.400000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830000 -4.800000 1002.390000 -0.400000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310000 -4.800000 1019.870000 -0.400000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250000 -4.800000 1037.810000 -0.400000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190000 -4.800000 1055.750000 -0.400000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130000 -4.800000 1073.690000 -0.400000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610000 -4.800000 1091.170000 -0.400000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550000 -4.800000 1109.110000 -0.400000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490000 -4.800000 1127.050000 -0.400000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430000 -4.800000 1144.990000 -0.400000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370000 -4.800000 1162.930000 -0.400000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290000 -4.800000 680.850000 -0.400000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850000 -4.800000 1180.410000 -0.400000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790000 -4.800000 1198.350000 -0.400000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730000 -4.800000 1216.290000 -0.400000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670000 -4.800000 1234.230000 -0.400000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610000 -4.800000 1252.170000 -0.400000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090000 -4.800000 1269.650000 -0.400000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030000 -4.800000 1287.590000 -0.400000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970000 -4.800000 1305.530000 -0.400000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910000 -4.800000 1323.470000 -0.400000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390000 -4.800000 1340.950000 -0.400000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230000 -4.800000 698.790000 -0.400000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330000 -4.800000 1358.890000 -0.400000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270000 -4.800000 1376.830000 -0.400000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210000 -4.800000 1394.770000 -0.400000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150000 -4.800000 1412.710000 -0.400000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630000 -4.800000 1430.190000 -0.400000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570000 -4.800000 1448.130000 -0.400000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510000 -4.800000 1466.070000 -0.400000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450000 -4.800000 1484.010000 -0.400000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390000 -4.800000 1501.950000 -0.400000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870000 -4.800000 1519.430000 -0.400000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170000 -4.800000 716.730000 -0.400000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810000 -4.800000 1537.370000 -0.400000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750000 -4.800000 1555.310000 -0.400000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690000 -4.800000 1573.250000 -0.400000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170000 -4.800000 1590.730000 -0.400000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110000 -4.800000 1608.670000 -0.400000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050000 -4.800000 1626.610000 -0.400000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990000 -4.800000 1644.550000 -0.400000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930000 -4.800000 1662.490000 -0.400000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410000 -4.800000 1679.970000 -0.400000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350000 -4.800000 1697.910000 -0.400000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110000 -4.800000 734.670000 -0.400000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290000 -4.800000 1715.850000 -0.400000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230000 -4.800000 1733.790000 -0.400000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170000 -4.800000 1751.730000 -0.400000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650000 -4.800000 1769.210000 -0.400000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590000 -4.800000 1787.150000 -0.400000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530000 -4.800000 1805.090000 -0.400000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470000 -4.800000 1823.030000 -0.400000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950000 -4.800000 1840.510000 -0.400000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890000 -4.800000 1858.450000 -0.400000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830000 -4.800000 1876.390000 -0.400000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050000 -4.800000 752.610000 -0.400000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770000 -4.800000 1894.330000 -0.400000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710000 -4.800000 1912.270000 -0.400000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190000 -4.800000 1929.750000 -0.400000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130000 -4.800000 1947.690000 -0.400000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070000 -4.800000 1965.630000 -0.400000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010000 -4.800000 1983.570000 -0.400000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950000 -4.800000 2001.510000 -0.400000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430000 -4.800000 2018.990000 -0.400000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370000 -4.800000 2036.930000 -0.400000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310000 -4.800000 2054.870000 -0.400000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530000 -4.800000 770.090000 -0.400000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250000 -4.800000 2072.810000 -0.400000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730000 -4.800000 2090.290000 -0.400000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670000 -4.800000 2108.230000 -0.400000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610000 -4.800000 2126.170000 -0.400000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550000 -4.800000 2144.110000 -0.400000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490000 -4.800000 2162.050000 -0.400000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970000 -4.800000 2179.530000 -0.400000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910000 -4.800000 2197.470000 -0.400000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850000 -4.800000 2215.410000 -0.400000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790000 -4.800000 2233.350000 -0.400000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470000 -4.800000 788.030000 -0.400000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730000 -4.800000 2251.290000 -0.400000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210000 -4.800000 2268.770000 -0.400000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150000 -4.800000 2286.710000 -0.400000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090000 -4.800000 2304.650000 -0.400000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030000 -4.800000 2322.590000 -0.400000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510000 -4.800000 2340.070000 -0.400000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450000 -4.800000 2358.010000 -0.400000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390000 -4.800000 2375.950000 -0.400000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330000 -4.800000 2393.890000 -0.400000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270000 -4.800000 2411.830000 -0.400000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410000 -4.800000 805.970000 -0.400000 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810000 -4.800000 2917.370000 -0.400000 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.710000 -4.800000 3.270000 -0.400000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.230000 -4.800000 8.790000 -0.400000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.210000 -4.800000 14.770000 -0.400000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.130000 -4.800000 38.690000 -0.400000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.530000 -4.800000 241.090000 -0.400000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.010000 -4.800000 258.570000 -0.400000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.950000 -4.800000 276.510000 -0.400000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.890000 -4.800000 294.450000 -0.400000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.830000 -4.800000 312.390000 -0.400000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.770000 -4.800000 330.330000 -0.400000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.250000 -4.800000 347.810000 -0.400000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.190000 -4.800000 365.750000 -0.400000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.130000 -4.800000 383.690000 -0.400000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.070000 -4.800000 401.630000 -0.400000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.050000 -4.800000 62.610000 -0.400000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.010000 -4.800000 419.570000 -0.400000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.490000 -4.800000 437.050000 -0.400000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.430000 -4.800000 454.990000 -0.400000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.370000 -4.800000 472.930000 -0.400000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.310000 -4.800000 490.870000 -0.400000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.790000 -4.800000 508.350000 -0.400000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.730000 -4.800000 526.290000 -0.400000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.670000 -4.800000 544.230000 -0.400000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.610000 -4.800000 562.170000 -0.400000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.550000 -4.800000 580.110000 -0.400000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.970000 -4.800000 86.530000 -0.400000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.030000 -4.800000 597.590000 -0.400000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 614.970000 -4.800000 615.530000 -0.400000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.430000 -4.800000 109.990000 -0.400000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.350000 -4.800000 133.910000 -0.400000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.290000 -4.800000 151.850000 -0.400000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.230000 -4.800000 169.790000 -0.400000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.710000 -4.800000 187.270000 -0.400000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.650000 -4.800000 205.210000 -0.400000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.590000 -4.800000 223.150000 -0.400000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.190000 -4.800000 20.750000 -0.400000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.110000 -4.800000 44.670000 -0.400000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.510000 -4.800000 247.070000 -0.400000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.990000 -4.800000 264.550000 -0.400000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.930000 -4.800000 282.490000 -0.400000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.870000 -4.800000 300.430000 -0.400000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.810000 -4.800000 318.370000 -0.400000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.750000 -4.800000 336.310000 -0.400000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.230000 -4.800000 353.790000 -0.400000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.170000 -4.800000 371.730000 -0.400000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.110000 -4.800000 389.670000 -0.400000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.050000 -4.800000 407.610000 -0.400000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.030000 -4.800000 68.590000 -0.400000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.530000 -4.800000 425.090000 -0.400000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.470000 -4.800000 443.030000 -0.400000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.410000 -4.800000 460.970000 -0.400000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.350000 -4.800000 478.910000 -0.400000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.290000 -4.800000 496.850000 -0.400000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.770000 -4.800000 514.330000 -0.400000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.710000 -4.800000 532.270000 -0.400000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.650000 -4.800000 550.210000 -0.400000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.590000 -4.800000 568.150000 -0.400000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.530000 -4.800000 586.090000 -0.400000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.490000 -4.800000 92.050000 -0.400000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.010000 -4.800000 603.570000 -0.400000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.950000 -4.800000 621.510000 -0.400000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.410000 -4.800000 115.970000 -0.400000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.330000 -4.800000 139.890000 -0.400000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.270000 -4.800000 157.830000 -0.400000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.750000 -4.800000 175.310000 -0.400000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.690000 -4.800000 193.250000 -0.400000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.630000 -4.800000 211.190000 -0.400000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.570000 -4.800000 229.130000 -0.400000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.090000 -4.800000 50.650000 -0.400000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.490000 -4.800000 253.050000 -0.400000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.970000 -4.800000 270.530000 -0.400000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.910000 -4.800000 288.470000 -0.400000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.850000 -4.800000 306.410000 -0.400000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.790000 -4.800000 324.350000 -0.400000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.270000 -4.800000 341.830000 -0.400000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.210000 -4.800000 359.770000 -0.400000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 377.150000 -4.800000 377.710000 -0.400000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.090000 -4.800000 395.650000 -0.400000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.030000 -4.800000 413.590000 -0.400000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.010000 -4.800000 74.570000 -0.400000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.510000 -4.800000 431.070000 -0.400000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.450000 -4.800000 449.010000 -0.400000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.390000 -4.800000 466.950000 -0.400000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.330000 -4.800000 484.890000 -0.400000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.270000 -4.800000 502.830000 -0.400000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.750000 -4.800000 520.310000 -0.400000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.690000 -4.800000 538.250000 -0.400000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.630000 -4.800000 556.190000 -0.400000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.570000 -4.800000 574.130000 -0.400000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 591.050000 -4.800000 591.610000 -0.400000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.470000 -4.800000 98.030000 -0.400000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 608.990000 -4.800000 609.550000 -0.400000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 626.930000 -4.800000 627.490000 -0.400000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390000 -4.800000 121.950000 -0.400000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.310000 -4.800000 145.870000 -0.400000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.250000 -4.800000 163.810000 -0.400000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.730000 -4.800000 181.290000 -0.400000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.670000 -4.800000 199.230000 -0.400000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.610000 -4.800000 217.170000 -0.400000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.550000 -4.800000 235.110000 -0.400000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.070000 -4.800000 56.630000 -0.400000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.990000 -4.800000 80.550000 -0.400000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.450000 -4.800000 104.010000 -0.400000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.370000 -4.800000 127.930000 -0.400000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.170000 -4.800000 26.730000 -0.400000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.150000 -4.800000 32.710000 -0.400000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980000 -4.620000 -6.980000 3524.300000 ;
        RECT 4.020000 3520.400000 7.020000 3529.000000 ;
        RECT 184.020000 3520.400000 187.020000 3529.000000 ;
        RECT 364.020000 3520.400000 367.020000 3529.000000 ;
        RECT 544.020000 3520.400000 547.020000 3529.000000 ;
        RECT 724.020000 3520.400000 727.020000 3529.000000 ;
        RECT 904.020000 3520.400000 907.020000 3529.000000 ;
        RECT 1084.020000 3520.400000 1087.020000 3529.000000 ;
        RECT 1264.020000 3520.400000 1267.020000 3529.000000 ;
        RECT 1444.020000 3520.400000 1447.020000 3529.000000 ;
        RECT 1624.020000 3520.400000 1627.020000 3529.000000 ;
        RECT 1804.020000 3520.400000 1807.020000 3529.000000 ;
        RECT 1984.020000 3520.400000 1987.020000 3529.000000 ;
        RECT 2164.020000 3520.400000 2167.020000 3529.000000 ;
        RECT 2344.020000 3520.400000 2347.020000 3529.000000 ;
        RECT 2524.020000 3520.400000 2527.020000 3529.000000 ;
        RECT 2704.020000 3520.400000 2707.020000 3529.000000 ;
        RECT 2884.020000 3520.400000 2887.020000 3529.000000 ;
        RECT 4.020000 -9.320000 7.020000 -0.400000 ;
        RECT 184.020000 -9.320000 187.020000 -0.400000 ;
        RECT 364.020000 -9.320000 367.020000 -0.400000 ;
        RECT 544.020000 -9.320000 547.020000 -0.400000 ;
        RECT 724.020000 -9.320000 727.020000 -0.400000 ;
        RECT 904.020000 -9.320000 907.020000 -0.400000 ;
        RECT 1084.020000 -9.320000 1087.020000 -0.400000 ;
        RECT 1264.020000 -9.320000 1267.020000 -0.400000 ;
        RECT 1444.020000 -9.320000 1447.020000 -0.400000 ;
        RECT 1624.020000 -9.320000 1627.020000 -0.400000 ;
        RECT 1804.020000 -9.320000 1807.020000 -0.400000 ;
        RECT 1984.020000 -9.320000 1987.020000 -0.400000 ;
        RECT 2164.020000 -9.320000 2167.020000 -0.400000 ;
        RECT 2344.020000 -9.320000 2347.020000 -0.400000 ;
        RECT 2524.020000 -9.320000 2527.020000 -0.400000 ;
        RECT 2704.020000 -9.320000 2707.020000 -0.400000 ;
        RECT 2884.020000 -9.320000 2887.020000 -0.400000 ;
        RECT 2926.600000 -4.620000 2929.600000 3524.300000 ;
      LAYER via4 ;
        RECT -9.070000 3523.010000 -7.890000 3524.190000 ;
        RECT -9.070000 3521.410000 -7.890000 3522.590000 ;
        RECT 4.930000 3523.010000 6.110000 3524.190000 ;
        RECT 4.930000 3521.410000 6.110000 3522.590000 ;
        RECT 184.930000 3523.010000 186.110000 3524.190000 ;
        RECT 184.930000 3521.410000 186.110000 3522.590000 ;
        RECT 364.930000 3523.010000 366.110000 3524.190000 ;
        RECT 364.930000 3521.410000 366.110000 3522.590000 ;
        RECT 544.930000 3523.010000 546.110000 3524.190000 ;
        RECT 544.930000 3521.410000 546.110000 3522.590000 ;
        RECT 724.930000 3523.010000 726.110000 3524.190000 ;
        RECT 724.930000 3521.410000 726.110000 3522.590000 ;
        RECT 904.930000 3523.010000 906.110000 3524.190000 ;
        RECT 904.930000 3521.410000 906.110000 3522.590000 ;
        RECT 1084.930000 3523.010000 1086.110000 3524.190000 ;
        RECT 1084.930000 3521.410000 1086.110000 3522.590000 ;
        RECT 1264.930000 3523.010000 1266.110000 3524.190000 ;
        RECT 1264.930000 3521.410000 1266.110000 3522.590000 ;
        RECT 1444.930000 3523.010000 1446.110000 3524.190000 ;
        RECT 1444.930000 3521.410000 1446.110000 3522.590000 ;
        RECT 1624.930000 3523.010000 1626.110000 3524.190000 ;
        RECT 1624.930000 3521.410000 1626.110000 3522.590000 ;
        RECT 1804.930000 3523.010000 1806.110000 3524.190000 ;
        RECT 1804.930000 3521.410000 1806.110000 3522.590000 ;
        RECT 1984.930000 3523.010000 1986.110000 3524.190000 ;
        RECT 1984.930000 3521.410000 1986.110000 3522.590000 ;
        RECT 2164.930000 3523.010000 2166.110000 3524.190000 ;
        RECT 2164.930000 3521.410000 2166.110000 3522.590000 ;
        RECT 2344.930000 3523.010000 2346.110000 3524.190000 ;
        RECT 2344.930000 3521.410000 2346.110000 3522.590000 ;
        RECT 2524.930000 3523.010000 2526.110000 3524.190000 ;
        RECT 2524.930000 3521.410000 2526.110000 3522.590000 ;
        RECT 2704.930000 3523.010000 2706.110000 3524.190000 ;
        RECT 2704.930000 3521.410000 2706.110000 3522.590000 ;
        RECT 2884.930000 3523.010000 2886.110000 3524.190000 ;
        RECT 2884.930000 3521.410000 2886.110000 3522.590000 ;
        RECT 2927.510000 3523.010000 2928.690000 3524.190000 ;
        RECT 2927.510000 3521.410000 2928.690000 3522.590000 ;
        RECT -9.070000 3431.090000 -7.890000 3432.270000 ;
        RECT -9.070000 3429.490000 -7.890000 3430.670000 ;
        RECT -9.070000 3251.090000 -7.890000 3252.270000 ;
        RECT -9.070000 3249.490000 -7.890000 3250.670000 ;
        RECT -9.070000 3071.090000 -7.890000 3072.270000 ;
        RECT -9.070000 3069.490000 -7.890000 3070.670000 ;
        RECT -9.070000 2891.090000 -7.890000 2892.270000 ;
        RECT -9.070000 2889.490000 -7.890000 2890.670000 ;
        RECT -9.070000 2711.090000 -7.890000 2712.270000 ;
        RECT -9.070000 2709.490000 -7.890000 2710.670000 ;
        RECT -9.070000 2531.090000 -7.890000 2532.270000 ;
        RECT -9.070000 2529.490000 -7.890000 2530.670000 ;
        RECT -9.070000 2351.090000 -7.890000 2352.270000 ;
        RECT -9.070000 2349.490000 -7.890000 2350.670000 ;
        RECT -9.070000 2171.090000 -7.890000 2172.270000 ;
        RECT -9.070000 2169.490000 -7.890000 2170.670000 ;
        RECT -9.070000 1991.090000 -7.890000 1992.270000 ;
        RECT -9.070000 1989.490000 -7.890000 1990.670000 ;
        RECT -9.070000 1811.090000 -7.890000 1812.270000 ;
        RECT -9.070000 1809.490000 -7.890000 1810.670000 ;
        RECT -9.070000 1631.090000 -7.890000 1632.270000 ;
        RECT -9.070000 1629.490000 -7.890000 1630.670000 ;
        RECT -9.070000 1451.090000 -7.890000 1452.270000 ;
        RECT -9.070000 1449.490000 -7.890000 1450.670000 ;
        RECT -9.070000 1271.090000 -7.890000 1272.270000 ;
        RECT -9.070000 1269.490000 -7.890000 1270.670000 ;
        RECT -9.070000 1091.090000 -7.890000 1092.270000 ;
        RECT -9.070000 1089.490000 -7.890000 1090.670000 ;
        RECT -9.070000 911.090000 -7.890000 912.270000 ;
        RECT -9.070000 909.490000 -7.890000 910.670000 ;
        RECT -9.070000 731.090000 -7.890000 732.270000 ;
        RECT -9.070000 729.490000 -7.890000 730.670000 ;
        RECT -9.070000 551.090000 -7.890000 552.270000 ;
        RECT -9.070000 549.490000 -7.890000 550.670000 ;
        RECT -9.070000 371.090000 -7.890000 372.270000 ;
        RECT -9.070000 369.490000 -7.890000 370.670000 ;
        RECT -9.070000 191.090000 -7.890000 192.270000 ;
        RECT -9.070000 189.490000 -7.890000 190.670000 ;
        RECT -9.070000 11.090000 -7.890000 12.270000 ;
        RECT -9.070000 9.490000 -7.890000 10.670000 ;
        RECT 2927.510000 3431.090000 2928.690000 3432.270000 ;
        RECT 2927.510000 3429.490000 2928.690000 3430.670000 ;
        RECT 2927.510000 3251.090000 2928.690000 3252.270000 ;
        RECT 2927.510000 3249.490000 2928.690000 3250.670000 ;
        RECT 2927.510000 3071.090000 2928.690000 3072.270000 ;
        RECT 2927.510000 3069.490000 2928.690000 3070.670000 ;
        RECT 2927.510000 2891.090000 2928.690000 2892.270000 ;
        RECT 2927.510000 2889.490000 2928.690000 2890.670000 ;
        RECT 2927.510000 2711.090000 2928.690000 2712.270000 ;
        RECT 2927.510000 2709.490000 2928.690000 2710.670000 ;
        RECT 2927.510000 2531.090000 2928.690000 2532.270000 ;
        RECT 2927.510000 2529.490000 2928.690000 2530.670000 ;
        RECT 2927.510000 2351.090000 2928.690000 2352.270000 ;
        RECT 2927.510000 2349.490000 2928.690000 2350.670000 ;
        RECT 2927.510000 2171.090000 2928.690000 2172.270000 ;
        RECT 2927.510000 2169.490000 2928.690000 2170.670000 ;
        RECT 2927.510000 1991.090000 2928.690000 1992.270000 ;
        RECT 2927.510000 1989.490000 2928.690000 1990.670000 ;
        RECT 2927.510000 1811.090000 2928.690000 1812.270000 ;
        RECT 2927.510000 1809.490000 2928.690000 1810.670000 ;
        RECT 2927.510000 1631.090000 2928.690000 1632.270000 ;
        RECT 2927.510000 1629.490000 2928.690000 1630.670000 ;
        RECT 2927.510000 1451.090000 2928.690000 1452.270000 ;
        RECT 2927.510000 1449.490000 2928.690000 1450.670000 ;
        RECT 2927.510000 1271.090000 2928.690000 1272.270000 ;
        RECT 2927.510000 1269.490000 2928.690000 1270.670000 ;
        RECT 2927.510000 1091.090000 2928.690000 1092.270000 ;
        RECT 2927.510000 1089.490000 2928.690000 1090.670000 ;
        RECT 2927.510000 911.090000 2928.690000 912.270000 ;
        RECT 2927.510000 909.490000 2928.690000 910.670000 ;
        RECT 2927.510000 731.090000 2928.690000 732.270000 ;
        RECT 2927.510000 729.490000 2928.690000 730.670000 ;
        RECT 2927.510000 551.090000 2928.690000 552.270000 ;
        RECT 2927.510000 549.490000 2928.690000 550.670000 ;
        RECT 2927.510000 371.090000 2928.690000 372.270000 ;
        RECT 2927.510000 369.490000 2928.690000 370.670000 ;
        RECT 2927.510000 191.090000 2928.690000 192.270000 ;
        RECT 2927.510000 189.490000 2928.690000 190.670000 ;
        RECT 2927.510000 11.090000 2928.690000 12.270000 ;
        RECT 2927.510000 9.490000 2928.690000 10.670000 ;
        RECT -9.070000 -2.910000 -7.890000 -1.730000 ;
        RECT -9.070000 -4.510000 -7.890000 -3.330000 ;
        RECT 4.930000 -2.910000 6.110000 -1.730000 ;
        RECT 4.930000 -4.510000 6.110000 -3.330000 ;
        RECT 184.930000 -2.910000 186.110000 -1.730000 ;
        RECT 184.930000 -4.510000 186.110000 -3.330000 ;
        RECT 364.930000 -2.910000 366.110000 -1.730000 ;
        RECT 364.930000 -4.510000 366.110000 -3.330000 ;
        RECT 544.930000 -2.910000 546.110000 -1.730000 ;
        RECT 544.930000 -4.510000 546.110000 -3.330000 ;
        RECT 724.930000 -2.910000 726.110000 -1.730000 ;
        RECT 724.930000 -4.510000 726.110000 -3.330000 ;
        RECT 904.930000 -2.910000 906.110000 -1.730000 ;
        RECT 904.930000 -4.510000 906.110000 -3.330000 ;
        RECT 1084.930000 -2.910000 1086.110000 -1.730000 ;
        RECT 1084.930000 -4.510000 1086.110000 -3.330000 ;
        RECT 1264.930000 -2.910000 1266.110000 -1.730000 ;
        RECT 1264.930000 -4.510000 1266.110000 -3.330000 ;
        RECT 1444.930000 -2.910000 1446.110000 -1.730000 ;
        RECT 1444.930000 -4.510000 1446.110000 -3.330000 ;
        RECT 1624.930000 -2.910000 1626.110000 -1.730000 ;
        RECT 1624.930000 -4.510000 1626.110000 -3.330000 ;
        RECT 1804.930000 -2.910000 1806.110000 -1.730000 ;
        RECT 1804.930000 -4.510000 1806.110000 -3.330000 ;
        RECT 1984.930000 -2.910000 1986.110000 -1.730000 ;
        RECT 1984.930000 -4.510000 1986.110000 -3.330000 ;
        RECT 2164.930000 -2.910000 2166.110000 -1.730000 ;
        RECT 2164.930000 -4.510000 2166.110000 -3.330000 ;
        RECT 2344.930000 -2.910000 2346.110000 -1.730000 ;
        RECT 2344.930000 -4.510000 2346.110000 -3.330000 ;
        RECT 2524.930000 -2.910000 2526.110000 -1.730000 ;
        RECT 2524.930000 -4.510000 2526.110000 -3.330000 ;
        RECT 2704.930000 -2.910000 2706.110000 -1.730000 ;
        RECT 2704.930000 -4.510000 2706.110000 -3.330000 ;
        RECT 2884.930000 -2.910000 2886.110000 -1.730000 ;
        RECT 2884.930000 -4.510000 2886.110000 -3.330000 ;
        RECT 2927.510000 -2.910000 2928.690000 -1.730000 ;
        RECT 2927.510000 -4.510000 2928.690000 -3.330000 ;
      LAYER met5 ;
        RECT -9.980000 3524.300000 -6.980000 3524.310000 ;
        RECT 4.020000 3524.300000 7.020000 3524.310000 ;
        RECT 184.020000 3524.300000 187.020000 3524.310000 ;
        RECT 364.020000 3524.300000 367.020000 3524.310000 ;
        RECT 544.020000 3524.300000 547.020000 3524.310000 ;
        RECT 724.020000 3524.300000 727.020000 3524.310000 ;
        RECT 904.020000 3524.300000 907.020000 3524.310000 ;
        RECT 1084.020000 3524.300000 1087.020000 3524.310000 ;
        RECT 1264.020000 3524.300000 1267.020000 3524.310000 ;
        RECT 1444.020000 3524.300000 1447.020000 3524.310000 ;
        RECT 1624.020000 3524.300000 1627.020000 3524.310000 ;
        RECT 1804.020000 3524.300000 1807.020000 3524.310000 ;
        RECT 1984.020000 3524.300000 1987.020000 3524.310000 ;
        RECT 2164.020000 3524.300000 2167.020000 3524.310000 ;
        RECT 2344.020000 3524.300000 2347.020000 3524.310000 ;
        RECT 2524.020000 3524.300000 2527.020000 3524.310000 ;
        RECT 2704.020000 3524.300000 2707.020000 3524.310000 ;
        RECT 2884.020000 3524.300000 2887.020000 3524.310000 ;
        RECT 2926.600000 3524.300000 2929.600000 3524.310000 ;
        RECT -9.980000 3521.300000 2929.600000 3524.300000 ;
        RECT -9.980000 3521.290000 -6.980000 3521.300000 ;
        RECT 4.020000 3521.290000 7.020000 3521.300000 ;
        RECT 184.020000 3521.290000 187.020000 3521.300000 ;
        RECT 364.020000 3521.290000 367.020000 3521.300000 ;
        RECT 544.020000 3521.290000 547.020000 3521.300000 ;
        RECT 724.020000 3521.290000 727.020000 3521.300000 ;
        RECT 904.020000 3521.290000 907.020000 3521.300000 ;
        RECT 1084.020000 3521.290000 1087.020000 3521.300000 ;
        RECT 1264.020000 3521.290000 1267.020000 3521.300000 ;
        RECT 1444.020000 3521.290000 1447.020000 3521.300000 ;
        RECT 1624.020000 3521.290000 1627.020000 3521.300000 ;
        RECT 1804.020000 3521.290000 1807.020000 3521.300000 ;
        RECT 1984.020000 3521.290000 1987.020000 3521.300000 ;
        RECT 2164.020000 3521.290000 2167.020000 3521.300000 ;
        RECT 2344.020000 3521.290000 2347.020000 3521.300000 ;
        RECT 2524.020000 3521.290000 2527.020000 3521.300000 ;
        RECT 2704.020000 3521.290000 2707.020000 3521.300000 ;
        RECT 2884.020000 3521.290000 2887.020000 3521.300000 ;
        RECT 2926.600000 3521.290000 2929.600000 3521.300000 ;
        RECT -9.980000 3432.380000 -6.980000 3432.390000 ;
        RECT 2926.600000 3432.380000 2929.600000 3432.390000 ;
        RECT -14.680000 3429.380000 -0.400000 3432.380000 ;
        RECT 2920.400000 3429.380000 2934.300000 3432.380000 ;
        RECT -9.980000 3429.370000 -6.980000 3429.380000 ;
        RECT 2926.600000 3429.370000 2929.600000 3429.380000 ;
        RECT -9.980000 3252.380000 -6.980000 3252.390000 ;
        RECT 2926.600000 3252.380000 2929.600000 3252.390000 ;
        RECT -14.680000 3249.380000 -0.400000 3252.380000 ;
        RECT 2920.400000 3249.380000 2934.300000 3252.380000 ;
        RECT -9.980000 3249.370000 -6.980000 3249.380000 ;
        RECT 2926.600000 3249.370000 2929.600000 3249.380000 ;
        RECT -9.980000 3072.380000 -6.980000 3072.390000 ;
        RECT 2926.600000 3072.380000 2929.600000 3072.390000 ;
        RECT -14.680000 3069.380000 -0.400000 3072.380000 ;
        RECT 2920.400000 3069.380000 2934.300000 3072.380000 ;
        RECT -9.980000 3069.370000 -6.980000 3069.380000 ;
        RECT 2926.600000 3069.370000 2929.600000 3069.380000 ;
        RECT -9.980000 2892.380000 -6.980000 2892.390000 ;
        RECT 2926.600000 2892.380000 2929.600000 2892.390000 ;
        RECT -14.680000 2889.380000 -0.400000 2892.380000 ;
        RECT 2920.400000 2889.380000 2934.300000 2892.380000 ;
        RECT -9.980000 2889.370000 -6.980000 2889.380000 ;
        RECT 2926.600000 2889.370000 2929.600000 2889.380000 ;
        RECT -9.980000 2712.380000 -6.980000 2712.390000 ;
        RECT 2926.600000 2712.380000 2929.600000 2712.390000 ;
        RECT -14.680000 2709.380000 -0.400000 2712.380000 ;
        RECT 2920.400000 2709.380000 2934.300000 2712.380000 ;
        RECT -9.980000 2709.370000 -6.980000 2709.380000 ;
        RECT 2926.600000 2709.370000 2929.600000 2709.380000 ;
        RECT -9.980000 2532.380000 -6.980000 2532.390000 ;
        RECT 2926.600000 2532.380000 2929.600000 2532.390000 ;
        RECT -14.680000 2529.380000 -0.400000 2532.380000 ;
        RECT 2920.400000 2529.380000 2934.300000 2532.380000 ;
        RECT -9.980000 2529.370000 -6.980000 2529.380000 ;
        RECT 2926.600000 2529.370000 2929.600000 2529.380000 ;
        RECT -9.980000 2352.380000 -6.980000 2352.390000 ;
        RECT 2926.600000 2352.380000 2929.600000 2352.390000 ;
        RECT -14.680000 2349.380000 -0.400000 2352.380000 ;
        RECT 2920.400000 2349.380000 2934.300000 2352.380000 ;
        RECT -9.980000 2349.370000 -6.980000 2349.380000 ;
        RECT 2926.600000 2349.370000 2929.600000 2349.380000 ;
        RECT -9.980000 2172.380000 -6.980000 2172.390000 ;
        RECT 2926.600000 2172.380000 2929.600000 2172.390000 ;
        RECT -14.680000 2169.380000 -0.400000 2172.380000 ;
        RECT 2920.400000 2169.380000 2934.300000 2172.380000 ;
        RECT -9.980000 2169.370000 -6.980000 2169.380000 ;
        RECT 2926.600000 2169.370000 2929.600000 2169.380000 ;
        RECT -9.980000 1992.380000 -6.980000 1992.390000 ;
        RECT 2926.600000 1992.380000 2929.600000 1992.390000 ;
        RECT -14.680000 1989.380000 -0.400000 1992.380000 ;
        RECT 2920.400000 1989.380000 2934.300000 1992.380000 ;
        RECT -9.980000 1989.370000 -6.980000 1989.380000 ;
        RECT 2926.600000 1989.370000 2929.600000 1989.380000 ;
        RECT -9.980000 1812.380000 -6.980000 1812.390000 ;
        RECT 2926.600000 1812.380000 2929.600000 1812.390000 ;
        RECT -14.680000 1809.380000 -0.400000 1812.380000 ;
        RECT 2920.400000 1809.380000 2934.300000 1812.380000 ;
        RECT -9.980000 1809.370000 -6.980000 1809.380000 ;
        RECT 2926.600000 1809.370000 2929.600000 1809.380000 ;
        RECT -9.980000 1632.380000 -6.980000 1632.390000 ;
        RECT 2926.600000 1632.380000 2929.600000 1632.390000 ;
        RECT -14.680000 1629.380000 -0.400000 1632.380000 ;
        RECT 2920.400000 1629.380000 2934.300000 1632.380000 ;
        RECT -9.980000 1629.370000 -6.980000 1629.380000 ;
        RECT 2926.600000 1629.370000 2929.600000 1629.380000 ;
        RECT -9.980000 1452.380000 -6.980000 1452.390000 ;
        RECT 2926.600000 1452.380000 2929.600000 1452.390000 ;
        RECT -14.680000 1449.380000 -0.400000 1452.380000 ;
        RECT 2920.400000 1449.380000 2934.300000 1452.380000 ;
        RECT -9.980000 1449.370000 -6.980000 1449.380000 ;
        RECT 2926.600000 1449.370000 2929.600000 1449.380000 ;
        RECT -9.980000 1272.380000 -6.980000 1272.390000 ;
        RECT 2926.600000 1272.380000 2929.600000 1272.390000 ;
        RECT -14.680000 1269.380000 -0.400000 1272.380000 ;
        RECT 2920.400000 1269.380000 2934.300000 1272.380000 ;
        RECT -9.980000 1269.370000 -6.980000 1269.380000 ;
        RECT 2926.600000 1269.370000 2929.600000 1269.380000 ;
        RECT -9.980000 1092.380000 -6.980000 1092.390000 ;
        RECT 2926.600000 1092.380000 2929.600000 1092.390000 ;
        RECT -14.680000 1089.380000 -0.400000 1092.380000 ;
        RECT 2920.400000 1089.380000 2934.300000 1092.380000 ;
        RECT -9.980000 1089.370000 -6.980000 1089.380000 ;
        RECT 2926.600000 1089.370000 2929.600000 1089.380000 ;
        RECT -9.980000 912.380000 -6.980000 912.390000 ;
        RECT 2926.600000 912.380000 2929.600000 912.390000 ;
        RECT -14.680000 909.380000 -0.400000 912.380000 ;
        RECT 2920.400000 909.380000 2934.300000 912.380000 ;
        RECT -9.980000 909.370000 -6.980000 909.380000 ;
        RECT 2926.600000 909.370000 2929.600000 909.380000 ;
        RECT -9.980000 732.380000 -6.980000 732.390000 ;
        RECT 2926.600000 732.380000 2929.600000 732.390000 ;
        RECT -14.680000 729.380000 -0.400000 732.380000 ;
        RECT 2920.400000 729.380000 2934.300000 732.380000 ;
        RECT -9.980000 729.370000 -6.980000 729.380000 ;
        RECT 2926.600000 729.370000 2929.600000 729.380000 ;
        RECT -9.980000 552.380000 -6.980000 552.390000 ;
        RECT 2926.600000 552.380000 2929.600000 552.390000 ;
        RECT -14.680000 549.380000 -0.400000 552.380000 ;
        RECT 2920.400000 549.380000 2934.300000 552.380000 ;
        RECT -9.980000 549.370000 -6.980000 549.380000 ;
        RECT 2926.600000 549.370000 2929.600000 549.380000 ;
        RECT -9.980000 372.380000 -6.980000 372.390000 ;
        RECT 2926.600000 372.380000 2929.600000 372.390000 ;
        RECT -14.680000 369.380000 -0.400000 372.380000 ;
        RECT 2920.400000 369.380000 2934.300000 372.380000 ;
        RECT -9.980000 369.370000 -6.980000 369.380000 ;
        RECT 2926.600000 369.370000 2929.600000 369.380000 ;
        RECT -9.980000 192.380000 -6.980000 192.390000 ;
        RECT 2926.600000 192.380000 2929.600000 192.390000 ;
        RECT -14.680000 189.380000 -0.400000 192.380000 ;
        RECT 2920.400000 189.380000 2934.300000 192.380000 ;
        RECT -9.980000 189.370000 -6.980000 189.380000 ;
        RECT 2926.600000 189.370000 2929.600000 189.380000 ;
        RECT -9.980000 12.380000 -6.980000 12.390000 ;
        RECT 2926.600000 12.380000 2929.600000 12.390000 ;
        RECT -14.680000 9.380000 -0.400000 12.380000 ;
        RECT 2920.400000 9.380000 2934.300000 12.380000 ;
        RECT -9.980000 9.370000 -6.980000 9.380000 ;
        RECT 2926.600000 9.370000 2929.600000 9.380000 ;
        RECT -9.980000 -1.620000 -6.980000 -1.610000 ;
        RECT 4.020000 -1.620000 7.020000 -1.610000 ;
        RECT 184.020000 -1.620000 187.020000 -1.610000 ;
        RECT 364.020000 -1.620000 367.020000 -1.610000 ;
        RECT 544.020000 -1.620000 547.020000 -1.610000 ;
        RECT 724.020000 -1.620000 727.020000 -1.610000 ;
        RECT 904.020000 -1.620000 907.020000 -1.610000 ;
        RECT 1084.020000 -1.620000 1087.020000 -1.610000 ;
        RECT 1264.020000 -1.620000 1267.020000 -1.610000 ;
        RECT 1444.020000 -1.620000 1447.020000 -1.610000 ;
        RECT 1624.020000 -1.620000 1627.020000 -1.610000 ;
        RECT 1804.020000 -1.620000 1807.020000 -1.610000 ;
        RECT 1984.020000 -1.620000 1987.020000 -1.610000 ;
        RECT 2164.020000 -1.620000 2167.020000 -1.610000 ;
        RECT 2344.020000 -1.620000 2347.020000 -1.610000 ;
        RECT 2524.020000 -1.620000 2527.020000 -1.610000 ;
        RECT 2704.020000 -1.620000 2707.020000 -1.610000 ;
        RECT 2884.020000 -1.620000 2887.020000 -1.610000 ;
        RECT 2926.600000 -1.620000 2929.600000 -1.610000 ;
        RECT -9.980000 -4.620000 2929.600000 -1.620000 ;
        RECT -9.980000 -4.630000 -6.980000 -4.620000 ;
        RECT 4.020000 -4.630000 7.020000 -4.620000 ;
        RECT 184.020000 -4.630000 187.020000 -4.620000 ;
        RECT 364.020000 -4.630000 367.020000 -4.620000 ;
        RECT 544.020000 -4.630000 547.020000 -4.620000 ;
        RECT 724.020000 -4.630000 727.020000 -4.620000 ;
        RECT 904.020000 -4.630000 907.020000 -4.620000 ;
        RECT 1084.020000 -4.630000 1087.020000 -4.620000 ;
        RECT 1264.020000 -4.630000 1267.020000 -4.620000 ;
        RECT 1444.020000 -4.630000 1447.020000 -4.620000 ;
        RECT 1624.020000 -4.630000 1627.020000 -4.620000 ;
        RECT 1804.020000 -4.630000 1807.020000 -4.620000 ;
        RECT 1984.020000 -4.630000 1987.020000 -4.620000 ;
        RECT 2164.020000 -4.630000 2167.020000 -4.620000 ;
        RECT 2344.020000 -4.630000 2347.020000 -4.620000 ;
        RECT 2524.020000 -4.630000 2527.020000 -4.620000 ;
        RECT 2704.020000 -4.630000 2707.020000 -4.620000 ;
        RECT 2884.020000 -4.630000 2887.020000 -4.620000 ;
        RECT 2926.600000 -4.630000 2929.600000 -4.620000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680000 -9.320000 -11.680000 3529.000000 ;
        RECT 94.020000 3520.400000 97.020000 3529.000000 ;
        RECT 274.020000 3520.400000 277.020000 3529.000000 ;
        RECT 454.020000 3520.400000 457.020000 3529.000000 ;
        RECT 634.020000 3520.400000 637.020000 3529.000000 ;
        RECT 814.020000 3520.400000 817.020000 3529.000000 ;
        RECT 994.020000 3520.400000 997.020000 3529.000000 ;
        RECT 1174.020000 3520.400000 1177.020000 3529.000000 ;
        RECT 1354.020000 3520.400000 1357.020000 3529.000000 ;
        RECT 1534.020000 3520.400000 1537.020000 3529.000000 ;
        RECT 1714.020000 3520.400000 1717.020000 3529.000000 ;
        RECT 1894.020000 3520.400000 1897.020000 3529.000000 ;
        RECT 2074.020000 3520.400000 2077.020000 3529.000000 ;
        RECT 2254.020000 3520.400000 2257.020000 3529.000000 ;
        RECT 2434.020000 3520.400000 2437.020000 3529.000000 ;
        RECT 2614.020000 3520.400000 2617.020000 3529.000000 ;
        RECT 2794.020000 3520.400000 2797.020000 3529.000000 ;
        RECT 94.020000 -9.320000 97.020000 -0.400000 ;
        RECT 274.020000 -9.320000 277.020000 -0.400000 ;
        RECT 454.020000 -9.320000 457.020000 -0.400000 ;
        RECT 634.020000 -9.320000 637.020000 -0.400000 ;
        RECT 814.020000 -9.320000 817.020000 -0.400000 ;
        RECT 994.020000 -9.320000 997.020000 -0.400000 ;
        RECT 1174.020000 -9.320000 1177.020000 -0.400000 ;
        RECT 1354.020000 -9.320000 1357.020000 -0.400000 ;
        RECT 1534.020000 -9.320000 1537.020000 -0.400000 ;
        RECT 1714.020000 -9.320000 1717.020000 -0.400000 ;
        RECT 1894.020000 -9.320000 1897.020000 -0.400000 ;
        RECT 2074.020000 -9.320000 2077.020000 -0.400000 ;
        RECT 2254.020000 -9.320000 2257.020000 -0.400000 ;
        RECT 2434.020000 -9.320000 2437.020000 -0.400000 ;
        RECT 2614.020000 -9.320000 2617.020000 -0.400000 ;
        RECT 2794.020000 -9.320000 2797.020000 -0.400000 ;
        RECT 2931.300000 -9.320000 2934.300000 3529.000000 ;
      LAYER via4 ;
        RECT -13.770000 3527.710000 -12.590000 3528.890000 ;
        RECT -13.770000 3526.110000 -12.590000 3527.290000 ;
        RECT 94.930000 3527.710000 96.110000 3528.890000 ;
        RECT 94.930000 3526.110000 96.110000 3527.290000 ;
        RECT 274.930000 3527.710000 276.110000 3528.890000 ;
        RECT 274.930000 3526.110000 276.110000 3527.290000 ;
        RECT 454.930000 3527.710000 456.110000 3528.890000 ;
        RECT 454.930000 3526.110000 456.110000 3527.290000 ;
        RECT 634.930000 3527.710000 636.110000 3528.890000 ;
        RECT 634.930000 3526.110000 636.110000 3527.290000 ;
        RECT 814.930000 3527.710000 816.110000 3528.890000 ;
        RECT 814.930000 3526.110000 816.110000 3527.290000 ;
        RECT 994.930000 3527.710000 996.110000 3528.890000 ;
        RECT 994.930000 3526.110000 996.110000 3527.290000 ;
        RECT 1174.930000 3527.710000 1176.110000 3528.890000 ;
        RECT 1174.930000 3526.110000 1176.110000 3527.290000 ;
        RECT 1354.930000 3527.710000 1356.110000 3528.890000 ;
        RECT 1354.930000 3526.110000 1356.110000 3527.290000 ;
        RECT 1534.930000 3527.710000 1536.110000 3528.890000 ;
        RECT 1534.930000 3526.110000 1536.110000 3527.290000 ;
        RECT 1714.930000 3527.710000 1716.110000 3528.890000 ;
        RECT 1714.930000 3526.110000 1716.110000 3527.290000 ;
        RECT 1894.930000 3527.710000 1896.110000 3528.890000 ;
        RECT 1894.930000 3526.110000 1896.110000 3527.290000 ;
        RECT 2074.930000 3527.710000 2076.110000 3528.890000 ;
        RECT 2074.930000 3526.110000 2076.110000 3527.290000 ;
        RECT 2254.930000 3527.710000 2256.110000 3528.890000 ;
        RECT 2254.930000 3526.110000 2256.110000 3527.290000 ;
        RECT 2434.930000 3527.710000 2436.110000 3528.890000 ;
        RECT 2434.930000 3526.110000 2436.110000 3527.290000 ;
        RECT 2614.930000 3527.710000 2616.110000 3528.890000 ;
        RECT 2614.930000 3526.110000 2616.110000 3527.290000 ;
        RECT 2794.930000 3527.710000 2796.110000 3528.890000 ;
        RECT 2794.930000 3526.110000 2796.110000 3527.290000 ;
        RECT 2932.210000 3527.710000 2933.390000 3528.890000 ;
        RECT 2932.210000 3526.110000 2933.390000 3527.290000 ;
        RECT -13.770000 3341.090000 -12.590000 3342.270000 ;
        RECT -13.770000 3339.490000 -12.590000 3340.670000 ;
        RECT -13.770000 3161.090000 -12.590000 3162.270000 ;
        RECT -13.770000 3159.490000 -12.590000 3160.670000 ;
        RECT -13.770000 2981.090000 -12.590000 2982.270000 ;
        RECT -13.770000 2979.490000 -12.590000 2980.670000 ;
        RECT -13.770000 2801.090000 -12.590000 2802.270000 ;
        RECT -13.770000 2799.490000 -12.590000 2800.670000 ;
        RECT -13.770000 2621.090000 -12.590000 2622.270000 ;
        RECT -13.770000 2619.490000 -12.590000 2620.670000 ;
        RECT -13.770000 2441.090000 -12.590000 2442.270000 ;
        RECT -13.770000 2439.490000 -12.590000 2440.670000 ;
        RECT -13.770000 2261.090000 -12.590000 2262.270000 ;
        RECT -13.770000 2259.490000 -12.590000 2260.670000 ;
        RECT -13.770000 2081.090000 -12.590000 2082.270000 ;
        RECT -13.770000 2079.490000 -12.590000 2080.670000 ;
        RECT -13.770000 1901.090000 -12.590000 1902.270000 ;
        RECT -13.770000 1899.490000 -12.590000 1900.670000 ;
        RECT -13.770000 1721.090000 -12.590000 1722.270000 ;
        RECT -13.770000 1719.490000 -12.590000 1720.670000 ;
        RECT -13.770000 1541.090000 -12.590000 1542.270000 ;
        RECT -13.770000 1539.490000 -12.590000 1540.670000 ;
        RECT -13.770000 1361.090000 -12.590000 1362.270000 ;
        RECT -13.770000 1359.490000 -12.590000 1360.670000 ;
        RECT -13.770000 1181.090000 -12.590000 1182.270000 ;
        RECT -13.770000 1179.490000 -12.590000 1180.670000 ;
        RECT -13.770000 1001.090000 -12.590000 1002.270000 ;
        RECT -13.770000 999.490000 -12.590000 1000.670000 ;
        RECT -13.770000 821.090000 -12.590000 822.270000 ;
        RECT -13.770000 819.490000 -12.590000 820.670000 ;
        RECT -13.770000 641.090000 -12.590000 642.270000 ;
        RECT -13.770000 639.490000 -12.590000 640.670000 ;
        RECT -13.770000 461.090000 -12.590000 462.270000 ;
        RECT -13.770000 459.490000 -12.590000 460.670000 ;
        RECT -13.770000 281.090000 -12.590000 282.270000 ;
        RECT -13.770000 279.490000 -12.590000 280.670000 ;
        RECT -13.770000 101.090000 -12.590000 102.270000 ;
        RECT -13.770000 99.490000 -12.590000 100.670000 ;
        RECT 2932.210000 3341.090000 2933.390000 3342.270000 ;
        RECT 2932.210000 3339.490000 2933.390000 3340.670000 ;
        RECT 2932.210000 3161.090000 2933.390000 3162.270000 ;
        RECT 2932.210000 3159.490000 2933.390000 3160.670000 ;
        RECT 2932.210000 2981.090000 2933.390000 2982.270000 ;
        RECT 2932.210000 2979.490000 2933.390000 2980.670000 ;
        RECT 2932.210000 2801.090000 2933.390000 2802.270000 ;
        RECT 2932.210000 2799.490000 2933.390000 2800.670000 ;
        RECT 2932.210000 2621.090000 2933.390000 2622.270000 ;
        RECT 2932.210000 2619.490000 2933.390000 2620.670000 ;
        RECT 2932.210000 2441.090000 2933.390000 2442.270000 ;
        RECT 2932.210000 2439.490000 2933.390000 2440.670000 ;
        RECT 2932.210000 2261.090000 2933.390000 2262.270000 ;
        RECT 2932.210000 2259.490000 2933.390000 2260.670000 ;
        RECT 2932.210000 2081.090000 2933.390000 2082.270000 ;
        RECT 2932.210000 2079.490000 2933.390000 2080.670000 ;
        RECT 2932.210000 1901.090000 2933.390000 1902.270000 ;
        RECT 2932.210000 1899.490000 2933.390000 1900.670000 ;
        RECT 2932.210000 1721.090000 2933.390000 1722.270000 ;
        RECT 2932.210000 1719.490000 2933.390000 1720.670000 ;
        RECT 2932.210000 1541.090000 2933.390000 1542.270000 ;
        RECT 2932.210000 1539.490000 2933.390000 1540.670000 ;
        RECT 2932.210000 1361.090000 2933.390000 1362.270000 ;
        RECT 2932.210000 1359.490000 2933.390000 1360.670000 ;
        RECT 2932.210000 1181.090000 2933.390000 1182.270000 ;
        RECT 2932.210000 1179.490000 2933.390000 1180.670000 ;
        RECT 2932.210000 1001.090000 2933.390000 1002.270000 ;
        RECT 2932.210000 999.490000 2933.390000 1000.670000 ;
        RECT 2932.210000 821.090000 2933.390000 822.270000 ;
        RECT 2932.210000 819.490000 2933.390000 820.670000 ;
        RECT 2932.210000 641.090000 2933.390000 642.270000 ;
        RECT 2932.210000 639.490000 2933.390000 640.670000 ;
        RECT 2932.210000 461.090000 2933.390000 462.270000 ;
        RECT 2932.210000 459.490000 2933.390000 460.670000 ;
        RECT 2932.210000 281.090000 2933.390000 282.270000 ;
        RECT 2932.210000 279.490000 2933.390000 280.670000 ;
        RECT 2932.210000 101.090000 2933.390000 102.270000 ;
        RECT 2932.210000 99.490000 2933.390000 100.670000 ;
        RECT -13.770000 -7.610000 -12.590000 -6.430000 ;
        RECT -13.770000 -9.210000 -12.590000 -8.030000 ;
        RECT 94.930000 -7.610000 96.110000 -6.430000 ;
        RECT 94.930000 -9.210000 96.110000 -8.030000 ;
        RECT 274.930000 -7.610000 276.110000 -6.430000 ;
        RECT 274.930000 -9.210000 276.110000 -8.030000 ;
        RECT 454.930000 -7.610000 456.110000 -6.430000 ;
        RECT 454.930000 -9.210000 456.110000 -8.030000 ;
        RECT 634.930000 -7.610000 636.110000 -6.430000 ;
        RECT 634.930000 -9.210000 636.110000 -8.030000 ;
        RECT 814.930000 -7.610000 816.110000 -6.430000 ;
        RECT 814.930000 -9.210000 816.110000 -8.030000 ;
        RECT 994.930000 -7.610000 996.110000 -6.430000 ;
        RECT 994.930000 -9.210000 996.110000 -8.030000 ;
        RECT 1174.930000 -7.610000 1176.110000 -6.430000 ;
        RECT 1174.930000 -9.210000 1176.110000 -8.030000 ;
        RECT 1354.930000 -7.610000 1356.110000 -6.430000 ;
        RECT 1354.930000 -9.210000 1356.110000 -8.030000 ;
        RECT 1534.930000 -7.610000 1536.110000 -6.430000 ;
        RECT 1534.930000 -9.210000 1536.110000 -8.030000 ;
        RECT 1714.930000 -7.610000 1716.110000 -6.430000 ;
        RECT 1714.930000 -9.210000 1716.110000 -8.030000 ;
        RECT 1894.930000 -7.610000 1896.110000 -6.430000 ;
        RECT 1894.930000 -9.210000 1896.110000 -8.030000 ;
        RECT 2074.930000 -7.610000 2076.110000 -6.430000 ;
        RECT 2074.930000 -9.210000 2076.110000 -8.030000 ;
        RECT 2254.930000 -7.610000 2256.110000 -6.430000 ;
        RECT 2254.930000 -9.210000 2256.110000 -8.030000 ;
        RECT 2434.930000 -7.610000 2436.110000 -6.430000 ;
        RECT 2434.930000 -9.210000 2436.110000 -8.030000 ;
        RECT 2614.930000 -7.610000 2616.110000 -6.430000 ;
        RECT 2614.930000 -9.210000 2616.110000 -8.030000 ;
        RECT 2794.930000 -7.610000 2796.110000 -6.430000 ;
        RECT 2794.930000 -9.210000 2796.110000 -8.030000 ;
        RECT 2932.210000 -7.610000 2933.390000 -6.430000 ;
        RECT 2932.210000 -9.210000 2933.390000 -8.030000 ;
      LAYER met5 ;
        RECT -14.680000 3529.000000 -11.680000 3529.010000 ;
        RECT 94.020000 3529.000000 97.020000 3529.010000 ;
        RECT 274.020000 3529.000000 277.020000 3529.010000 ;
        RECT 454.020000 3529.000000 457.020000 3529.010000 ;
        RECT 634.020000 3529.000000 637.020000 3529.010000 ;
        RECT 814.020000 3529.000000 817.020000 3529.010000 ;
        RECT 994.020000 3529.000000 997.020000 3529.010000 ;
        RECT 1174.020000 3529.000000 1177.020000 3529.010000 ;
        RECT 1354.020000 3529.000000 1357.020000 3529.010000 ;
        RECT 1534.020000 3529.000000 1537.020000 3529.010000 ;
        RECT 1714.020000 3529.000000 1717.020000 3529.010000 ;
        RECT 1894.020000 3529.000000 1897.020000 3529.010000 ;
        RECT 2074.020000 3529.000000 2077.020000 3529.010000 ;
        RECT 2254.020000 3529.000000 2257.020000 3529.010000 ;
        RECT 2434.020000 3529.000000 2437.020000 3529.010000 ;
        RECT 2614.020000 3529.000000 2617.020000 3529.010000 ;
        RECT 2794.020000 3529.000000 2797.020000 3529.010000 ;
        RECT 2931.300000 3529.000000 2934.300000 3529.010000 ;
        RECT -14.680000 3526.000000 2934.300000 3529.000000 ;
        RECT -14.680000 3525.990000 -11.680000 3526.000000 ;
        RECT 94.020000 3525.990000 97.020000 3526.000000 ;
        RECT 274.020000 3525.990000 277.020000 3526.000000 ;
        RECT 454.020000 3525.990000 457.020000 3526.000000 ;
        RECT 634.020000 3525.990000 637.020000 3526.000000 ;
        RECT 814.020000 3525.990000 817.020000 3526.000000 ;
        RECT 994.020000 3525.990000 997.020000 3526.000000 ;
        RECT 1174.020000 3525.990000 1177.020000 3526.000000 ;
        RECT 1354.020000 3525.990000 1357.020000 3526.000000 ;
        RECT 1534.020000 3525.990000 1537.020000 3526.000000 ;
        RECT 1714.020000 3525.990000 1717.020000 3526.000000 ;
        RECT 1894.020000 3525.990000 1897.020000 3526.000000 ;
        RECT 2074.020000 3525.990000 2077.020000 3526.000000 ;
        RECT 2254.020000 3525.990000 2257.020000 3526.000000 ;
        RECT 2434.020000 3525.990000 2437.020000 3526.000000 ;
        RECT 2614.020000 3525.990000 2617.020000 3526.000000 ;
        RECT 2794.020000 3525.990000 2797.020000 3526.000000 ;
        RECT 2931.300000 3525.990000 2934.300000 3526.000000 ;
        RECT -14.680000 3342.380000 -11.680000 3342.390000 ;
        RECT 2931.300000 3342.380000 2934.300000 3342.390000 ;
        RECT -14.680000 3339.380000 -0.400000 3342.380000 ;
        RECT 2920.400000 3339.380000 2934.300000 3342.380000 ;
        RECT -14.680000 3339.370000 -11.680000 3339.380000 ;
        RECT 2931.300000 3339.370000 2934.300000 3339.380000 ;
        RECT -14.680000 3162.380000 -11.680000 3162.390000 ;
        RECT 2931.300000 3162.380000 2934.300000 3162.390000 ;
        RECT -14.680000 3159.380000 -0.400000 3162.380000 ;
        RECT 2920.400000 3159.380000 2934.300000 3162.380000 ;
        RECT -14.680000 3159.370000 -11.680000 3159.380000 ;
        RECT 2931.300000 3159.370000 2934.300000 3159.380000 ;
        RECT -14.680000 2982.380000 -11.680000 2982.390000 ;
        RECT 2931.300000 2982.380000 2934.300000 2982.390000 ;
        RECT -14.680000 2979.380000 -0.400000 2982.380000 ;
        RECT 2920.400000 2979.380000 2934.300000 2982.380000 ;
        RECT -14.680000 2979.370000 -11.680000 2979.380000 ;
        RECT 2931.300000 2979.370000 2934.300000 2979.380000 ;
        RECT -14.680000 2802.380000 -11.680000 2802.390000 ;
        RECT 2931.300000 2802.380000 2934.300000 2802.390000 ;
        RECT -14.680000 2799.380000 -0.400000 2802.380000 ;
        RECT 2920.400000 2799.380000 2934.300000 2802.380000 ;
        RECT -14.680000 2799.370000 -11.680000 2799.380000 ;
        RECT 2931.300000 2799.370000 2934.300000 2799.380000 ;
        RECT -14.680000 2622.380000 -11.680000 2622.390000 ;
        RECT 2931.300000 2622.380000 2934.300000 2622.390000 ;
        RECT -14.680000 2619.380000 -0.400000 2622.380000 ;
        RECT 2920.400000 2619.380000 2934.300000 2622.380000 ;
        RECT -14.680000 2619.370000 -11.680000 2619.380000 ;
        RECT 2931.300000 2619.370000 2934.300000 2619.380000 ;
        RECT -14.680000 2442.380000 -11.680000 2442.390000 ;
        RECT 2931.300000 2442.380000 2934.300000 2442.390000 ;
        RECT -14.680000 2439.380000 -0.400000 2442.380000 ;
        RECT 2920.400000 2439.380000 2934.300000 2442.380000 ;
        RECT -14.680000 2439.370000 -11.680000 2439.380000 ;
        RECT 2931.300000 2439.370000 2934.300000 2439.380000 ;
        RECT -14.680000 2262.380000 -11.680000 2262.390000 ;
        RECT 2931.300000 2262.380000 2934.300000 2262.390000 ;
        RECT -14.680000 2259.380000 -0.400000 2262.380000 ;
        RECT 2920.400000 2259.380000 2934.300000 2262.380000 ;
        RECT -14.680000 2259.370000 -11.680000 2259.380000 ;
        RECT 2931.300000 2259.370000 2934.300000 2259.380000 ;
        RECT -14.680000 2082.380000 -11.680000 2082.390000 ;
        RECT 2931.300000 2082.380000 2934.300000 2082.390000 ;
        RECT -14.680000 2079.380000 -0.400000 2082.380000 ;
        RECT 2920.400000 2079.380000 2934.300000 2082.380000 ;
        RECT -14.680000 2079.370000 -11.680000 2079.380000 ;
        RECT 2931.300000 2079.370000 2934.300000 2079.380000 ;
        RECT -14.680000 1902.380000 -11.680000 1902.390000 ;
        RECT 2931.300000 1902.380000 2934.300000 1902.390000 ;
        RECT -14.680000 1899.380000 -0.400000 1902.380000 ;
        RECT 2920.400000 1899.380000 2934.300000 1902.380000 ;
        RECT -14.680000 1899.370000 -11.680000 1899.380000 ;
        RECT 2931.300000 1899.370000 2934.300000 1899.380000 ;
        RECT -14.680000 1722.380000 -11.680000 1722.390000 ;
        RECT 2931.300000 1722.380000 2934.300000 1722.390000 ;
        RECT -14.680000 1719.380000 -0.400000 1722.380000 ;
        RECT 2920.400000 1719.380000 2934.300000 1722.380000 ;
        RECT -14.680000 1719.370000 -11.680000 1719.380000 ;
        RECT 2931.300000 1719.370000 2934.300000 1719.380000 ;
        RECT -14.680000 1542.380000 -11.680000 1542.390000 ;
        RECT 2931.300000 1542.380000 2934.300000 1542.390000 ;
        RECT -14.680000 1539.380000 -0.400000 1542.380000 ;
        RECT 2920.400000 1539.380000 2934.300000 1542.380000 ;
        RECT -14.680000 1539.370000 -11.680000 1539.380000 ;
        RECT 2931.300000 1539.370000 2934.300000 1539.380000 ;
        RECT -14.680000 1362.380000 -11.680000 1362.390000 ;
        RECT 2931.300000 1362.380000 2934.300000 1362.390000 ;
        RECT -14.680000 1359.380000 -0.400000 1362.380000 ;
        RECT 2920.400000 1359.380000 2934.300000 1362.380000 ;
        RECT -14.680000 1359.370000 -11.680000 1359.380000 ;
        RECT 2931.300000 1359.370000 2934.300000 1359.380000 ;
        RECT -14.680000 1182.380000 -11.680000 1182.390000 ;
        RECT 2931.300000 1182.380000 2934.300000 1182.390000 ;
        RECT -14.680000 1179.380000 -0.400000 1182.380000 ;
        RECT 2920.400000 1179.380000 2934.300000 1182.380000 ;
        RECT -14.680000 1179.370000 -11.680000 1179.380000 ;
        RECT 2931.300000 1179.370000 2934.300000 1179.380000 ;
        RECT -14.680000 1002.380000 -11.680000 1002.390000 ;
        RECT 2931.300000 1002.380000 2934.300000 1002.390000 ;
        RECT -14.680000 999.380000 -0.400000 1002.380000 ;
        RECT 2920.400000 999.380000 2934.300000 1002.380000 ;
        RECT -14.680000 999.370000 -11.680000 999.380000 ;
        RECT 2931.300000 999.370000 2934.300000 999.380000 ;
        RECT -14.680000 822.380000 -11.680000 822.390000 ;
        RECT 2931.300000 822.380000 2934.300000 822.390000 ;
        RECT -14.680000 819.380000 -0.400000 822.380000 ;
        RECT 2920.400000 819.380000 2934.300000 822.380000 ;
        RECT -14.680000 819.370000 -11.680000 819.380000 ;
        RECT 2931.300000 819.370000 2934.300000 819.380000 ;
        RECT -14.680000 642.380000 -11.680000 642.390000 ;
        RECT 2931.300000 642.380000 2934.300000 642.390000 ;
        RECT -14.680000 639.380000 -0.400000 642.380000 ;
        RECT 2920.400000 639.380000 2934.300000 642.380000 ;
        RECT -14.680000 639.370000 -11.680000 639.380000 ;
        RECT 2931.300000 639.370000 2934.300000 639.380000 ;
        RECT -14.680000 462.380000 -11.680000 462.390000 ;
        RECT 2931.300000 462.380000 2934.300000 462.390000 ;
        RECT -14.680000 459.380000 -0.400000 462.380000 ;
        RECT 2920.400000 459.380000 2934.300000 462.380000 ;
        RECT -14.680000 459.370000 -11.680000 459.380000 ;
        RECT 2931.300000 459.370000 2934.300000 459.380000 ;
        RECT -14.680000 282.380000 -11.680000 282.390000 ;
        RECT 2931.300000 282.380000 2934.300000 282.390000 ;
        RECT -14.680000 279.380000 -0.400000 282.380000 ;
        RECT 2920.400000 279.380000 2934.300000 282.380000 ;
        RECT -14.680000 279.370000 -11.680000 279.380000 ;
        RECT 2931.300000 279.370000 2934.300000 279.380000 ;
        RECT -14.680000 102.380000 -11.680000 102.390000 ;
        RECT 2931.300000 102.380000 2934.300000 102.390000 ;
        RECT -14.680000 99.380000 -0.400000 102.380000 ;
        RECT 2920.400000 99.380000 2934.300000 102.380000 ;
        RECT -14.680000 99.370000 -11.680000 99.380000 ;
        RECT 2931.300000 99.370000 2934.300000 99.380000 ;
        RECT -14.680000 -6.320000 -11.680000 -6.310000 ;
        RECT 94.020000 -6.320000 97.020000 -6.310000 ;
        RECT 274.020000 -6.320000 277.020000 -6.310000 ;
        RECT 454.020000 -6.320000 457.020000 -6.310000 ;
        RECT 634.020000 -6.320000 637.020000 -6.310000 ;
        RECT 814.020000 -6.320000 817.020000 -6.310000 ;
        RECT 994.020000 -6.320000 997.020000 -6.310000 ;
        RECT 1174.020000 -6.320000 1177.020000 -6.310000 ;
        RECT 1354.020000 -6.320000 1357.020000 -6.310000 ;
        RECT 1534.020000 -6.320000 1537.020000 -6.310000 ;
        RECT 1714.020000 -6.320000 1717.020000 -6.310000 ;
        RECT 1894.020000 -6.320000 1897.020000 -6.310000 ;
        RECT 2074.020000 -6.320000 2077.020000 -6.310000 ;
        RECT 2254.020000 -6.320000 2257.020000 -6.310000 ;
        RECT 2434.020000 -6.320000 2437.020000 -6.310000 ;
        RECT 2614.020000 -6.320000 2617.020000 -6.310000 ;
        RECT 2794.020000 -6.320000 2797.020000 -6.310000 ;
        RECT 2931.300000 -6.320000 2934.300000 -6.310000 ;
        RECT -14.680000 -9.320000 2934.300000 -6.320000 ;
        RECT -14.680000 -9.330000 -11.680000 -9.320000 ;
        RECT 94.020000 -9.330000 97.020000 -9.320000 ;
        RECT 274.020000 -9.330000 277.020000 -9.320000 ;
        RECT 454.020000 -9.330000 457.020000 -9.320000 ;
        RECT 634.020000 -9.330000 637.020000 -9.320000 ;
        RECT 814.020000 -9.330000 817.020000 -9.320000 ;
        RECT 994.020000 -9.330000 997.020000 -9.320000 ;
        RECT 1174.020000 -9.330000 1177.020000 -9.320000 ;
        RECT 1354.020000 -9.330000 1357.020000 -9.320000 ;
        RECT 1534.020000 -9.330000 1537.020000 -9.320000 ;
        RECT 1714.020000 -9.330000 1717.020000 -9.320000 ;
        RECT 1894.020000 -9.330000 1897.020000 -9.320000 ;
        RECT 2074.020000 -9.330000 2077.020000 -9.320000 ;
        RECT 2254.020000 -9.330000 2257.020000 -9.320000 ;
        RECT 2434.020000 -9.330000 2437.020000 -9.320000 ;
        RECT 2614.020000 -9.330000 2617.020000 -9.320000 ;
        RECT 2794.020000 -9.330000 2797.020000 -9.320000 ;
        RECT 2931.300000 -9.330000 2934.300000 -9.320000 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380000 -14.020000 -16.380000 3533.700000 ;
        RECT 22.020000 3520.400000 25.020000 3538.400000 ;
        RECT 202.020000 3520.400000 205.020000 3538.400000 ;
        RECT 382.020000 3520.400000 385.020000 3538.400000 ;
        RECT 562.020000 3520.400000 565.020000 3538.400000 ;
        RECT 742.020000 3520.400000 745.020000 3538.400000 ;
        RECT 922.020000 3520.400000 925.020000 3538.400000 ;
        RECT 1102.020000 3520.400000 1105.020000 3538.400000 ;
        RECT 1282.020000 3520.400000 1285.020000 3538.400000 ;
        RECT 1462.020000 3520.400000 1465.020000 3538.400000 ;
        RECT 1642.020000 3520.400000 1645.020000 3538.400000 ;
        RECT 1822.020000 3520.400000 1825.020000 3538.400000 ;
        RECT 2002.020000 3520.400000 2005.020000 3538.400000 ;
        RECT 2182.020000 3520.400000 2185.020000 3538.400000 ;
        RECT 2362.020000 3520.400000 2365.020000 3538.400000 ;
        RECT 2542.020000 3520.400000 2545.020000 3538.400000 ;
        RECT 2722.020000 3520.400000 2725.020000 3538.400000 ;
        RECT 2902.020000 3520.400000 2905.020000 3538.400000 ;
        RECT 22.020000 -18.720000 25.020000 -0.400000 ;
        RECT 202.020000 -18.720000 205.020000 -0.400000 ;
        RECT 382.020000 -18.720000 385.020000 -0.400000 ;
        RECT 562.020000 -18.720000 565.020000 -0.400000 ;
        RECT 742.020000 -18.720000 745.020000 -0.400000 ;
        RECT 922.020000 -18.720000 925.020000 -0.400000 ;
        RECT 1102.020000 -18.720000 1105.020000 -0.400000 ;
        RECT 1282.020000 -18.720000 1285.020000 -0.400000 ;
        RECT 1462.020000 -18.720000 1465.020000 -0.400000 ;
        RECT 1642.020000 -18.720000 1645.020000 -0.400000 ;
        RECT 1822.020000 -18.720000 1825.020000 -0.400000 ;
        RECT 2002.020000 -18.720000 2005.020000 -0.400000 ;
        RECT 2182.020000 -18.720000 2185.020000 -0.400000 ;
        RECT 2362.020000 -18.720000 2365.020000 -0.400000 ;
        RECT 2542.020000 -18.720000 2545.020000 -0.400000 ;
        RECT 2722.020000 -18.720000 2725.020000 -0.400000 ;
        RECT 2902.020000 -18.720000 2905.020000 -0.400000 ;
        RECT 2936.000000 -14.020000 2939.000000 3533.700000 ;
      LAYER via4 ;
        RECT -18.470000 3532.410000 -17.290000 3533.590000 ;
        RECT -18.470000 3530.810000 -17.290000 3531.990000 ;
        RECT 22.930000 3532.410000 24.110000 3533.590000 ;
        RECT 22.930000 3530.810000 24.110000 3531.990000 ;
        RECT 202.930000 3532.410000 204.110000 3533.590000 ;
        RECT 202.930000 3530.810000 204.110000 3531.990000 ;
        RECT 382.930000 3532.410000 384.110000 3533.590000 ;
        RECT 382.930000 3530.810000 384.110000 3531.990000 ;
        RECT 562.930000 3532.410000 564.110000 3533.590000 ;
        RECT 562.930000 3530.810000 564.110000 3531.990000 ;
        RECT 742.930000 3532.410000 744.110000 3533.590000 ;
        RECT 742.930000 3530.810000 744.110000 3531.990000 ;
        RECT 922.930000 3532.410000 924.110000 3533.590000 ;
        RECT 922.930000 3530.810000 924.110000 3531.990000 ;
        RECT 1102.930000 3532.410000 1104.110000 3533.590000 ;
        RECT 1102.930000 3530.810000 1104.110000 3531.990000 ;
        RECT 1282.930000 3532.410000 1284.110000 3533.590000 ;
        RECT 1282.930000 3530.810000 1284.110000 3531.990000 ;
        RECT 1462.930000 3532.410000 1464.110000 3533.590000 ;
        RECT 1462.930000 3530.810000 1464.110000 3531.990000 ;
        RECT 1642.930000 3532.410000 1644.110000 3533.590000 ;
        RECT 1642.930000 3530.810000 1644.110000 3531.990000 ;
        RECT 1822.930000 3532.410000 1824.110000 3533.590000 ;
        RECT 1822.930000 3530.810000 1824.110000 3531.990000 ;
        RECT 2002.930000 3532.410000 2004.110000 3533.590000 ;
        RECT 2002.930000 3530.810000 2004.110000 3531.990000 ;
        RECT 2182.930000 3532.410000 2184.110000 3533.590000 ;
        RECT 2182.930000 3530.810000 2184.110000 3531.990000 ;
        RECT 2362.930000 3532.410000 2364.110000 3533.590000 ;
        RECT 2362.930000 3530.810000 2364.110000 3531.990000 ;
        RECT 2542.930000 3532.410000 2544.110000 3533.590000 ;
        RECT 2542.930000 3530.810000 2544.110000 3531.990000 ;
        RECT 2722.930000 3532.410000 2724.110000 3533.590000 ;
        RECT 2722.930000 3530.810000 2724.110000 3531.990000 ;
        RECT 2902.930000 3532.410000 2904.110000 3533.590000 ;
        RECT 2902.930000 3530.810000 2904.110000 3531.990000 ;
        RECT 2936.910000 3532.410000 2938.090000 3533.590000 ;
        RECT 2936.910000 3530.810000 2938.090000 3531.990000 ;
        RECT -18.470000 3449.090000 -17.290000 3450.270000 ;
        RECT -18.470000 3447.490000 -17.290000 3448.670000 ;
        RECT -18.470000 3269.090000 -17.290000 3270.270000 ;
        RECT -18.470000 3267.490000 -17.290000 3268.670000 ;
        RECT -18.470000 3089.090000 -17.290000 3090.270000 ;
        RECT -18.470000 3087.490000 -17.290000 3088.670000 ;
        RECT -18.470000 2909.090000 -17.290000 2910.270000 ;
        RECT -18.470000 2907.490000 -17.290000 2908.670000 ;
        RECT -18.470000 2729.090000 -17.290000 2730.270000 ;
        RECT -18.470000 2727.490000 -17.290000 2728.670000 ;
        RECT -18.470000 2549.090000 -17.290000 2550.270000 ;
        RECT -18.470000 2547.490000 -17.290000 2548.670000 ;
        RECT -18.470000 2369.090000 -17.290000 2370.270000 ;
        RECT -18.470000 2367.490000 -17.290000 2368.670000 ;
        RECT -18.470000 2189.090000 -17.290000 2190.270000 ;
        RECT -18.470000 2187.490000 -17.290000 2188.670000 ;
        RECT -18.470000 2009.090000 -17.290000 2010.270000 ;
        RECT -18.470000 2007.490000 -17.290000 2008.670000 ;
        RECT -18.470000 1829.090000 -17.290000 1830.270000 ;
        RECT -18.470000 1827.490000 -17.290000 1828.670000 ;
        RECT -18.470000 1649.090000 -17.290000 1650.270000 ;
        RECT -18.470000 1647.490000 -17.290000 1648.670000 ;
        RECT -18.470000 1469.090000 -17.290000 1470.270000 ;
        RECT -18.470000 1467.490000 -17.290000 1468.670000 ;
        RECT -18.470000 1289.090000 -17.290000 1290.270000 ;
        RECT -18.470000 1287.490000 -17.290000 1288.670000 ;
        RECT -18.470000 1109.090000 -17.290000 1110.270000 ;
        RECT -18.470000 1107.490000 -17.290000 1108.670000 ;
        RECT -18.470000 929.090000 -17.290000 930.270000 ;
        RECT -18.470000 927.490000 -17.290000 928.670000 ;
        RECT -18.470000 749.090000 -17.290000 750.270000 ;
        RECT -18.470000 747.490000 -17.290000 748.670000 ;
        RECT -18.470000 569.090000 -17.290000 570.270000 ;
        RECT -18.470000 567.490000 -17.290000 568.670000 ;
        RECT -18.470000 389.090000 -17.290000 390.270000 ;
        RECT -18.470000 387.490000 -17.290000 388.670000 ;
        RECT -18.470000 209.090000 -17.290000 210.270000 ;
        RECT -18.470000 207.490000 -17.290000 208.670000 ;
        RECT -18.470000 29.090000 -17.290000 30.270000 ;
        RECT -18.470000 27.490000 -17.290000 28.670000 ;
        RECT 2936.910000 3449.090000 2938.090000 3450.270000 ;
        RECT 2936.910000 3447.490000 2938.090000 3448.670000 ;
        RECT 2936.910000 3269.090000 2938.090000 3270.270000 ;
        RECT 2936.910000 3267.490000 2938.090000 3268.670000 ;
        RECT 2936.910000 3089.090000 2938.090000 3090.270000 ;
        RECT 2936.910000 3087.490000 2938.090000 3088.670000 ;
        RECT 2936.910000 2909.090000 2938.090000 2910.270000 ;
        RECT 2936.910000 2907.490000 2938.090000 2908.670000 ;
        RECT 2936.910000 2729.090000 2938.090000 2730.270000 ;
        RECT 2936.910000 2727.490000 2938.090000 2728.670000 ;
        RECT 2936.910000 2549.090000 2938.090000 2550.270000 ;
        RECT 2936.910000 2547.490000 2938.090000 2548.670000 ;
        RECT 2936.910000 2369.090000 2938.090000 2370.270000 ;
        RECT 2936.910000 2367.490000 2938.090000 2368.670000 ;
        RECT 2936.910000 2189.090000 2938.090000 2190.270000 ;
        RECT 2936.910000 2187.490000 2938.090000 2188.670000 ;
        RECT 2936.910000 2009.090000 2938.090000 2010.270000 ;
        RECT 2936.910000 2007.490000 2938.090000 2008.670000 ;
        RECT 2936.910000 1829.090000 2938.090000 1830.270000 ;
        RECT 2936.910000 1827.490000 2938.090000 1828.670000 ;
        RECT 2936.910000 1649.090000 2938.090000 1650.270000 ;
        RECT 2936.910000 1647.490000 2938.090000 1648.670000 ;
        RECT 2936.910000 1469.090000 2938.090000 1470.270000 ;
        RECT 2936.910000 1467.490000 2938.090000 1468.670000 ;
        RECT 2936.910000 1289.090000 2938.090000 1290.270000 ;
        RECT 2936.910000 1287.490000 2938.090000 1288.670000 ;
        RECT 2936.910000 1109.090000 2938.090000 1110.270000 ;
        RECT 2936.910000 1107.490000 2938.090000 1108.670000 ;
        RECT 2936.910000 929.090000 2938.090000 930.270000 ;
        RECT 2936.910000 927.490000 2938.090000 928.670000 ;
        RECT 2936.910000 749.090000 2938.090000 750.270000 ;
        RECT 2936.910000 747.490000 2938.090000 748.670000 ;
        RECT 2936.910000 569.090000 2938.090000 570.270000 ;
        RECT 2936.910000 567.490000 2938.090000 568.670000 ;
        RECT 2936.910000 389.090000 2938.090000 390.270000 ;
        RECT 2936.910000 387.490000 2938.090000 388.670000 ;
        RECT 2936.910000 209.090000 2938.090000 210.270000 ;
        RECT 2936.910000 207.490000 2938.090000 208.670000 ;
        RECT 2936.910000 29.090000 2938.090000 30.270000 ;
        RECT 2936.910000 27.490000 2938.090000 28.670000 ;
        RECT -18.470000 -12.310000 -17.290000 -11.130000 ;
        RECT -18.470000 -13.910000 -17.290000 -12.730000 ;
        RECT 22.930000 -12.310000 24.110000 -11.130000 ;
        RECT 22.930000 -13.910000 24.110000 -12.730000 ;
        RECT 202.930000 -12.310000 204.110000 -11.130000 ;
        RECT 202.930000 -13.910000 204.110000 -12.730000 ;
        RECT 382.930000 -12.310000 384.110000 -11.130000 ;
        RECT 382.930000 -13.910000 384.110000 -12.730000 ;
        RECT 562.930000 -12.310000 564.110000 -11.130000 ;
        RECT 562.930000 -13.910000 564.110000 -12.730000 ;
        RECT 742.930000 -12.310000 744.110000 -11.130000 ;
        RECT 742.930000 -13.910000 744.110000 -12.730000 ;
        RECT 922.930000 -12.310000 924.110000 -11.130000 ;
        RECT 922.930000 -13.910000 924.110000 -12.730000 ;
        RECT 1102.930000 -12.310000 1104.110000 -11.130000 ;
        RECT 1102.930000 -13.910000 1104.110000 -12.730000 ;
        RECT 1282.930000 -12.310000 1284.110000 -11.130000 ;
        RECT 1282.930000 -13.910000 1284.110000 -12.730000 ;
        RECT 1462.930000 -12.310000 1464.110000 -11.130000 ;
        RECT 1462.930000 -13.910000 1464.110000 -12.730000 ;
        RECT 1642.930000 -12.310000 1644.110000 -11.130000 ;
        RECT 1642.930000 -13.910000 1644.110000 -12.730000 ;
        RECT 1822.930000 -12.310000 1824.110000 -11.130000 ;
        RECT 1822.930000 -13.910000 1824.110000 -12.730000 ;
        RECT 2002.930000 -12.310000 2004.110000 -11.130000 ;
        RECT 2002.930000 -13.910000 2004.110000 -12.730000 ;
        RECT 2182.930000 -12.310000 2184.110000 -11.130000 ;
        RECT 2182.930000 -13.910000 2184.110000 -12.730000 ;
        RECT 2362.930000 -12.310000 2364.110000 -11.130000 ;
        RECT 2362.930000 -13.910000 2364.110000 -12.730000 ;
        RECT 2542.930000 -12.310000 2544.110000 -11.130000 ;
        RECT 2542.930000 -13.910000 2544.110000 -12.730000 ;
        RECT 2722.930000 -12.310000 2724.110000 -11.130000 ;
        RECT 2722.930000 -13.910000 2724.110000 -12.730000 ;
        RECT 2902.930000 -12.310000 2904.110000 -11.130000 ;
        RECT 2902.930000 -13.910000 2904.110000 -12.730000 ;
        RECT 2936.910000 -12.310000 2938.090000 -11.130000 ;
        RECT 2936.910000 -13.910000 2938.090000 -12.730000 ;
      LAYER met5 ;
        RECT -19.380000 3533.700000 -16.380000 3533.710000 ;
        RECT 22.020000 3533.700000 25.020000 3533.710000 ;
        RECT 202.020000 3533.700000 205.020000 3533.710000 ;
        RECT 382.020000 3533.700000 385.020000 3533.710000 ;
        RECT 562.020000 3533.700000 565.020000 3533.710000 ;
        RECT 742.020000 3533.700000 745.020000 3533.710000 ;
        RECT 922.020000 3533.700000 925.020000 3533.710000 ;
        RECT 1102.020000 3533.700000 1105.020000 3533.710000 ;
        RECT 1282.020000 3533.700000 1285.020000 3533.710000 ;
        RECT 1462.020000 3533.700000 1465.020000 3533.710000 ;
        RECT 1642.020000 3533.700000 1645.020000 3533.710000 ;
        RECT 1822.020000 3533.700000 1825.020000 3533.710000 ;
        RECT 2002.020000 3533.700000 2005.020000 3533.710000 ;
        RECT 2182.020000 3533.700000 2185.020000 3533.710000 ;
        RECT 2362.020000 3533.700000 2365.020000 3533.710000 ;
        RECT 2542.020000 3533.700000 2545.020000 3533.710000 ;
        RECT 2722.020000 3533.700000 2725.020000 3533.710000 ;
        RECT 2902.020000 3533.700000 2905.020000 3533.710000 ;
        RECT 2936.000000 3533.700000 2939.000000 3533.710000 ;
        RECT -19.380000 3530.700000 2939.000000 3533.700000 ;
        RECT -19.380000 3530.690000 -16.380000 3530.700000 ;
        RECT 22.020000 3530.690000 25.020000 3530.700000 ;
        RECT 202.020000 3530.690000 205.020000 3530.700000 ;
        RECT 382.020000 3530.690000 385.020000 3530.700000 ;
        RECT 562.020000 3530.690000 565.020000 3530.700000 ;
        RECT 742.020000 3530.690000 745.020000 3530.700000 ;
        RECT 922.020000 3530.690000 925.020000 3530.700000 ;
        RECT 1102.020000 3530.690000 1105.020000 3530.700000 ;
        RECT 1282.020000 3530.690000 1285.020000 3530.700000 ;
        RECT 1462.020000 3530.690000 1465.020000 3530.700000 ;
        RECT 1642.020000 3530.690000 1645.020000 3530.700000 ;
        RECT 1822.020000 3530.690000 1825.020000 3530.700000 ;
        RECT 2002.020000 3530.690000 2005.020000 3530.700000 ;
        RECT 2182.020000 3530.690000 2185.020000 3530.700000 ;
        RECT 2362.020000 3530.690000 2365.020000 3530.700000 ;
        RECT 2542.020000 3530.690000 2545.020000 3530.700000 ;
        RECT 2722.020000 3530.690000 2725.020000 3530.700000 ;
        RECT 2902.020000 3530.690000 2905.020000 3530.700000 ;
        RECT 2936.000000 3530.690000 2939.000000 3530.700000 ;
        RECT -19.380000 3450.380000 -16.380000 3450.390000 ;
        RECT 2936.000000 3450.380000 2939.000000 3450.390000 ;
        RECT -24.080000 3447.380000 -0.400000 3450.380000 ;
        RECT 2920.400000 3447.380000 2943.700000 3450.380000 ;
        RECT -19.380000 3447.370000 -16.380000 3447.380000 ;
        RECT 2936.000000 3447.370000 2939.000000 3447.380000 ;
        RECT -19.380000 3270.380000 -16.380000 3270.390000 ;
        RECT 2936.000000 3270.380000 2939.000000 3270.390000 ;
        RECT -24.080000 3267.380000 -0.400000 3270.380000 ;
        RECT 2920.400000 3267.380000 2943.700000 3270.380000 ;
        RECT -19.380000 3267.370000 -16.380000 3267.380000 ;
        RECT 2936.000000 3267.370000 2939.000000 3267.380000 ;
        RECT -19.380000 3090.380000 -16.380000 3090.390000 ;
        RECT 2936.000000 3090.380000 2939.000000 3090.390000 ;
        RECT -24.080000 3087.380000 -0.400000 3090.380000 ;
        RECT 2920.400000 3087.380000 2943.700000 3090.380000 ;
        RECT -19.380000 3087.370000 -16.380000 3087.380000 ;
        RECT 2936.000000 3087.370000 2939.000000 3087.380000 ;
        RECT -19.380000 2910.380000 -16.380000 2910.390000 ;
        RECT 2936.000000 2910.380000 2939.000000 2910.390000 ;
        RECT -24.080000 2907.380000 -0.400000 2910.380000 ;
        RECT 2920.400000 2907.380000 2943.700000 2910.380000 ;
        RECT -19.380000 2907.370000 -16.380000 2907.380000 ;
        RECT 2936.000000 2907.370000 2939.000000 2907.380000 ;
        RECT -19.380000 2730.380000 -16.380000 2730.390000 ;
        RECT 2936.000000 2730.380000 2939.000000 2730.390000 ;
        RECT -24.080000 2727.380000 -0.400000 2730.380000 ;
        RECT 2920.400000 2727.380000 2943.700000 2730.380000 ;
        RECT -19.380000 2727.370000 -16.380000 2727.380000 ;
        RECT 2936.000000 2727.370000 2939.000000 2727.380000 ;
        RECT -19.380000 2550.380000 -16.380000 2550.390000 ;
        RECT 2936.000000 2550.380000 2939.000000 2550.390000 ;
        RECT -24.080000 2547.380000 -0.400000 2550.380000 ;
        RECT 2920.400000 2547.380000 2943.700000 2550.380000 ;
        RECT -19.380000 2547.370000 -16.380000 2547.380000 ;
        RECT 2936.000000 2547.370000 2939.000000 2547.380000 ;
        RECT -19.380000 2370.380000 -16.380000 2370.390000 ;
        RECT 2936.000000 2370.380000 2939.000000 2370.390000 ;
        RECT -24.080000 2367.380000 -0.400000 2370.380000 ;
        RECT 2920.400000 2367.380000 2943.700000 2370.380000 ;
        RECT -19.380000 2367.370000 -16.380000 2367.380000 ;
        RECT 2936.000000 2367.370000 2939.000000 2367.380000 ;
        RECT -19.380000 2190.380000 -16.380000 2190.390000 ;
        RECT 2936.000000 2190.380000 2939.000000 2190.390000 ;
        RECT -24.080000 2187.380000 -0.400000 2190.380000 ;
        RECT 2920.400000 2187.380000 2943.700000 2190.380000 ;
        RECT -19.380000 2187.370000 -16.380000 2187.380000 ;
        RECT 2936.000000 2187.370000 2939.000000 2187.380000 ;
        RECT -19.380000 2010.380000 -16.380000 2010.390000 ;
        RECT 2936.000000 2010.380000 2939.000000 2010.390000 ;
        RECT -24.080000 2007.380000 -0.400000 2010.380000 ;
        RECT 2920.400000 2007.380000 2943.700000 2010.380000 ;
        RECT -19.380000 2007.370000 -16.380000 2007.380000 ;
        RECT 2936.000000 2007.370000 2939.000000 2007.380000 ;
        RECT -19.380000 1830.380000 -16.380000 1830.390000 ;
        RECT 2936.000000 1830.380000 2939.000000 1830.390000 ;
        RECT -24.080000 1827.380000 -0.400000 1830.380000 ;
        RECT 2920.400000 1827.380000 2943.700000 1830.380000 ;
        RECT -19.380000 1827.370000 -16.380000 1827.380000 ;
        RECT 2936.000000 1827.370000 2939.000000 1827.380000 ;
        RECT -19.380000 1650.380000 -16.380000 1650.390000 ;
        RECT 2936.000000 1650.380000 2939.000000 1650.390000 ;
        RECT -24.080000 1647.380000 -0.400000 1650.380000 ;
        RECT 2920.400000 1647.380000 2943.700000 1650.380000 ;
        RECT -19.380000 1647.370000 -16.380000 1647.380000 ;
        RECT 2936.000000 1647.370000 2939.000000 1647.380000 ;
        RECT -19.380000 1470.380000 -16.380000 1470.390000 ;
        RECT 2936.000000 1470.380000 2939.000000 1470.390000 ;
        RECT -24.080000 1467.380000 -0.400000 1470.380000 ;
        RECT 2920.400000 1467.380000 2943.700000 1470.380000 ;
        RECT -19.380000 1467.370000 -16.380000 1467.380000 ;
        RECT 2936.000000 1467.370000 2939.000000 1467.380000 ;
        RECT -19.380000 1290.380000 -16.380000 1290.390000 ;
        RECT 2936.000000 1290.380000 2939.000000 1290.390000 ;
        RECT -24.080000 1287.380000 -0.400000 1290.380000 ;
        RECT 2920.400000 1287.380000 2943.700000 1290.380000 ;
        RECT -19.380000 1287.370000 -16.380000 1287.380000 ;
        RECT 2936.000000 1287.370000 2939.000000 1287.380000 ;
        RECT -19.380000 1110.380000 -16.380000 1110.390000 ;
        RECT 2936.000000 1110.380000 2939.000000 1110.390000 ;
        RECT -24.080000 1107.380000 -0.400000 1110.380000 ;
        RECT 2920.400000 1107.380000 2943.700000 1110.380000 ;
        RECT -19.380000 1107.370000 -16.380000 1107.380000 ;
        RECT 2936.000000 1107.370000 2939.000000 1107.380000 ;
        RECT -19.380000 930.380000 -16.380000 930.390000 ;
        RECT 2936.000000 930.380000 2939.000000 930.390000 ;
        RECT -24.080000 927.380000 -0.400000 930.380000 ;
        RECT 2920.400000 927.380000 2943.700000 930.380000 ;
        RECT -19.380000 927.370000 -16.380000 927.380000 ;
        RECT 2936.000000 927.370000 2939.000000 927.380000 ;
        RECT -19.380000 750.380000 -16.380000 750.390000 ;
        RECT 2936.000000 750.380000 2939.000000 750.390000 ;
        RECT -24.080000 747.380000 -0.400000 750.380000 ;
        RECT 2920.400000 747.380000 2943.700000 750.380000 ;
        RECT -19.380000 747.370000 -16.380000 747.380000 ;
        RECT 2936.000000 747.370000 2939.000000 747.380000 ;
        RECT -19.380000 570.380000 -16.380000 570.390000 ;
        RECT 2936.000000 570.380000 2939.000000 570.390000 ;
        RECT -24.080000 567.380000 -0.400000 570.380000 ;
        RECT 2920.400000 567.380000 2943.700000 570.380000 ;
        RECT -19.380000 567.370000 -16.380000 567.380000 ;
        RECT 2936.000000 567.370000 2939.000000 567.380000 ;
        RECT -19.380000 390.380000 -16.380000 390.390000 ;
        RECT 2936.000000 390.380000 2939.000000 390.390000 ;
        RECT -24.080000 387.380000 -0.400000 390.380000 ;
        RECT 2920.400000 387.380000 2943.700000 390.380000 ;
        RECT -19.380000 387.370000 -16.380000 387.380000 ;
        RECT 2936.000000 387.370000 2939.000000 387.380000 ;
        RECT -19.380000 210.380000 -16.380000 210.390000 ;
        RECT 2936.000000 210.380000 2939.000000 210.390000 ;
        RECT -24.080000 207.380000 -0.400000 210.380000 ;
        RECT 2920.400000 207.380000 2943.700000 210.380000 ;
        RECT -19.380000 207.370000 -16.380000 207.380000 ;
        RECT 2936.000000 207.370000 2939.000000 207.380000 ;
        RECT -19.380000 30.380000 -16.380000 30.390000 ;
        RECT 2936.000000 30.380000 2939.000000 30.390000 ;
        RECT -24.080000 27.380000 -0.400000 30.380000 ;
        RECT 2920.400000 27.380000 2943.700000 30.380000 ;
        RECT -19.380000 27.370000 -16.380000 27.380000 ;
        RECT 2936.000000 27.370000 2939.000000 27.380000 ;
        RECT -19.380000 -11.020000 -16.380000 -11.010000 ;
        RECT 22.020000 -11.020000 25.020000 -11.010000 ;
        RECT 202.020000 -11.020000 205.020000 -11.010000 ;
        RECT 382.020000 -11.020000 385.020000 -11.010000 ;
        RECT 562.020000 -11.020000 565.020000 -11.010000 ;
        RECT 742.020000 -11.020000 745.020000 -11.010000 ;
        RECT 922.020000 -11.020000 925.020000 -11.010000 ;
        RECT 1102.020000 -11.020000 1105.020000 -11.010000 ;
        RECT 1282.020000 -11.020000 1285.020000 -11.010000 ;
        RECT 1462.020000 -11.020000 1465.020000 -11.010000 ;
        RECT 1642.020000 -11.020000 1645.020000 -11.010000 ;
        RECT 1822.020000 -11.020000 1825.020000 -11.010000 ;
        RECT 2002.020000 -11.020000 2005.020000 -11.010000 ;
        RECT 2182.020000 -11.020000 2185.020000 -11.010000 ;
        RECT 2362.020000 -11.020000 2365.020000 -11.010000 ;
        RECT 2542.020000 -11.020000 2545.020000 -11.010000 ;
        RECT 2722.020000 -11.020000 2725.020000 -11.010000 ;
        RECT 2902.020000 -11.020000 2905.020000 -11.010000 ;
        RECT 2936.000000 -11.020000 2939.000000 -11.010000 ;
        RECT -19.380000 -14.020000 2939.000000 -11.020000 ;
        RECT -19.380000 -14.030000 -16.380000 -14.020000 ;
        RECT 22.020000 -14.030000 25.020000 -14.020000 ;
        RECT 202.020000 -14.030000 205.020000 -14.020000 ;
        RECT 382.020000 -14.030000 385.020000 -14.020000 ;
        RECT 562.020000 -14.030000 565.020000 -14.020000 ;
        RECT 742.020000 -14.030000 745.020000 -14.020000 ;
        RECT 922.020000 -14.030000 925.020000 -14.020000 ;
        RECT 1102.020000 -14.030000 1105.020000 -14.020000 ;
        RECT 1282.020000 -14.030000 1285.020000 -14.020000 ;
        RECT 1462.020000 -14.030000 1465.020000 -14.020000 ;
        RECT 1642.020000 -14.030000 1645.020000 -14.020000 ;
        RECT 1822.020000 -14.030000 1825.020000 -14.020000 ;
        RECT 2002.020000 -14.030000 2005.020000 -14.020000 ;
        RECT 2182.020000 -14.030000 2185.020000 -14.020000 ;
        RECT 2362.020000 -14.030000 2365.020000 -14.020000 ;
        RECT 2542.020000 -14.030000 2545.020000 -14.020000 ;
        RECT 2722.020000 -14.030000 2725.020000 -14.020000 ;
        RECT 2902.020000 -14.030000 2905.020000 -14.020000 ;
        RECT 2936.000000 -14.030000 2939.000000 -14.020000 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080000 -18.720000 -21.080000 3538.400000 ;
        RECT 112.020000 3520.400000 115.020000 3538.400000 ;
        RECT 292.020000 3520.400000 295.020000 3538.400000 ;
        RECT 472.020000 3520.400000 475.020000 3538.400000 ;
        RECT 652.020000 3520.400000 655.020000 3538.400000 ;
        RECT 832.020000 3520.400000 835.020000 3538.400000 ;
        RECT 1012.020000 3520.400000 1015.020000 3538.400000 ;
        RECT 1192.020000 3520.400000 1195.020000 3538.400000 ;
        RECT 1372.020000 3520.400000 1375.020000 3538.400000 ;
        RECT 1552.020000 3520.400000 1555.020000 3538.400000 ;
        RECT 1732.020000 3520.400000 1735.020000 3538.400000 ;
        RECT 1912.020000 3520.400000 1915.020000 3538.400000 ;
        RECT 2092.020000 3520.400000 2095.020000 3538.400000 ;
        RECT 2272.020000 3520.400000 2275.020000 3538.400000 ;
        RECT 2452.020000 3520.400000 2455.020000 3538.400000 ;
        RECT 2632.020000 3520.400000 2635.020000 3538.400000 ;
        RECT 2812.020000 3520.400000 2815.020000 3538.400000 ;
        RECT 112.020000 -18.720000 115.020000 -0.400000 ;
        RECT 292.020000 -18.720000 295.020000 -0.400000 ;
        RECT 472.020000 -18.720000 475.020000 -0.400000 ;
        RECT 652.020000 -18.720000 655.020000 -0.400000 ;
        RECT 832.020000 -18.720000 835.020000 -0.400000 ;
        RECT 1012.020000 -18.720000 1015.020000 -0.400000 ;
        RECT 1192.020000 -18.720000 1195.020000 -0.400000 ;
        RECT 1372.020000 -18.720000 1375.020000 -0.400000 ;
        RECT 1552.020000 -18.720000 1555.020000 -0.400000 ;
        RECT 1732.020000 -18.720000 1735.020000 -0.400000 ;
        RECT 1912.020000 -18.720000 1915.020000 -0.400000 ;
        RECT 2092.020000 -18.720000 2095.020000 -0.400000 ;
        RECT 2272.020000 -18.720000 2275.020000 -0.400000 ;
        RECT 2452.020000 -18.720000 2455.020000 -0.400000 ;
        RECT 2632.020000 -18.720000 2635.020000 -0.400000 ;
        RECT 2812.020000 -18.720000 2815.020000 -0.400000 ;
        RECT 2940.700000 -18.720000 2943.700000 3538.400000 ;
      LAYER via4 ;
        RECT -23.170000 3537.110000 -21.990000 3538.290000 ;
        RECT -23.170000 3535.510000 -21.990000 3536.690000 ;
        RECT 112.930000 3537.110000 114.110000 3538.290000 ;
        RECT 112.930000 3535.510000 114.110000 3536.690000 ;
        RECT 292.930000 3537.110000 294.110000 3538.290000 ;
        RECT 292.930000 3535.510000 294.110000 3536.690000 ;
        RECT 472.930000 3537.110000 474.110000 3538.290000 ;
        RECT 472.930000 3535.510000 474.110000 3536.690000 ;
        RECT 652.930000 3537.110000 654.110000 3538.290000 ;
        RECT 652.930000 3535.510000 654.110000 3536.690000 ;
        RECT 832.930000 3537.110000 834.110000 3538.290000 ;
        RECT 832.930000 3535.510000 834.110000 3536.690000 ;
        RECT 1012.930000 3537.110000 1014.110000 3538.290000 ;
        RECT 1012.930000 3535.510000 1014.110000 3536.690000 ;
        RECT 1192.930000 3537.110000 1194.110000 3538.290000 ;
        RECT 1192.930000 3535.510000 1194.110000 3536.690000 ;
        RECT 1372.930000 3537.110000 1374.110000 3538.290000 ;
        RECT 1372.930000 3535.510000 1374.110000 3536.690000 ;
        RECT 1552.930000 3537.110000 1554.110000 3538.290000 ;
        RECT 1552.930000 3535.510000 1554.110000 3536.690000 ;
        RECT 1732.930000 3537.110000 1734.110000 3538.290000 ;
        RECT 1732.930000 3535.510000 1734.110000 3536.690000 ;
        RECT 1912.930000 3537.110000 1914.110000 3538.290000 ;
        RECT 1912.930000 3535.510000 1914.110000 3536.690000 ;
        RECT 2092.930000 3537.110000 2094.110000 3538.290000 ;
        RECT 2092.930000 3535.510000 2094.110000 3536.690000 ;
        RECT 2272.930000 3537.110000 2274.110000 3538.290000 ;
        RECT 2272.930000 3535.510000 2274.110000 3536.690000 ;
        RECT 2452.930000 3537.110000 2454.110000 3538.290000 ;
        RECT 2452.930000 3535.510000 2454.110000 3536.690000 ;
        RECT 2632.930000 3537.110000 2634.110000 3538.290000 ;
        RECT 2632.930000 3535.510000 2634.110000 3536.690000 ;
        RECT 2812.930000 3537.110000 2814.110000 3538.290000 ;
        RECT 2812.930000 3535.510000 2814.110000 3536.690000 ;
        RECT 2941.610000 3537.110000 2942.790000 3538.290000 ;
        RECT 2941.610000 3535.510000 2942.790000 3536.690000 ;
        RECT -23.170000 3359.090000 -21.990000 3360.270000 ;
        RECT -23.170000 3357.490000 -21.990000 3358.670000 ;
        RECT -23.170000 3179.090000 -21.990000 3180.270000 ;
        RECT -23.170000 3177.490000 -21.990000 3178.670000 ;
        RECT -23.170000 2999.090000 -21.990000 3000.270000 ;
        RECT -23.170000 2997.490000 -21.990000 2998.670000 ;
        RECT -23.170000 2819.090000 -21.990000 2820.270000 ;
        RECT -23.170000 2817.490000 -21.990000 2818.670000 ;
        RECT -23.170000 2639.090000 -21.990000 2640.270000 ;
        RECT -23.170000 2637.490000 -21.990000 2638.670000 ;
        RECT -23.170000 2459.090000 -21.990000 2460.270000 ;
        RECT -23.170000 2457.490000 -21.990000 2458.670000 ;
        RECT -23.170000 2279.090000 -21.990000 2280.270000 ;
        RECT -23.170000 2277.490000 -21.990000 2278.670000 ;
        RECT -23.170000 2099.090000 -21.990000 2100.270000 ;
        RECT -23.170000 2097.490000 -21.990000 2098.670000 ;
        RECT -23.170000 1919.090000 -21.990000 1920.270000 ;
        RECT -23.170000 1917.490000 -21.990000 1918.670000 ;
        RECT -23.170000 1739.090000 -21.990000 1740.270000 ;
        RECT -23.170000 1737.490000 -21.990000 1738.670000 ;
        RECT -23.170000 1559.090000 -21.990000 1560.270000 ;
        RECT -23.170000 1557.490000 -21.990000 1558.670000 ;
        RECT -23.170000 1379.090000 -21.990000 1380.270000 ;
        RECT -23.170000 1377.490000 -21.990000 1378.670000 ;
        RECT -23.170000 1199.090000 -21.990000 1200.270000 ;
        RECT -23.170000 1197.490000 -21.990000 1198.670000 ;
        RECT -23.170000 1019.090000 -21.990000 1020.270000 ;
        RECT -23.170000 1017.490000 -21.990000 1018.670000 ;
        RECT -23.170000 839.090000 -21.990000 840.270000 ;
        RECT -23.170000 837.490000 -21.990000 838.670000 ;
        RECT -23.170000 659.090000 -21.990000 660.270000 ;
        RECT -23.170000 657.490000 -21.990000 658.670000 ;
        RECT -23.170000 479.090000 -21.990000 480.270000 ;
        RECT -23.170000 477.490000 -21.990000 478.670000 ;
        RECT -23.170000 299.090000 -21.990000 300.270000 ;
        RECT -23.170000 297.490000 -21.990000 298.670000 ;
        RECT -23.170000 119.090000 -21.990000 120.270000 ;
        RECT -23.170000 117.490000 -21.990000 118.670000 ;
        RECT 2941.610000 3359.090000 2942.790000 3360.270000 ;
        RECT 2941.610000 3357.490000 2942.790000 3358.670000 ;
        RECT 2941.610000 3179.090000 2942.790000 3180.270000 ;
        RECT 2941.610000 3177.490000 2942.790000 3178.670000 ;
        RECT 2941.610000 2999.090000 2942.790000 3000.270000 ;
        RECT 2941.610000 2997.490000 2942.790000 2998.670000 ;
        RECT 2941.610000 2819.090000 2942.790000 2820.270000 ;
        RECT 2941.610000 2817.490000 2942.790000 2818.670000 ;
        RECT 2941.610000 2639.090000 2942.790000 2640.270000 ;
        RECT 2941.610000 2637.490000 2942.790000 2638.670000 ;
        RECT 2941.610000 2459.090000 2942.790000 2460.270000 ;
        RECT 2941.610000 2457.490000 2942.790000 2458.670000 ;
        RECT 2941.610000 2279.090000 2942.790000 2280.270000 ;
        RECT 2941.610000 2277.490000 2942.790000 2278.670000 ;
        RECT 2941.610000 2099.090000 2942.790000 2100.270000 ;
        RECT 2941.610000 2097.490000 2942.790000 2098.670000 ;
        RECT 2941.610000 1919.090000 2942.790000 1920.270000 ;
        RECT 2941.610000 1917.490000 2942.790000 1918.670000 ;
        RECT 2941.610000 1739.090000 2942.790000 1740.270000 ;
        RECT 2941.610000 1737.490000 2942.790000 1738.670000 ;
        RECT 2941.610000 1559.090000 2942.790000 1560.270000 ;
        RECT 2941.610000 1557.490000 2942.790000 1558.670000 ;
        RECT 2941.610000 1379.090000 2942.790000 1380.270000 ;
        RECT 2941.610000 1377.490000 2942.790000 1378.670000 ;
        RECT 2941.610000 1199.090000 2942.790000 1200.270000 ;
        RECT 2941.610000 1197.490000 2942.790000 1198.670000 ;
        RECT 2941.610000 1019.090000 2942.790000 1020.270000 ;
        RECT 2941.610000 1017.490000 2942.790000 1018.670000 ;
        RECT 2941.610000 839.090000 2942.790000 840.270000 ;
        RECT 2941.610000 837.490000 2942.790000 838.670000 ;
        RECT 2941.610000 659.090000 2942.790000 660.270000 ;
        RECT 2941.610000 657.490000 2942.790000 658.670000 ;
        RECT 2941.610000 479.090000 2942.790000 480.270000 ;
        RECT 2941.610000 477.490000 2942.790000 478.670000 ;
        RECT 2941.610000 299.090000 2942.790000 300.270000 ;
        RECT 2941.610000 297.490000 2942.790000 298.670000 ;
        RECT 2941.610000 119.090000 2942.790000 120.270000 ;
        RECT 2941.610000 117.490000 2942.790000 118.670000 ;
        RECT -23.170000 -17.010000 -21.990000 -15.830000 ;
        RECT -23.170000 -18.610000 -21.990000 -17.430000 ;
        RECT 112.930000 -17.010000 114.110000 -15.830000 ;
        RECT 112.930000 -18.610000 114.110000 -17.430000 ;
        RECT 292.930000 -17.010000 294.110000 -15.830000 ;
        RECT 292.930000 -18.610000 294.110000 -17.430000 ;
        RECT 472.930000 -17.010000 474.110000 -15.830000 ;
        RECT 472.930000 -18.610000 474.110000 -17.430000 ;
        RECT 652.930000 -17.010000 654.110000 -15.830000 ;
        RECT 652.930000 -18.610000 654.110000 -17.430000 ;
        RECT 832.930000 -17.010000 834.110000 -15.830000 ;
        RECT 832.930000 -18.610000 834.110000 -17.430000 ;
        RECT 1012.930000 -17.010000 1014.110000 -15.830000 ;
        RECT 1012.930000 -18.610000 1014.110000 -17.430000 ;
        RECT 1192.930000 -17.010000 1194.110000 -15.830000 ;
        RECT 1192.930000 -18.610000 1194.110000 -17.430000 ;
        RECT 1372.930000 -17.010000 1374.110000 -15.830000 ;
        RECT 1372.930000 -18.610000 1374.110000 -17.430000 ;
        RECT 1552.930000 -17.010000 1554.110000 -15.830000 ;
        RECT 1552.930000 -18.610000 1554.110000 -17.430000 ;
        RECT 1732.930000 -17.010000 1734.110000 -15.830000 ;
        RECT 1732.930000 -18.610000 1734.110000 -17.430000 ;
        RECT 1912.930000 -17.010000 1914.110000 -15.830000 ;
        RECT 1912.930000 -18.610000 1914.110000 -17.430000 ;
        RECT 2092.930000 -17.010000 2094.110000 -15.830000 ;
        RECT 2092.930000 -18.610000 2094.110000 -17.430000 ;
        RECT 2272.930000 -17.010000 2274.110000 -15.830000 ;
        RECT 2272.930000 -18.610000 2274.110000 -17.430000 ;
        RECT 2452.930000 -17.010000 2454.110000 -15.830000 ;
        RECT 2452.930000 -18.610000 2454.110000 -17.430000 ;
        RECT 2632.930000 -17.010000 2634.110000 -15.830000 ;
        RECT 2632.930000 -18.610000 2634.110000 -17.430000 ;
        RECT 2812.930000 -17.010000 2814.110000 -15.830000 ;
        RECT 2812.930000 -18.610000 2814.110000 -17.430000 ;
        RECT 2941.610000 -17.010000 2942.790000 -15.830000 ;
        RECT 2941.610000 -18.610000 2942.790000 -17.430000 ;
      LAYER met5 ;
        RECT -24.080000 3538.400000 -21.080000 3538.410000 ;
        RECT 112.020000 3538.400000 115.020000 3538.410000 ;
        RECT 292.020000 3538.400000 295.020000 3538.410000 ;
        RECT 472.020000 3538.400000 475.020000 3538.410000 ;
        RECT 652.020000 3538.400000 655.020000 3538.410000 ;
        RECT 832.020000 3538.400000 835.020000 3538.410000 ;
        RECT 1012.020000 3538.400000 1015.020000 3538.410000 ;
        RECT 1192.020000 3538.400000 1195.020000 3538.410000 ;
        RECT 1372.020000 3538.400000 1375.020000 3538.410000 ;
        RECT 1552.020000 3538.400000 1555.020000 3538.410000 ;
        RECT 1732.020000 3538.400000 1735.020000 3538.410000 ;
        RECT 1912.020000 3538.400000 1915.020000 3538.410000 ;
        RECT 2092.020000 3538.400000 2095.020000 3538.410000 ;
        RECT 2272.020000 3538.400000 2275.020000 3538.410000 ;
        RECT 2452.020000 3538.400000 2455.020000 3538.410000 ;
        RECT 2632.020000 3538.400000 2635.020000 3538.410000 ;
        RECT 2812.020000 3538.400000 2815.020000 3538.410000 ;
        RECT 2940.700000 3538.400000 2943.700000 3538.410000 ;
        RECT -24.080000 3535.400000 2943.700000 3538.400000 ;
        RECT -24.080000 3535.390000 -21.080000 3535.400000 ;
        RECT 112.020000 3535.390000 115.020000 3535.400000 ;
        RECT 292.020000 3535.390000 295.020000 3535.400000 ;
        RECT 472.020000 3535.390000 475.020000 3535.400000 ;
        RECT 652.020000 3535.390000 655.020000 3535.400000 ;
        RECT 832.020000 3535.390000 835.020000 3535.400000 ;
        RECT 1012.020000 3535.390000 1015.020000 3535.400000 ;
        RECT 1192.020000 3535.390000 1195.020000 3535.400000 ;
        RECT 1372.020000 3535.390000 1375.020000 3535.400000 ;
        RECT 1552.020000 3535.390000 1555.020000 3535.400000 ;
        RECT 1732.020000 3535.390000 1735.020000 3535.400000 ;
        RECT 1912.020000 3535.390000 1915.020000 3535.400000 ;
        RECT 2092.020000 3535.390000 2095.020000 3535.400000 ;
        RECT 2272.020000 3535.390000 2275.020000 3535.400000 ;
        RECT 2452.020000 3535.390000 2455.020000 3535.400000 ;
        RECT 2632.020000 3535.390000 2635.020000 3535.400000 ;
        RECT 2812.020000 3535.390000 2815.020000 3535.400000 ;
        RECT 2940.700000 3535.390000 2943.700000 3535.400000 ;
        RECT -24.080000 3360.380000 -21.080000 3360.390000 ;
        RECT 2940.700000 3360.380000 2943.700000 3360.390000 ;
        RECT -24.080000 3357.380000 -0.400000 3360.380000 ;
        RECT 2920.400000 3357.380000 2943.700000 3360.380000 ;
        RECT -24.080000 3357.370000 -21.080000 3357.380000 ;
        RECT 2940.700000 3357.370000 2943.700000 3357.380000 ;
        RECT -24.080000 3180.380000 -21.080000 3180.390000 ;
        RECT 2940.700000 3180.380000 2943.700000 3180.390000 ;
        RECT -24.080000 3177.380000 -0.400000 3180.380000 ;
        RECT 2920.400000 3177.380000 2943.700000 3180.380000 ;
        RECT -24.080000 3177.370000 -21.080000 3177.380000 ;
        RECT 2940.700000 3177.370000 2943.700000 3177.380000 ;
        RECT -24.080000 3000.380000 -21.080000 3000.390000 ;
        RECT 2940.700000 3000.380000 2943.700000 3000.390000 ;
        RECT -24.080000 2997.380000 -0.400000 3000.380000 ;
        RECT 2920.400000 2997.380000 2943.700000 3000.380000 ;
        RECT -24.080000 2997.370000 -21.080000 2997.380000 ;
        RECT 2940.700000 2997.370000 2943.700000 2997.380000 ;
        RECT -24.080000 2820.380000 -21.080000 2820.390000 ;
        RECT 2940.700000 2820.380000 2943.700000 2820.390000 ;
        RECT -24.080000 2817.380000 -0.400000 2820.380000 ;
        RECT 2920.400000 2817.380000 2943.700000 2820.380000 ;
        RECT -24.080000 2817.370000 -21.080000 2817.380000 ;
        RECT 2940.700000 2817.370000 2943.700000 2817.380000 ;
        RECT -24.080000 2640.380000 -21.080000 2640.390000 ;
        RECT 2940.700000 2640.380000 2943.700000 2640.390000 ;
        RECT -24.080000 2637.380000 -0.400000 2640.380000 ;
        RECT 2920.400000 2637.380000 2943.700000 2640.380000 ;
        RECT -24.080000 2637.370000 -21.080000 2637.380000 ;
        RECT 2940.700000 2637.370000 2943.700000 2637.380000 ;
        RECT -24.080000 2460.380000 -21.080000 2460.390000 ;
        RECT 2940.700000 2460.380000 2943.700000 2460.390000 ;
        RECT -24.080000 2457.380000 -0.400000 2460.380000 ;
        RECT 2920.400000 2457.380000 2943.700000 2460.380000 ;
        RECT -24.080000 2457.370000 -21.080000 2457.380000 ;
        RECT 2940.700000 2457.370000 2943.700000 2457.380000 ;
        RECT -24.080000 2280.380000 -21.080000 2280.390000 ;
        RECT 2940.700000 2280.380000 2943.700000 2280.390000 ;
        RECT -24.080000 2277.380000 -0.400000 2280.380000 ;
        RECT 2920.400000 2277.380000 2943.700000 2280.380000 ;
        RECT -24.080000 2277.370000 -21.080000 2277.380000 ;
        RECT 2940.700000 2277.370000 2943.700000 2277.380000 ;
        RECT -24.080000 2100.380000 -21.080000 2100.390000 ;
        RECT 2940.700000 2100.380000 2943.700000 2100.390000 ;
        RECT -24.080000 2097.380000 -0.400000 2100.380000 ;
        RECT 2920.400000 2097.380000 2943.700000 2100.380000 ;
        RECT -24.080000 2097.370000 -21.080000 2097.380000 ;
        RECT 2940.700000 2097.370000 2943.700000 2097.380000 ;
        RECT -24.080000 1920.380000 -21.080000 1920.390000 ;
        RECT 2940.700000 1920.380000 2943.700000 1920.390000 ;
        RECT -24.080000 1917.380000 -0.400000 1920.380000 ;
        RECT 2920.400000 1917.380000 2943.700000 1920.380000 ;
        RECT -24.080000 1917.370000 -21.080000 1917.380000 ;
        RECT 2940.700000 1917.370000 2943.700000 1917.380000 ;
        RECT -24.080000 1740.380000 -21.080000 1740.390000 ;
        RECT 2940.700000 1740.380000 2943.700000 1740.390000 ;
        RECT -24.080000 1737.380000 -0.400000 1740.380000 ;
        RECT 2920.400000 1737.380000 2943.700000 1740.380000 ;
        RECT -24.080000 1737.370000 -21.080000 1737.380000 ;
        RECT 2940.700000 1737.370000 2943.700000 1737.380000 ;
        RECT -24.080000 1560.380000 -21.080000 1560.390000 ;
        RECT 2940.700000 1560.380000 2943.700000 1560.390000 ;
        RECT -24.080000 1557.380000 -0.400000 1560.380000 ;
        RECT 2920.400000 1557.380000 2943.700000 1560.380000 ;
        RECT -24.080000 1557.370000 -21.080000 1557.380000 ;
        RECT 2940.700000 1557.370000 2943.700000 1557.380000 ;
        RECT -24.080000 1380.380000 -21.080000 1380.390000 ;
        RECT 2940.700000 1380.380000 2943.700000 1380.390000 ;
        RECT -24.080000 1377.380000 -0.400000 1380.380000 ;
        RECT 2920.400000 1377.380000 2943.700000 1380.380000 ;
        RECT -24.080000 1377.370000 -21.080000 1377.380000 ;
        RECT 2940.700000 1377.370000 2943.700000 1377.380000 ;
        RECT -24.080000 1200.380000 -21.080000 1200.390000 ;
        RECT 2940.700000 1200.380000 2943.700000 1200.390000 ;
        RECT -24.080000 1197.380000 -0.400000 1200.380000 ;
        RECT 2920.400000 1197.380000 2943.700000 1200.380000 ;
        RECT -24.080000 1197.370000 -21.080000 1197.380000 ;
        RECT 2940.700000 1197.370000 2943.700000 1197.380000 ;
        RECT -24.080000 1020.380000 -21.080000 1020.390000 ;
        RECT 2940.700000 1020.380000 2943.700000 1020.390000 ;
        RECT -24.080000 1017.380000 -0.400000 1020.380000 ;
        RECT 2920.400000 1017.380000 2943.700000 1020.380000 ;
        RECT -24.080000 1017.370000 -21.080000 1017.380000 ;
        RECT 2940.700000 1017.370000 2943.700000 1017.380000 ;
        RECT -24.080000 840.380000 -21.080000 840.390000 ;
        RECT 2940.700000 840.380000 2943.700000 840.390000 ;
        RECT -24.080000 837.380000 -0.400000 840.380000 ;
        RECT 2920.400000 837.380000 2943.700000 840.380000 ;
        RECT -24.080000 837.370000 -21.080000 837.380000 ;
        RECT 2940.700000 837.370000 2943.700000 837.380000 ;
        RECT -24.080000 660.380000 -21.080000 660.390000 ;
        RECT 2940.700000 660.380000 2943.700000 660.390000 ;
        RECT -24.080000 657.380000 -0.400000 660.380000 ;
        RECT 2920.400000 657.380000 2943.700000 660.380000 ;
        RECT -24.080000 657.370000 -21.080000 657.380000 ;
        RECT 2940.700000 657.370000 2943.700000 657.380000 ;
        RECT -24.080000 480.380000 -21.080000 480.390000 ;
        RECT 2940.700000 480.380000 2943.700000 480.390000 ;
        RECT -24.080000 477.380000 -0.400000 480.380000 ;
        RECT 2920.400000 477.380000 2943.700000 480.380000 ;
        RECT -24.080000 477.370000 -21.080000 477.380000 ;
        RECT 2940.700000 477.370000 2943.700000 477.380000 ;
        RECT -24.080000 300.380000 -21.080000 300.390000 ;
        RECT 2940.700000 300.380000 2943.700000 300.390000 ;
        RECT -24.080000 297.380000 -0.400000 300.380000 ;
        RECT 2920.400000 297.380000 2943.700000 300.380000 ;
        RECT -24.080000 297.370000 -21.080000 297.380000 ;
        RECT 2940.700000 297.370000 2943.700000 297.380000 ;
        RECT -24.080000 120.380000 -21.080000 120.390000 ;
        RECT 2940.700000 120.380000 2943.700000 120.390000 ;
        RECT -24.080000 117.380000 -0.400000 120.380000 ;
        RECT 2920.400000 117.380000 2943.700000 120.380000 ;
        RECT -24.080000 117.370000 -21.080000 117.380000 ;
        RECT 2940.700000 117.370000 2943.700000 117.380000 ;
        RECT -24.080000 -15.720000 -21.080000 -15.710000 ;
        RECT 112.020000 -15.720000 115.020000 -15.710000 ;
        RECT 292.020000 -15.720000 295.020000 -15.710000 ;
        RECT 472.020000 -15.720000 475.020000 -15.710000 ;
        RECT 652.020000 -15.720000 655.020000 -15.710000 ;
        RECT 832.020000 -15.720000 835.020000 -15.710000 ;
        RECT 1012.020000 -15.720000 1015.020000 -15.710000 ;
        RECT 1192.020000 -15.720000 1195.020000 -15.710000 ;
        RECT 1372.020000 -15.720000 1375.020000 -15.710000 ;
        RECT 1552.020000 -15.720000 1555.020000 -15.710000 ;
        RECT 1732.020000 -15.720000 1735.020000 -15.710000 ;
        RECT 1912.020000 -15.720000 1915.020000 -15.710000 ;
        RECT 2092.020000 -15.720000 2095.020000 -15.710000 ;
        RECT 2272.020000 -15.720000 2275.020000 -15.710000 ;
        RECT 2452.020000 -15.720000 2455.020000 -15.710000 ;
        RECT 2632.020000 -15.720000 2635.020000 -15.710000 ;
        RECT 2812.020000 -15.720000 2815.020000 -15.710000 ;
        RECT 2940.700000 -15.720000 2943.700000 -15.710000 ;
        RECT -24.080000 -18.720000 2943.700000 -15.720000 ;
        RECT -24.080000 -18.730000 -21.080000 -18.720000 ;
        RECT 112.020000 -18.730000 115.020000 -18.720000 ;
        RECT 292.020000 -18.730000 295.020000 -18.720000 ;
        RECT 472.020000 -18.730000 475.020000 -18.720000 ;
        RECT 652.020000 -18.730000 655.020000 -18.720000 ;
        RECT 832.020000 -18.730000 835.020000 -18.720000 ;
        RECT 1012.020000 -18.730000 1015.020000 -18.720000 ;
        RECT 1192.020000 -18.730000 1195.020000 -18.720000 ;
        RECT 1372.020000 -18.730000 1375.020000 -18.720000 ;
        RECT 1552.020000 -18.730000 1555.020000 -18.720000 ;
        RECT 1732.020000 -18.730000 1735.020000 -18.720000 ;
        RECT 1912.020000 -18.730000 1915.020000 -18.720000 ;
        RECT 2092.020000 -18.730000 2095.020000 -18.720000 ;
        RECT 2272.020000 -18.730000 2275.020000 -18.720000 ;
        RECT 2452.020000 -18.730000 2455.020000 -18.720000 ;
        RECT 2632.020000 -18.730000 2635.020000 -18.720000 ;
        RECT 2812.020000 -18.730000 2815.020000 -18.720000 ;
        RECT 2940.700000 -18.730000 2943.700000 -18.720000 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780000 -23.420000 -25.780000 3543.100000 ;
        RECT 40.020000 3520.400000 43.020000 3547.800000 ;
        RECT 220.020000 3520.400000 223.020000 3547.800000 ;
        RECT 400.020000 3520.400000 403.020000 3547.800000 ;
        RECT 580.020000 3520.400000 583.020000 3547.800000 ;
        RECT 760.020000 3520.400000 763.020000 3547.800000 ;
        RECT 940.020000 3520.400000 943.020000 3547.800000 ;
        RECT 1120.020000 3520.400000 1123.020000 3547.800000 ;
        RECT 1300.020000 3520.400000 1303.020000 3547.800000 ;
        RECT 1480.020000 3520.400000 1483.020000 3547.800000 ;
        RECT 1660.020000 3520.400000 1663.020000 3547.800000 ;
        RECT 1840.020000 3520.400000 1843.020000 3547.800000 ;
        RECT 2020.020000 3520.400000 2023.020000 3547.800000 ;
        RECT 2200.020000 3520.400000 2203.020000 3547.800000 ;
        RECT 2380.020000 3520.400000 2383.020000 3547.800000 ;
        RECT 2560.020000 3520.400000 2563.020000 3547.800000 ;
        RECT 2740.020000 3520.400000 2743.020000 3547.800000 ;
        RECT 40.020000 -28.120000 43.020000 -0.400000 ;
        RECT 220.020000 -28.120000 223.020000 -0.400000 ;
        RECT 400.020000 -28.120000 403.020000 -0.400000 ;
        RECT 580.020000 -28.120000 583.020000 -0.400000 ;
        RECT 760.020000 -28.120000 763.020000 -0.400000 ;
        RECT 940.020000 -28.120000 943.020000 -0.400000 ;
        RECT 1120.020000 -28.120000 1123.020000 -0.400000 ;
        RECT 1300.020000 -28.120000 1303.020000 -0.400000 ;
        RECT 1480.020000 -28.120000 1483.020000 -0.400000 ;
        RECT 1660.020000 -28.120000 1663.020000 -0.400000 ;
        RECT 1840.020000 -28.120000 1843.020000 -0.400000 ;
        RECT 2020.020000 -28.120000 2023.020000 -0.400000 ;
        RECT 2200.020000 -28.120000 2203.020000 -0.400000 ;
        RECT 2380.020000 -28.120000 2383.020000 -0.400000 ;
        RECT 2560.020000 -28.120000 2563.020000 -0.400000 ;
        RECT 2740.020000 -28.120000 2743.020000 -0.400000 ;
        RECT 2945.400000 -23.420000 2948.400000 3543.100000 ;
      LAYER via4 ;
        RECT -27.870000 3541.810000 -26.690000 3542.990000 ;
        RECT -27.870000 3540.210000 -26.690000 3541.390000 ;
        RECT 40.930000 3541.810000 42.110000 3542.990000 ;
        RECT 40.930000 3540.210000 42.110000 3541.390000 ;
        RECT 220.930000 3541.810000 222.110000 3542.990000 ;
        RECT 220.930000 3540.210000 222.110000 3541.390000 ;
        RECT 400.930000 3541.810000 402.110000 3542.990000 ;
        RECT 400.930000 3540.210000 402.110000 3541.390000 ;
        RECT 580.930000 3541.810000 582.110000 3542.990000 ;
        RECT 580.930000 3540.210000 582.110000 3541.390000 ;
        RECT 760.930000 3541.810000 762.110000 3542.990000 ;
        RECT 760.930000 3540.210000 762.110000 3541.390000 ;
        RECT 940.930000 3541.810000 942.110000 3542.990000 ;
        RECT 940.930000 3540.210000 942.110000 3541.390000 ;
        RECT 1120.930000 3541.810000 1122.110000 3542.990000 ;
        RECT 1120.930000 3540.210000 1122.110000 3541.390000 ;
        RECT 1300.930000 3541.810000 1302.110000 3542.990000 ;
        RECT 1300.930000 3540.210000 1302.110000 3541.390000 ;
        RECT 1480.930000 3541.810000 1482.110000 3542.990000 ;
        RECT 1480.930000 3540.210000 1482.110000 3541.390000 ;
        RECT 1660.930000 3541.810000 1662.110000 3542.990000 ;
        RECT 1660.930000 3540.210000 1662.110000 3541.390000 ;
        RECT 1840.930000 3541.810000 1842.110000 3542.990000 ;
        RECT 1840.930000 3540.210000 1842.110000 3541.390000 ;
        RECT 2020.930000 3541.810000 2022.110000 3542.990000 ;
        RECT 2020.930000 3540.210000 2022.110000 3541.390000 ;
        RECT 2200.930000 3541.810000 2202.110000 3542.990000 ;
        RECT 2200.930000 3540.210000 2202.110000 3541.390000 ;
        RECT 2380.930000 3541.810000 2382.110000 3542.990000 ;
        RECT 2380.930000 3540.210000 2382.110000 3541.390000 ;
        RECT 2560.930000 3541.810000 2562.110000 3542.990000 ;
        RECT 2560.930000 3540.210000 2562.110000 3541.390000 ;
        RECT 2740.930000 3541.810000 2742.110000 3542.990000 ;
        RECT 2740.930000 3540.210000 2742.110000 3541.390000 ;
        RECT 2946.310000 3541.810000 2947.490000 3542.990000 ;
        RECT 2946.310000 3540.210000 2947.490000 3541.390000 ;
        RECT -27.870000 3467.090000 -26.690000 3468.270000 ;
        RECT -27.870000 3465.490000 -26.690000 3466.670000 ;
        RECT -27.870000 3287.090000 -26.690000 3288.270000 ;
        RECT -27.870000 3285.490000 -26.690000 3286.670000 ;
        RECT -27.870000 3107.090000 -26.690000 3108.270000 ;
        RECT -27.870000 3105.490000 -26.690000 3106.670000 ;
        RECT -27.870000 2927.090000 -26.690000 2928.270000 ;
        RECT -27.870000 2925.490000 -26.690000 2926.670000 ;
        RECT -27.870000 2747.090000 -26.690000 2748.270000 ;
        RECT -27.870000 2745.490000 -26.690000 2746.670000 ;
        RECT -27.870000 2567.090000 -26.690000 2568.270000 ;
        RECT -27.870000 2565.490000 -26.690000 2566.670000 ;
        RECT -27.870000 2387.090000 -26.690000 2388.270000 ;
        RECT -27.870000 2385.490000 -26.690000 2386.670000 ;
        RECT -27.870000 2207.090000 -26.690000 2208.270000 ;
        RECT -27.870000 2205.490000 -26.690000 2206.670000 ;
        RECT -27.870000 2027.090000 -26.690000 2028.270000 ;
        RECT -27.870000 2025.490000 -26.690000 2026.670000 ;
        RECT -27.870000 1847.090000 -26.690000 1848.270000 ;
        RECT -27.870000 1845.490000 -26.690000 1846.670000 ;
        RECT -27.870000 1667.090000 -26.690000 1668.270000 ;
        RECT -27.870000 1665.490000 -26.690000 1666.670000 ;
        RECT -27.870000 1487.090000 -26.690000 1488.270000 ;
        RECT -27.870000 1485.490000 -26.690000 1486.670000 ;
        RECT -27.870000 1307.090000 -26.690000 1308.270000 ;
        RECT -27.870000 1305.490000 -26.690000 1306.670000 ;
        RECT -27.870000 1127.090000 -26.690000 1128.270000 ;
        RECT -27.870000 1125.490000 -26.690000 1126.670000 ;
        RECT -27.870000 947.090000 -26.690000 948.270000 ;
        RECT -27.870000 945.490000 -26.690000 946.670000 ;
        RECT -27.870000 767.090000 -26.690000 768.270000 ;
        RECT -27.870000 765.490000 -26.690000 766.670000 ;
        RECT -27.870000 587.090000 -26.690000 588.270000 ;
        RECT -27.870000 585.490000 -26.690000 586.670000 ;
        RECT -27.870000 407.090000 -26.690000 408.270000 ;
        RECT -27.870000 405.490000 -26.690000 406.670000 ;
        RECT -27.870000 227.090000 -26.690000 228.270000 ;
        RECT -27.870000 225.490000 -26.690000 226.670000 ;
        RECT -27.870000 47.090000 -26.690000 48.270000 ;
        RECT -27.870000 45.490000 -26.690000 46.670000 ;
        RECT 2946.310000 3467.090000 2947.490000 3468.270000 ;
        RECT 2946.310000 3465.490000 2947.490000 3466.670000 ;
        RECT 2946.310000 3287.090000 2947.490000 3288.270000 ;
        RECT 2946.310000 3285.490000 2947.490000 3286.670000 ;
        RECT 2946.310000 3107.090000 2947.490000 3108.270000 ;
        RECT 2946.310000 3105.490000 2947.490000 3106.670000 ;
        RECT 2946.310000 2927.090000 2947.490000 2928.270000 ;
        RECT 2946.310000 2925.490000 2947.490000 2926.670000 ;
        RECT 2946.310000 2747.090000 2947.490000 2748.270000 ;
        RECT 2946.310000 2745.490000 2947.490000 2746.670000 ;
        RECT 2946.310000 2567.090000 2947.490000 2568.270000 ;
        RECT 2946.310000 2565.490000 2947.490000 2566.670000 ;
        RECT 2946.310000 2387.090000 2947.490000 2388.270000 ;
        RECT 2946.310000 2385.490000 2947.490000 2386.670000 ;
        RECT 2946.310000 2207.090000 2947.490000 2208.270000 ;
        RECT 2946.310000 2205.490000 2947.490000 2206.670000 ;
        RECT 2946.310000 2027.090000 2947.490000 2028.270000 ;
        RECT 2946.310000 2025.490000 2947.490000 2026.670000 ;
        RECT 2946.310000 1847.090000 2947.490000 1848.270000 ;
        RECT 2946.310000 1845.490000 2947.490000 1846.670000 ;
        RECT 2946.310000 1667.090000 2947.490000 1668.270000 ;
        RECT 2946.310000 1665.490000 2947.490000 1666.670000 ;
        RECT 2946.310000 1487.090000 2947.490000 1488.270000 ;
        RECT 2946.310000 1485.490000 2947.490000 1486.670000 ;
        RECT 2946.310000 1307.090000 2947.490000 1308.270000 ;
        RECT 2946.310000 1305.490000 2947.490000 1306.670000 ;
        RECT 2946.310000 1127.090000 2947.490000 1128.270000 ;
        RECT 2946.310000 1125.490000 2947.490000 1126.670000 ;
        RECT 2946.310000 947.090000 2947.490000 948.270000 ;
        RECT 2946.310000 945.490000 2947.490000 946.670000 ;
        RECT 2946.310000 767.090000 2947.490000 768.270000 ;
        RECT 2946.310000 765.490000 2947.490000 766.670000 ;
        RECT 2946.310000 587.090000 2947.490000 588.270000 ;
        RECT 2946.310000 585.490000 2947.490000 586.670000 ;
        RECT 2946.310000 407.090000 2947.490000 408.270000 ;
        RECT 2946.310000 405.490000 2947.490000 406.670000 ;
        RECT 2946.310000 227.090000 2947.490000 228.270000 ;
        RECT 2946.310000 225.490000 2947.490000 226.670000 ;
        RECT 2946.310000 47.090000 2947.490000 48.270000 ;
        RECT 2946.310000 45.490000 2947.490000 46.670000 ;
        RECT -27.870000 -21.710000 -26.690000 -20.530000 ;
        RECT -27.870000 -23.310000 -26.690000 -22.130000 ;
        RECT 40.930000 -21.710000 42.110000 -20.530000 ;
        RECT 40.930000 -23.310000 42.110000 -22.130000 ;
        RECT 220.930000 -21.710000 222.110000 -20.530000 ;
        RECT 220.930000 -23.310000 222.110000 -22.130000 ;
        RECT 400.930000 -21.710000 402.110000 -20.530000 ;
        RECT 400.930000 -23.310000 402.110000 -22.130000 ;
        RECT 580.930000 -21.710000 582.110000 -20.530000 ;
        RECT 580.930000 -23.310000 582.110000 -22.130000 ;
        RECT 760.930000 -21.710000 762.110000 -20.530000 ;
        RECT 760.930000 -23.310000 762.110000 -22.130000 ;
        RECT 940.930000 -21.710000 942.110000 -20.530000 ;
        RECT 940.930000 -23.310000 942.110000 -22.130000 ;
        RECT 1120.930000 -21.710000 1122.110000 -20.530000 ;
        RECT 1120.930000 -23.310000 1122.110000 -22.130000 ;
        RECT 1300.930000 -21.710000 1302.110000 -20.530000 ;
        RECT 1300.930000 -23.310000 1302.110000 -22.130000 ;
        RECT 1480.930000 -21.710000 1482.110000 -20.530000 ;
        RECT 1480.930000 -23.310000 1482.110000 -22.130000 ;
        RECT 1660.930000 -21.710000 1662.110000 -20.530000 ;
        RECT 1660.930000 -23.310000 1662.110000 -22.130000 ;
        RECT 1840.930000 -21.710000 1842.110000 -20.530000 ;
        RECT 1840.930000 -23.310000 1842.110000 -22.130000 ;
        RECT 2020.930000 -21.710000 2022.110000 -20.530000 ;
        RECT 2020.930000 -23.310000 2022.110000 -22.130000 ;
        RECT 2200.930000 -21.710000 2202.110000 -20.530000 ;
        RECT 2200.930000 -23.310000 2202.110000 -22.130000 ;
        RECT 2380.930000 -21.710000 2382.110000 -20.530000 ;
        RECT 2380.930000 -23.310000 2382.110000 -22.130000 ;
        RECT 2560.930000 -21.710000 2562.110000 -20.530000 ;
        RECT 2560.930000 -23.310000 2562.110000 -22.130000 ;
        RECT 2740.930000 -21.710000 2742.110000 -20.530000 ;
        RECT 2740.930000 -23.310000 2742.110000 -22.130000 ;
        RECT 2946.310000 -21.710000 2947.490000 -20.530000 ;
        RECT 2946.310000 -23.310000 2947.490000 -22.130000 ;
      LAYER met5 ;
        RECT -28.780000 3543.100000 -25.780000 3543.110000 ;
        RECT 40.020000 3543.100000 43.020000 3543.110000 ;
        RECT 220.020000 3543.100000 223.020000 3543.110000 ;
        RECT 400.020000 3543.100000 403.020000 3543.110000 ;
        RECT 580.020000 3543.100000 583.020000 3543.110000 ;
        RECT 760.020000 3543.100000 763.020000 3543.110000 ;
        RECT 940.020000 3543.100000 943.020000 3543.110000 ;
        RECT 1120.020000 3543.100000 1123.020000 3543.110000 ;
        RECT 1300.020000 3543.100000 1303.020000 3543.110000 ;
        RECT 1480.020000 3543.100000 1483.020000 3543.110000 ;
        RECT 1660.020000 3543.100000 1663.020000 3543.110000 ;
        RECT 1840.020000 3543.100000 1843.020000 3543.110000 ;
        RECT 2020.020000 3543.100000 2023.020000 3543.110000 ;
        RECT 2200.020000 3543.100000 2203.020000 3543.110000 ;
        RECT 2380.020000 3543.100000 2383.020000 3543.110000 ;
        RECT 2560.020000 3543.100000 2563.020000 3543.110000 ;
        RECT 2740.020000 3543.100000 2743.020000 3543.110000 ;
        RECT 2945.400000 3543.100000 2948.400000 3543.110000 ;
        RECT -28.780000 3540.100000 2948.400000 3543.100000 ;
        RECT -28.780000 3540.090000 -25.780000 3540.100000 ;
        RECT 40.020000 3540.090000 43.020000 3540.100000 ;
        RECT 220.020000 3540.090000 223.020000 3540.100000 ;
        RECT 400.020000 3540.090000 403.020000 3540.100000 ;
        RECT 580.020000 3540.090000 583.020000 3540.100000 ;
        RECT 760.020000 3540.090000 763.020000 3540.100000 ;
        RECT 940.020000 3540.090000 943.020000 3540.100000 ;
        RECT 1120.020000 3540.090000 1123.020000 3540.100000 ;
        RECT 1300.020000 3540.090000 1303.020000 3540.100000 ;
        RECT 1480.020000 3540.090000 1483.020000 3540.100000 ;
        RECT 1660.020000 3540.090000 1663.020000 3540.100000 ;
        RECT 1840.020000 3540.090000 1843.020000 3540.100000 ;
        RECT 2020.020000 3540.090000 2023.020000 3540.100000 ;
        RECT 2200.020000 3540.090000 2203.020000 3540.100000 ;
        RECT 2380.020000 3540.090000 2383.020000 3540.100000 ;
        RECT 2560.020000 3540.090000 2563.020000 3540.100000 ;
        RECT 2740.020000 3540.090000 2743.020000 3540.100000 ;
        RECT 2945.400000 3540.090000 2948.400000 3540.100000 ;
        RECT -28.780000 3468.380000 -25.780000 3468.390000 ;
        RECT 2945.400000 3468.380000 2948.400000 3468.390000 ;
        RECT -33.480000 3465.380000 -0.400000 3468.380000 ;
        RECT 2920.400000 3465.380000 2953.100000 3468.380000 ;
        RECT -28.780000 3465.370000 -25.780000 3465.380000 ;
        RECT 2945.400000 3465.370000 2948.400000 3465.380000 ;
        RECT -28.780000 3288.380000 -25.780000 3288.390000 ;
        RECT 2945.400000 3288.380000 2948.400000 3288.390000 ;
        RECT -33.480000 3285.380000 -0.400000 3288.380000 ;
        RECT 2920.400000 3285.380000 2953.100000 3288.380000 ;
        RECT -28.780000 3285.370000 -25.780000 3285.380000 ;
        RECT 2945.400000 3285.370000 2948.400000 3285.380000 ;
        RECT -28.780000 3108.380000 -25.780000 3108.390000 ;
        RECT 2945.400000 3108.380000 2948.400000 3108.390000 ;
        RECT -33.480000 3105.380000 -0.400000 3108.380000 ;
        RECT 2920.400000 3105.380000 2953.100000 3108.380000 ;
        RECT -28.780000 3105.370000 -25.780000 3105.380000 ;
        RECT 2945.400000 3105.370000 2948.400000 3105.380000 ;
        RECT -28.780000 2928.380000 -25.780000 2928.390000 ;
        RECT 2945.400000 2928.380000 2948.400000 2928.390000 ;
        RECT -33.480000 2925.380000 -0.400000 2928.380000 ;
        RECT 2920.400000 2925.380000 2953.100000 2928.380000 ;
        RECT -28.780000 2925.370000 -25.780000 2925.380000 ;
        RECT 2945.400000 2925.370000 2948.400000 2925.380000 ;
        RECT -28.780000 2748.380000 -25.780000 2748.390000 ;
        RECT 2945.400000 2748.380000 2948.400000 2748.390000 ;
        RECT -33.480000 2745.380000 -0.400000 2748.380000 ;
        RECT 2920.400000 2745.380000 2953.100000 2748.380000 ;
        RECT -28.780000 2745.370000 -25.780000 2745.380000 ;
        RECT 2945.400000 2745.370000 2948.400000 2745.380000 ;
        RECT -28.780000 2568.380000 -25.780000 2568.390000 ;
        RECT 2945.400000 2568.380000 2948.400000 2568.390000 ;
        RECT -33.480000 2565.380000 -0.400000 2568.380000 ;
        RECT 2920.400000 2565.380000 2953.100000 2568.380000 ;
        RECT -28.780000 2565.370000 -25.780000 2565.380000 ;
        RECT 2945.400000 2565.370000 2948.400000 2565.380000 ;
        RECT -28.780000 2388.380000 -25.780000 2388.390000 ;
        RECT 2945.400000 2388.380000 2948.400000 2388.390000 ;
        RECT -33.480000 2385.380000 -0.400000 2388.380000 ;
        RECT 2920.400000 2385.380000 2953.100000 2388.380000 ;
        RECT -28.780000 2385.370000 -25.780000 2385.380000 ;
        RECT 2945.400000 2385.370000 2948.400000 2385.380000 ;
        RECT -28.780000 2208.380000 -25.780000 2208.390000 ;
        RECT 2945.400000 2208.380000 2948.400000 2208.390000 ;
        RECT -33.480000 2205.380000 -0.400000 2208.380000 ;
        RECT 2920.400000 2205.380000 2953.100000 2208.380000 ;
        RECT -28.780000 2205.370000 -25.780000 2205.380000 ;
        RECT 2945.400000 2205.370000 2948.400000 2205.380000 ;
        RECT -28.780000 2028.380000 -25.780000 2028.390000 ;
        RECT 2945.400000 2028.380000 2948.400000 2028.390000 ;
        RECT -33.480000 2025.380000 -0.400000 2028.380000 ;
        RECT 2920.400000 2025.380000 2953.100000 2028.380000 ;
        RECT -28.780000 2025.370000 -25.780000 2025.380000 ;
        RECT 2945.400000 2025.370000 2948.400000 2025.380000 ;
        RECT -28.780000 1848.380000 -25.780000 1848.390000 ;
        RECT 2945.400000 1848.380000 2948.400000 1848.390000 ;
        RECT -33.480000 1845.380000 -0.400000 1848.380000 ;
        RECT 2920.400000 1845.380000 2953.100000 1848.380000 ;
        RECT -28.780000 1845.370000 -25.780000 1845.380000 ;
        RECT 2945.400000 1845.370000 2948.400000 1845.380000 ;
        RECT -28.780000 1668.380000 -25.780000 1668.390000 ;
        RECT 2945.400000 1668.380000 2948.400000 1668.390000 ;
        RECT -33.480000 1665.380000 -0.400000 1668.380000 ;
        RECT 2920.400000 1665.380000 2953.100000 1668.380000 ;
        RECT -28.780000 1665.370000 -25.780000 1665.380000 ;
        RECT 2945.400000 1665.370000 2948.400000 1665.380000 ;
        RECT -28.780000 1488.380000 -25.780000 1488.390000 ;
        RECT 2945.400000 1488.380000 2948.400000 1488.390000 ;
        RECT -33.480000 1485.380000 -0.400000 1488.380000 ;
        RECT 2920.400000 1485.380000 2953.100000 1488.380000 ;
        RECT -28.780000 1485.370000 -25.780000 1485.380000 ;
        RECT 2945.400000 1485.370000 2948.400000 1485.380000 ;
        RECT -28.780000 1308.380000 -25.780000 1308.390000 ;
        RECT 2945.400000 1308.380000 2948.400000 1308.390000 ;
        RECT -33.480000 1305.380000 -0.400000 1308.380000 ;
        RECT 2920.400000 1305.380000 2953.100000 1308.380000 ;
        RECT -28.780000 1305.370000 -25.780000 1305.380000 ;
        RECT 2945.400000 1305.370000 2948.400000 1305.380000 ;
        RECT -28.780000 1128.380000 -25.780000 1128.390000 ;
        RECT 2945.400000 1128.380000 2948.400000 1128.390000 ;
        RECT -33.480000 1125.380000 -0.400000 1128.380000 ;
        RECT 2920.400000 1125.380000 2953.100000 1128.380000 ;
        RECT -28.780000 1125.370000 -25.780000 1125.380000 ;
        RECT 2945.400000 1125.370000 2948.400000 1125.380000 ;
        RECT -28.780000 948.380000 -25.780000 948.390000 ;
        RECT 2945.400000 948.380000 2948.400000 948.390000 ;
        RECT -33.480000 945.380000 -0.400000 948.380000 ;
        RECT 2920.400000 945.380000 2953.100000 948.380000 ;
        RECT -28.780000 945.370000 -25.780000 945.380000 ;
        RECT 2945.400000 945.370000 2948.400000 945.380000 ;
        RECT -28.780000 768.380000 -25.780000 768.390000 ;
        RECT 2945.400000 768.380000 2948.400000 768.390000 ;
        RECT -33.480000 765.380000 -0.400000 768.380000 ;
        RECT 2920.400000 765.380000 2953.100000 768.380000 ;
        RECT -28.780000 765.370000 -25.780000 765.380000 ;
        RECT 2945.400000 765.370000 2948.400000 765.380000 ;
        RECT -28.780000 588.380000 -25.780000 588.390000 ;
        RECT 2945.400000 588.380000 2948.400000 588.390000 ;
        RECT -33.480000 585.380000 -0.400000 588.380000 ;
        RECT 2920.400000 585.380000 2953.100000 588.380000 ;
        RECT -28.780000 585.370000 -25.780000 585.380000 ;
        RECT 2945.400000 585.370000 2948.400000 585.380000 ;
        RECT -28.780000 408.380000 -25.780000 408.390000 ;
        RECT 2945.400000 408.380000 2948.400000 408.390000 ;
        RECT -33.480000 405.380000 -0.400000 408.380000 ;
        RECT 2920.400000 405.380000 2953.100000 408.380000 ;
        RECT -28.780000 405.370000 -25.780000 405.380000 ;
        RECT 2945.400000 405.370000 2948.400000 405.380000 ;
        RECT -28.780000 228.380000 -25.780000 228.390000 ;
        RECT 2945.400000 228.380000 2948.400000 228.390000 ;
        RECT -33.480000 225.380000 -0.400000 228.380000 ;
        RECT 2920.400000 225.380000 2953.100000 228.380000 ;
        RECT -28.780000 225.370000 -25.780000 225.380000 ;
        RECT 2945.400000 225.370000 2948.400000 225.380000 ;
        RECT -28.780000 48.380000 -25.780000 48.390000 ;
        RECT 2945.400000 48.380000 2948.400000 48.390000 ;
        RECT -33.480000 45.380000 -0.400000 48.380000 ;
        RECT 2920.400000 45.380000 2953.100000 48.380000 ;
        RECT -28.780000 45.370000 -25.780000 45.380000 ;
        RECT 2945.400000 45.370000 2948.400000 45.380000 ;
        RECT -28.780000 -20.420000 -25.780000 -20.410000 ;
        RECT 40.020000 -20.420000 43.020000 -20.410000 ;
        RECT 220.020000 -20.420000 223.020000 -20.410000 ;
        RECT 400.020000 -20.420000 403.020000 -20.410000 ;
        RECT 580.020000 -20.420000 583.020000 -20.410000 ;
        RECT 760.020000 -20.420000 763.020000 -20.410000 ;
        RECT 940.020000 -20.420000 943.020000 -20.410000 ;
        RECT 1120.020000 -20.420000 1123.020000 -20.410000 ;
        RECT 1300.020000 -20.420000 1303.020000 -20.410000 ;
        RECT 1480.020000 -20.420000 1483.020000 -20.410000 ;
        RECT 1660.020000 -20.420000 1663.020000 -20.410000 ;
        RECT 1840.020000 -20.420000 1843.020000 -20.410000 ;
        RECT 2020.020000 -20.420000 2023.020000 -20.410000 ;
        RECT 2200.020000 -20.420000 2203.020000 -20.410000 ;
        RECT 2380.020000 -20.420000 2383.020000 -20.410000 ;
        RECT 2560.020000 -20.420000 2563.020000 -20.410000 ;
        RECT 2740.020000 -20.420000 2743.020000 -20.410000 ;
        RECT 2945.400000 -20.420000 2948.400000 -20.410000 ;
        RECT -28.780000 -23.420000 2948.400000 -20.420000 ;
        RECT -28.780000 -23.430000 -25.780000 -23.420000 ;
        RECT 40.020000 -23.430000 43.020000 -23.420000 ;
        RECT 220.020000 -23.430000 223.020000 -23.420000 ;
        RECT 400.020000 -23.430000 403.020000 -23.420000 ;
        RECT 580.020000 -23.430000 583.020000 -23.420000 ;
        RECT 760.020000 -23.430000 763.020000 -23.420000 ;
        RECT 940.020000 -23.430000 943.020000 -23.420000 ;
        RECT 1120.020000 -23.430000 1123.020000 -23.420000 ;
        RECT 1300.020000 -23.430000 1303.020000 -23.420000 ;
        RECT 1480.020000 -23.430000 1483.020000 -23.420000 ;
        RECT 1660.020000 -23.430000 1663.020000 -23.420000 ;
        RECT 1840.020000 -23.430000 1843.020000 -23.420000 ;
        RECT 2020.020000 -23.430000 2023.020000 -23.420000 ;
        RECT 2200.020000 -23.430000 2203.020000 -23.420000 ;
        RECT 2380.020000 -23.430000 2383.020000 -23.420000 ;
        RECT 2560.020000 -23.430000 2563.020000 -23.420000 ;
        RECT 2740.020000 -23.430000 2743.020000 -23.420000 ;
        RECT 2945.400000 -23.430000 2948.400000 -23.420000 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480000 -28.120000 -30.480000 3547.800000 ;
        RECT 130.020000 3520.400000 133.020000 3547.800000 ;
        RECT 310.020000 3520.400000 313.020000 3547.800000 ;
        RECT 490.020000 3520.400000 493.020000 3547.800000 ;
        RECT 670.020000 3520.400000 673.020000 3547.800000 ;
        RECT 850.020000 3520.400000 853.020000 3547.800000 ;
        RECT 1030.020000 3520.400000 1033.020000 3547.800000 ;
        RECT 1210.020000 3520.400000 1213.020000 3547.800000 ;
        RECT 1390.020000 3520.400000 1393.020000 3547.800000 ;
        RECT 1570.020000 3520.400000 1573.020000 3547.800000 ;
        RECT 1750.020000 3520.400000 1753.020000 3547.800000 ;
        RECT 1930.020000 3520.400000 1933.020000 3547.800000 ;
        RECT 2110.020000 3520.400000 2113.020000 3547.800000 ;
        RECT 2290.020000 3520.400000 2293.020000 3547.800000 ;
        RECT 2470.020000 3520.400000 2473.020000 3547.800000 ;
        RECT 2650.020000 3520.400000 2653.020000 3547.800000 ;
        RECT 2830.020000 3520.400000 2833.020000 3547.800000 ;
        RECT 130.020000 -28.120000 133.020000 -0.400000 ;
        RECT 310.020000 -28.120000 313.020000 -0.400000 ;
        RECT 490.020000 -28.120000 493.020000 -0.400000 ;
        RECT 670.020000 -28.120000 673.020000 -0.400000 ;
        RECT 850.020000 -28.120000 853.020000 -0.400000 ;
        RECT 1030.020000 -28.120000 1033.020000 -0.400000 ;
        RECT 1210.020000 -28.120000 1213.020000 -0.400000 ;
        RECT 1390.020000 -28.120000 1393.020000 -0.400000 ;
        RECT 1570.020000 -28.120000 1573.020000 -0.400000 ;
        RECT 1750.020000 -28.120000 1753.020000 -0.400000 ;
        RECT 1930.020000 -28.120000 1933.020000 -0.400000 ;
        RECT 2110.020000 -28.120000 2113.020000 -0.400000 ;
        RECT 2290.020000 -28.120000 2293.020000 -0.400000 ;
        RECT 2470.020000 -28.120000 2473.020000 -0.400000 ;
        RECT 2650.020000 -28.120000 2653.020000 -0.400000 ;
        RECT 2830.020000 -28.120000 2833.020000 -0.400000 ;
        RECT 2950.100000 -28.120000 2953.100000 3547.800000 ;
      LAYER via4 ;
        RECT -32.570000 3546.510000 -31.390000 3547.690000 ;
        RECT -32.570000 3544.910000 -31.390000 3546.090000 ;
        RECT 130.930000 3546.510000 132.110000 3547.690000 ;
        RECT 130.930000 3544.910000 132.110000 3546.090000 ;
        RECT 310.930000 3546.510000 312.110000 3547.690000 ;
        RECT 310.930000 3544.910000 312.110000 3546.090000 ;
        RECT 490.930000 3546.510000 492.110000 3547.690000 ;
        RECT 490.930000 3544.910000 492.110000 3546.090000 ;
        RECT 670.930000 3546.510000 672.110000 3547.690000 ;
        RECT 670.930000 3544.910000 672.110000 3546.090000 ;
        RECT 850.930000 3546.510000 852.110000 3547.690000 ;
        RECT 850.930000 3544.910000 852.110000 3546.090000 ;
        RECT 1030.930000 3546.510000 1032.110000 3547.690000 ;
        RECT 1030.930000 3544.910000 1032.110000 3546.090000 ;
        RECT 1210.930000 3546.510000 1212.110000 3547.690000 ;
        RECT 1210.930000 3544.910000 1212.110000 3546.090000 ;
        RECT 1390.930000 3546.510000 1392.110000 3547.690000 ;
        RECT 1390.930000 3544.910000 1392.110000 3546.090000 ;
        RECT 1570.930000 3546.510000 1572.110000 3547.690000 ;
        RECT 1570.930000 3544.910000 1572.110000 3546.090000 ;
        RECT 1750.930000 3546.510000 1752.110000 3547.690000 ;
        RECT 1750.930000 3544.910000 1752.110000 3546.090000 ;
        RECT 1930.930000 3546.510000 1932.110000 3547.690000 ;
        RECT 1930.930000 3544.910000 1932.110000 3546.090000 ;
        RECT 2110.930000 3546.510000 2112.110000 3547.690000 ;
        RECT 2110.930000 3544.910000 2112.110000 3546.090000 ;
        RECT 2290.930000 3546.510000 2292.110000 3547.690000 ;
        RECT 2290.930000 3544.910000 2292.110000 3546.090000 ;
        RECT 2470.930000 3546.510000 2472.110000 3547.690000 ;
        RECT 2470.930000 3544.910000 2472.110000 3546.090000 ;
        RECT 2650.930000 3546.510000 2652.110000 3547.690000 ;
        RECT 2650.930000 3544.910000 2652.110000 3546.090000 ;
        RECT 2830.930000 3546.510000 2832.110000 3547.690000 ;
        RECT 2830.930000 3544.910000 2832.110000 3546.090000 ;
        RECT 2951.010000 3546.510000 2952.190000 3547.690000 ;
        RECT 2951.010000 3544.910000 2952.190000 3546.090000 ;
        RECT -32.570000 3377.090000 -31.390000 3378.270000 ;
        RECT -32.570000 3375.490000 -31.390000 3376.670000 ;
        RECT -32.570000 3197.090000 -31.390000 3198.270000 ;
        RECT -32.570000 3195.490000 -31.390000 3196.670000 ;
        RECT -32.570000 3017.090000 -31.390000 3018.270000 ;
        RECT -32.570000 3015.490000 -31.390000 3016.670000 ;
        RECT -32.570000 2837.090000 -31.390000 2838.270000 ;
        RECT -32.570000 2835.490000 -31.390000 2836.670000 ;
        RECT -32.570000 2657.090000 -31.390000 2658.270000 ;
        RECT -32.570000 2655.490000 -31.390000 2656.670000 ;
        RECT -32.570000 2477.090000 -31.390000 2478.270000 ;
        RECT -32.570000 2475.490000 -31.390000 2476.670000 ;
        RECT -32.570000 2297.090000 -31.390000 2298.270000 ;
        RECT -32.570000 2295.490000 -31.390000 2296.670000 ;
        RECT -32.570000 2117.090000 -31.390000 2118.270000 ;
        RECT -32.570000 2115.490000 -31.390000 2116.670000 ;
        RECT -32.570000 1937.090000 -31.390000 1938.270000 ;
        RECT -32.570000 1935.490000 -31.390000 1936.670000 ;
        RECT -32.570000 1757.090000 -31.390000 1758.270000 ;
        RECT -32.570000 1755.490000 -31.390000 1756.670000 ;
        RECT -32.570000 1577.090000 -31.390000 1578.270000 ;
        RECT -32.570000 1575.490000 -31.390000 1576.670000 ;
        RECT -32.570000 1397.090000 -31.390000 1398.270000 ;
        RECT -32.570000 1395.490000 -31.390000 1396.670000 ;
        RECT -32.570000 1217.090000 -31.390000 1218.270000 ;
        RECT -32.570000 1215.490000 -31.390000 1216.670000 ;
        RECT -32.570000 1037.090000 -31.390000 1038.270000 ;
        RECT -32.570000 1035.490000 -31.390000 1036.670000 ;
        RECT -32.570000 857.090000 -31.390000 858.270000 ;
        RECT -32.570000 855.490000 -31.390000 856.670000 ;
        RECT -32.570000 677.090000 -31.390000 678.270000 ;
        RECT -32.570000 675.490000 -31.390000 676.670000 ;
        RECT -32.570000 497.090000 -31.390000 498.270000 ;
        RECT -32.570000 495.490000 -31.390000 496.670000 ;
        RECT -32.570000 317.090000 -31.390000 318.270000 ;
        RECT -32.570000 315.490000 -31.390000 316.670000 ;
        RECT -32.570000 137.090000 -31.390000 138.270000 ;
        RECT -32.570000 135.490000 -31.390000 136.670000 ;
        RECT 2951.010000 3377.090000 2952.190000 3378.270000 ;
        RECT 2951.010000 3375.490000 2952.190000 3376.670000 ;
        RECT 2951.010000 3197.090000 2952.190000 3198.270000 ;
        RECT 2951.010000 3195.490000 2952.190000 3196.670000 ;
        RECT 2951.010000 3017.090000 2952.190000 3018.270000 ;
        RECT 2951.010000 3015.490000 2952.190000 3016.670000 ;
        RECT 2951.010000 2837.090000 2952.190000 2838.270000 ;
        RECT 2951.010000 2835.490000 2952.190000 2836.670000 ;
        RECT 2951.010000 2657.090000 2952.190000 2658.270000 ;
        RECT 2951.010000 2655.490000 2952.190000 2656.670000 ;
        RECT 2951.010000 2477.090000 2952.190000 2478.270000 ;
        RECT 2951.010000 2475.490000 2952.190000 2476.670000 ;
        RECT 2951.010000 2297.090000 2952.190000 2298.270000 ;
        RECT 2951.010000 2295.490000 2952.190000 2296.670000 ;
        RECT 2951.010000 2117.090000 2952.190000 2118.270000 ;
        RECT 2951.010000 2115.490000 2952.190000 2116.670000 ;
        RECT 2951.010000 1937.090000 2952.190000 1938.270000 ;
        RECT 2951.010000 1935.490000 2952.190000 1936.670000 ;
        RECT 2951.010000 1757.090000 2952.190000 1758.270000 ;
        RECT 2951.010000 1755.490000 2952.190000 1756.670000 ;
        RECT 2951.010000 1577.090000 2952.190000 1578.270000 ;
        RECT 2951.010000 1575.490000 2952.190000 1576.670000 ;
        RECT 2951.010000 1397.090000 2952.190000 1398.270000 ;
        RECT 2951.010000 1395.490000 2952.190000 1396.670000 ;
        RECT 2951.010000 1217.090000 2952.190000 1218.270000 ;
        RECT 2951.010000 1215.490000 2952.190000 1216.670000 ;
        RECT 2951.010000 1037.090000 2952.190000 1038.270000 ;
        RECT 2951.010000 1035.490000 2952.190000 1036.670000 ;
        RECT 2951.010000 857.090000 2952.190000 858.270000 ;
        RECT 2951.010000 855.490000 2952.190000 856.670000 ;
        RECT 2951.010000 677.090000 2952.190000 678.270000 ;
        RECT 2951.010000 675.490000 2952.190000 676.670000 ;
        RECT 2951.010000 497.090000 2952.190000 498.270000 ;
        RECT 2951.010000 495.490000 2952.190000 496.670000 ;
        RECT 2951.010000 317.090000 2952.190000 318.270000 ;
        RECT 2951.010000 315.490000 2952.190000 316.670000 ;
        RECT 2951.010000 137.090000 2952.190000 138.270000 ;
        RECT 2951.010000 135.490000 2952.190000 136.670000 ;
        RECT -32.570000 -26.410000 -31.390000 -25.230000 ;
        RECT -32.570000 -28.010000 -31.390000 -26.830000 ;
        RECT 130.930000 -26.410000 132.110000 -25.230000 ;
        RECT 130.930000 -28.010000 132.110000 -26.830000 ;
        RECT 310.930000 -26.410000 312.110000 -25.230000 ;
        RECT 310.930000 -28.010000 312.110000 -26.830000 ;
        RECT 490.930000 -26.410000 492.110000 -25.230000 ;
        RECT 490.930000 -28.010000 492.110000 -26.830000 ;
        RECT 670.930000 -26.410000 672.110000 -25.230000 ;
        RECT 670.930000 -28.010000 672.110000 -26.830000 ;
        RECT 850.930000 -26.410000 852.110000 -25.230000 ;
        RECT 850.930000 -28.010000 852.110000 -26.830000 ;
        RECT 1030.930000 -26.410000 1032.110000 -25.230000 ;
        RECT 1030.930000 -28.010000 1032.110000 -26.830000 ;
        RECT 1210.930000 -26.410000 1212.110000 -25.230000 ;
        RECT 1210.930000 -28.010000 1212.110000 -26.830000 ;
        RECT 1390.930000 -26.410000 1392.110000 -25.230000 ;
        RECT 1390.930000 -28.010000 1392.110000 -26.830000 ;
        RECT 1570.930000 -26.410000 1572.110000 -25.230000 ;
        RECT 1570.930000 -28.010000 1572.110000 -26.830000 ;
        RECT 1750.930000 -26.410000 1752.110000 -25.230000 ;
        RECT 1750.930000 -28.010000 1752.110000 -26.830000 ;
        RECT 1930.930000 -26.410000 1932.110000 -25.230000 ;
        RECT 1930.930000 -28.010000 1932.110000 -26.830000 ;
        RECT 2110.930000 -26.410000 2112.110000 -25.230000 ;
        RECT 2110.930000 -28.010000 2112.110000 -26.830000 ;
        RECT 2290.930000 -26.410000 2292.110000 -25.230000 ;
        RECT 2290.930000 -28.010000 2292.110000 -26.830000 ;
        RECT 2470.930000 -26.410000 2472.110000 -25.230000 ;
        RECT 2470.930000 -28.010000 2472.110000 -26.830000 ;
        RECT 2650.930000 -26.410000 2652.110000 -25.230000 ;
        RECT 2650.930000 -28.010000 2652.110000 -26.830000 ;
        RECT 2830.930000 -26.410000 2832.110000 -25.230000 ;
        RECT 2830.930000 -28.010000 2832.110000 -26.830000 ;
        RECT 2951.010000 -26.410000 2952.190000 -25.230000 ;
        RECT 2951.010000 -28.010000 2952.190000 -26.830000 ;
      LAYER met5 ;
        RECT -33.480000 3547.800000 -30.480000 3547.810000 ;
        RECT 130.020000 3547.800000 133.020000 3547.810000 ;
        RECT 310.020000 3547.800000 313.020000 3547.810000 ;
        RECT 490.020000 3547.800000 493.020000 3547.810000 ;
        RECT 670.020000 3547.800000 673.020000 3547.810000 ;
        RECT 850.020000 3547.800000 853.020000 3547.810000 ;
        RECT 1030.020000 3547.800000 1033.020000 3547.810000 ;
        RECT 1210.020000 3547.800000 1213.020000 3547.810000 ;
        RECT 1390.020000 3547.800000 1393.020000 3547.810000 ;
        RECT 1570.020000 3547.800000 1573.020000 3547.810000 ;
        RECT 1750.020000 3547.800000 1753.020000 3547.810000 ;
        RECT 1930.020000 3547.800000 1933.020000 3547.810000 ;
        RECT 2110.020000 3547.800000 2113.020000 3547.810000 ;
        RECT 2290.020000 3547.800000 2293.020000 3547.810000 ;
        RECT 2470.020000 3547.800000 2473.020000 3547.810000 ;
        RECT 2650.020000 3547.800000 2653.020000 3547.810000 ;
        RECT 2830.020000 3547.800000 2833.020000 3547.810000 ;
        RECT 2950.100000 3547.800000 2953.100000 3547.810000 ;
        RECT -33.480000 3544.800000 2953.100000 3547.800000 ;
        RECT -33.480000 3544.790000 -30.480000 3544.800000 ;
        RECT 130.020000 3544.790000 133.020000 3544.800000 ;
        RECT 310.020000 3544.790000 313.020000 3544.800000 ;
        RECT 490.020000 3544.790000 493.020000 3544.800000 ;
        RECT 670.020000 3544.790000 673.020000 3544.800000 ;
        RECT 850.020000 3544.790000 853.020000 3544.800000 ;
        RECT 1030.020000 3544.790000 1033.020000 3544.800000 ;
        RECT 1210.020000 3544.790000 1213.020000 3544.800000 ;
        RECT 1390.020000 3544.790000 1393.020000 3544.800000 ;
        RECT 1570.020000 3544.790000 1573.020000 3544.800000 ;
        RECT 1750.020000 3544.790000 1753.020000 3544.800000 ;
        RECT 1930.020000 3544.790000 1933.020000 3544.800000 ;
        RECT 2110.020000 3544.790000 2113.020000 3544.800000 ;
        RECT 2290.020000 3544.790000 2293.020000 3544.800000 ;
        RECT 2470.020000 3544.790000 2473.020000 3544.800000 ;
        RECT 2650.020000 3544.790000 2653.020000 3544.800000 ;
        RECT 2830.020000 3544.790000 2833.020000 3544.800000 ;
        RECT 2950.100000 3544.790000 2953.100000 3544.800000 ;
        RECT -33.480000 3378.380000 -30.480000 3378.390000 ;
        RECT 2950.100000 3378.380000 2953.100000 3378.390000 ;
        RECT -33.480000 3375.380000 -0.400000 3378.380000 ;
        RECT 2920.400000 3375.380000 2953.100000 3378.380000 ;
        RECT -33.480000 3375.370000 -30.480000 3375.380000 ;
        RECT 2950.100000 3375.370000 2953.100000 3375.380000 ;
        RECT -33.480000 3198.380000 -30.480000 3198.390000 ;
        RECT 2950.100000 3198.380000 2953.100000 3198.390000 ;
        RECT -33.480000 3195.380000 -0.400000 3198.380000 ;
        RECT 2920.400000 3195.380000 2953.100000 3198.380000 ;
        RECT -33.480000 3195.370000 -30.480000 3195.380000 ;
        RECT 2950.100000 3195.370000 2953.100000 3195.380000 ;
        RECT -33.480000 3018.380000 -30.480000 3018.390000 ;
        RECT 2950.100000 3018.380000 2953.100000 3018.390000 ;
        RECT -33.480000 3015.380000 -0.400000 3018.380000 ;
        RECT 2920.400000 3015.380000 2953.100000 3018.380000 ;
        RECT -33.480000 3015.370000 -30.480000 3015.380000 ;
        RECT 2950.100000 3015.370000 2953.100000 3015.380000 ;
        RECT -33.480000 2838.380000 -30.480000 2838.390000 ;
        RECT 2950.100000 2838.380000 2953.100000 2838.390000 ;
        RECT -33.480000 2835.380000 -0.400000 2838.380000 ;
        RECT 2920.400000 2835.380000 2953.100000 2838.380000 ;
        RECT -33.480000 2835.370000 -30.480000 2835.380000 ;
        RECT 2950.100000 2835.370000 2953.100000 2835.380000 ;
        RECT -33.480000 2658.380000 -30.480000 2658.390000 ;
        RECT 2950.100000 2658.380000 2953.100000 2658.390000 ;
        RECT -33.480000 2655.380000 -0.400000 2658.380000 ;
        RECT 2920.400000 2655.380000 2953.100000 2658.380000 ;
        RECT -33.480000 2655.370000 -30.480000 2655.380000 ;
        RECT 2950.100000 2655.370000 2953.100000 2655.380000 ;
        RECT -33.480000 2478.380000 -30.480000 2478.390000 ;
        RECT 2950.100000 2478.380000 2953.100000 2478.390000 ;
        RECT -33.480000 2475.380000 -0.400000 2478.380000 ;
        RECT 2920.400000 2475.380000 2953.100000 2478.380000 ;
        RECT -33.480000 2475.370000 -30.480000 2475.380000 ;
        RECT 2950.100000 2475.370000 2953.100000 2475.380000 ;
        RECT -33.480000 2298.380000 -30.480000 2298.390000 ;
        RECT 2950.100000 2298.380000 2953.100000 2298.390000 ;
        RECT -33.480000 2295.380000 -0.400000 2298.380000 ;
        RECT 2920.400000 2295.380000 2953.100000 2298.380000 ;
        RECT -33.480000 2295.370000 -30.480000 2295.380000 ;
        RECT 2950.100000 2295.370000 2953.100000 2295.380000 ;
        RECT -33.480000 2118.380000 -30.480000 2118.390000 ;
        RECT 2950.100000 2118.380000 2953.100000 2118.390000 ;
        RECT -33.480000 2115.380000 -0.400000 2118.380000 ;
        RECT 2920.400000 2115.380000 2953.100000 2118.380000 ;
        RECT -33.480000 2115.370000 -30.480000 2115.380000 ;
        RECT 2950.100000 2115.370000 2953.100000 2115.380000 ;
        RECT -33.480000 1938.380000 -30.480000 1938.390000 ;
        RECT 2950.100000 1938.380000 2953.100000 1938.390000 ;
        RECT -33.480000 1935.380000 -0.400000 1938.380000 ;
        RECT 2920.400000 1935.380000 2953.100000 1938.380000 ;
        RECT -33.480000 1935.370000 -30.480000 1935.380000 ;
        RECT 2950.100000 1935.370000 2953.100000 1935.380000 ;
        RECT -33.480000 1758.380000 -30.480000 1758.390000 ;
        RECT 2950.100000 1758.380000 2953.100000 1758.390000 ;
        RECT -33.480000 1755.380000 -0.400000 1758.380000 ;
        RECT 2920.400000 1755.380000 2953.100000 1758.380000 ;
        RECT -33.480000 1755.370000 -30.480000 1755.380000 ;
        RECT 2950.100000 1755.370000 2953.100000 1755.380000 ;
        RECT -33.480000 1578.380000 -30.480000 1578.390000 ;
        RECT 2950.100000 1578.380000 2953.100000 1578.390000 ;
        RECT -33.480000 1575.380000 -0.400000 1578.380000 ;
        RECT 2920.400000 1575.380000 2953.100000 1578.380000 ;
        RECT -33.480000 1575.370000 -30.480000 1575.380000 ;
        RECT 2950.100000 1575.370000 2953.100000 1575.380000 ;
        RECT -33.480000 1398.380000 -30.480000 1398.390000 ;
        RECT 2950.100000 1398.380000 2953.100000 1398.390000 ;
        RECT -33.480000 1395.380000 -0.400000 1398.380000 ;
        RECT 2920.400000 1395.380000 2953.100000 1398.380000 ;
        RECT -33.480000 1395.370000 -30.480000 1395.380000 ;
        RECT 2950.100000 1395.370000 2953.100000 1395.380000 ;
        RECT -33.480000 1218.380000 -30.480000 1218.390000 ;
        RECT 2950.100000 1218.380000 2953.100000 1218.390000 ;
        RECT -33.480000 1215.380000 -0.400000 1218.380000 ;
        RECT 2920.400000 1215.380000 2953.100000 1218.380000 ;
        RECT -33.480000 1215.370000 -30.480000 1215.380000 ;
        RECT 2950.100000 1215.370000 2953.100000 1215.380000 ;
        RECT -33.480000 1038.380000 -30.480000 1038.390000 ;
        RECT 2950.100000 1038.380000 2953.100000 1038.390000 ;
        RECT -33.480000 1035.380000 -0.400000 1038.380000 ;
        RECT 2920.400000 1035.380000 2953.100000 1038.380000 ;
        RECT -33.480000 1035.370000 -30.480000 1035.380000 ;
        RECT 2950.100000 1035.370000 2953.100000 1035.380000 ;
        RECT -33.480000 858.380000 -30.480000 858.390000 ;
        RECT 2950.100000 858.380000 2953.100000 858.390000 ;
        RECT -33.480000 855.380000 -0.400000 858.380000 ;
        RECT 2920.400000 855.380000 2953.100000 858.380000 ;
        RECT -33.480000 855.370000 -30.480000 855.380000 ;
        RECT 2950.100000 855.370000 2953.100000 855.380000 ;
        RECT -33.480000 678.380000 -30.480000 678.390000 ;
        RECT 2950.100000 678.380000 2953.100000 678.390000 ;
        RECT -33.480000 675.380000 -0.400000 678.380000 ;
        RECT 2920.400000 675.380000 2953.100000 678.380000 ;
        RECT -33.480000 675.370000 -30.480000 675.380000 ;
        RECT 2950.100000 675.370000 2953.100000 675.380000 ;
        RECT -33.480000 498.380000 -30.480000 498.390000 ;
        RECT 2950.100000 498.380000 2953.100000 498.390000 ;
        RECT -33.480000 495.380000 -0.400000 498.380000 ;
        RECT 2920.400000 495.380000 2953.100000 498.380000 ;
        RECT -33.480000 495.370000 -30.480000 495.380000 ;
        RECT 2950.100000 495.370000 2953.100000 495.380000 ;
        RECT -33.480000 318.380000 -30.480000 318.390000 ;
        RECT 2950.100000 318.380000 2953.100000 318.390000 ;
        RECT -33.480000 315.380000 -0.400000 318.380000 ;
        RECT 2920.400000 315.380000 2953.100000 318.380000 ;
        RECT -33.480000 315.370000 -30.480000 315.380000 ;
        RECT 2950.100000 315.370000 2953.100000 315.380000 ;
        RECT -33.480000 138.380000 -30.480000 138.390000 ;
        RECT 2950.100000 138.380000 2953.100000 138.390000 ;
        RECT -33.480000 135.380000 -0.400000 138.380000 ;
        RECT 2920.400000 135.380000 2953.100000 138.380000 ;
        RECT -33.480000 135.370000 -30.480000 135.380000 ;
        RECT 2950.100000 135.370000 2953.100000 135.380000 ;
        RECT -33.480000 -25.120000 -30.480000 -25.110000 ;
        RECT 130.020000 -25.120000 133.020000 -25.110000 ;
        RECT 310.020000 -25.120000 313.020000 -25.110000 ;
        RECT 490.020000 -25.120000 493.020000 -25.110000 ;
        RECT 670.020000 -25.120000 673.020000 -25.110000 ;
        RECT 850.020000 -25.120000 853.020000 -25.110000 ;
        RECT 1030.020000 -25.120000 1033.020000 -25.110000 ;
        RECT 1210.020000 -25.120000 1213.020000 -25.110000 ;
        RECT 1390.020000 -25.120000 1393.020000 -25.110000 ;
        RECT 1570.020000 -25.120000 1573.020000 -25.110000 ;
        RECT 1750.020000 -25.120000 1753.020000 -25.110000 ;
        RECT 1930.020000 -25.120000 1933.020000 -25.110000 ;
        RECT 2110.020000 -25.120000 2113.020000 -25.110000 ;
        RECT 2290.020000 -25.120000 2293.020000 -25.110000 ;
        RECT 2470.020000 -25.120000 2473.020000 -25.110000 ;
        RECT 2650.020000 -25.120000 2653.020000 -25.110000 ;
        RECT 2830.020000 -25.120000 2833.020000 -25.110000 ;
        RECT 2950.100000 -25.120000 2953.100000 -25.110000 ;
        RECT -33.480000 -28.120000 2953.100000 -25.120000 ;
        RECT -33.480000 -28.130000 -30.480000 -28.120000 ;
        RECT 130.020000 -28.130000 133.020000 -28.120000 ;
        RECT 310.020000 -28.130000 313.020000 -28.120000 ;
        RECT 490.020000 -28.130000 493.020000 -28.120000 ;
        RECT 670.020000 -28.130000 673.020000 -28.120000 ;
        RECT 850.020000 -28.130000 853.020000 -28.120000 ;
        RECT 1030.020000 -28.130000 1033.020000 -28.120000 ;
        RECT 1210.020000 -28.130000 1213.020000 -28.120000 ;
        RECT 1390.020000 -28.130000 1393.020000 -28.120000 ;
        RECT 1570.020000 -28.130000 1573.020000 -28.120000 ;
        RECT 1750.020000 -28.130000 1753.020000 -28.120000 ;
        RECT 1930.020000 -28.130000 1933.020000 -28.120000 ;
        RECT 2110.020000 -28.130000 2113.020000 -28.120000 ;
        RECT 2290.020000 -28.130000 2293.020000 -28.120000 ;
        RECT 2470.020000 -28.130000 2473.020000 -28.120000 ;
        RECT 2650.020000 -28.130000 2653.020000 -28.120000 ;
        RECT 2830.020000 -28.130000 2833.020000 -28.120000 ;
        RECT 2950.100000 -28.130000 2953.100000 -28.120000 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180000 -32.820000 -35.180000 3552.500000 ;
        RECT 58.020000 3520.400000 61.020000 3557.200000 ;
        RECT 238.020000 3520.400000 241.020000 3557.200000 ;
        RECT 418.020000 3520.400000 421.020000 3557.200000 ;
        RECT 598.020000 3520.400000 601.020000 3557.200000 ;
        RECT 778.020000 3520.400000 781.020000 3557.200000 ;
        RECT 958.020000 3520.400000 961.020000 3557.200000 ;
        RECT 1138.020000 3520.400000 1141.020000 3557.200000 ;
        RECT 1318.020000 3520.400000 1321.020000 3557.200000 ;
        RECT 1498.020000 3520.400000 1501.020000 3557.200000 ;
        RECT 1678.020000 3520.400000 1681.020000 3557.200000 ;
        RECT 1858.020000 3520.400000 1861.020000 3557.200000 ;
        RECT 2038.020000 3520.400000 2041.020000 3557.200000 ;
        RECT 2218.020000 3520.400000 2221.020000 3557.200000 ;
        RECT 2398.020000 3520.400000 2401.020000 3557.200000 ;
        RECT 2578.020000 3520.400000 2581.020000 3557.200000 ;
        RECT 2758.020000 3520.400000 2761.020000 3557.200000 ;
        RECT 58.020000 -37.520000 61.020000 -0.400000 ;
        RECT 238.020000 -37.520000 241.020000 -0.400000 ;
        RECT 418.020000 -37.520000 421.020000 -0.400000 ;
        RECT 598.020000 -37.520000 601.020000 -0.400000 ;
        RECT 778.020000 -37.520000 781.020000 -0.400000 ;
        RECT 958.020000 -37.520000 961.020000 -0.400000 ;
        RECT 1138.020000 -37.520000 1141.020000 -0.400000 ;
        RECT 1318.020000 -37.520000 1321.020000 -0.400000 ;
        RECT 1498.020000 -37.520000 1501.020000 -0.400000 ;
        RECT 1678.020000 -37.520000 1681.020000 -0.400000 ;
        RECT 1858.020000 -37.520000 1861.020000 -0.400000 ;
        RECT 2038.020000 -37.520000 2041.020000 -0.400000 ;
        RECT 2218.020000 -37.520000 2221.020000 -0.400000 ;
        RECT 2398.020000 -37.520000 2401.020000 -0.400000 ;
        RECT 2578.020000 -37.520000 2581.020000 -0.400000 ;
        RECT 2758.020000 -37.520000 2761.020000 -0.400000 ;
        RECT 2954.800000 -32.820000 2957.800000 3552.500000 ;
      LAYER via4 ;
        RECT -37.270000 3551.210000 -36.090000 3552.390000 ;
        RECT -37.270000 3549.610000 -36.090000 3550.790000 ;
        RECT 58.930000 3551.210000 60.110000 3552.390000 ;
        RECT 58.930000 3549.610000 60.110000 3550.790000 ;
        RECT 238.930000 3551.210000 240.110000 3552.390000 ;
        RECT 238.930000 3549.610000 240.110000 3550.790000 ;
        RECT 418.930000 3551.210000 420.110000 3552.390000 ;
        RECT 418.930000 3549.610000 420.110000 3550.790000 ;
        RECT 598.930000 3551.210000 600.110000 3552.390000 ;
        RECT 598.930000 3549.610000 600.110000 3550.790000 ;
        RECT 778.930000 3551.210000 780.110000 3552.390000 ;
        RECT 778.930000 3549.610000 780.110000 3550.790000 ;
        RECT 958.930000 3551.210000 960.110000 3552.390000 ;
        RECT 958.930000 3549.610000 960.110000 3550.790000 ;
        RECT 1138.930000 3551.210000 1140.110000 3552.390000 ;
        RECT 1138.930000 3549.610000 1140.110000 3550.790000 ;
        RECT 1318.930000 3551.210000 1320.110000 3552.390000 ;
        RECT 1318.930000 3549.610000 1320.110000 3550.790000 ;
        RECT 1498.930000 3551.210000 1500.110000 3552.390000 ;
        RECT 1498.930000 3549.610000 1500.110000 3550.790000 ;
        RECT 1678.930000 3551.210000 1680.110000 3552.390000 ;
        RECT 1678.930000 3549.610000 1680.110000 3550.790000 ;
        RECT 1858.930000 3551.210000 1860.110000 3552.390000 ;
        RECT 1858.930000 3549.610000 1860.110000 3550.790000 ;
        RECT 2038.930000 3551.210000 2040.110000 3552.390000 ;
        RECT 2038.930000 3549.610000 2040.110000 3550.790000 ;
        RECT 2218.930000 3551.210000 2220.110000 3552.390000 ;
        RECT 2218.930000 3549.610000 2220.110000 3550.790000 ;
        RECT 2398.930000 3551.210000 2400.110000 3552.390000 ;
        RECT 2398.930000 3549.610000 2400.110000 3550.790000 ;
        RECT 2578.930000 3551.210000 2580.110000 3552.390000 ;
        RECT 2578.930000 3549.610000 2580.110000 3550.790000 ;
        RECT 2758.930000 3551.210000 2760.110000 3552.390000 ;
        RECT 2758.930000 3549.610000 2760.110000 3550.790000 ;
        RECT 2955.710000 3551.210000 2956.890000 3552.390000 ;
        RECT 2955.710000 3549.610000 2956.890000 3550.790000 ;
        RECT -37.270000 3485.090000 -36.090000 3486.270000 ;
        RECT -37.270000 3483.490000 -36.090000 3484.670000 ;
        RECT -37.270000 3305.090000 -36.090000 3306.270000 ;
        RECT -37.270000 3303.490000 -36.090000 3304.670000 ;
        RECT -37.270000 3125.090000 -36.090000 3126.270000 ;
        RECT -37.270000 3123.490000 -36.090000 3124.670000 ;
        RECT -37.270000 2945.090000 -36.090000 2946.270000 ;
        RECT -37.270000 2943.490000 -36.090000 2944.670000 ;
        RECT -37.270000 2765.090000 -36.090000 2766.270000 ;
        RECT -37.270000 2763.490000 -36.090000 2764.670000 ;
        RECT -37.270000 2585.090000 -36.090000 2586.270000 ;
        RECT -37.270000 2583.490000 -36.090000 2584.670000 ;
        RECT -37.270000 2405.090000 -36.090000 2406.270000 ;
        RECT -37.270000 2403.490000 -36.090000 2404.670000 ;
        RECT -37.270000 2225.090000 -36.090000 2226.270000 ;
        RECT -37.270000 2223.490000 -36.090000 2224.670000 ;
        RECT -37.270000 2045.090000 -36.090000 2046.270000 ;
        RECT -37.270000 2043.490000 -36.090000 2044.670000 ;
        RECT -37.270000 1865.090000 -36.090000 1866.270000 ;
        RECT -37.270000 1863.490000 -36.090000 1864.670000 ;
        RECT -37.270000 1685.090000 -36.090000 1686.270000 ;
        RECT -37.270000 1683.490000 -36.090000 1684.670000 ;
        RECT -37.270000 1505.090000 -36.090000 1506.270000 ;
        RECT -37.270000 1503.490000 -36.090000 1504.670000 ;
        RECT -37.270000 1325.090000 -36.090000 1326.270000 ;
        RECT -37.270000 1323.490000 -36.090000 1324.670000 ;
        RECT -37.270000 1145.090000 -36.090000 1146.270000 ;
        RECT -37.270000 1143.490000 -36.090000 1144.670000 ;
        RECT -37.270000 965.090000 -36.090000 966.270000 ;
        RECT -37.270000 963.490000 -36.090000 964.670000 ;
        RECT -37.270000 785.090000 -36.090000 786.270000 ;
        RECT -37.270000 783.490000 -36.090000 784.670000 ;
        RECT -37.270000 605.090000 -36.090000 606.270000 ;
        RECT -37.270000 603.490000 -36.090000 604.670000 ;
        RECT -37.270000 425.090000 -36.090000 426.270000 ;
        RECT -37.270000 423.490000 -36.090000 424.670000 ;
        RECT -37.270000 245.090000 -36.090000 246.270000 ;
        RECT -37.270000 243.490000 -36.090000 244.670000 ;
        RECT -37.270000 65.090000 -36.090000 66.270000 ;
        RECT -37.270000 63.490000 -36.090000 64.670000 ;
        RECT 2955.710000 3485.090000 2956.890000 3486.270000 ;
        RECT 2955.710000 3483.490000 2956.890000 3484.670000 ;
        RECT 2955.710000 3305.090000 2956.890000 3306.270000 ;
        RECT 2955.710000 3303.490000 2956.890000 3304.670000 ;
        RECT 2955.710000 3125.090000 2956.890000 3126.270000 ;
        RECT 2955.710000 3123.490000 2956.890000 3124.670000 ;
        RECT 2955.710000 2945.090000 2956.890000 2946.270000 ;
        RECT 2955.710000 2943.490000 2956.890000 2944.670000 ;
        RECT 2955.710000 2765.090000 2956.890000 2766.270000 ;
        RECT 2955.710000 2763.490000 2956.890000 2764.670000 ;
        RECT 2955.710000 2585.090000 2956.890000 2586.270000 ;
        RECT 2955.710000 2583.490000 2956.890000 2584.670000 ;
        RECT 2955.710000 2405.090000 2956.890000 2406.270000 ;
        RECT 2955.710000 2403.490000 2956.890000 2404.670000 ;
        RECT 2955.710000 2225.090000 2956.890000 2226.270000 ;
        RECT 2955.710000 2223.490000 2956.890000 2224.670000 ;
        RECT 2955.710000 2045.090000 2956.890000 2046.270000 ;
        RECT 2955.710000 2043.490000 2956.890000 2044.670000 ;
        RECT 2955.710000 1865.090000 2956.890000 1866.270000 ;
        RECT 2955.710000 1863.490000 2956.890000 1864.670000 ;
        RECT 2955.710000 1685.090000 2956.890000 1686.270000 ;
        RECT 2955.710000 1683.490000 2956.890000 1684.670000 ;
        RECT 2955.710000 1505.090000 2956.890000 1506.270000 ;
        RECT 2955.710000 1503.490000 2956.890000 1504.670000 ;
        RECT 2955.710000 1325.090000 2956.890000 1326.270000 ;
        RECT 2955.710000 1323.490000 2956.890000 1324.670000 ;
        RECT 2955.710000 1145.090000 2956.890000 1146.270000 ;
        RECT 2955.710000 1143.490000 2956.890000 1144.670000 ;
        RECT 2955.710000 965.090000 2956.890000 966.270000 ;
        RECT 2955.710000 963.490000 2956.890000 964.670000 ;
        RECT 2955.710000 785.090000 2956.890000 786.270000 ;
        RECT 2955.710000 783.490000 2956.890000 784.670000 ;
        RECT 2955.710000 605.090000 2956.890000 606.270000 ;
        RECT 2955.710000 603.490000 2956.890000 604.670000 ;
        RECT 2955.710000 425.090000 2956.890000 426.270000 ;
        RECT 2955.710000 423.490000 2956.890000 424.670000 ;
        RECT 2955.710000 245.090000 2956.890000 246.270000 ;
        RECT 2955.710000 243.490000 2956.890000 244.670000 ;
        RECT 2955.710000 65.090000 2956.890000 66.270000 ;
        RECT 2955.710000 63.490000 2956.890000 64.670000 ;
        RECT -37.270000 -31.110000 -36.090000 -29.930000 ;
        RECT -37.270000 -32.710000 -36.090000 -31.530000 ;
        RECT 58.930000 -31.110000 60.110000 -29.930000 ;
        RECT 58.930000 -32.710000 60.110000 -31.530000 ;
        RECT 238.930000 -31.110000 240.110000 -29.930000 ;
        RECT 238.930000 -32.710000 240.110000 -31.530000 ;
        RECT 418.930000 -31.110000 420.110000 -29.930000 ;
        RECT 418.930000 -32.710000 420.110000 -31.530000 ;
        RECT 598.930000 -31.110000 600.110000 -29.930000 ;
        RECT 598.930000 -32.710000 600.110000 -31.530000 ;
        RECT 778.930000 -31.110000 780.110000 -29.930000 ;
        RECT 778.930000 -32.710000 780.110000 -31.530000 ;
        RECT 958.930000 -31.110000 960.110000 -29.930000 ;
        RECT 958.930000 -32.710000 960.110000 -31.530000 ;
        RECT 1138.930000 -31.110000 1140.110000 -29.930000 ;
        RECT 1138.930000 -32.710000 1140.110000 -31.530000 ;
        RECT 1318.930000 -31.110000 1320.110000 -29.930000 ;
        RECT 1318.930000 -32.710000 1320.110000 -31.530000 ;
        RECT 1498.930000 -31.110000 1500.110000 -29.930000 ;
        RECT 1498.930000 -32.710000 1500.110000 -31.530000 ;
        RECT 1678.930000 -31.110000 1680.110000 -29.930000 ;
        RECT 1678.930000 -32.710000 1680.110000 -31.530000 ;
        RECT 1858.930000 -31.110000 1860.110000 -29.930000 ;
        RECT 1858.930000 -32.710000 1860.110000 -31.530000 ;
        RECT 2038.930000 -31.110000 2040.110000 -29.930000 ;
        RECT 2038.930000 -32.710000 2040.110000 -31.530000 ;
        RECT 2218.930000 -31.110000 2220.110000 -29.930000 ;
        RECT 2218.930000 -32.710000 2220.110000 -31.530000 ;
        RECT 2398.930000 -31.110000 2400.110000 -29.930000 ;
        RECT 2398.930000 -32.710000 2400.110000 -31.530000 ;
        RECT 2578.930000 -31.110000 2580.110000 -29.930000 ;
        RECT 2578.930000 -32.710000 2580.110000 -31.530000 ;
        RECT 2758.930000 -31.110000 2760.110000 -29.930000 ;
        RECT 2758.930000 -32.710000 2760.110000 -31.530000 ;
        RECT 2955.710000 -31.110000 2956.890000 -29.930000 ;
        RECT 2955.710000 -32.710000 2956.890000 -31.530000 ;
      LAYER met5 ;
        RECT -38.180000 3552.500000 -35.180000 3552.510000 ;
        RECT 58.020000 3552.500000 61.020000 3552.510000 ;
        RECT 238.020000 3552.500000 241.020000 3552.510000 ;
        RECT 418.020000 3552.500000 421.020000 3552.510000 ;
        RECT 598.020000 3552.500000 601.020000 3552.510000 ;
        RECT 778.020000 3552.500000 781.020000 3552.510000 ;
        RECT 958.020000 3552.500000 961.020000 3552.510000 ;
        RECT 1138.020000 3552.500000 1141.020000 3552.510000 ;
        RECT 1318.020000 3552.500000 1321.020000 3552.510000 ;
        RECT 1498.020000 3552.500000 1501.020000 3552.510000 ;
        RECT 1678.020000 3552.500000 1681.020000 3552.510000 ;
        RECT 1858.020000 3552.500000 1861.020000 3552.510000 ;
        RECT 2038.020000 3552.500000 2041.020000 3552.510000 ;
        RECT 2218.020000 3552.500000 2221.020000 3552.510000 ;
        RECT 2398.020000 3552.500000 2401.020000 3552.510000 ;
        RECT 2578.020000 3552.500000 2581.020000 3552.510000 ;
        RECT 2758.020000 3552.500000 2761.020000 3552.510000 ;
        RECT 2954.800000 3552.500000 2957.800000 3552.510000 ;
        RECT -38.180000 3549.500000 2957.800000 3552.500000 ;
        RECT -38.180000 3549.490000 -35.180000 3549.500000 ;
        RECT 58.020000 3549.490000 61.020000 3549.500000 ;
        RECT 238.020000 3549.490000 241.020000 3549.500000 ;
        RECT 418.020000 3549.490000 421.020000 3549.500000 ;
        RECT 598.020000 3549.490000 601.020000 3549.500000 ;
        RECT 778.020000 3549.490000 781.020000 3549.500000 ;
        RECT 958.020000 3549.490000 961.020000 3549.500000 ;
        RECT 1138.020000 3549.490000 1141.020000 3549.500000 ;
        RECT 1318.020000 3549.490000 1321.020000 3549.500000 ;
        RECT 1498.020000 3549.490000 1501.020000 3549.500000 ;
        RECT 1678.020000 3549.490000 1681.020000 3549.500000 ;
        RECT 1858.020000 3549.490000 1861.020000 3549.500000 ;
        RECT 2038.020000 3549.490000 2041.020000 3549.500000 ;
        RECT 2218.020000 3549.490000 2221.020000 3549.500000 ;
        RECT 2398.020000 3549.490000 2401.020000 3549.500000 ;
        RECT 2578.020000 3549.490000 2581.020000 3549.500000 ;
        RECT 2758.020000 3549.490000 2761.020000 3549.500000 ;
        RECT 2954.800000 3549.490000 2957.800000 3549.500000 ;
        RECT -38.180000 3486.380000 -35.180000 3486.390000 ;
        RECT 2954.800000 3486.380000 2957.800000 3486.390000 ;
        RECT -42.880000 3483.380000 -0.400000 3486.380000 ;
        RECT 2920.400000 3483.380000 2962.500000 3486.380000 ;
        RECT -38.180000 3483.370000 -35.180000 3483.380000 ;
        RECT 2954.800000 3483.370000 2957.800000 3483.380000 ;
        RECT -38.180000 3306.380000 -35.180000 3306.390000 ;
        RECT 2954.800000 3306.380000 2957.800000 3306.390000 ;
        RECT -42.880000 3303.380000 -0.400000 3306.380000 ;
        RECT 2920.400000 3303.380000 2962.500000 3306.380000 ;
        RECT -38.180000 3303.370000 -35.180000 3303.380000 ;
        RECT 2954.800000 3303.370000 2957.800000 3303.380000 ;
        RECT -38.180000 3126.380000 -35.180000 3126.390000 ;
        RECT 2954.800000 3126.380000 2957.800000 3126.390000 ;
        RECT -42.880000 3123.380000 -0.400000 3126.380000 ;
        RECT 2920.400000 3123.380000 2962.500000 3126.380000 ;
        RECT -38.180000 3123.370000 -35.180000 3123.380000 ;
        RECT 2954.800000 3123.370000 2957.800000 3123.380000 ;
        RECT -38.180000 2946.380000 -35.180000 2946.390000 ;
        RECT 2954.800000 2946.380000 2957.800000 2946.390000 ;
        RECT -42.880000 2943.380000 -0.400000 2946.380000 ;
        RECT 2920.400000 2943.380000 2962.500000 2946.380000 ;
        RECT -38.180000 2943.370000 -35.180000 2943.380000 ;
        RECT 2954.800000 2943.370000 2957.800000 2943.380000 ;
        RECT -38.180000 2766.380000 -35.180000 2766.390000 ;
        RECT 2954.800000 2766.380000 2957.800000 2766.390000 ;
        RECT -42.880000 2763.380000 -0.400000 2766.380000 ;
        RECT 2920.400000 2763.380000 2962.500000 2766.380000 ;
        RECT -38.180000 2763.370000 -35.180000 2763.380000 ;
        RECT 2954.800000 2763.370000 2957.800000 2763.380000 ;
        RECT -38.180000 2586.380000 -35.180000 2586.390000 ;
        RECT 2954.800000 2586.380000 2957.800000 2586.390000 ;
        RECT -42.880000 2583.380000 -0.400000 2586.380000 ;
        RECT 2920.400000 2583.380000 2962.500000 2586.380000 ;
        RECT -38.180000 2583.370000 -35.180000 2583.380000 ;
        RECT 2954.800000 2583.370000 2957.800000 2583.380000 ;
        RECT -38.180000 2406.380000 -35.180000 2406.390000 ;
        RECT 2954.800000 2406.380000 2957.800000 2406.390000 ;
        RECT -42.880000 2403.380000 -0.400000 2406.380000 ;
        RECT 2920.400000 2403.380000 2962.500000 2406.380000 ;
        RECT -38.180000 2403.370000 -35.180000 2403.380000 ;
        RECT 2954.800000 2403.370000 2957.800000 2403.380000 ;
        RECT -38.180000 2226.380000 -35.180000 2226.390000 ;
        RECT 2954.800000 2226.380000 2957.800000 2226.390000 ;
        RECT -42.880000 2223.380000 -0.400000 2226.380000 ;
        RECT 2920.400000 2223.380000 2962.500000 2226.380000 ;
        RECT -38.180000 2223.370000 -35.180000 2223.380000 ;
        RECT 2954.800000 2223.370000 2957.800000 2223.380000 ;
        RECT -38.180000 2046.380000 -35.180000 2046.390000 ;
        RECT 2954.800000 2046.380000 2957.800000 2046.390000 ;
        RECT -42.880000 2043.380000 -0.400000 2046.380000 ;
        RECT 2920.400000 2043.380000 2962.500000 2046.380000 ;
        RECT -38.180000 2043.370000 -35.180000 2043.380000 ;
        RECT 2954.800000 2043.370000 2957.800000 2043.380000 ;
        RECT -38.180000 1866.380000 -35.180000 1866.390000 ;
        RECT 2954.800000 1866.380000 2957.800000 1866.390000 ;
        RECT -42.880000 1863.380000 -0.400000 1866.380000 ;
        RECT 2920.400000 1863.380000 2962.500000 1866.380000 ;
        RECT -38.180000 1863.370000 -35.180000 1863.380000 ;
        RECT 2954.800000 1863.370000 2957.800000 1863.380000 ;
        RECT -38.180000 1686.380000 -35.180000 1686.390000 ;
        RECT 2954.800000 1686.380000 2957.800000 1686.390000 ;
        RECT -42.880000 1683.380000 -0.400000 1686.380000 ;
        RECT 2920.400000 1683.380000 2962.500000 1686.380000 ;
        RECT -38.180000 1683.370000 -35.180000 1683.380000 ;
        RECT 2954.800000 1683.370000 2957.800000 1683.380000 ;
        RECT -38.180000 1506.380000 -35.180000 1506.390000 ;
        RECT 2954.800000 1506.380000 2957.800000 1506.390000 ;
        RECT -42.880000 1503.380000 -0.400000 1506.380000 ;
        RECT 2920.400000 1503.380000 2962.500000 1506.380000 ;
        RECT -38.180000 1503.370000 -35.180000 1503.380000 ;
        RECT 2954.800000 1503.370000 2957.800000 1503.380000 ;
        RECT -38.180000 1326.380000 -35.180000 1326.390000 ;
        RECT 2954.800000 1326.380000 2957.800000 1326.390000 ;
        RECT -42.880000 1323.380000 -0.400000 1326.380000 ;
        RECT 2920.400000 1323.380000 2962.500000 1326.380000 ;
        RECT -38.180000 1323.370000 -35.180000 1323.380000 ;
        RECT 2954.800000 1323.370000 2957.800000 1323.380000 ;
        RECT -38.180000 1146.380000 -35.180000 1146.390000 ;
        RECT 2954.800000 1146.380000 2957.800000 1146.390000 ;
        RECT -42.880000 1143.380000 -0.400000 1146.380000 ;
        RECT 2920.400000 1143.380000 2962.500000 1146.380000 ;
        RECT -38.180000 1143.370000 -35.180000 1143.380000 ;
        RECT 2954.800000 1143.370000 2957.800000 1143.380000 ;
        RECT -38.180000 966.380000 -35.180000 966.390000 ;
        RECT 2954.800000 966.380000 2957.800000 966.390000 ;
        RECT -42.880000 963.380000 -0.400000 966.380000 ;
        RECT 2920.400000 963.380000 2962.500000 966.380000 ;
        RECT -38.180000 963.370000 -35.180000 963.380000 ;
        RECT 2954.800000 963.370000 2957.800000 963.380000 ;
        RECT -38.180000 786.380000 -35.180000 786.390000 ;
        RECT 2954.800000 786.380000 2957.800000 786.390000 ;
        RECT -42.880000 783.380000 -0.400000 786.380000 ;
        RECT 2920.400000 783.380000 2962.500000 786.380000 ;
        RECT -38.180000 783.370000 -35.180000 783.380000 ;
        RECT 2954.800000 783.370000 2957.800000 783.380000 ;
        RECT -38.180000 606.380000 -35.180000 606.390000 ;
        RECT 2954.800000 606.380000 2957.800000 606.390000 ;
        RECT -42.880000 603.380000 -0.400000 606.380000 ;
        RECT 2920.400000 603.380000 2962.500000 606.380000 ;
        RECT -38.180000 603.370000 -35.180000 603.380000 ;
        RECT 2954.800000 603.370000 2957.800000 603.380000 ;
        RECT -38.180000 426.380000 -35.180000 426.390000 ;
        RECT 2954.800000 426.380000 2957.800000 426.390000 ;
        RECT -42.880000 423.380000 -0.400000 426.380000 ;
        RECT 2920.400000 423.380000 2962.500000 426.380000 ;
        RECT -38.180000 423.370000 -35.180000 423.380000 ;
        RECT 2954.800000 423.370000 2957.800000 423.380000 ;
        RECT -38.180000 246.380000 -35.180000 246.390000 ;
        RECT 2954.800000 246.380000 2957.800000 246.390000 ;
        RECT -42.880000 243.380000 -0.400000 246.380000 ;
        RECT 2920.400000 243.380000 2962.500000 246.380000 ;
        RECT -38.180000 243.370000 -35.180000 243.380000 ;
        RECT 2954.800000 243.370000 2957.800000 243.380000 ;
        RECT -38.180000 66.380000 -35.180000 66.390000 ;
        RECT 2954.800000 66.380000 2957.800000 66.390000 ;
        RECT -42.880000 63.380000 -0.400000 66.380000 ;
        RECT 2920.400000 63.380000 2962.500000 66.380000 ;
        RECT -38.180000 63.370000 -35.180000 63.380000 ;
        RECT 2954.800000 63.370000 2957.800000 63.380000 ;
        RECT -38.180000 -29.820000 -35.180000 -29.810000 ;
        RECT 58.020000 -29.820000 61.020000 -29.810000 ;
        RECT 238.020000 -29.820000 241.020000 -29.810000 ;
        RECT 418.020000 -29.820000 421.020000 -29.810000 ;
        RECT 598.020000 -29.820000 601.020000 -29.810000 ;
        RECT 778.020000 -29.820000 781.020000 -29.810000 ;
        RECT 958.020000 -29.820000 961.020000 -29.810000 ;
        RECT 1138.020000 -29.820000 1141.020000 -29.810000 ;
        RECT 1318.020000 -29.820000 1321.020000 -29.810000 ;
        RECT 1498.020000 -29.820000 1501.020000 -29.810000 ;
        RECT 1678.020000 -29.820000 1681.020000 -29.810000 ;
        RECT 1858.020000 -29.820000 1861.020000 -29.810000 ;
        RECT 2038.020000 -29.820000 2041.020000 -29.810000 ;
        RECT 2218.020000 -29.820000 2221.020000 -29.810000 ;
        RECT 2398.020000 -29.820000 2401.020000 -29.810000 ;
        RECT 2578.020000 -29.820000 2581.020000 -29.810000 ;
        RECT 2758.020000 -29.820000 2761.020000 -29.810000 ;
        RECT 2954.800000 -29.820000 2957.800000 -29.810000 ;
        RECT -38.180000 -32.820000 2957.800000 -29.820000 ;
        RECT -38.180000 -32.830000 -35.180000 -32.820000 ;
        RECT 58.020000 -32.830000 61.020000 -32.820000 ;
        RECT 238.020000 -32.830000 241.020000 -32.820000 ;
        RECT 418.020000 -32.830000 421.020000 -32.820000 ;
        RECT 598.020000 -32.830000 601.020000 -32.820000 ;
        RECT 778.020000 -32.830000 781.020000 -32.820000 ;
        RECT 958.020000 -32.830000 961.020000 -32.820000 ;
        RECT 1138.020000 -32.830000 1141.020000 -32.820000 ;
        RECT 1318.020000 -32.830000 1321.020000 -32.820000 ;
        RECT 1498.020000 -32.830000 1501.020000 -32.820000 ;
        RECT 1678.020000 -32.830000 1681.020000 -32.820000 ;
        RECT 1858.020000 -32.830000 1861.020000 -32.820000 ;
        RECT 2038.020000 -32.830000 2041.020000 -32.820000 ;
        RECT 2218.020000 -32.830000 2221.020000 -32.820000 ;
        RECT 2398.020000 -32.830000 2401.020000 -32.820000 ;
        RECT 2578.020000 -32.830000 2581.020000 -32.820000 ;
        RECT 2758.020000 -32.830000 2761.020000 -32.820000 ;
        RECT 2954.800000 -32.830000 2957.800000 -32.820000 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880000 -37.520000 -39.880000 3557.200000 ;
        RECT 148.020000 3520.400000 151.020000 3557.200000 ;
        RECT 328.020000 3520.400000 331.020000 3557.200000 ;
        RECT 508.020000 3520.400000 511.020000 3557.200000 ;
        RECT 688.020000 3520.400000 691.020000 3557.200000 ;
        RECT 868.020000 3520.400000 871.020000 3557.200000 ;
        RECT 1048.020000 3520.400000 1051.020000 3557.200000 ;
        RECT 1228.020000 3520.400000 1231.020000 3557.200000 ;
        RECT 1408.020000 3520.400000 1411.020000 3557.200000 ;
        RECT 1588.020000 3520.400000 1591.020000 3557.200000 ;
        RECT 1768.020000 3520.400000 1771.020000 3557.200000 ;
        RECT 1948.020000 3520.400000 1951.020000 3557.200000 ;
        RECT 2128.020000 3520.400000 2131.020000 3557.200000 ;
        RECT 2308.020000 3520.400000 2311.020000 3557.200000 ;
        RECT 2488.020000 3520.400000 2491.020000 3557.200000 ;
        RECT 2668.020000 3520.400000 2671.020000 3557.200000 ;
        RECT 2848.020000 3520.400000 2851.020000 3557.200000 ;
        RECT 148.020000 -37.520000 151.020000 -0.400000 ;
        RECT 328.020000 -37.520000 331.020000 -0.400000 ;
        RECT 508.020000 -37.520000 511.020000 -0.400000 ;
        RECT 688.020000 -37.520000 691.020000 -0.400000 ;
        RECT 868.020000 -37.520000 871.020000 -0.400000 ;
        RECT 1048.020000 -37.520000 1051.020000 -0.400000 ;
        RECT 1228.020000 -37.520000 1231.020000 -0.400000 ;
        RECT 1408.020000 -37.520000 1411.020000 -0.400000 ;
        RECT 1588.020000 -37.520000 1591.020000 -0.400000 ;
        RECT 1768.020000 -37.520000 1771.020000 -0.400000 ;
        RECT 1948.020000 -37.520000 1951.020000 -0.400000 ;
        RECT 2128.020000 -37.520000 2131.020000 -0.400000 ;
        RECT 2308.020000 -37.520000 2311.020000 -0.400000 ;
        RECT 2488.020000 -37.520000 2491.020000 -0.400000 ;
        RECT 2668.020000 -37.520000 2671.020000 -0.400000 ;
        RECT 2848.020000 -37.520000 2851.020000 -0.400000 ;
        RECT 2959.500000 -37.520000 2962.500000 3557.200000 ;
      LAYER via4 ;
        RECT -41.970000 3555.910000 -40.790000 3557.090000 ;
        RECT -41.970000 3554.310000 -40.790000 3555.490000 ;
        RECT 148.930000 3555.910000 150.110000 3557.090000 ;
        RECT 148.930000 3554.310000 150.110000 3555.490000 ;
        RECT 328.930000 3555.910000 330.110000 3557.090000 ;
        RECT 328.930000 3554.310000 330.110000 3555.490000 ;
        RECT 508.930000 3555.910000 510.110000 3557.090000 ;
        RECT 508.930000 3554.310000 510.110000 3555.490000 ;
        RECT 688.930000 3555.910000 690.110000 3557.090000 ;
        RECT 688.930000 3554.310000 690.110000 3555.490000 ;
        RECT 868.930000 3555.910000 870.110000 3557.090000 ;
        RECT 868.930000 3554.310000 870.110000 3555.490000 ;
        RECT 1048.930000 3555.910000 1050.110000 3557.090000 ;
        RECT 1048.930000 3554.310000 1050.110000 3555.490000 ;
        RECT 1228.930000 3555.910000 1230.110000 3557.090000 ;
        RECT 1228.930000 3554.310000 1230.110000 3555.490000 ;
        RECT 1408.930000 3555.910000 1410.110000 3557.090000 ;
        RECT 1408.930000 3554.310000 1410.110000 3555.490000 ;
        RECT 1588.930000 3555.910000 1590.110000 3557.090000 ;
        RECT 1588.930000 3554.310000 1590.110000 3555.490000 ;
        RECT 1768.930000 3555.910000 1770.110000 3557.090000 ;
        RECT 1768.930000 3554.310000 1770.110000 3555.490000 ;
        RECT 1948.930000 3555.910000 1950.110000 3557.090000 ;
        RECT 1948.930000 3554.310000 1950.110000 3555.490000 ;
        RECT 2128.930000 3555.910000 2130.110000 3557.090000 ;
        RECT 2128.930000 3554.310000 2130.110000 3555.490000 ;
        RECT 2308.930000 3555.910000 2310.110000 3557.090000 ;
        RECT 2308.930000 3554.310000 2310.110000 3555.490000 ;
        RECT 2488.930000 3555.910000 2490.110000 3557.090000 ;
        RECT 2488.930000 3554.310000 2490.110000 3555.490000 ;
        RECT 2668.930000 3555.910000 2670.110000 3557.090000 ;
        RECT 2668.930000 3554.310000 2670.110000 3555.490000 ;
        RECT 2848.930000 3555.910000 2850.110000 3557.090000 ;
        RECT 2848.930000 3554.310000 2850.110000 3555.490000 ;
        RECT 2960.410000 3555.910000 2961.590000 3557.090000 ;
        RECT 2960.410000 3554.310000 2961.590000 3555.490000 ;
        RECT -41.970000 3395.090000 -40.790000 3396.270000 ;
        RECT -41.970000 3393.490000 -40.790000 3394.670000 ;
        RECT -41.970000 3215.090000 -40.790000 3216.270000 ;
        RECT -41.970000 3213.490000 -40.790000 3214.670000 ;
        RECT -41.970000 3035.090000 -40.790000 3036.270000 ;
        RECT -41.970000 3033.490000 -40.790000 3034.670000 ;
        RECT -41.970000 2855.090000 -40.790000 2856.270000 ;
        RECT -41.970000 2853.490000 -40.790000 2854.670000 ;
        RECT -41.970000 2675.090000 -40.790000 2676.270000 ;
        RECT -41.970000 2673.490000 -40.790000 2674.670000 ;
        RECT -41.970000 2495.090000 -40.790000 2496.270000 ;
        RECT -41.970000 2493.490000 -40.790000 2494.670000 ;
        RECT -41.970000 2315.090000 -40.790000 2316.270000 ;
        RECT -41.970000 2313.490000 -40.790000 2314.670000 ;
        RECT -41.970000 2135.090000 -40.790000 2136.270000 ;
        RECT -41.970000 2133.490000 -40.790000 2134.670000 ;
        RECT -41.970000 1955.090000 -40.790000 1956.270000 ;
        RECT -41.970000 1953.490000 -40.790000 1954.670000 ;
        RECT -41.970000 1775.090000 -40.790000 1776.270000 ;
        RECT -41.970000 1773.490000 -40.790000 1774.670000 ;
        RECT -41.970000 1595.090000 -40.790000 1596.270000 ;
        RECT -41.970000 1593.490000 -40.790000 1594.670000 ;
        RECT -41.970000 1415.090000 -40.790000 1416.270000 ;
        RECT -41.970000 1413.490000 -40.790000 1414.670000 ;
        RECT -41.970000 1235.090000 -40.790000 1236.270000 ;
        RECT -41.970000 1233.490000 -40.790000 1234.670000 ;
        RECT -41.970000 1055.090000 -40.790000 1056.270000 ;
        RECT -41.970000 1053.490000 -40.790000 1054.670000 ;
        RECT -41.970000 875.090000 -40.790000 876.270000 ;
        RECT -41.970000 873.490000 -40.790000 874.670000 ;
        RECT -41.970000 695.090000 -40.790000 696.270000 ;
        RECT -41.970000 693.490000 -40.790000 694.670000 ;
        RECT -41.970000 515.090000 -40.790000 516.270000 ;
        RECT -41.970000 513.490000 -40.790000 514.670000 ;
        RECT -41.970000 335.090000 -40.790000 336.270000 ;
        RECT -41.970000 333.490000 -40.790000 334.670000 ;
        RECT -41.970000 155.090000 -40.790000 156.270000 ;
        RECT -41.970000 153.490000 -40.790000 154.670000 ;
        RECT 2960.410000 3395.090000 2961.590000 3396.270000 ;
        RECT 2960.410000 3393.490000 2961.590000 3394.670000 ;
        RECT 2960.410000 3215.090000 2961.590000 3216.270000 ;
        RECT 2960.410000 3213.490000 2961.590000 3214.670000 ;
        RECT 2960.410000 3035.090000 2961.590000 3036.270000 ;
        RECT 2960.410000 3033.490000 2961.590000 3034.670000 ;
        RECT 2960.410000 2855.090000 2961.590000 2856.270000 ;
        RECT 2960.410000 2853.490000 2961.590000 2854.670000 ;
        RECT 2960.410000 2675.090000 2961.590000 2676.270000 ;
        RECT 2960.410000 2673.490000 2961.590000 2674.670000 ;
        RECT 2960.410000 2495.090000 2961.590000 2496.270000 ;
        RECT 2960.410000 2493.490000 2961.590000 2494.670000 ;
        RECT 2960.410000 2315.090000 2961.590000 2316.270000 ;
        RECT 2960.410000 2313.490000 2961.590000 2314.670000 ;
        RECT 2960.410000 2135.090000 2961.590000 2136.270000 ;
        RECT 2960.410000 2133.490000 2961.590000 2134.670000 ;
        RECT 2960.410000 1955.090000 2961.590000 1956.270000 ;
        RECT 2960.410000 1953.490000 2961.590000 1954.670000 ;
        RECT 2960.410000 1775.090000 2961.590000 1776.270000 ;
        RECT 2960.410000 1773.490000 2961.590000 1774.670000 ;
        RECT 2960.410000 1595.090000 2961.590000 1596.270000 ;
        RECT 2960.410000 1593.490000 2961.590000 1594.670000 ;
        RECT 2960.410000 1415.090000 2961.590000 1416.270000 ;
        RECT 2960.410000 1413.490000 2961.590000 1414.670000 ;
        RECT 2960.410000 1235.090000 2961.590000 1236.270000 ;
        RECT 2960.410000 1233.490000 2961.590000 1234.670000 ;
        RECT 2960.410000 1055.090000 2961.590000 1056.270000 ;
        RECT 2960.410000 1053.490000 2961.590000 1054.670000 ;
        RECT 2960.410000 875.090000 2961.590000 876.270000 ;
        RECT 2960.410000 873.490000 2961.590000 874.670000 ;
        RECT 2960.410000 695.090000 2961.590000 696.270000 ;
        RECT 2960.410000 693.490000 2961.590000 694.670000 ;
        RECT 2960.410000 515.090000 2961.590000 516.270000 ;
        RECT 2960.410000 513.490000 2961.590000 514.670000 ;
        RECT 2960.410000 335.090000 2961.590000 336.270000 ;
        RECT 2960.410000 333.490000 2961.590000 334.670000 ;
        RECT 2960.410000 155.090000 2961.590000 156.270000 ;
        RECT 2960.410000 153.490000 2961.590000 154.670000 ;
        RECT -41.970000 -35.810000 -40.790000 -34.630000 ;
        RECT -41.970000 -37.410000 -40.790000 -36.230000 ;
        RECT 148.930000 -35.810000 150.110000 -34.630000 ;
        RECT 148.930000 -37.410000 150.110000 -36.230000 ;
        RECT 328.930000 -35.810000 330.110000 -34.630000 ;
        RECT 328.930000 -37.410000 330.110000 -36.230000 ;
        RECT 508.930000 -35.810000 510.110000 -34.630000 ;
        RECT 508.930000 -37.410000 510.110000 -36.230000 ;
        RECT 688.930000 -35.810000 690.110000 -34.630000 ;
        RECT 688.930000 -37.410000 690.110000 -36.230000 ;
        RECT 868.930000 -35.810000 870.110000 -34.630000 ;
        RECT 868.930000 -37.410000 870.110000 -36.230000 ;
        RECT 1048.930000 -35.810000 1050.110000 -34.630000 ;
        RECT 1048.930000 -37.410000 1050.110000 -36.230000 ;
        RECT 1228.930000 -35.810000 1230.110000 -34.630000 ;
        RECT 1228.930000 -37.410000 1230.110000 -36.230000 ;
        RECT 1408.930000 -35.810000 1410.110000 -34.630000 ;
        RECT 1408.930000 -37.410000 1410.110000 -36.230000 ;
        RECT 1588.930000 -35.810000 1590.110000 -34.630000 ;
        RECT 1588.930000 -37.410000 1590.110000 -36.230000 ;
        RECT 1768.930000 -35.810000 1770.110000 -34.630000 ;
        RECT 1768.930000 -37.410000 1770.110000 -36.230000 ;
        RECT 1948.930000 -35.810000 1950.110000 -34.630000 ;
        RECT 1948.930000 -37.410000 1950.110000 -36.230000 ;
        RECT 2128.930000 -35.810000 2130.110000 -34.630000 ;
        RECT 2128.930000 -37.410000 2130.110000 -36.230000 ;
        RECT 2308.930000 -35.810000 2310.110000 -34.630000 ;
        RECT 2308.930000 -37.410000 2310.110000 -36.230000 ;
        RECT 2488.930000 -35.810000 2490.110000 -34.630000 ;
        RECT 2488.930000 -37.410000 2490.110000 -36.230000 ;
        RECT 2668.930000 -35.810000 2670.110000 -34.630000 ;
        RECT 2668.930000 -37.410000 2670.110000 -36.230000 ;
        RECT 2848.930000 -35.810000 2850.110000 -34.630000 ;
        RECT 2848.930000 -37.410000 2850.110000 -36.230000 ;
        RECT 2960.410000 -35.810000 2961.590000 -34.630000 ;
        RECT 2960.410000 -37.410000 2961.590000 -36.230000 ;
      LAYER met5 ;
        RECT -42.880000 3557.200000 -39.880000 3557.210000 ;
        RECT 148.020000 3557.200000 151.020000 3557.210000 ;
        RECT 328.020000 3557.200000 331.020000 3557.210000 ;
        RECT 508.020000 3557.200000 511.020000 3557.210000 ;
        RECT 688.020000 3557.200000 691.020000 3557.210000 ;
        RECT 868.020000 3557.200000 871.020000 3557.210000 ;
        RECT 1048.020000 3557.200000 1051.020000 3557.210000 ;
        RECT 1228.020000 3557.200000 1231.020000 3557.210000 ;
        RECT 1408.020000 3557.200000 1411.020000 3557.210000 ;
        RECT 1588.020000 3557.200000 1591.020000 3557.210000 ;
        RECT 1768.020000 3557.200000 1771.020000 3557.210000 ;
        RECT 1948.020000 3557.200000 1951.020000 3557.210000 ;
        RECT 2128.020000 3557.200000 2131.020000 3557.210000 ;
        RECT 2308.020000 3557.200000 2311.020000 3557.210000 ;
        RECT 2488.020000 3557.200000 2491.020000 3557.210000 ;
        RECT 2668.020000 3557.200000 2671.020000 3557.210000 ;
        RECT 2848.020000 3557.200000 2851.020000 3557.210000 ;
        RECT 2959.500000 3557.200000 2962.500000 3557.210000 ;
        RECT -42.880000 3554.200000 2962.500000 3557.200000 ;
        RECT -42.880000 3554.190000 -39.880000 3554.200000 ;
        RECT 148.020000 3554.190000 151.020000 3554.200000 ;
        RECT 328.020000 3554.190000 331.020000 3554.200000 ;
        RECT 508.020000 3554.190000 511.020000 3554.200000 ;
        RECT 688.020000 3554.190000 691.020000 3554.200000 ;
        RECT 868.020000 3554.190000 871.020000 3554.200000 ;
        RECT 1048.020000 3554.190000 1051.020000 3554.200000 ;
        RECT 1228.020000 3554.190000 1231.020000 3554.200000 ;
        RECT 1408.020000 3554.190000 1411.020000 3554.200000 ;
        RECT 1588.020000 3554.190000 1591.020000 3554.200000 ;
        RECT 1768.020000 3554.190000 1771.020000 3554.200000 ;
        RECT 1948.020000 3554.190000 1951.020000 3554.200000 ;
        RECT 2128.020000 3554.190000 2131.020000 3554.200000 ;
        RECT 2308.020000 3554.190000 2311.020000 3554.200000 ;
        RECT 2488.020000 3554.190000 2491.020000 3554.200000 ;
        RECT 2668.020000 3554.190000 2671.020000 3554.200000 ;
        RECT 2848.020000 3554.190000 2851.020000 3554.200000 ;
        RECT 2959.500000 3554.190000 2962.500000 3554.200000 ;
        RECT -42.880000 3396.380000 -39.880000 3396.390000 ;
        RECT 2959.500000 3396.380000 2962.500000 3396.390000 ;
        RECT -42.880000 3393.380000 -0.400000 3396.380000 ;
        RECT 2920.400000 3393.380000 2962.500000 3396.380000 ;
        RECT -42.880000 3393.370000 -39.880000 3393.380000 ;
        RECT 2959.500000 3393.370000 2962.500000 3393.380000 ;
        RECT -42.880000 3216.380000 -39.880000 3216.390000 ;
        RECT 2959.500000 3216.380000 2962.500000 3216.390000 ;
        RECT -42.880000 3213.380000 -0.400000 3216.380000 ;
        RECT 2920.400000 3213.380000 2962.500000 3216.380000 ;
        RECT -42.880000 3213.370000 -39.880000 3213.380000 ;
        RECT 2959.500000 3213.370000 2962.500000 3213.380000 ;
        RECT -42.880000 3036.380000 -39.880000 3036.390000 ;
        RECT 2959.500000 3036.380000 2962.500000 3036.390000 ;
        RECT -42.880000 3033.380000 -0.400000 3036.380000 ;
        RECT 2920.400000 3033.380000 2962.500000 3036.380000 ;
        RECT -42.880000 3033.370000 -39.880000 3033.380000 ;
        RECT 2959.500000 3033.370000 2962.500000 3033.380000 ;
        RECT -42.880000 2856.380000 -39.880000 2856.390000 ;
        RECT 2959.500000 2856.380000 2962.500000 2856.390000 ;
        RECT -42.880000 2853.380000 -0.400000 2856.380000 ;
        RECT 2920.400000 2853.380000 2962.500000 2856.380000 ;
        RECT -42.880000 2853.370000 -39.880000 2853.380000 ;
        RECT 2959.500000 2853.370000 2962.500000 2853.380000 ;
        RECT -42.880000 2676.380000 -39.880000 2676.390000 ;
        RECT 2959.500000 2676.380000 2962.500000 2676.390000 ;
        RECT -42.880000 2673.380000 -0.400000 2676.380000 ;
        RECT 2920.400000 2673.380000 2962.500000 2676.380000 ;
        RECT -42.880000 2673.370000 -39.880000 2673.380000 ;
        RECT 2959.500000 2673.370000 2962.500000 2673.380000 ;
        RECT -42.880000 2496.380000 -39.880000 2496.390000 ;
        RECT 2959.500000 2496.380000 2962.500000 2496.390000 ;
        RECT -42.880000 2493.380000 -0.400000 2496.380000 ;
        RECT 2920.400000 2493.380000 2962.500000 2496.380000 ;
        RECT -42.880000 2493.370000 -39.880000 2493.380000 ;
        RECT 2959.500000 2493.370000 2962.500000 2493.380000 ;
        RECT -42.880000 2316.380000 -39.880000 2316.390000 ;
        RECT 2959.500000 2316.380000 2962.500000 2316.390000 ;
        RECT -42.880000 2313.380000 -0.400000 2316.380000 ;
        RECT 2920.400000 2313.380000 2962.500000 2316.380000 ;
        RECT -42.880000 2313.370000 -39.880000 2313.380000 ;
        RECT 2959.500000 2313.370000 2962.500000 2313.380000 ;
        RECT -42.880000 2136.380000 -39.880000 2136.390000 ;
        RECT 2959.500000 2136.380000 2962.500000 2136.390000 ;
        RECT -42.880000 2133.380000 -0.400000 2136.380000 ;
        RECT 2920.400000 2133.380000 2962.500000 2136.380000 ;
        RECT -42.880000 2133.370000 -39.880000 2133.380000 ;
        RECT 2959.500000 2133.370000 2962.500000 2133.380000 ;
        RECT -42.880000 1956.380000 -39.880000 1956.390000 ;
        RECT 2959.500000 1956.380000 2962.500000 1956.390000 ;
        RECT -42.880000 1953.380000 -0.400000 1956.380000 ;
        RECT 2920.400000 1953.380000 2962.500000 1956.380000 ;
        RECT -42.880000 1953.370000 -39.880000 1953.380000 ;
        RECT 2959.500000 1953.370000 2962.500000 1953.380000 ;
        RECT -42.880000 1776.380000 -39.880000 1776.390000 ;
        RECT 2959.500000 1776.380000 2962.500000 1776.390000 ;
        RECT -42.880000 1773.380000 -0.400000 1776.380000 ;
        RECT 2920.400000 1773.380000 2962.500000 1776.380000 ;
        RECT -42.880000 1773.370000 -39.880000 1773.380000 ;
        RECT 2959.500000 1773.370000 2962.500000 1773.380000 ;
        RECT -42.880000 1596.380000 -39.880000 1596.390000 ;
        RECT 2959.500000 1596.380000 2962.500000 1596.390000 ;
        RECT -42.880000 1593.380000 -0.400000 1596.380000 ;
        RECT 2920.400000 1593.380000 2962.500000 1596.380000 ;
        RECT -42.880000 1593.370000 -39.880000 1593.380000 ;
        RECT 2959.500000 1593.370000 2962.500000 1593.380000 ;
        RECT -42.880000 1416.380000 -39.880000 1416.390000 ;
        RECT 2959.500000 1416.380000 2962.500000 1416.390000 ;
        RECT -42.880000 1413.380000 -0.400000 1416.380000 ;
        RECT 2920.400000 1413.380000 2962.500000 1416.380000 ;
        RECT -42.880000 1413.370000 -39.880000 1413.380000 ;
        RECT 2959.500000 1413.370000 2962.500000 1413.380000 ;
        RECT -42.880000 1236.380000 -39.880000 1236.390000 ;
        RECT 2959.500000 1236.380000 2962.500000 1236.390000 ;
        RECT -42.880000 1233.380000 -0.400000 1236.380000 ;
        RECT 2920.400000 1233.380000 2962.500000 1236.380000 ;
        RECT -42.880000 1233.370000 -39.880000 1233.380000 ;
        RECT 2959.500000 1233.370000 2962.500000 1233.380000 ;
        RECT -42.880000 1056.380000 -39.880000 1056.390000 ;
        RECT 2959.500000 1056.380000 2962.500000 1056.390000 ;
        RECT -42.880000 1053.380000 -0.400000 1056.380000 ;
        RECT 2920.400000 1053.380000 2962.500000 1056.380000 ;
        RECT -42.880000 1053.370000 -39.880000 1053.380000 ;
        RECT 2959.500000 1053.370000 2962.500000 1053.380000 ;
        RECT -42.880000 876.380000 -39.880000 876.390000 ;
        RECT 2959.500000 876.380000 2962.500000 876.390000 ;
        RECT -42.880000 873.380000 -0.400000 876.380000 ;
        RECT 2920.400000 873.380000 2962.500000 876.380000 ;
        RECT -42.880000 873.370000 -39.880000 873.380000 ;
        RECT 2959.500000 873.370000 2962.500000 873.380000 ;
        RECT -42.880000 696.380000 -39.880000 696.390000 ;
        RECT 2959.500000 696.380000 2962.500000 696.390000 ;
        RECT -42.880000 693.380000 -0.400000 696.380000 ;
        RECT 2920.400000 693.380000 2962.500000 696.380000 ;
        RECT -42.880000 693.370000 -39.880000 693.380000 ;
        RECT 2959.500000 693.370000 2962.500000 693.380000 ;
        RECT -42.880000 516.380000 -39.880000 516.390000 ;
        RECT 2959.500000 516.380000 2962.500000 516.390000 ;
        RECT -42.880000 513.380000 -0.400000 516.380000 ;
        RECT 2920.400000 513.380000 2962.500000 516.380000 ;
        RECT -42.880000 513.370000 -39.880000 513.380000 ;
        RECT 2959.500000 513.370000 2962.500000 513.380000 ;
        RECT -42.880000 336.380000 -39.880000 336.390000 ;
        RECT 2959.500000 336.380000 2962.500000 336.390000 ;
        RECT -42.880000 333.380000 -0.400000 336.380000 ;
        RECT 2920.400000 333.380000 2962.500000 336.380000 ;
        RECT -42.880000 333.370000 -39.880000 333.380000 ;
        RECT 2959.500000 333.370000 2962.500000 333.380000 ;
        RECT -42.880000 156.380000 -39.880000 156.390000 ;
        RECT 2959.500000 156.380000 2962.500000 156.390000 ;
        RECT -42.880000 153.380000 -0.400000 156.380000 ;
        RECT 2920.400000 153.380000 2962.500000 156.380000 ;
        RECT -42.880000 153.370000 -39.880000 153.380000 ;
        RECT 2959.500000 153.370000 2962.500000 153.380000 ;
        RECT -42.880000 -34.520000 -39.880000 -34.510000 ;
        RECT 148.020000 -34.520000 151.020000 -34.510000 ;
        RECT 328.020000 -34.520000 331.020000 -34.510000 ;
        RECT 508.020000 -34.520000 511.020000 -34.510000 ;
        RECT 688.020000 -34.520000 691.020000 -34.510000 ;
        RECT 868.020000 -34.520000 871.020000 -34.510000 ;
        RECT 1048.020000 -34.520000 1051.020000 -34.510000 ;
        RECT 1228.020000 -34.520000 1231.020000 -34.510000 ;
        RECT 1408.020000 -34.520000 1411.020000 -34.510000 ;
        RECT 1588.020000 -34.520000 1591.020000 -34.510000 ;
        RECT 1768.020000 -34.520000 1771.020000 -34.510000 ;
        RECT 1948.020000 -34.520000 1951.020000 -34.510000 ;
        RECT 2128.020000 -34.520000 2131.020000 -34.510000 ;
        RECT 2308.020000 -34.520000 2311.020000 -34.510000 ;
        RECT 2488.020000 -34.520000 2491.020000 -34.510000 ;
        RECT 2668.020000 -34.520000 2671.020000 -34.510000 ;
        RECT 2848.020000 -34.520000 2851.020000 -34.510000 ;
        RECT 2959.500000 -34.520000 2962.500000 -34.510000 ;
        RECT -42.880000 -37.520000 2962.500000 -34.520000 ;
        RECT -42.880000 -37.530000 -39.880000 -37.520000 ;
        RECT 148.020000 -37.530000 151.020000 -37.520000 ;
        RECT 328.020000 -37.530000 331.020000 -37.520000 ;
        RECT 508.020000 -37.530000 511.020000 -37.520000 ;
        RECT 688.020000 -37.530000 691.020000 -37.520000 ;
        RECT 868.020000 -37.530000 871.020000 -37.520000 ;
        RECT 1048.020000 -37.530000 1051.020000 -37.520000 ;
        RECT 1228.020000 -37.530000 1231.020000 -37.520000 ;
        RECT 1408.020000 -37.530000 1411.020000 -37.520000 ;
        RECT 1588.020000 -37.530000 1591.020000 -37.520000 ;
        RECT 1768.020000 -37.530000 1771.020000 -37.520000 ;
        RECT 1948.020000 -37.530000 1951.020000 -37.520000 ;
        RECT 2128.020000 -37.530000 2131.020000 -37.520000 ;
        RECT 2308.020000 -37.530000 2311.020000 -37.520000 ;
        RECT 2488.020000 -37.530000 2491.020000 -37.520000 ;
        RECT 2668.020000 -37.530000 2671.020000 -37.520000 ;
        RECT 2848.020000 -37.530000 2851.020000 -37.520000 ;
        RECT 2959.500000 -37.530000 2962.500000 -37.520000 ;
    END
  END vssa2
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 2920.0 3520.0 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 2920.0 3520.0 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 2920.0 3520.0 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 2920.0 3520.0 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 2920.0 3520.0 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 2920.0 3520.0 ;
   END
END user_project_wrapper
END LIBRARY
