magic
tech sky130A
magscale 12 1
timestamp 1598786935
<< metal5 >>
rect 30 90 45 105
rect 25 75 45 90
rect 20 70 45 75
rect 20 65 40 70
rect 15 60 40 65
rect 15 55 35 60
rect 10 50 35 55
rect 10 45 30 50
rect 5 40 30 45
rect 5 35 25 40
rect 0 30 25 35
rect 0 15 20 30
rect 0 0 15 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
