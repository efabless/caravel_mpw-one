magic
tech sky130A
magscale 1 2
timestamp 1621458646
<< locali >>
rect 6193 5015 6227 5185
<< viali >>
rect 5641 11305 5675 11339
rect 6193 11305 6227 11339
rect 6745 11305 6779 11339
rect 7205 11237 7239 11271
rect 9321 11237 9355 11271
rect 5457 11169 5491 11203
rect 5917 11169 5951 11203
rect 6009 11169 6043 11203
rect 6561 11169 6595 11203
rect 7021 11169 7055 11203
rect 7573 11169 7607 11203
rect 7849 11169 7883 11203
rect 8677 11169 8711 11203
rect 7941 11101 7975 11135
rect 5733 11033 5767 11067
rect 6377 11033 6411 11067
rect 7665 11033 7699 11067
rect 8585 11033 8619 11067
rect 9505 11033 9539 11067
rect 8861 10965 8895 10999
rect 6009 10761 6043 10795
rect 9137 10761 9171 10795
rect 8769 10693 8803 10727
rect 6745 10625 6779 10659
rect 5825 10557 5859 10591
rect 6469 10557 6503 10591
rect 8953 10557 8987 10591
rect 9321 10557 9355 10591
rect 8585 10489 8619 10523
rect 8217 10421 8251 10455
rect 9505 10421 9539 10455
rect 5825 10217 5859 10251
rect 6929 10149 6963 10183
rect 5365 10081 5399 10115
rect 5641 10081 5675 10115
rect 5917 10081 5951 10115
rect 6285 10081 6319 10115
rect 7021 10081 7055 10115
rect 7205 10081 7239 10115
rect 7481 10081 7515 10115
rect 7849 10013 7883 10047
rect 5549 9945 5583 9979
rect 6101 9877 6135 9911
rect 7297 9877 7331 9911
rect 9275 9877 9309 9911
rect 4905 9673 4939 9707
rect 5917 9673 5951 9707
rect 5825 9537 5859 9571
rect 6561 9537 6595 9571
rect 6929 9537 6963 9571
rect 9505 9537 9539 9571
rect 4721 9469 4755 9503
rect 4997 9469 5031 9503
rect 5273 9469 5307 9503
rect 6653 9469 6687 9503
rect 9045 9469 9079 9503
rect 8585 9401 8619 9435
rect 8769 9401 8803 9435
rect 5181 9333 5215 9367
rect 5457 9333 5491 9367
rect 8401 9333 8435 9367
rect 9045 9333 9079 9367
rect 5089 9129 5123 9163
rect 5733 9129 5767 9163
rect 9505 9129 9539 9163
rect 5825 9061 5859 9095
rect 7389 9061 7423 9095
rect 8033 9061 8067 9095
rect 5273 8993 5307 9027
rect 6285 8993 6319 9027
rect 6653 8993 6687 9027
rect 7297 8993 7331 9027
rect 7757 8993 7791 9027
rect 6009 8925 6043 8959
rect 7481 8925 7515 8959
rect 6837 8857 6871 8891
rect 5365 8789 5399 8823
rect 6469 8789 6503 8823
rect 6929 8789 6963 8823
rect 8309 8585 8343 8619
rect 9137 8585 9171 8619
rect 4629 8517 4663 8551
rect 8769 8517 8803 8551
rect 6469 8449 6503 8483
rect 6837 8449 6871 8483
rect 4445 8381 4479 8415
rect 4721 8381 4755 8415
rect 6561 8381 6595 8415
rect 8585 8381 8619 8415
rect 8953 8381 8987 8415
rect 9321 8381 9355 8415
rect 4997 8313 5031 8347
rect 9505 8313 9539 8347
rect 4353 7973 4387 8007
rect 6561 7973 6595 8007
rect 8769 7973 8803 8007
rect 4077 7905 4111 7939
rect 6285 7905 6319 7939
rect 8861 7905 8895 7939
rect 9321 7905 9355 7939
rect 8125 7837 8159 7871
rect 4261 7769 4295 7803
rect 9505 7769 9539 7803
rect 5641 7701 5675 7735
rect 8033 7701 8067 7735
rect 9321 7497 9355 7531
rect 4721 7361 4755 7395
rect 6193 7361 6227 7395
rect 6653 7361 6687 7395
rect 4169 7293 4203 7327
rect 4445 7293 4479 7327
rect 6377 7293 6411 7327
rect 8217 7293 8251 7327
rect 9045 7293 9079 7327
rect 9137 7293 9171 7327
rect 8585 7225 8619 7259
rect 8769 7225 8803 7259
rect 4353 7157 4387 7191
rect 8125 7157 8159 7191
rect 8401 7157 8435 7191
rect 4261 6953 4295 6987
rect 8815 6885 8849 6919
rect 3525 6817 3559 6851
rect 3801 6817 3835 6851
rect 4077 6817 4111 6851
rect 6285 6817 6319 6851
rect 6561 6817 6595 6851
rect 7021 6817 7055 6851
rect 8953 6817 8987 6851
rect 9046 6817 9080 6851
rect 4353 6749 4387 6783
rect 4629 6749 4663 6783
rect 7389 6749 7423 6783
rect 3709 6681 3743 6715
rect 6469 6681 6503 6715
rect 3433 6613 3467 6647
rect 3985 6613 4019 6647
rect 6101 6613 6135 6647
rect 6745 6613 6779 6647
rect 9137 6613 9171 6647
rect 8125 6409 8159 6443
rect 6653 6273 6687 6307
rect 8769 6273 8803 6307
rect 4261 6205 4295 6239
rect 4537 6205 4571 6239
rect 6377 6205 6411 6239
rect 8217 6205 8251 6239
rect 8953 6205 8987 6239
rect 9321 6205 9355 6239
rect 4813 6137 4847 6171
rect 8585 6137 8619 6171
rect 9505 6137 9539 6171
rect 4353 6069 4387 6103
rect 6285 6069 6319 6103
rect 8401 6069 8435 6103
rect 9137 6069 9171 6103
rect 4261 5865 4295 5899
rect 7389 5797 7423 5831
rect 3801 5729 3835 5763
rect 4077 5729 4111 5763
rect 6285 5729 6319 5763
rect 6745 5729 6779 5763
rect 7021 5729 7055 5763
rect 7573 5729 7607 5763
rect 4353 5661 4387 5695
rect 4629 5661 4663 5695
rect 7665 5661 7699 5695
rect 8033 5661 8067 5695
rect 3985 5525 4019 5559
rect 6101 5525 6135 5559
rect 6469 5525 6503 5559
rect 6929 5525 6963 5559
rect 7205 5525 7239 5559
rect 9459 5525 9493 5559
rect 6101 5253 6135 5287
rect 4629 5185 4663 5219
rect 6193 5185 6227 5219
rect 6837 5185 6871 5219
rect 8861 5185 8895 5219
rect 4261 5117 4295 5151
rect 4353 5117 4387 5151
rect 6377 5117 6411 5151
rect 9321 5117 9355 5151
rect 7113 5049 7147 5083
rect 9505 5049 9539 5083
rect 4077 4981 4111 5015
rect 6193 4981 6227 5015
rect 6561 4981 6595 5015
rect 8355 4777 8389 4811
rect 8769 4709 8803 4743
rect 4353 4641 4387 4675
rect 6193 4641 6227 4675
rect 4629 4573 4663 4607
rect 6561 4573 6595 4607
rect 6929 4573 6963 4607
rect 8677 4573 8711 4607
rect 9045 4573 9079 4607
rect 6101 4437 6135 4471
rect 6377 4437 6411 4471
rect 4340 4233 4374 4267
rect 4077 4097 4111 4131
rect 6929 4097 6963 4131
rect 8677 4097 8711 4131
rect 6009 4029 6043 4063
rect 6377 4029 6411 4063
rect 6653 4029 6687 4063
rect 8769 4029 8803 4063
rect 8862 4029 8896 4063
rect 9321 3961 9355 3995
rect 9505 3961 9539 3995
rect 5825 3893 5859 3927
rect 6193 3893 6227 3927
rect 6561 3893 6595 3927
rect 9137 3893 9171 3927
rect 8585 3689 8619 3723
rect 4629 3621 4663 3655
rect 6469 3621 6503 3655
rect 8401 3621 8435 3655
rect 4353 3553 4387 3587
rect 8217 3553 8251 3587
rect 8953 3553 8987 3587
rect 6101 3485 6135 3519
rect 6193 3485 6227 3519
rect 7941 3485 7975 3519
rect 9045 3485 9079 3519
rect 9137 3485 9171 3519
rect 5825 3145 5859 3179
rect 8585 3145 8619 3179
rect 4077 3009 4111 3043
rect 4353 3009 4387 3043
rect 6285 3009 6319 3043
rect 9137 3009 9171 3043
rect 6009 2941 6043 2975
rect 9045 2941 9079 2975
rect 6561 2873 6595 2907
rect 8309 2873 8343 2907
rect 8493 2873 8527 2907
rect 6193 2805 6227 2839
rect 8033 2805 8067 2839
rect 8953 2805 8987 2839
rect 4445 2601 4479 2635
rect 5733 2601 5767 2635
rect 8493 2601 8527 2635
rect 5365 2533 5399 2567
rect 7021 2533 7055 2567
rect 9321 2533 9355 2567
rect 4629 2465 4663 2499
rect 5089 2465 5123 2499
rect 5641 2465 5675 2499
rect 6101 2465 6135 2499
rect 6469 2465 6503 2499
rect 6745 2465 6779 2499
rect 8953 2465 8987 2499
rect 5549 2397 5583 2431
rect 9505 2397 9539 2431
rect 6653 2329 6687 2363
rect 9137 2329 9171 2363
rect 4997 2261 5031 2295
rect 5273 2261 5307 2295
rect 6285 2261 6319 2295
<< metal1 >>
rect 7190 12588 7196 12640
rect 7248 12628 7254 12640
rect 14366 12628 14372 12640
rect 7248 12600 14372 12628
rect 7248 12588 7254 12600
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 6730 12520 6736 12572
rect 6788 12560 6794 12572
rect 14274 12560 14280 12572
rect 6788 12532 14280 12560
rect 6788 12520 6794 12532
rect 14274 12520 14280 12532
rect 14332 12520 14338 12572
rect 5902 12452 5908 12504
rect 5960 12492 5966 12504
rect 14182 12492 14188 12504
rect 5960 12464 14188 12492
rect 5960 12452 5966 12464
rect 14182 12452 14188 12464
rect 14240 12452 14246 12504
rect 5626 11500 5632 11552
rect 5684 11540 5690 11552
rect 14274 11540 14280 11552
rect 5684 11512 14280 11540
rect 5684 11500 5690 11512
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 920 11450 9844 11472
rect 920 11398 2898 11450
rect 2950 11398 2962 11450
rect 3014 11398 3026 11450
rect 3078 11398 3090 11450
rect 3142 11398 6098 11450
rect 6150 11398 6162 11450
rect 6214 11398 6226 11450
rect 6278 11398 6290 11450
rect 6342 11398 9298 11450
rect 9350 11398 9362 11450
rect 9414 11398 9426 11450
rect 9478 11398 9490 11450
rect 9542 11398 9844 11450
rect 920 11376 9844 11398
rect 5626 11336 5632 11348
rect 5587 11308 5632 11336
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 6181 11339 6239 11345
rect 6181 11305 6193 11339
rect 6227 11305 6239 11339
rect 6730 11336 6736 11348
rect 6691 11308 6736 11336
rect 6181 11299 6239 11305
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11169 5503 11203
rect 5902 11200 5908 11212
rect 5863 11172 5908 11200
rect 5445 11163 5503 11169
rect 5460 11132 5488 11163
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 5994 11160 6000 11212
rect 6052 11200 6058 11212
rect 6052 11172 6097 11200
rect 6052 11160 6058 11172
rect 6196 11132 6224 11299
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 6840 11308 9352 11336
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11200 6607 11203
rect 6748 11200 6776 11296
rect 6595 11172 6776 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 6840 11132 6868 11308
rect 7190 11268 7196 11280
rect 7151 11240 7196 11268
rect 7190 11228 7196 11240
rect 7248 11228 7254 11280
rect 8754 11268 8760 11280
rect 7484 11240 8760 11268
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 7484 11200 7512 11240
rect 8754 11228 8760 11240
rect 8812 11228 8818 11280
rect 9324 11277 9352 11308
rect 9309 11271 9367 11277
rect 9309 11237 9321 11271
rect 9355 11237 9367 11271
rect 9309 11231 9367 11237
rect 7055 11172 7512 11200
rect 7561 11203 7619 11209
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 7561 11169 7573 11203
rect 7607 11200 7619 11203
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 7607 11172 7849 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 7837 11169 7849 11172
rect 7883 11200 7895 11203
rect 8665 11203 8723 11209
rect 7883 11172 8616 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 5460 11104 5856 11132
rect 6196 11104 6868 11132
rect 5718 11064 5724 11076
rect 5679 11036 5724 11064
rect 5718 11024 5724 11036
rect 5776 11024 5782 11076
rect 5828 10996 5856 11104
rect 6914 11092 6920 11144
rect 6972 11132 6978 11144
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 6972 11104 7941 11132
rect 6972 11092 6978 11104
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 8588 11132 8616 11172
rect 8665 11169 8677 11203
rect 8711 11200 8723 11203
rect 9122 11200 9128 11212
rect 8711 11172 9128 11200
rect 8711 11169 8723 11172
rect 8665 11163 8723 11169
rect 9122 11160 9128 11172
rect 9180 11160 9186 11212
rect 14182 11160 14188 11212
rect 14240 11160 14246 11212
rect 14200 11132 14228 11160
rect 8588 11104 14228 11132
rect 7929 11095 7987 11101
rect 5902 11024 5908 11076
rect 5960 11064 5966 11076
rect 6365 11067 6423 11073
rect 6365 11064 6377 11067
rect 5960 11036 6377 11064
rect 5960 11024 5966 11036
rect 6365 11033 6377 11036
rect 6411 11033 6423 11067
rect 6365 11027 6423 11033
rect 7098 11024 7104 11076
rect 7156 11064 7162 11076
rect 7653 11067 7711 11073
rect 7653 11064 7665 11067
rect 7156 11036 7665 11064
rect 7156 11024 7162 11036
rect 7653 11033 7665 11036
rect 7699 11033 7711 11067
rect 7653 11027 7711 11033
rect 8573 11067 8631 11073
rect 8573 11033 8585 11067
rect 8619 11064 8631 11067
rect 9030 11064 9036 11076
rect 8619 11036 9036 11064
rect 8619 11033 8631 11036
rect 8573 11027 8631 11033
rect 9030 11024 9036 11036
rect 9088 11024 9094 11076
rect 9493 11067 9551 11073
rect 9493 11033 9505 11067
rect 9539 11064 9551 11067
rect 14182 11064 14188 11076
rect 9539 11036 14188 11064
rect 9539 11033 9551 11036
rect 9493 11027 9551 11033
rect 14182 11024 14188 11036
rect 14240 11024 14246 11076
rect 8202 10996 8208 11008
rect 5828 10968 8208 10996
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 8846 10996 8852 11008
rect 8807 10968 8852 10996
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 920 10906 9844 10928
rect 920 10854 1298 10906
rect 1350 10854 1362 10906
rect 1414 10854 1426 10906
rect 1478 10854 1490 10906
rect 1542 10854 4498 10906
rect 4550 10854 4562 10906
rect 4614 10854 4626 10906
rect 4678 10854 4690 10906
rect 4742 10854 7698 10906
rect 7750 10854 7762 10906
rect 7814 10854 7826 10906
rect 7878 10854 7890 10906
rect 7942 10854 9844 10906
rect 920 10832 9844 10854
rect 5994 10792 6000 10804
rect 5955 10764 6000 10792
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 8202 10752 8208 10804
rect 8260 10792 8266 10804
rect 9125 10795 9183 10801
rect 9125 10792 9137 10795
rect 8260 10764 9137 10792
rect 8260 10752 8266 10764
rect 9125 10761 9137 10764
rect 9171 10761 9183 10795
rect 9125 10755 9183 10761
rect 8757 10727 8815 10733
rect 8757 10693 8769 10727
rect 8803 10724 8815 10727
rect 14366 10724 14372 10736
rect 8803 10696 14372 10724
rect 8803 10693 8815 10696
rect 8757 10687 8815 10693
rect 14366 10684 14372 10696
rect 14424 10684 14430 10736
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 7098 10656 7104 10668
rect 6779 10628 7104 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 8036 10628 9168 10656
rect 5810 10588 5816 10600
rect 5771 10560 5816 10588
rect 5810 10548 5816 10560
rect 5868 10548 5874 10600
rect 6457 10591 6515 10597
rect 6457 10557 6469 10591
rect 6503 10557 6515 10591
rect 6457 10551 6515 10557
rect 6472 10520 6500 10551
rect 6638 10520 6644 10532
rect 6472 10492 6644 10520
rect 6638 10480 6644 10492
rect 6696 10480 6702 10532
rect 7190 10480 7196 10532
rect 7248 10480 7254 10532
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 8036 10452 8064 10628
rect 9140 10600 9168 10628
rect 8938 10588 8944 10600
rect 8899 10560 8944 10588
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 9122 10548 9128 10600
rect 9180 10588 9186 10600
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 9180 10560 9321 10588
rect 9180 10548 9186 10560
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 8386 10480 8392 10532
rect 8444 10520 8450 10532
rect 8573 10523 8631 10529
rect 8573 10520 8585 10523
rect 8444 10492 8585 10520
rect 8444 10480 8450 10492
rect 8573 10489 8585 10492
rect 8619 10489 8631 10523
rect 8573 10483 8631 10489
rect 8202 10452 8208 10464
rect 5408 10424 8064 10452
rect 8163 10424 8208 10452
rect 5408 10412 5414 10424
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 9493 10455 9551 10461
rect 9493 10421 9505 10455
rect 9539 10452 9551 10455
rect 9582 10452 9588 10464
rect 9539 10424 9588 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 920 10362 9844 10384
rect 920 10310 2898 10362
rect 2950 10310 2962 10362
rect 3014 10310 3026 10362
rect 3078 10310 3090 10362
rect 3142 10310 6098 10362
rect 6150 10310 6162 10362
rect 6214 10310 6226 10362
rect 6278 10310 6290 10362
rect 6342 10310 9298 10362
rect 9350 10310 9362 10362
rect 9414 10310 9426 10362
rect 9478 10310 9490 10362
rect 9542 10310 9844 10362
rect 920 10288 9844 10310
rect 5813 10251 5871 10257
rect 5813 10217 5825 10251
rect 5859 10248 5871 10251
rect 7190 10248 7196 10260
rect 5859 10220 7196 10248
rect 5859 10217 5871 10220
rect 5813 10211 5871 10217
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 7300 10220 8984 10248
rect 6730 10180 6736 10192
rect 5920 10152 6736 10180
rect 5350 10112 5356 10124
rect 5311 10084 5356 10112
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 5920 10121 5948 10152
rect 6730 10140 6736 10152
rect 6788 10140 6794 10192
rect 6914 10180 6920 10192
rect 6875 10152 6920 10180
rect 6914 10140 6920 10152
rect 6972 10140 6978 10192
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10112 5687 10115
rect 5905 10115 5963 10121
rect 5905 10112 5917 10115
rect 5675 10084 5917 10112
rect 5675 10081 5687 10084
rect 5629 10075 5687 10081
rect 5905 10081 5917 10084
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6273 10115 6331 10121
rect 6273 10112 6285 10115
rect 6052 10084 6285 10112
rect 6052 10072 6058 10084
rect 6273 10081 6285 10084
rect 6319 10112 6331 10115
rect 7009 10115 7067 10121
rect 7009 10112 7021 10115
rect 6319 10084 7021 10112
rect 6319 10081 6331 10084
rect 6273 10075 6331 10081
rect 7009 10081 7021 10084
rect 7055 10081 7067 10115
rect 7009 10075 7067 10081
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10112 7251 10115
rect 7300 10112 7328 10220
rect 8846 10140 8852 10192
rect 8904 10140 8910 10192
rect 7239 10084 7328 10112
rect 7469 10115 7527 10121
rect 7239 10081 7251 10084
rect 7193 10075 7251 10081
rect 7469 10081 7481 10115
rect 7515 10112 7527 10115
rect 7558 10112 7564 10124
rect 7515 10084 7564 10112
rect 7515 10081 7527 10084
rect 7469 10075 7527 10081
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 7208 10044 7236 10075
rect 6696 10016 7236 10044
rect 6696 10004 6702 10016
rect 7282 10004 7288 10056
rect 7340 10044 7346 10056
rect 7484 10044 7512 10075
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 8956 10056 8984 10220
rect 7340 10016 7512 10044
rect 7837 10047 7895 10053
rect 7340 10004 7346 10016
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 8202 10044 8208 10056
rect 7883 10016 8208 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8938 10004 8944 10056
rect 8996 10004 9002 10056
rect 5537 9979 5595 9985
rect 5537 9945 5549 9979
rect 5583 9976 5595 9979
rect 6730 9976 6736 9988
rect 5583 9948 6736 9976
rect 5583 9945 5595 9948
rect 5537 9939 5595 9945
rect 6730 9936 6736 9948
rect 6788 9936 6794 9988
rect 6089 9911 6147 9917
rect 6089 9877 6101 9911
rect 6135 9908 6147 9911
rect 6454 9908 6460 9920
rect 6135 9880 6460 9908
rect 6135 9877 6147 9880
rect 6089 9871 6147 9877
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 6546 9868 6552 9920
rect 6604 9908 6610 9920
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 6604 9880 7297 9908
rect 6604 9868 6610 9880
rect 7285 9877 7297 9880
rect 7331 9877 7343 9911
rect 7285 9871 7343 9877
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 9263 9911 9321 9917
rect 9263 9908 9275 9911
rect 7524 9880 9275 9908
rect 7524 9868 7530 9880
rect 9263 9877 9275 9880
rect 9309 9877 9321 9911
rect 14274 9908 14280 9920
rect 9263 9871 9321 9877
rect 12406 9880 14280 9908
rect 920 9818 9844 9840
rect 920 9766 1298 9818
rect 1350 9766 1362 9818
rect 1414 9766 1426 9818
rect 1478 9766 1490 9818
rect 1542 9766 4498 9818
rect 4550 9766 4562 9818
rect 4614 9766 4626 9818
rect 4678 9766 4690 9818
rect 4742 9766 7698 9818
rect 7750 9766 7762 9818
rect 7814 9766 7826 9818
rect 7878 9766 7890 9818
rect 7942 9766 9844 9818
rect 920 9744 9844 9766
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 4893 9707 4951 9713
rect 4893 9704 4905 9707
rect 4396 9676 4905 9704
rect 4396 9664 4402 9676
rect 4893 9673 4905 9676
rect 4939 9704 4951 9707
rect 5350 9704 5356 9716
rect 4939 9676 5356 9704
rect 4939 9673 4951 9676
rect 4893 9667 4951 9673
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 5905 9707 5963 9713
rect 5905 9704 5917 9707
rect 5868 9676 5917 9704
rect 5868 9664 5874 9676
rect 5905 9673 5917 9676
rect 5951 9673 5963 9707
rect 5905 9667 5963 9673
rect 6546 9664 6552 9716
rect 6604 9664 6610 9716
rect 6748 9676 7972 9704
rect 6564 9636 6592 9664
rect 4724 9608 6592 9636
rect 4724 9509 4752 9608
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 5859 9540 6561 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 6549 9537 6561 9540
rect 6595 9568 6607 9571
rect 6748 9568 6776 9676
rect 7944 9636 7972 9676
rect 8018 9664 8024 9716
rect 8076 9704 8082 9716
rect 12406 9704 12434 9880
rect 14274 9868 14280 9880
rect 14332 9868 14338 9920
rect 8076 9676 12434 9704
rect 8076 9664 8082 9676
rect 7944 9608 12434 9636
rect 6595 9540 6776 9568
rect 6917 9571 6975 9577
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 6917 9537 6929 9571
rect 6963 9568 6975 9571
rect 8202 9568 8208 9580
rect 6963 9540 8208 9568
rect 6963 9537 6975 9540
rect 6917 9531 6975 9537
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 8938 9528 8944 9580
rect 8996 9568 9002 9580
rect 9493 9571 9551 9577
rect 9493 9568 9505 9571
rect 8996 9540 9505 9568
rect 8996 9528 9002 9540
rect 9493 9537 9505 9540
rect 9539 9537 9551 9571
rect 12406 9568 12434 9608
rect 14182 9568 14188 9580
rect 12406 9540 14188 9568
rect 9493 9531 9551 9537
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 4985 9503 5043 9509
rect 4985 9469 4997 9503
rect 5031 9500 5043 9503
rect 5074 9500 5080 9512
rect 5031 9472 5080 9500
rect 5031 9469 5043 9472
rect 4985 9463 5043 9469
rect 5074 9460 5080 9472
rect 5132 9500 5138 9512
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 5132 9472 5273 9500
rect 5132 9460 5138 9472
rect 5261 9469 5273 9472
rect 5307 9469 5319 9503
rect 5261 9463 5319 9469
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 6638 9500 6644 9512
rect 5592 9472 6644 9500
rect 5592 9460 5598 9472
rect 6638 9460 6644 9472
rect 6696 9460 6702 9512
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 7006 9432 7012 9444
rect 5460 9404 7012 9432
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5258 9364 5264 9376
rect 5215 9336 5264 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5460 9373 5488 9404
rect 7006 9392 7012 9404
rect 7064 9392 7070 9444
rect 5445 9367 5503 9373
rect 5445 9333 5457 9367
rect 5491 9333 5503 9367
rect 5445 9327 5503 9333
rect 6454 9324 6460 9376
rect 6512 9364 6518 9376
rect 7392 9364 7420 9418
rect 8294 9392 8300 9444
rect 8352 9432 8358 9444
rect 8573 9435 8631 9441
rect 8573 9432 8585 9435
rect 8352 9404 8585 9432
rect 8352 9392 8358 9404
rect 8573 9401 8585 9404
rect 8619 9401 8631 9435
rect 8573 9395 8631 9401
rect 8757 9435 8815 9441
rect 8757 9401 8769 9435
rect 8803 9432 8815 9435
rect 14274 9432 14280 9444
rect 8803 9404 14280 9432
rect 8803 9401 8815 9404
rect 8757 9395 8815 9401
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 6512 9336 7420 9364
rect 6512 9324 6518 9336
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 7616 9336 8401 9364
rect 7616 9324 7622 9336
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 8389 9327 8447 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 920 9274 9844 9296
rect 920 9222 2898 9274
rect 2950 9222 2962 9274
rect 3014 9222 3026 9274
rect 3078 9222 3090 9274
rect 3142 9222 6098 9274
rect 6150 9222 6162 9274
rect 6214 9222 6226 9274
rect 6278 9222 6290 9274
rect 6342 9222 9298 9274
rect 9350 9222 9362 9274
rect 9414 9222 9426 9274
rect 9478 9222 9490 9274
rect 9542 9222 9844 9274
rect 920 9200 9844 9222
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 5077 9163 5135 9169
rect 5077 9160 5089 9163
rect 4856 9132 5089 9160
rect 4856 9120 4862 9132
rect 5077 9129 5089 9132
rect 5123 9160 5135 9163
rect 5534 9160 5540 9172
rect 5123 9132 5540 9160
rect 5123 9129 5135 9132
rect 5077 9123 5135 9129
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 5721 9163 5779 9169
rect 5721 9129 5733 9163
rect 5767 9160 5779 9163
rect 5902 9160 5908 9172
rect 5767 9132 5908 9160
rect 5767 9129 5779 9132
rect 5721 9123 5779 9129
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 9493 9163 9551 9169
rect 9493 9160 9505 9163
rect 7116 9132 9505 9160
rect 5813 9095 5871 9101
rect 5813 9061 5825 9095
rect 5859 9092 5871 9095
rect 6454 9092 6460 9104
rect 5859 9064 6460 9092
rect 5859 9061 5871 9064
rect 5813 9055 5871 9061
rect 6454 9052 6460 9064
rect 6512 9052 6518 9104
rect 5166 8984 5172 9036
rect 5224 9024 5230 9036
rect 5261 9027 5319 9033
rect 5261 9024 5273 9027
rect 5224 8996 5273 9024
rect 5224 8984 5230 8996
rect 5261 8993 5273 8996
rect 5307 8993 5319 9027
rect 5261 8987 5319 8993
rect 6273 9027 6331 9033
rect 6273 8993 6285 9027
rect 6319 9024 6331 9027
rect 6362 9024 6368 9036
rect 6319 8996 6368 9024
rect 6319 8993 6331 8996
rect 6273 8987 6331 8993
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 6641 9027 6699 9033
rect 6641 8993 6653 9027
rect 6687 9024 6699 9027
rect 7116 9024 7144 9132
rect 9493 9129 9505 9132
rect 9539 9129 9551 9163
rect 14182 9160 14188 9172
rect 9493 9123 9551 9129
rect 12406 9132 14188 9160
rect 7377 9095 7435 9101
rect 7377 9061 7389 9095
rect 7423 9092 7435 9095
rect 7650 9092 7656 9104
rect 7423 9064 7656 9092
rect 7423 9061 7435 9064
rect 7377 9055 7435 9061
rect 7650 9052 7656 9064
rect 7708 9052 7714 9104
rect 8021 9095 8079 9101
rect 8021 9061 8033 9095
rect 8067 9092 8079 9095
rect 8110 9092 8116 9104
rect 8067 9064 8116 9092
rect 8067 9061 8079 9064
rect 8021 9055 8079 9061
rect 8110 9052 8116 9064
rect 8168 9052 8174 9104
rect 9582 9092 9588 9104
rect 9246 9064 9588 9092
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 6687 8996 7144 9024
rect 6687 8993 6699 8996
rect 6641 8987 6699 8993
rect 7190 8984 7196 9036
rect 7248 9024 7254 9036
rect 7285 9027 7343 9033
rect 7285 9024 7297 9027
rect 7248 8996 7297 9024
rect 7248 8984 7254 8996
rect 7285 8993 7297 8996
rect 7331 8993 7343 9027
rect 7742 9024 7748 9036
rect 7703 8996 7748 9024
rect 7285 8987 7343 8993
rect 7742 8984 7748 8996
rect 7800 8984 7806 9036
rect 5994 8956 6000 8968
rect 5955 8928 6000 8956
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 7466 8956 7472 8968
rect 7427 8928 7472 8956
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 12406 8956 12434 9132
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 7852 8928 12434 8956
rect 6825 8891 6883 8897
rect 6825 8857 6837 8891
rect 6871 8888 6883 8891
rect 7852 8888 7880 8928
rect 6871 8860 7880 8888
rect 6871 8857 6883 8860
rect 6825 8851 6883 8857
rect 5350 8820 5356 8832
rect 5311 8792 5356 8820
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 6457 8823 6515 8829
rect 6457 8820 6469 8823
rect 5960 8792 6469 8820
rect 5960 8780 5966 8792
rect 6457 8789 6469 8792
rect 6503 8789 6515 8823
rect 6457 8783 6515 8789
rect 6917 8823 6975 8829
rect 6917 8789 6929 8823
rect 6963 8820 6975 8823
rect 8570 8820 8576 8832
rect 6963 8792 8576 8820
rect 6963 8789 6975 8792
rect 6917 8783 6975 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 920 8730 9844 8752
rect 920 8678 1298 8730
rect 1350 8678 1362 8730
rect 1414 8678 1426 8730
rect 1478 8678 1490 8730
rect 1542 8678 4498 8730
rect 4550 8678 4562 8730
rect 4614 8678 4626 8730
rect 4678 8678 4690 8730
rect 4742 8678 7698 8730
rect 7750 8678 7762 8730
rect 7814 8678 7826 8730
rect 7878 8678 7890 8730
rect 7942 8678 9844 8730
rect 920 8656 9844 8678
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 8294 8616 8300 8628
rect 5408 8588 8156 8616
rect 8255 8588 8300 8616
rect 5408 8576 5414 8588
rect 4617 8551 4675 8557
rect 4617 8517 4629 8551
rect 4663 8517 4675 8551
rect 4617 8511 4675 8517
rect 4632 8480 4660 8511
rect 6454 8480 6460 8492
rect 4632 8452 6316 8480
rect 6367 8452 6460 8480
rect 4154 8372 4160 8424
rect 4212 8412 4218 8424
rect 4338 8412 4344 8424
rect 4212 8384 4344 8412
rect 4212 8372 4218 8384
rect 4338 8372 4344 8384
rect 4396 8412 4402 8424
rect 4433 8415 4491 8421
rect 4433 8412 4445 8415
rect 4396 8384 4445 8412
rect 4396 8372 4402 8384
rect 4433 8381 4445 8384
rect 4479 8381 4491 8415
rect 4706 8412 4712 8424
rect 4667 8384 4712 8412
rect 4433 8375 4491 8381
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 4982 8344 4988 8356
rect 4943 8316 4988 8344
rect 4982 8304 4988 8316
rect 5040 8304 5046 8356
rect 5258 8304 5264 8356
rect 5316 8344 5322 8356
rect 6288 8344 6316 8452
rect 6454 8440 6460 8452
rect 6512 8480 6518 8492
rect 6825 8483 6883 8489
rect 6825 8480 6837 8483
rect 6512 8452 6837 8480
rect 6512 8440 6518 8452
rect 6825 8449 6837 8452
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 8128 8480 8156 8588
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 9125 8619 9183 8625
rect 9125 8616 9137 8619
rect 8404 8588 9137 8616
rect 8202 8508 8208 8560
rect 8260 8548 8266 8560
rect 8404 8548 8432 8588
rect 9125 8585 9137 8588
rect 9171 8585 9183 8619
rect 9125 8579 9183 8585
rect 8260 8520 8432 8548
rect 8757 8551 8815 8557
rect 8260 8508 8266 8520
rect 8757 8517 8769 8551
rect 8803 8548 8815 8551
rect 14182 8548 14188 8560
rect 8803 8520 14188 8548
rect 8803 8517 8815 8520
rect 8757 8511 8815 8517
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 6972 8452 8064 8480
rect 8128 8452 9352 8480
rect 6972 8440 6978 8452
rect 6546 8412 6552 8424
rect 6507 8384 6552 8412
rect 6546 8372 6552 8384
rect 6604 8372 6610 8424
rect 8036 8412 8064 8452
rect 8570 8412 8576 8424
rect 8036 8384 8432 8412
rect 8531 8384 8576 8412
rect 5316 8316 5474 8344
rect 6288 8316 6684 8344
rect 5316 8304 5322 8316
rect 6656 8276 6684 8316
rect 6730 8304 6736 8356
rect 6788 8344 6794 8356
rect 8404 8344 8432 8384
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 9324 8421 9352 8452
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 8956 8344 8984 8375
rect 6788 8316 7314 8344
rect 8404 8316 8984 8344
rect 9493 8347 9551 8353
rect 6788 8304 6794 8316
rect 9493 8313 9505 8347
rect 9539 8344 9551 8347
rect 14274 8344 14280 8356
rect 9539 8316 14280 8344
rect 9539 8313 9551 8316
rect 9493 8307 9551 8313
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 6914 8276 6920 8288
rect 6656 8248 6920 8276
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 920 8186 9844 8208
rect 920 8134 2898 8186
rect 2950 8134 2962 8186
rect 3014 8134 3026 8186
rect 3078 8134 3090 8186
rect 3142 8134 6098 8186
rect 6150 8134 6162 8186
rect 6214 8134 6226 8186
rect 6278 8134 6290 8186
rect 6342 8134 9298 8186
rect 9350 8134 9362 8186
rect 9414 8134 9426 8186
rect 9478 8134 9490 8186
rect 9542 8134 9844 8186
rect 920 8112 9844 8134
rect 8018 8072 8024 8084
rect 4356 8044 8024 8072
rect 4356 8013 4384 8044
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 4341 8007 4399 8013
rect 4341 7973 4353 8007
rect 4387 7973 4399 8007
rect 4341 7967 4399 7973
rect 6454 7964 6460 8016
rect 6512 8004 6518 8016
rect 6549 8007 6607 8013
rect 6549 8004 6561 8007
rect 6512 7976 6561 8004
rect 6512 7964 6518 7976
rect 6549 7973 6561 7976
rect 6595 7973 6607 8007
rect 6549 7967 6607 7973
rect 7006 7964 7012 8016
rect 7064 7964 7070 8016
rect 8754 8004 8760 8016
rect 8715 7976 8760 8004
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 3786 7896 3792 7948
rect 3844 7936 3850 7948
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 3844 7908 4077 7936
rect 3844 7896 3850 7908
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 4080 7868 4108 7899
rect 5534 7896 5540 7948
rect 5592 7936 5598 7948
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 5592 7908 6285 7936
rect 5592 7896 5598 7908
rect 6273 7905 6285 7908
rect 6319 7905 6331 7939
rect 8849 7939 8907 7945
rect 8849 7936 8861 7939
rect 6273 7899 6331 7905
rect 7760 7908 8861 7936
rect 5902 7868 5908 7880
rect 4080 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 7760 7868 7788 7908
rect 8849 7905 8861 7908
rect 8895 7905 8907 7939
rect 8849 7899 8907 7905
rect 9309 7939 9367 7945
rect 9309 7905 9321 7939
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 6380 7840 7788 7868
rect 4249 7803 4307 7809
rect 4249 7769 4261 7803
rect 4295 7800 4307 7803
rect 5074 7800 5080 7812
rect 4295 7772 5080 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 5074 7760 5080 7772
rect 5132 7760 5138 7812
rect 5534 7760 5540 7812
rect 5592 7800 5598 7812
rect 6380 7800 6408 7840
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 8076 7840 8125 7868
rect 8076 7828 8082 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 9324 7868 9352 7899
rect 8260 7840 9352 7868
rect 8260 7828 8266 7840
rect 5592 7772 6408 7800
rect 9493 7803 9551 7809
rect 5592 7760 5598 7772
rect 9493 7769 9505 7803
rect 9539 7800 9551 7803
rect 13998 7800 14004 7812
rect 9539 7772 14004 7800
rect 9539 7769 9551 7772
rect 9493 7763 9551 7769
rect 13998 7760 14004 7772
rect 14056 7760 14062 7812
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 5166 7732 5172 7744
rect 4396 7704 5172 7732
rect 4396 7692 4402 7704
rect 5166 7692 5172 7704
rect 5224 7732 5230 7744
rect 5629 7735 5687 7741
rect 5629 7732 5641 7735
rect 5224 7704 5641 7732
rect 5224 7692 5230 7704
rect 5629 7701 5641 7704
rect 5675 7701 5687 7735
rect 5629 7695 5687 7701
rect 7190 7692 7196 7744
rect 7248 7732 7254 7744
rect 8021 7735 8079 7741
rect 8021 7732 8033 7735
rect 7248 7704 8033 7732
rect 7248 7692 7254 7704
rect 8021 7701 8033 7704
rect 8067 7732 8079 7735
rect 8110 7732 8116 7744
rect 8067 7704 8116 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 920 7642 9844 7664
rect 920 7590 1298 7642
rect 1350 7590 1362 7642
rect 1414 7590 1426 7642
rect 1478 7590 1490 7642
rect 1542 7590 4498 7642
rect 4550 7590 4562 7642
rect 4614 7590 4626 7642
rect 4678 7590 4690 7642
rect 4742 7590 7698 7642
rect 7750 7590 7762 7642
rect 7814 7590 7826 7642
rect 7878 7590 7890 7642
rect 7942 7590 9844 7642
rect 920 7568 9844 7590
rect 7282 7528 7288 7540
rect 5736 7500 7288 7528
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7392 4767 7395
rect 5736 7392 5764 7500
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 9309 7531 9367 7537
rect 9309 7528 9321 7531
rect 9180 7500 9321 7528
rect 9180 7488 9186 7500
rect 9309 7497 9321 7500
rect 9355 7497 9367 7531
rect 9309 7491 9367 7497
rect 4755 7364 5764 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 6181 7395 6239 7401
rect 6181 7392 6193 7395
rect 6052 7364 6193 7392
rect 6052 7352 6058 7364
rect 6181 7361 6193 7364
rect 6227 7392 6239 7395
rect 6641 7395 6699 7401
rect 6641 7392 6653 7395
rect 6227 7364 6653 7392
rect 6227 7361 6239 7364
rect 6181 7355 6239 7361
rect 6641 7361 6653 7364
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 4154 7324 4160 7336
rect 4115 7296 4160 7324
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 4338 7284 4344 7336
rect 4396 7324 4402 7336
rect 4433 7327 4491 7333
rect 4433 7324 4445 7327
rect 4396 7296 4445 7324
rect 4396 7284 4402 7296
rect 4433 7293 4445 7296
rect 4479 7293 4491 7327
rect 4433 7287 4491 7293
rect 6365 7327 6423 7333
rect 6365 7293 6377 7327
rect 6411 7293 6423 7327
rect 6365 7287 6423 7293
rect 5166 7216 5172 7268
rect 5224 7216 5230 7268
rect 6380 7256 6408 7287
rect 8110 7284 8116 7336
rect 8168 7324 8174 7336
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 8168 7296 8217 7324
rect 8168 7284 8174 7296
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 9030 7324 9036 7336
rect 8991 7296 9036 7324
rect 8205 7287 8263 7293
rect 9030 7284 9036 7296
rect 9088 7284 9094 7336
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 9180 7296 9225 7324
rect 9180 7284 9186 7296
rect 6546 7256 6552 7268
rect 6012 7228 6316 7256
rect 6380 7228 6552 7256
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 6012 7188 6040 7228
rect 4387 7160 6040 7188
rect 6288 7188 6316 7228
rect 6546 7216 6552 7228
rect 6604 7216 6610 7268
rect 8573 7259 8631 7265
rect 7116 7188 7144 7242
rect 8573 7225 8585 7259
rect 8619 7225 8631 7259
rect 8573 7219 8631 7225
rect 8757 7259 8815 7265
rect 8757 7225 8769 7259
rect 8803 7256 8815 7259
rect 14182 7256 14188 7268
rect 8803 7228 14188 7256
rect 8803 7225 8815 7228
rect 8757 7219 8815 7225
rect 6288 7160 7144 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 7374 7148 7380 7200
rect 7432 7188 7438 7200
rect 8113 7191 8171 7197
rect 8113 7188 8125 7191
rect 7432 7160 8125 7188
rect 7432 7148 7438 7160
rect 8113 7157 8125 7160
rect 8159 7157 8171 7191
rect 8386 7188 8392 7200
rect 8347 7160 8392 7188
rect 8113 7151 8171 7157
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 8588 7188 8616 7219
rect 14182 7216 14188 7228
rect 14240 7216 14246 7268
rect 8938 7188 8944 7200
rect 8588 7160 8944 7188
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 920 7098 9844 7120
rect 920 7046 2898 7098
rect 2950 7046 2962 7098
rect 3014 7046 3026 7098
rect 3078 7046 3090 7098
rect 3142 7046 6098 7098
rect 6150 7046 6162 7098
rect 6214 7046 6226 7098
rect 6278 7046 6290 7098
rect 6342 7046 9298 7098
rect 9350 7046 9362 7098
rect 9414 7046 9426 7098
rect 9478 7046 9490 7098
rect 9542 7046 9844 7098
rect 920 7024 9844 7046
rect 4249 6987 4307 6993
rect 4249 6953 4261 6987
rect 4295 6953 4307 6987
rect 4249 6947 4307 6953
rect 4264 6916 4292 6947
rect 6546 6944 6552 6996
rect 6604 6984 6610 6996
rect 6604 6956 7052 6984
rect 6604 6944 6610 6956
rect 6730 6916 6736 6928
rect 4264 6888 5106 6916
rect 6380 6888 6736 6916
rect 3513 6851 3571 6857
rect 3513 6848 3525 6851
rect 3436 6820 3525 6848
rect 3436 6656 3464 6820
rect 3513 6817 3525 6820
rect 3559 6817 3571 6851
rect 3513 6811 3571 6817
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6848 3847 6851
rect 4062 6848 4068 6860
rect 3835 6820 4068 6848
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 5902 6808 5908 6860
rect 5960 6848 5966 6860
rect 6273 6851 6331 6857
rect 6273 6848 6285 6851
rect 5960 6820 6285 6848
rect 5960 6808 5966 6820
rect 6273 6817 6285 6820
rect 6319 6848 6331 6851
rect 6380 6848 6408 6888
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 7024 6857 7052 6956
rect 7466 6944 7472 6996
rect 7524 6984 7530 6996
rect 8018 6984 8024 6996
rect 7524 6956 8024 6984
rect 7524 6944 7530 6956
rect 8018 6944 8024 6956
rect 8076 6944 8082 6996
rect 8386 6876 8392 6928
rect 8444 6876 8450 6928
rect 8803 6919 8861 6925
rect 8803 6885 8815 6919
rect 8849 6916 8861 6919
rect 8849 6888 9076 6916
rect 8849 6885 8861 6888
rect 8803 6879 8861 6885
rect 9048 6860 9076 6888
rect 6549 6851 6607 6857
rect 6549 6848 6561 6851
rect 6319 6820 6408 6848
rect 6472 6820 6561 6848
rect 6319 6817 6331 6820
rect 6273 6811 6331 6817
rect 4338 6780 4344 6792
rect 4299 6752 4344 6780
rect 4338 6740 4344 6752
rect 4396 6740 4402 6792
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6780 4675 6783
rect 5994 6780 6000 6792
rect 4663 6752 6000 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 3697 6715 3755 6721
rect 3697 6681 3709 6715
rect 3743 6712 3755 6715
rect 4154 6712 4160 6724
rect 3743 6684 4160 6712
rect 3743 6681 3755 6684
rect 3697 6675 3755 6681
rect 4154 6672 4160 6684
rect 4212 6672 4218 6724
rect 5810 6672 5816 6724
rect 5868 6712 5874 6724
rect 6472 6721 6500 6820
rect 6549 6817 6561 6820
rect 6595 6817 6607 6851
rect 6549 6811 6607 6817
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6817 7067 6851
rect 8938 6848 8944 6860
rect 8899 6820 8944 6848
rect 7009 6811 7067 6817
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 9030 6808 9036 6860
rect 9088 6848 9094 6860
rect 9088 6820 9133 6848
rect 9088 6808 9094 6820
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 7558 6780 7564 6792
rect 7423 6752 7564 6780
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 6457 6715 6515 6721
rect 6457 6712 6469 6715
rect 5868 6684 6469 6712
rect 5868 6672 5874 6684
rect 6457 6681 6469 6684
rect 6503 6681 6515 6715
rect 6457 6675 6515 6681
rect 3418 6644 3424 6656
rect 3379 6616 3424 6644
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3973 6647 4031 6653
rect 3973 6613 3985 6647
rect 4019 6644 4031 6647
rect 5166 6644 5172 6656
rect 4019 6616 5172 6644
rect 4019 6613 4031 6616
rect 3973 6607 4031 6613
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 5994 6604 6000 6656
rect 6052 6644 6058 6656
rect 6089 6647 6147 6653
rect 6089 6644 6101 6647
rect 6052 6616 6101 6644
rect 6052 6604 6058 6616
rect 6089 6613 6101 6616
rect 6135 6613 6147 6647
rect 6089 6607 6147 6613
rect 6546 6604 6552 6656
rect 6604 6644 6610 6656
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 6604 6616 6745 6644
rect 6604 6604 6610 6616
rect 6733 6613 6745 6616
rect 6779 6613 6791 6647
rect 6733 6607 6791 6613
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 8812 6616 9137 6644
rect 8812 6604 8818 6616
rect 9125 6613 9137 6616
rect 9171 6613 9183 6647
rect 9125 6607 9183 6613
rect 920 6554 9844 6576
rect 920 6502 1298 6554
rect 1350 6502 1362 6554
rect 1414 6502 1426 6554
rect 1478 6502 1490 6554
rect 1542 6502 4498 6554
rect 4550 6502 4562 6554
rect 4614 6502 4626 6554
rect 4678 6502 4690 6554
rect 4742 6502 7698 6554
rect 7750 6502 7762 6554
rect 7814 6502 7826 6554
rect 7878 6502 7890 6554
rect 7942 6502 9844 6554
rect 920 6480 9844 6502
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 8113 6443 8171 6449
rect 3476 6412 7696 6440
rect 3476 6400 3482 6412
rect 7668 6372 7696 6412
rect 8113 6409 8125 6443
rect 8159 6440 8171 6443
rect 8938 6440 8944 6452
rect 8159 6412 8944 6440
rect 8159 6409 8171 6412
rect 8113 6403 8171 6409
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 14182 6440 14188 6452
rect 12406 6412 14188 6440
rect 12406 6372 12434 6412
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 7668 6344 12434 6372
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 5810 6304 5816 6316
rect 4120 6276 5816 6304
rect 4120 6264 4126 6276
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 6052 6276 6653 6304
rect 6052 6264 6058 6276
rect 6641 6273 6653 6276
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 8757 6307 8815 6313
rect 6788 6276 8248 6304
rect 6788 6264 6794 6276
rect 4154 6196 4160 6248
rect 4212 6236 4218 6248
rect 4249 6239 4307 6245
rect 4249 6236 4261 6239
rect 4212 6208 4261 6236
rect 4212 6196 4218 6208
rect 4249 6205 4261 6208
rect 4295 6205 4307 6239
rect 4522 6236 4528 6248
rect 4483 6208 4528 6236
rect 4249 6199 4307 6205
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 6362 6236 6368 6248
rect 6323 6208 6368 6236
rect 6362 6196 6368 6208
rect 6420 6196 6426 6248
rect 8220 6245 8248 6276
rect 8757 6273 8769 6307
rect 8803 6304 8815 6307
rect 14274 6304 14280 6316
rect 8803 6276 14280 6304
rect 8803 6273 8815 6276
rect 8757 6267 8815 6273
rect 14274 6264 14280 6276
rect 14332 6264 14338 6316
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6205 8263 6239
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8205 6199 8263 6205
rect 8404 6208 8953 6236
rect 4798 6168 4804 6180
rect 4759 6140 4804 6168
rect 4798 6128 4804 6140
rect 4856 6128 4862 6180
rect 4890 6128 4896 6180
rect 4948 6168 4954 6180
rect 4948 6140 5290 6168
rect 4948 6128 4954 6140
rect 6914 6128 6920 6180
rect 6972 6168 6978 6180
rect 6972 6140 7130 6168
rect 6972 6128 6978 6140
rect 8110 6128 8116 6180
rect 8168 6168 8174 6180
rect 8404 6168 8432 6208
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 9122 6196 9128 6248
rect 9180 6196 9186 6248
rect 9309 6239 9367 6245
rect 9309 6205 9321 6239
rect 9355 6236 9367 6239
rect 9582 6236 9588 6248
rect 9355 6208 9588 6236
rect 9355 6205 9367 6208
rect 9309 6199 9367 6205
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 8168 6140 8432 6168
rect 8168 6128 8174 6140
rect 4341 6103 4399 6109
rect 4341 6069 4353 6103
rect 4387 6100 4399 6103
rect 5534 6100 5540 6112
rect 4387 6072 5540 6100
rect 4387 6069 4399 6072
rect 4341 6063 4399 6069
rect 5534 6060 5540 6072
rect 5592 6060 5598 6112
rect 6273 6103 6331 6109
rect 6273 6069 6285 6103
rect 6319 6100 6331 6103
rect 8202 6100 8208 6112
rect 6319 6072 8208 6100
rect 6319 6069 6331 6072
rect 6273 6063 6331 6069
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 8404 6109 8432 6140
rect 8573 6171 8631 6177
rect 8573 6137 8585 6171
rect 8619 6168 8631 6171
rect 9140 6168 9168 6196
rect 8619 6140 9168 6168
rect 9493 6171 9551 6177
rect 8619 6137 8631 6140
rect 8573 6131 8631 6137
rect 9493 6137 9505 6171
rect 9539 6168 9551 6171
rect 14366 6168 14372 6180
rect 9539 6140 14372 6168
rect 9539 6137 9551 6140
rect 9493 6131 9551 6137
rect 14366 6128 14372 6140
rect 14424 6128 14430 6180
rect 8389 6103 8447 6109
rect 8389 6069 8401 6103
rect 8435 6069 8447 6103
rect 8389 6063 8447 6069
rect 9030 6060 9036 6112
rect 9088 6100 9094 6112
rect 9125 6103 9183 6109
rect 9125 6100 9137 6103
rect 9088 6072 9137 6100
rect 9088 6060 9094 6072
rect 9125 6069 9137 6072
rect 9171 6069 9183 6103
rect 9125 6063 9183 6069
rect 920 6010 9844 6032
rect 920 5958 2898 6010
rect 2950 5958 2962 6010
rect 3014 5958 3026 6010
rect 3078 5958 3090 6010
rect 3142 5958 6098 6010
rect 6150 5958 6162 6010
rect 6214 5958 6226 6010
rect 6278 5958 6290 6010
rect 6342 5958 9298 6010
rect 9350 5958 9362 6010
rect 9414 5958 9426 6010
rect 9478 5958 9490 6010
rect 9542 5958 9844 6010
rect 920 5936 9844 5958
rect 4249 5899 4307 5905
rect 4249 5865 4261 5899
rect 4295 5896 4307 5899
rect 4890 5896 4896 5908
rect 4295 5868 4896 5896
rect 4295 5865 4307 5868
rect 4249 5859 4307 5865
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 8110 5896 8116 5908
rect 5000 5868 8116 5896
rect 5000 5828 5028 5868
rect 6546 5828 6552 5840
rect 4080 5800 5028 5828
rect 5842 5800 6552 5828
rect 3786 5760 3792 5772
rect 3747 5732 3792 5760
rect 3786 5720 3792 5732
rect 3844 5720 3850 5772
rect 4080 5769 4108 5800
rect 6546 5788 6552 5800
rect 6604 5788 6610 5840
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 6270 5760 6276 5772
rect 5960 5732 6276 5760
rect 5960 5720 5966 5732
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 6748 5769 6776 5868
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 7374 5828 7380 5840
rect 7335 5800 7380 5828
rect 7374 5788 7380 5800
rect 7432 5788 7438 5840
rect 9030 5788 9036 5840
rect 9088 5788 9094 5840
rect 6733 5763 6791 5769
rect 6733 5729 6745 5763
rect 6779 5760 6791 5763
rect 7009 5763 7067 5769
rect 7009 5760 7021 5763
rect 6779 5732 7021 5760
rect 6779 5729 6791 5732
rect 6733 5723 6791 5729
rect 7009 5729 7021 5732
rect 7055 5729 7067 5763
rect 7009 5723 7067 5729
rect 7561 5763 7619 5769
rect 7561 5729 7573 5763
rect 7607 5760 7619 5763
rect 7607 5732 8156 5760
rect 7607 5729 7619 5732
rect 7561 5723 7619 5729
rect 4338 5692 4344 5704
rect 4251 5664 4344 5692
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5692 4675 5695
rect 5994 5692 6000 5704
rect 4663 5664 6000 5692
rect 4663 5661 4675 5664
rect 4617 5655 4675 5661
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 6454 5652 6460 5704
rect 6512 5692 6518 5704
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 6512 5664 7665 5692
rect 6512 5652 6518 5664
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 4356 5624 4384 5652
rect 6748 5636 6776 5664
rect 7653 5661 7665 5664
rect 7699 5661 7711 5695
rect 8018 5692 8024 5704
rect 7979 5664 8024 5692
rect 7653 5655 7711 5661
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 8128 5692 8156 5732
rect 14182 5692 14188 5704
rect 8128 5664 14188 5692
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 4120 5596 4384 5624
rect 4120 5584 4126 5596
rect 6730 5584 6736 5636
rect 6788 5584 6794 5636
rect 3973 5559 4031 5565
rect 3973 5525 3985 5559
rect 4019 5556 4031 5559
rect 4338 5556 4344 5568
rect 4019 5528 4344 5556
rect 4019 5525 4031 5528
rect 3973 5519 4031 5525
rect 4338 5516 4344 5528
rect 4396 5516 4402 5568
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 6089 5559 6147 5565
rect 6089 5556 6101 5559
rect 4856 5528 6101 5556
rect 4856 5516 4862 5528
rect 6089 5525 6101 5528
rect 6135 5525 6147 5559
rect 6454 5556 6460 5568
rect 6415 5528 6460 5556
rect 6089 5519 6147 5525
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 6917 5559 6975 5565
rect 6917 5525 6929 5559
rect 6963 5556 6975 5559
rect 7006 5556 7012 5568
rect 6963 5528 7012 5556
rect 6963 5525 6975 5528
rect 6917 5519 6975 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7193 5559 7251 5565
rect 7193 5525 7205 5559
rect 7239 5556 7251 5559
rect 7282 5556 7288 5568
rect 7239 5528 7288 5556
rect 7239 5525 7251 5528
rect 7193 5519 7251 5525
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 9447 5559 9505 5565
rect 9447 5556 9459 5559
rect 9180 5528 9459 5556
rect 9180 5516 9186 5528
rect 9447 5525 9459 5528
rect 9493 5525 9505 5559
rect 9447 5519 9505 5525
rect 920 5466 9844 5488
rect 920 5414 1298 5466
rect 1350 5414 1362 5466
rect 1414 5414 1426 5466
rect 1478 5414 1490 5466
rect 1542 5414 4498 5466
rect 4550 5414 4562 5466
rect 4614 5414 4626 5466
rect 4678 5414 4690 5466
rect 4742 5414 7698 5466
rect 7750 5414 7762 5466
rect 7814 5414 7826 5466
rect 7878 5414 7890 5466
rect 7942 5414 9844 5466
rect 920 5392 9844 5414
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 4396 5324 8248 5352
rect 4396 5312 4402 5324
rect 5718 5244 5724 5296
rect 5776 5284 5782 5296
rect 6089 5287 6147 5293
rect 6089 5284 6101 5287
rect 5776 5256 6101 5284
rect 5776 5244 5782 5256
rect 6089 5253 6101 5256
rect 6135 5253 6147 5287
rect 6089 5247 6147 5253
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 4706 5216 4712 5228
rect 4663 5188 4712 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6227 5188 6837 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 4246 5148 4252 5160
rect 4207 5120 4252 5148
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 4356 5024 4384 5111
rect 6270 5108 6276 5160
rect 6328 5148 6334 5160
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 6328 5120 6377 5148
rect 6328 5108 6334 5120
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 8220 5134 8248 5324
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 8849 5219 8907 5225
rect 8849 5216 8861 5219
rect 8352 5188 8861 5216
rect 8352 5176 8358 5188
rect 8849 5185 8861 5188
rect 8895 5185 8907 5219
rect 8849 5179 8907 5185
rect 6365 5111 6423 5117
rect 8662 5108 8668 5160
rect 8720 5148 8726 5160
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 8720 5120 9321 5148
rect 8720 5108 8726 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9309 5111 9367 5117
rect 6454 5080 6460 5092
rect 5842 5052 6460 5080
rect 6454 5040 6460 5052
rect 6512 5040 6518 5092
rect 7098 5080 7104 5092
rect 7059 5052 7104 5080
rect 7098 5040 7104 5052
rect 7156 5040 7162 5092
rect 9493 5083 9551 5089
rect 9493 5049 9505 5083
rect 9539 5080 9551 5083
rect 14182 5080 14188 5092
rect 9539 5052 14188 5080
rect 9539 5049 9551 5052
rect 9493 5043 9551 5049
rect 14182 5040 14188 5052
rect 14240 5040 14246 5092
rect 4062 5012 4068 5024
rect 3975 4984 4068 5012
rect 4062 4972 4068 4984
rect 4120 5012 4126 5024
rect 4338 5012 4344 5024
rect 4120 4984 4344 5012
rect 4120 4972 4126 4984
rect 4338 4972 4344 4984
rect 4396 5012 4402 5024
rect 6181 5015 6239 5021
rect 6181 5012 6193 5015
rect 4396 4984 6193 5012
rect 4396 4972 4402 4984
rect 6181 4981 6193 4984
rect 6227 4981 6239 5015
rect 6546 5012 6552 5024
rect 6507 4984 6552 5012
rect 6181 4975 6239 4981
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 920 4922 9844 4944
rect 920 4870 2898 4922
rect 2950 4870 2962 4922
rect 3014 4870 3026 4922
rect 3078 4870 3090 4922
rect 3142 4870 6098 4922
rect 6150 4870 6162 4922
rect 6214 4870 6226 4922
rect 6278 4870 6290 4922
rect 6342 4870 9298 4922
rect 9350 4870 9362 4922
rect 9414 4870 9426 4922
rect 9478 4870 9490 4922
rect 9542 4870 9844 4922
rect 920 4848 9844 4870
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 8343 4811 8401 4817
rect 4212 4780 8156 4808
rect 4212 4768 4218 4780
rect 6546 4740 6552 4752
rect 5842 4712 6552 4740
rect 6546 4700 6552 4712
rect 6604 4700 6610 4752
rect 7282 4700 7288 4752
rect 7340 4700 7346 4752
rect 4338 4672 4344 4684
rect 4299 4644 4344 4672
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 6178 4672 6184 4684
rect 6139 4644 6184 4672
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4604 4675 4607
rect 6549 4607 6607 4613
rect 4663 4576 5764 4604
rect 4663 4573 4675 4576
rect 4617 4567 4675 4573
rect 5736 4548 5764 4576
rect 6549 4573 6561 4607
rect 6595 4604 6607 4607
rect 6730 4604 6736 4616
rect 6595 4576 6736 4604
rect 6595 4573 6607 4576
rect 6549 4567 6607 4573
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 6914 4604 6920 4616
rect 6875 4576 6920 4604
rect 6914 4564 6920 4576
rect 6972 4604 6978 4616
rect 7098 4604 7104 4616
rect 6972 4576 7104 4604
rect 6972 4564 6978 4576
rect 7098 4564 7104 4576
rect 7156 4564 7162 4616
rect 8128 4604 8156 4780
rect 8343 4777 8355 4811
rect 8389 4808 8401 4811
rect 8846 4808 8852 4820
rect 8389 4780 8852 4808
rect 8389 4777 8401 4780
rect 8343 4771 8401 4777
rect 8846 4768 8852 4780
rect 8904 4808 8910 4820
rect 9582 4808 9588 4820
rect 8904 4780 9588 4808
rect 8904 4768 8910 4780
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 8754 4740 8760 4752
rect 8715 4712 8760 4740
rect 8754 4700 8760 4712
rect 8812 4700 8818 4752
rect 8665 4607 8723 4613
rect 8665 4604 8677 4607
rect 8128 4576 8677 4604
rect 8665 4573 8677 4576
rect 8711 4573 8723 4607
rect 9030 4604 9036 4616
rect 8991 4576 9036 4604
rect 8665 4567 8723 4573
rect 9030 4564 9036 4576
rect 9088 4564 9094 4616
rect 5718 4496 5724 4548
rect 5776 4496 5782 4548
rect 5994 4428 6000 4480
rect 6052 4468 6058 4480
rect 6089 4471 6147 4477
rect 6089 4468 6101 4471
rect 6052 4440 6101 4468
rect 6052 4428 6058 4440
rect 6089 4437 6101 4440
rect 6135 4437 6147 4471
rect 6089 4431 6147 4437
rect 6270 4428 6276 4480
rect 6328 4468 6334 4480
rect 6365 4471 6423 4477
rect 6365 4468 6377 4471
rect 6328 4440 6377 4468
rect 6328 4428 6334 4440
rect 6365 4437 6377 4440
rect 6411 4437 6423 4471
rect 6365 4431 6423 4437
rect 3220 4378 9844 4400
rect 3220 4326 4498 4378
rect 4550 4326 4562 4378
rect 4614 4326 4626 4378
rect 4678 4326 4690 4378
rect 4742 4326 7698 4378
rect 7750 4326 7762 4378
rect 7814 4326 7826 4378
rect 7878 4326 7890 4378
rect 7942 4326 9844 4378
rect 3220 4304 9844 4326
rect 4328 4267 4386 4273
rect 4328 4233 4340 4267
rect 4374 4264 4386 4267
rect 7098 4264 7104 4276
rect 4374 4236 7104 4264
rect 4374 4233 4386 4236
rect 4328 4227 4386 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4128 4123 4131
rect 4338 4128 4344 4140
rect 4111 4100 4344 4128
rect 4111 4097 4123 4100
rect 4065 4091 4123 4097
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 5074 4088 5080 4140
rect 5132 4128 5138 4140
rect 5132 4100 5580 4128
rect 5132 4088 5138 4100
rect 5552 4060 5580 4100
rect 5810 4088 5816 4140
rect 5868 4128 5874 4140
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 5868 4100 6929 4128
rect 5868 4088 5874 4100
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 8662 4128 8668 4140
rect 8623 4100 8668 4128
rect 6917 4091 6975 4097
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 9122 4128 9128 4140
rect 8772 4100 9128 4128
rect 5997 4063 6055 4069
rect 5997 4060 6009 4063
rect 5552 4032 6009 4060
rect 5997 4029 6009 4032
rect 6043 4060 6055 4063
rect 6178 4060 6184 4072
rect 6043 4032 6184 4060
rect 6043 4029 6055 4032
rect 5997 4023 6055 4029
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 6365 4063 6423 4069
rect 6365 4029 6377 4063
rect 6411 4060 6423 4063
rect 6546 4060 6552 4072
rect 6411 4032 6552 4060
rect 6411 4029 6423 4032
rect 6365 4023 6423 4029
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 8772 4069 8800 4100
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4029 6699 4063
rect 6641 4023 6699 4029
rect 8757 4063 8815 4069
rect 8757 4029 8769 4063
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 6270 3992 6276 4004
rect 5566 3964 6276 3992
rect 6270 3952 6276 3964
rect 6328 3952 6334 4004
rect 6454 3952 6460 4004
rect 6512 3992 6518 4004
rect 6656 3992 6684 4023
rect 8846 4020 8852 4072
rect 8904 4060 8910 4072
rect 8904 4032 8949 4060
rect 8904 4020 8910 4032
rect 6512 3964 6776 3992
rect 6512 3952 6518 3964
rect 6748 3936 6776 3964
rect 7006 3952 7012 4004
rect 7064 3992 7070 4004
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 7064 3964 7406 3992
rect 8772 3964 9321 3992
rect 7064 3952 7070 3964
rect 8772 3936 8800 3964
rect 9309 3961 9321 3964
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 9493 3995 9551 4001
rect 9493 3961 9505 3995
rect 9539 3992 9551 3995
rect 14182 3992 14188 4004
rect 9539 3964 14188 3992
rect 9539 3961 9551 3964
rect 9493 3955 9551 3961
rect 14182 3952 14188 3964
rect 14240 3952 14246 4004
rect 5810 3924 5816 3936
rect 5771 3896 5816 3924
rect 5810 3884 5816 3896
rect 5868 3884 5874 3936
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 6181 3927 6239 3933
rect 6181 3924 6193 3927
rect 5960 3896 6193 3924
rect 5960 3884 5966 3896
rect 6181 3893 6193 3896
rect 6227 3893 6239 3927
rect 6546 3924 6552 3936
rect 6507 3896 6552 3924
rect 6181 3887 6239 3893
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 6730 3884 6736 3936
rect 6788 3884 6794 3936
rect 8754 3884 8760 3936
rect 8812 3884 8818 3936
rect 9122 3924 9128 3936
rect 9083 3896 9128 3924
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 3220 3834 9844 3856
rect 3220 3782 6098 3834
rect 6150 3782 6162 3834
rect 6214 3782 6226 3834
rect 6278 3782 6290 3834
rect 6342 3782 9298 3834
rect 9350 3782 9362 3834
rect 9414 3782 9426 3834
rect 9478 3782 9490 3834
rect 9542 3782 9844 3834
rect 3220 3760 9844 3782
rect 5994 3720 6000 3732
rect 4632 3692 6000 3720
rect 4632 3661 4660 3692
rect 5994 3680 6000 3692
rect 6052 3720 6058 3732
rect 6052 3692 6500 3720
rect 6052 3680 6058 3692
rect 4617 3655 4675 3661
rect 4617 3621 4629 3655
rect 4663 3621 4675 3655
rect 5902 3652 5908 3664
rect 5842 3624 5908 3652
rect 4617 3615 4675 3621
rect 5902 3612 5908 3624
rect 5960 3612 5966 3664
rect 6472 3661 6500 3692
rect 8478 3680 8484 3732
rect 8536 3720 8542 3732
rect 8573 3723 8631 3729
rect 8573 3720 8585 3723
rect 8536 3692 8585 3720
rect 8536 3680 8542 3692
rect 8573 3689 8585 3692
rect 8619 3689 8631 3723
rect 8573 3683 8631 3689
rect 6457 3655 6515 3661
rect 6457 3621 6469 3655
rect 6503 3621 6515 3655
rect 6457 3615 6515 3621
rect 6546 3612 6552 3664
rect 6604 3652 6610 3664
rect 8389 3655 8447 3661
rect 6604 3624 6946 3652
rect 6604 3612 6610 3624
rect 8389 3621 8401 3655
rect 8435 3652 8447 3655
rect 14274 3652 14280 3664
rect 8435 3624 14280 3652
rect 8435 3621 8447 3624
rect 8389 3615 8447 3621
rect 14274 3612 14280 3624
rect 14332 3612 14338 3664
rect 4338 3584 4344 3596
rect 4299 3556 4344 3584
rect 4338 3544 4344 3556
rect 4396 3544 4402 3596
rect 8205 3587 8263 3593
rect 8205 3584 8217 3587
rect 7944 3556 8217 3584
rect 4982 3476 4988 3528
rect 5040 3516 5046 3528
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 5040 3488 6101 3516
rect 5040 3476 5046 3488
rect 6012 3380 6040 3488
rect 6089 3485 6101 3488
rect 6135 3485 6147 3519
rect 6089 3479 6147 3485
rect 6178 3476 6184 3528
rect 6236 3516 6242 3528
rect 6454 3516 6460 3528
rect 6236 3488 6460 3516
rect 6236 3476 6242 3488
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 7944 3525 7972 3556
rect 8205 3553 8217 3556
rect 8251 3553 8263 3587
rect 8938 3584 8944 3596
rect 8899 3556 8944 3584
rect 8205 3547 8263 3553
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 8570 3476 8576 3528
rect 8628 3516 8634 3528
rect 9033 3519 9091 3525
rect 9033 3516 9045 3519
rect 8628 3488 9045 3516
rect 8628 3476 8634 3488
rect 9033 3485 9045 3488
rect 9079 3485 9091 3519
rect 9033 3479 9091 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 8846 3408 8852 3460
rect 8904 3448 8910 3460
rect 9140 3448 9168 3479
rect 9582 3448 9588 3460
rect 8904 3420 9588 3448
rect 8904 3408 8910 3420
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 7006 3380 7012 3392
rect 6012 3352 7012 3380
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 3220 3290 9844 3312
rect 3220 3238 4498 3290
rect 4550 3238 4562 3290
rect 4614 3238 4626 3290
rect 4678 3238 4690 3290
rect 4742 3238 7698 3290
rect 7750 3238 7762 3290
rect 7814 3238 7826 3290
rect 7878 3238 7890 3290
rect 7942 3238 9844 3290
rect 3220 3216 9844 3238
rect 4338 3176 4344 3188
rect 4172 3148 4344 3176
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3040 4123 3043
rect 4172 3040 4200 3148
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 6914 3176 6920 3188
rect 5859 3148 6920 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 8570 3176 8576 3188
rect 8531 3148 8576 3176
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 4111 3012 4200 3040
rect 4341 3043 4399 3049
rect 4111 3009 4123 3012
rect 4065 3003 4123 3009
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 5810 3040 5816 3052
rect 4387 3012 5816 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 6086 3000 6092 3052
rect 6144 3040 6150 3052
rect 6273 3043 6331 3049
rect 6273 3040 6285 3043
rect 6144 3012 6285 3040
rect 6144 3000 6150 3012
rect 6273 3009 6285 3012
rect 6319 3009 6331 3043
rect 6273 3003 6331 3009
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 9122 3040 9128 3052
rect 7156 3012 8432 3040
rect 9083 3012 9128 3040
rect 7156 3000 7162 3012
rect 5994 2972 6000 2984
rect 5907 2944 6000 2972
rect 5994 2932 6000 2944
rect 6052 2972 6058 2984
rect 6178 2972 6184 2984
rect 6052 2944 6184 2972
rect 6052 2932 6058 2944
rect 6178 2932 6184 2944
rect 6236 2932 6242 2984
rect 5074 2864 5080 2916
rect 5132 2864 5138 2916
rect 5718 2864 5724 2916
rect 5776 2904 5782 2916
rect 6549 2907 6607 2913
rect 6549 2904 6561 2907
rect 5776 2876 6561 2904
rect 5776 2864 5782 2876
rect 6549 2873 6561 2876
rect 6595 2873 6607 2907
rect 6549 2867 6607 2873
rect 7006 2864 7012 2916
rect 7064 2864 7070 2916
rect 8297 2907 8355 2913
rect 8297 2873 8309 2907
rect 8343 2873 8355 2907
rect 8297 2867 8355 2873
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 6638 2836 6644 2848
rect 6227 2808 6644 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 8021 2839 8079 2845
rect 8021 2805 8033 2839
rect 8067 2836 8079 2839
rect 8312 2836 8340 2867
rect 8067 2808 8340 2836
rect 8404 2836 8432 3012
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 8996 2944 9045 2972
rect 8996 2932 9002 2944
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 8481 2907 8539 2913
rect 8481 2873 8493 2907
rect 8527 2904 8539 2907
rect 14182 2904 14188 2916
rect 8527 2876 14188 2904
rect 8527 2873 8539 2876
rect 8481 2867 8539 2873
rect 14182 2864 14188 2876
rect 14240 2864 14246 2916
rect 8941 2839 8999 2845
rect 8941 2836 8953 2839
rect 8404 2808 8953 2836
rect 8067 2805 8079 2808
rect 8021 2799 8079 2805
rect 8941 2805 8953 2808
rect 8987 2805 8999 2839
rect 8941 2799 8999 2805
rect 3220 2746 9844 2768
rect 3220 2694 6098 2746
rect 6150 2694 6162 2746
rect 6214 2694 6226 2746
rect 6278 2694 6290 2746
rect 6342 2694 9298 2746
rect 9350 2694 9362 2746
rect 9414 2694 9426 2746
rect 9478 2694 9490 2746
rect 9542 2694 9844 2746
rect 3220 2672 9844 2694
rect 4430 2632 4436 2644
rect 4391 2604 4436 2632
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 5721 2635 5779 2641
rect 5721 2601 5733 2635
rect 5767 2632 5779 2635
rect 6546 2632 6552 2644
rect 5767 2604 6552 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 6638 2592 6644 2644
rect 6696 2632 6702 2644
rect 8481 2635 8539 2641
rect 6696 2604 7512 2632
rect 6696 2592 6702 2604
rect 5353 2567 5411 2573
rect 5353 2533 5365 2567
rect 5399 2564 5411 2567
rect 5399 2536 6592 2564
rect 5399 2533 5411 2536
rect 5353 2527 5411 2533
rect 4617 2499 4675 2505
rect 4617 2465 4629 2499
rect 4663 2496 4675 2499
rect 4890 2496 4896 2508
rect 4663 2468 4896 2496
rect 4663 2465 4675 2468
rect 4617 2459 4675 2465
rect 4890 2456 4896 2468
rect 4948 2456 4954 2508
rect 5077 2499 5135 2505
rect 5077 2496 5089 2499
rect 5000 2468 5089 2496
rect 5000 2304 5028 2468
rect 5077 2465 5089 2468
rect 5123 2465 5135 2499
rect 5626 2496 5632 2508
rect 5587 2468 5632 2496
rect 5077 2459 5135 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6089 2499 6147 2505
rect 6089 2496 6101 2499
rect 6052 2468 6101 2496
rect 6052 2456 6058 2468
rect 6089 2465 6101 2468
rect 6135 2465 6147 2499
rect 6089 2459 6147 2465
rect 6457 2499 6515 2505
rect 6457 2465 6469 2499
rect 6503 2465 6515 2499
rect 6457 2459 6515 2465
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2428 5595 2431
rect 6472 2428 6500 2459
rect 5583 2400 6500 2428
rect 6564 2428 6592 2536
rect 6914 2524 6920 2576
rect 6972 2564 6978 2576
rect 7009 2567 7067 2573
rect 7009 2564 7021 2567
rect 6972 2536 7021 2564
rect 6972 2524 6978 2536
rect 7009 2533 7021 2536
rect 7055 2533 7067 2567
rect 7484 2550 7512 2604
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 8754 2632 8760 2644
rect 8527 2604 8760 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 7009 2527 7067 2533
rect 9030 2524 9036 2576
rect 9088 2564 9094 2576
rect 9309 2567 9367 2573
rect 9309 2564 9321 2567
rect 9088 2536 9321 2564
rect 9088 2524 9094 2536
rect 9309 2533 9321 2536
rect 9355 2533 9367 2567
rect 9309 2527 9367 2533
rect 6730 2496 6736 2508
rect 6691 2468 6736 2496
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 8941 2499 8999 2505
rect 8941 2465 8953 2499
rect 8987 2465 8999 2499
rect 8941 2459 8999 2465
rect 8956 2428 8984 2459
rect 6564 2400 8984 2428
rect 9493 2431 9551 2437
rect 5583 2397 5595 2400
rect 5537 2391 5595 2397
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 9539 2400 12434 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 6638 2360 6644 2372
rect 6599 2332 6644 2360
rect 6638 2320 6644 2332
rect 6696 2320 6702 2372
rect 9125 2363 9183 2369
rect 9125 2329 9137 2363
rect 9171 2360 9183 2363
rect 12406 2360 12434 2400
rect 14182 2360 14188 2372
rect 9171 2332 11008 2360
rect 12406 2332 14188 2360
rect 9171 2329 9183 2332
rect 9125 2323 9183 2329
rect 4982 2292 4988 2304
rect 4943 2264 4988 2292
rect 4982 2252 4988 2264
rect 5040 2252 5046 2304
rect 5258 2292 5264 2304
rect 5219 2264 5264 2292
rect 5258 2252 5264 2264
rect 5316 2252 5322 2304
rect 6273 2295 6331 2301
rect 6273 2261 6285 2295
rect 6319 2292 6331 2295
rect 7006 2292 7012 2304
rect 6319 2264 7012 2292
rect 6319 2261 6331 2264
rect 6273 2255 6331 2261
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 10980 2292 11008 2332
rect 14182 2320 14188 2332
rect 14240 2320 14246 2372
rect 14366 2292 14372 2304
rect 10980 2264 14372 2292
rect 14366 2252 14372 2264
rect 14424 2252 14430 2304
rect 3220 2202 9844 2224
rect 3220 2150 4498 2202
rect 4550 2150 4562 2202
rect 4614 2150 4626 2202
rect 4678 2150 4690 2202
rect 4742 2150 7698 2202
rect 7750 2150 7762 2202
rect 7814 2150 7826 2202
rect 7878 2150 7890 2202
rect 7942 2150 9844 2202
rect 3220 2128 9844 2150
rect 5626 2048 5632 2100
rect 5684 2088 5690 2100
rect 8662 2088 8668 2100
rect 5684 2060 8668 2088
rect 5684 2048 5690 2060
rect 8662 2048 8668 2060
rect 8720 2048 8726 2100
rect 4982 1980 4988 2032
rect 5040 2020 5046 2032
rect 14090 2020 14096 2032
rect 5040 1992 14096 2020
rect 5040 1980 5046 1992
rect 14090 1980 14096 1992
rect 14148 1980 14154 2032
rect 4890 1844 4896 1896
rect 4948 1884 4954 1896
rect 14274 1884 14280 1896
rect 4948 1856 14280 1884
rect 4948 1844 4954 1856
rect 14274 1844 14280 1856
rect 14332 1844 14338 1896
rect 5258 1776 5264 1828
rect 5316 1816 5322 1828
rect 9582 1816 9588 1828
rect 5316 1788 9588 1816
rect 5316 1776 5322 1788
rect 9582 1776 9588 1788
rect 9640 1776 9646 1828
rect 6638 8 6644 60
rect 6696 48 6702 60
rect 14182 48 14188 60
rect 6696 20 14188 48
rect 6696 8 6702 20
rect 14182 8 14188 20
rect 14240 8 14246 60
<< via1 >>
rect 7196 12588 7248 12640
rect 14372 12588 14424 12640
rect 6736 12520 6788 12572
rect 14280 12520 14332 12572
rect 5908 12452 5960 12504
rect 14188 12452 14240 12504
rect 5632 11500 5684 11552
rect 14280 11500 14332 11552
rect 2898 11398 2950 11450
rect 2962 11398 3014 11450
rect 3026 11398 3078 11450
rect 3090 11398 3142 11450
rect 6098 11398 6150 11450
rect 6162 11398 6214 11450
rect 6226 11398 6278 11450
rect 6290 11398 6342 11450
rect 9298 11398 9350 11450
rect 9362 11398 9414 11450
rect 9426 11398 9478 11450
rect 9490 11398 9542 11450
rect 5632 11339 5684 11348
rect 5632 11305 5641 11339
rect 5641 11305 5675 11339
rect 5675 11305 5684 11339
rect 5632 11296 5684 11305
rect 6736 11339 6788 11348
rect 5908 11203 5960 11212
rect 5908 11169 5917 11203
rect 5917 11169 5951 11203
rect 5951 11169 5960 11203
rect 5908 11160 5960 11169
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 6736 11305 6745 11339
rect 6745 11305 6779 11339
rect 6779 11305 6788 11339
rect 6736 11296 6788 11305
rect 7196 11271 7248 11280
rect 7196 11237 7205 11271
rect 7205 11237 7239 11271
rect 7239 11237 7248 11271
rect 7196 11228 7248 11237
rect 8760 11228 8812 11280
rect 5724 11067 5776 11076
rect 5724 11033 5733 11067
rect 5733 11033 5767 11067
rect 5767 11033 5776 11067
rect 5724 11024 5776 11033
rect 6920 11092 6972 11144
rect 9128 11160 9180 11212
rect 14188 11160 14240 11212
rect 5908 11024 5960 11076
rect 7104 11024 7156 11076
rect 9036 11024 9088 11076
rect 14188 11024 14240 11076
rect 8208 10956 8260 11008
rect 8852 10999 8904 11008
rect 8852 10965 8861 10999
rect 8861 10965 8895 10999
rect 8895 10965 8904 10999
rect 8852 10956 8904 10965
rect 1298 10854 1350 10906
rect 1362 10854 1414 10906
rect 1426 10854 1478 10906
rect 1490 10854 1542 10906
rect 4498 10854 4550 10906
rect 4562 10854 4614 10906
rect 4626 10854 4678 10906
rect 4690 10854 4742 10906
rect 7698 10854 7750 10906
rect 7762 10854 7814 10906
rect 7826 10854 7878 10906
rect 7890 10854 7942 10906
rect 6000 10795 6052 10804
rect 6000 10761 6009 10795
rect 6009 10761 6043 10795
rect 6043 10761 6052 10795
rect 6000 10752 6052 10761
rect 8208 10752 8260 10804
rect 14372 10684 14424 10736
rect 7104 10616 7156 10668
rect 5816 10591 5868 10600
rect 5816 10557 5825 10591
rect 5825 10557 5859 10591
rect 5859 10557 5868 10591
rect 5816 10548 5868 10557
rect 6644 10480 6696 10532
rect 7196 10480 7248 10532
rect 5356 10412 5408 10464
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 9128 10548 9180 10600
rect 8392 10480 8444 10532
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 9588 10412 9640 10464
rect 2898 10310 2950 10362
rect 2962 10310 3014 10362
rect 3026 10310 3078 10362
rect 3090 10310 3142 10362
rect 6098 10310 6150 10362
rect 6162 10310 6214 10362
rect 6226 10310 6278 10362
rect 6290 10310 6342 10362
rect 9298 10310 9350 10362
rect 9362 10310 9414 10362
rect 9426 10310 9478 10362
rect 9490 10310 9542 10362
rect 7196 10208 7248 10260
rect 5356 10115 5408 10124
rect 5356 10081 5365 10115
rect 5365 10081 5399 10115
rect 5399 10081 5408 10115
rect 5356 10072 5408 10081
rect 6736 10140 6788 10192
rect 6920 10183 6972 10192
rect 6920 10149 6929 10183
rect 6929 10149 6963 10183
rect 6963 10149 6972 10183
rect 6920 10140 6972 10149
rect 6000 10072 6052 10124
rect 8852 10140 8904 10192
rect 6644 10004 6696 10056
rect 7288 10004 7340 10056
rect 7564 10072 7616 10124
rect 8208 10004 8260 10056
rect 8944 10004 8996 10056
rect 6736 9936 6788 9988
rect 6460 9868 6512 9920
rect 6552 9868 6604 9920
rect 7472 9868 7524 9920
rect 1298 9766 1350 9818
rect 1362 9766 1414 9818
rect 1426 9766 1478 9818
rect 1490 9766 1542 9818
rect 4498 9766 4550 9818
rect 4562 9766 4614 9818
rect 4626 9766 4678 9818
rect 4690 9766 4742 9818
rect 7698 9766 7750 9818
rect 7762 9766 7814 9818
rect 7826 9766 7878 9818
rect 7890 9766 7942 9818
rect 4344 9664 4396 9716
rect 5356 9664 5408 9716
rect 5816 9664 5868 9716
rect 6552 9664 6604 9716
rect 8024 9664 8076 9716
rect 14280 9868 14332 9920
rect 8208 9528 8260 9580
rect 8944 9528 8996 9580
rect 14188 9528 14240 9580
rect 5080 9460 5132 9512
rect 5540 9460 5592 9512
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 5264 9324 5316 9376
rect 7012 9392 7064 9444
rect 6460 9324 6512 9376
rect 8300 9392 8352 9444
rect 14280 9392 14332 9444
rect 7564 9324 7616 9376
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 2898 9222 2950 9274
rect 2962 9222 3014 9274
rect 3026 9222 3078 9274
rect 3090 9222 3142 9274
rect 6098 9222 6150 9274
rect 6162 9222 6214 9274
rect 6226 9222 6278 9274
rect 6290 9222 6342 9274
rect 9298 9222 9350 9274
rect 9362 9222 9414 9274
rect 9426 9222 9478 9274
rect 9490 9222 9542 9274
rect 4804 9120 4856 9172
rect 5540 9120 5592 9172
rect 5908 9120 5960 9172
rect 6460 9052 6512 9104
rect 5172 8984 5224 9036
rect 6368 8984 6420 9036
rect 7656 9052 7708 9104
rect 8116 9052 8168 9104
rect 9588 9052 9640 9104
rect 7196 8984 7248 9036
rect 7748 9027 7800 9036
rect 7748 8993 7757 9027
rect 7757 8993 7791 9027
rect 7791 8993 7800 9027
rect 7748 8984 7800 8993
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 14188 9120 14240 9172
rect 5356 8823 5408 8832
rect 5356 8789 5365 8823
rect 5365 8789 5399 8823
rect 5399 8789 5408 8823
rect 5356 8780 5408 8789
rect 5908 8780 5960 8832
rect 8576 8780 8628 8832
rect 1298 8678 1350 8730
rect 1362 8678 1414 8730
rect 1426 8678 1478 8730
rect 1490 8678 1542 8730
rect 4498 8678 4550 8730
rect 4562 8678 4614 8730
rect 4626 8678 4678 8730
rect 4690 8678 4742 8730
rect 7698 8678 7750 8730
rect 7762 8678 7814 8730
rect 7826 8678 7878 8730
rect 7890 8678 7942 8730
rect 5356 8576 5408 8628
rect 8300 8619 8352 8628
rect 6460 8483 6512 8492
rect 4160 8372 4212 8424
rect 4344 8372 4396 8424
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 4988 8347 5040 8356
rect 4988 8313 4997 8347
rect 4997 8313 5031 8347
rect 5031 8313 5040 8347
rect 4988 8304 5040 8313
rect 5264 8304 5316 8356
rect 6460 8449 6469 8483
rect 6469 8449 6503 8483
rect 6503 8449 6512 8483
rect 6460 8440 6512 8449
rect 6920 8440 6972 8492
rect 8300 8585 8309 8619
rect 8309 8585 8343 8619
rect 8343 8585 8352 8619
rect 8300 8576 8352 8585
rect 8208 8508 8260 8560
rect 14188 8508 14240 8560
rect 6552 8415 6604 8424
rect 6552 8381 6561 8415
rect 6561 8381 6595 8415
rect 6595 8381 6604 8415
rect 6552 8372 6604 8381
rect 8576 8415 8628 8424
rect 6736 8304 6788 8356
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 14280 8304 14332 8356
rect 6920 8236 6972 8288
rect 2898 8134 2950 8186
rect 2962 8134 3014 8186
rect 3026 8134 3078 8186
rect 3090 8134 3142 8186
rect 6098 8134 6150 8186
rect 6162 8134 6214 8186
rect 6226 8134 6278 8186
rect 6290 8134 6342 8186
rect 9298 8134 9350 8186
rect 9362 8134 9414 8186
rect 9426 8134 9478 8186
rect 9490 8134 9542 8186
rect 8024 8032 8076 8084
rect 6460 7964 6512 8016
rect 7012 7964 7064 8016
rect 8760 8007 8812 8016
rect 8760 7973 8769 8007
rect 8769 7973 8803 8007
rect 8803 7973 8812 8007
rect 8760 7964 8812 7973
rect 3792 7896 3844 7948
rect 5540 7896 5592 7948
rect 5908 7828 5960 7880
rect 5080 7760 5132 7812
rect 5540 7760 5592 7812
rect 8024 7828 8076 7880
rect 8208 7828 8260 7880
rect 14004 7760 14056 7812
rect 4344 7692 4396 7744
rect 5172 7692 5224 7744
rect 7196 7692 7248 7744
rect 8116 7692 8168 7744
rect 1298 7590 1350 7642
rect 1362 7590 1414 7642
rect 1426 7590 1478 7642
rect 1490 7590 1542 7642
rect 4498 7590 4550 7642
rect 4562 7590 4614 7642
rect 4626 7590 4678 7642
rect 4690 7590 4742 7642
rect 7698 7590 7750 7642
rect 7762 7590 7814 7642
rect 7826 7590 7878 7642
rect 7890 7590 7942 7642
rect 7288 7488 7340 7540
rect 9128 7488 9180 7540
rect 6000 7352 6052 7404
rect 4160 7327 4212 7336
rect 4160 7293 4169 7327
rect 4169 7293 4203 7327
rect 4203 7293 4212 7327
rect 4160 7284 4212 7293
rect 4344 7284 4396 7336
rect 5172 7216 5224 7268
rect 8116 7284 8168 7336
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 6552 7216 6604 7268
rect 7380 7148 7432 7200
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 14188 7216 14240 7268
rect 8944 7148 8996 7200
rect 2898 7046 2950 7098
rect 2962 7046 3014 7098
rect 3026 7046 3078 7098
rect 3090 7046 3142 7098
rect 6098 7046 6150 7098
rect 6162 7046 6214 7098
rect 6226 7046 6278 7098
rect 6290 7046 6342 7098
rect 9298 7046 9350 7098
rect 9362 7046 9414 7098
rect 9426 7046 9478 7098
rect 9490 7046 9542 7098
rect 6552 6944 6604 6996
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 5908 6808 5960 6860
rect 6736 6876 6788 6928
rect 7472 6944 7524 6996
rect 8024 6944 8076 6996
rect 8392 6876 8444 6928
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 6000 6740 6052 6792
rect 4160 6672 4212 6724
rect 5816 6672 5868 6724
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 9036 6851 9088 6860
rect 9036 6817 9046 6851
rect 9046 6817 9080 6851
rect 9080 6817 9088 6851
rect 9036 6808 9088 6817
rect 7564 6740 7616 6792
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 5172 6604 5224 6656
rect 6000 6604 6052 6656
rect 6552 6604 6604 6656
rect 8760 6604 8812 6656
rect 1298 6502 1350 6554
rect 1362 6502 1414 6554
rect 1426 6502 1478 6554
rect 1490 6502 1542 6554
rect 4498 6502 4550 6554
rect 4562 6502 4614 6554
rect 4626 6502 4678 6554
rect 4690 6502 4742 6554
rect 7698 6502 7750 6554
rect 7762 6502 7814 6554
rect 7826 6502 7878 6554
rect 7890 6502 7942 6554
rect 3424 6400 3476 6452
rect 8944 6400 8996 6452
rect 14188 6400 14240 6452
rect 4068 6264 4120 6316
rect 5816 6264 5868 6316
rect 6000 6264 6052 6316
rect 6736 6264 6788 6316
rect 4160 6196 4212 6248
rect 4528 6239 4580 6248
rect 4528 6205 4537 6239
rect 4537 6205 4571 6239
rect 4571 6205 4580 6239
rect 4528 6196 4580 6205
rect 6368 6239 6420 6248
rect 6368 6205 6377 6239
rect 6377 6205 6411 6239
rect 6411 6205 6420 6239
rect 6368 6196 6420 6205
rect 14280 6264 14332 6316
rect 4804 6171 4856 6180
rect 4804 6137 4813 6171
rect 4813 6137 4847 6171
rect 4847 6137 4856 6171
rect 4804 6128 4856 6137
rect 4896 6128 4948 6180
rect 6920 6128 6972 6180
rect 8116 6128 8168 6180
rect 9128 6196 9180 6248
rect 9588 6196 9640 6248
rect 5540 6060 5592 6112
rect 8208 6060 8260 6112
rect 14372 6128 14424 6180
rect 9036 6060 9088 6112
rect 2898 5958 2950 6010
rect 2962 5958 3014 6010
rect 3026 5958 3078 6010
rect 3090 5958 3142 6010
rect 6098 5958 6150 6010
rect 6162 5958 6214 6010
rect 6226 5958 6278 6010
rect 6290 5958 6342 6010
rect 9298 5958 9350 6010
rect 9362 5958 9414 6010
rect 9426 5958 9478 6010
rect 9490 5958 9542 6010
rect 4896 5856 4948 5908
rect 3792 5763 3844 5772
rect 3792 5729 3801 5763
rect 3801 5729 3835 5763
rect 3835 5729 3844 5763
rect 3792 5720 3844 5729
rect 6552 5788 6604 5840
rect 5908 5720 5960 5772
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 8116 5856 8168 5908
rect 7380 5831 7432 5840
rect 7380 5797 7389 5831
rect 7389 5797 7423 5831
rect 7423 5797 7432 5831
rect 7380 5788 7432 5797
rect 9036 5788 9088 5840
rect 4344 5695 4396 5704
rect 4344 5661 4353 5695
rect 4353 5661 4387 5695
rect 4387 5661 4396 5695
rect 4344 5652 4396 5661
rect 6000 5652 6052 5704
rect 6460 5652 6512 5704
rect 4068 5584 4120 5636
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 14188 5652 14240 5704
rect 6736 5584 6788 5636
rect 4344 5516 4396 5568
rect 4804 5516 4856 5568
rect 6460 5559 6512 5568
rect 6460 5525 6469 5559
rect 6469 5525 6503 5559
rect 6503 5525 6512 5559
rect 6460 5516 6512 5525
rect 7012 5516 7064 5568
rect 7288 5516 7340 5568
rect 9128 5516 9180 5568
rect 1298 5414 1350 5466
rect 1362 5414 1414 5466
rect 1426 5414 1478 5466
rect 1490 5414 1542 5466
rect 4498 5414 4550 5466
rect 4562 5414 4614 5466
rect 4626 5414 4678 5466
rect 4690 5414 4742 5466
rect 7698 5414 7750 5466
rect 7762 5414 7814 5466
rect 7826 5414 7878 5466
rect 7890 5414 7942 5466
rect 4344 5312 4396 5364
rect 5724 5244 5776 5296
rect 4712 5176 4764 5228
rect 4252 5151 4304 5160
rect 4252 5117 4261 5151
rect 4261 5117 4295 5151
rect 4295 5117 4304 5151
rect 4252 5108 4304 5117
rect 6276 5108 6328 5160
rect 8300 5176 8352 5228
rect 8668 5108 8720 5160
rect 6460 5040 6512 5092
rect 7104 5083 7156 5092
rect 7104 5049 7113 5083
rect 7113 5049 7147 5083
rect 7147 5049 7156 5083
rect 7104 5040 7156 5049
rect 14188 5040 14240 5092
rect 4068 5015 4120 5024
rect 4068 4981 4077 5015
rect 4077 4981 4111 5015
rect 4111 4981 4120 5015
rect 4068 4972 4120 4981
rect 4344 4972 4396 5024
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 2898 4870 2950 4922
rect 2962 4870 3014 4922
rect 3026 4870 3078 4922
rect 3090 4870 3142 4922
rect 6098 4870 6150 4922
rect 6162 4870 6214 4922
rect 6226 4870 6278 4922
rect 6290 4870 6342 4922
rect 9298 4870 9350 4922
rect 9362 4870 9414 4922
rect 9426 4870 9478 4922
rect 9490 4870 9542 4922
rect 4160 4768 4212 4820
rect 6552 4700 6604 4752
rect 7288 4700 7340 4752
rect 4344 4675 4396 4684
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 6736 4564 6788 4616
rect 6920 4607 6972 4616
rect 6920 4573 6929 4607
rect 6929 4573 6963 4607
rect 6963 4573 6972 4607
rect 6920 4564 6972 4573
rect 7104 4564 7156 4616
rect 8852 4768 8904 4820
rect 9588 4768 9640 4820
rect 8760 4743 8812 4752
rect 8760 4709 8769 4743
rect 8769 4709 8803 4743
rect 8803 4709 8812 4743
rect 8760 4700 8812 4709
rect 9036 4607 9088 4616
rect 9036 4573 9045 4607
rect 9045 4573 9079 4607
rect 9079 4573 9088 4607
rect 9036 4564 9088 4573
rect 5724 4496 5776 4548
rect 6000 4428 6052 4480
rect 6276 4428 6328 4480
rect 4498 4326 4550 4378
rect 4562 4326 4614 4378
rect 4626 4326 4678 4378
rect 4690 4326 4742 4378
rect 7698 4326 7750 4378
rect 7762 4326 7814 4378
rect 7826 4326 7878 4378
rect 7890 4326 7942 4378
rect 7104 4224 7156 4276
rect 4344 4088 4396 4140
rect 5080 4088 5132 4140
rect 5816 4088 5868 4140
rect 8668 4131 8720 4140
rect 8668 4097 8677 4131
rect 8677 4097 8711 4131
rect 8711 4097 8720 4131
rect 8668 4088 8720 4097
rect 6184 4020 6236 4072
rect 6552 4020 6604 4072
rect 9128 4088 9180 4140
rect 6276 3952 6328 4004
rect 6460 3952 6512 4004
rect 8852 4063 8904 4072
rect 8852 4029 8862 4063
rect 8862 4029 8896 4063
rect 8896 4029 8904 4063
rect 8852 4020 8904 4029
rect 7012 3952 7064 4004
rect 14188 3952 14240 4004
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 5908 3884 5960 3936
rect 6552 3927 6604 3936
rect 6552 3893 6561 3927
rect 6561 3893 6595 3927
rect 6595 3893 6604 3927
rect 6552 3884 6604 3893
rect 6736 3884 6788 3936
rect 8760 3884 8812 3936
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 6098 3782 6150 3834
rect 6162 3782 6214 3834
rect 6226 3782 6278 3834
rect 6290 3782 6342 3834
rect 9298 3782 9350 3834
rect 9362 3782 9414 3834
rect 9426 3782 9478 3834
rect 9490 3782 9542 3834
rect 6000 3680 6052 3732
rect 5908 3612 5960 3664
rect 8484 3680 8536 3732
rect 6552 3612 6604 3664
rect 14280 3612 14332 3664
rect 4344 3587 4396 3596
rect 4344 3553 4353 3587
rect 4353 3553 4387 3587
rect 4387 3553 4396 3587
rect 4344 3544 4396 3553
rect 4988 3476 5040 3528
rect 6184 3519 6236 3528
rect 6184 3485 6193 3519
rect 6193 3485 6227 3519
rect 6227 3485 6236 3519
rect 6184 3476 6236 3485
rect 6460 3476 6512 3528
rect 8944 3587 8996 3596
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 8576 3476 8628 3528
rect 8852 3408 8904 3460
rect 9588 3408 9640 3460
rect 7012 3340 7064 3392
rect 4498 3238 4550 3290
rect 4562 3238 4614 3290
rect 4626 3238 4678 3290
rect 4690 3238 4742 3290
rect 7698 3238 7750 3290
rect 7762 3238 7814 3290
rect 7826 3238 7878 3290
rect 7890 3238 7942 3290
rect 4344 3136 4396 3188
rect 6920 3136 6972 3188
rect 8576 3179 8628 3188
rect 8576 3145 8585 3179
rect 8585 3145 8619 3179
rect 8619 3145 8628 3179
rect 8576 3136 8628 3145
rect 5816 3000 5868 3052
rect 6092 3000 6144 3052
rect 7104 3000 7156 3052
rect 9128 3043 9180 3052
rect 6000 2975 6052 2984
rect 6000 2941 6009 2975
rect 6009 2941 6043 2975
rect 6043 2941 6052 2975
rect 6000 2932 6052 2941
rect 6184 2932 6236 2984
rect 5080 2864 5132 2916
rect 5724 2864 5776 2916
rect 7012 2864 7064 2916
rect 6644 2796 6696 2848
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 8944 2932 8996 2984
rect 14188 2864 14240 2916
rect 6098 2694 6150 2746
rect 6162 2694 6214 2746
rect 6226 2694 6278 2746
rect 6290 2694 6342 2746
rect 9298 2694 9350 2746
rect 9362 2694 9414 2746
rect 9426 2694 9478 2746
rect 9490 2694 9542 2746
rect 4436 2635 4488 2644
rect 4436 2601 4445 2635
rect 4445 2601 4479 2635
rect 4479 2601 4488 2635
rect 4436 2592 4488 2601
rect 6552 2592 6604 2644
rect 6644 2592 6696 2644
rect 4896 2456 4948 2508
rect 5632 2499 5684 2508
rect 5632 2465 5641 2499
rect 5641 2465 5675 2499
rect 5675 2465 5684 2499
rect 5632 2456 5684 2465
rect 6000 2456 6052 2508
rect 6920 2524 6972 2576
rect 8760 2592 8812 2644
rect 9036 2524 9088 2576
rect 6736 2499 6788 2508
rect 6736 2465 6745 2499
rect 6745 2465 6779 2499
rect 6779 2465 6788 2499
rect 6736 2456 6788 2465
rect 6644 2363 6696 2372
rect 6644 2329 6653 2363
rect 6653 2329 6687 2363
rect 6687 2329 6696 2363
rect 6644 2320 6696 2329
rect 4988 2295 5040 2304
rect 4988 2261 4997 2295
rect 4997 2261 5031 2295
rect 5031 2261 5040 2295
rect 4988 2252 5040 2261
rect 5264 2295 5316 2304
rect 5264 2261 5273 2295
rect 5273 2261 5307 2295
rect 5307 2261 5316 2295
rect 5264 2252 5316 2261
rect 7012 2252 7064 2304
rect 14188 2320 14240 2372
rect 14372 2252 14424 2304
rect 4498 2150 4550 2202
rect 4562 2150 4614 2202
rect 4626 2150 4678 2202
rect 4690 2150 4742 2202
rect 7698 2150 7750 2202
rect 7762 2150 7814 2202
rect 7826 2150 7878 2202
rect 7890 2150 7942 2202
rect 5632 2048 5684 2100
rect 8668 2048 8720 2100
rect 4988 1980 5040 2032
rect 14096 1980 14148 2032
rect 4896 1844 4948 1896
rect 14280 1844 14332 1896
rect 5264 1776 5316 1828
rect 9588 1776 9640 1828
rect 6644 8 6696 60
rect 14188 8 14240 60
<< metal2 >>
rect 14278 13696 14334 13705
rect 14278 13631 14334 13640
rect 14186 13152 14242 13161
rect 14186 13087 14242 13096
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 6736 12572 6788 12578
rect 6736 12514 6788 12520
rect 5908 12504 5960 12510
rect 5908 12446 5960 12452
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 2872 11452 3168 11472
rect 2928 11450 2952 11452
rect 3008 11450 3032 11452
rect 3088 11450 3112 11452
rect 2950 11398 2952 11450
rect 3014 11398 3026 11450
rect 3088 11398 3090 11450
rect 2928 11396 2952 11398
rect 3008 11396 3032 11398
rect 3088 11396 3112 11398
rect 2872 11376 3168 11396
rect 5644 11354 5672 11494
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5920 11218 5948 12446
rect 6072 11452 6368 11472
rect 6128 11450 6152 11452
rect 6208 11450 6232 11452
rect 6288 11450 6312 11452
rect 6150 11398 6152 11450
rect 6214 11398 6226 11450
rect 6288 11398 6290 11450
rect 6128 11396 6152 11398
rect 6208 11396 6232 11398
rect 6288 11396 6312 11398
rect 6072 11376 6368 11396
rect 6748 11354 6776 12514
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 7208 11286 7236 12582
rect 14200 12510 14228 13087
rect 14292 12578 14320 13631
rect 14372 12640 14424 12646
rect 14370 12608 14372 12617
rect 14424 12608 14426 12617
rect 14280 12572 14332 12578
rect 14370 12543 14426 12552
rect 14280 12514 14332 12520
rect 14188 12504 14240 12510
rect 14188 12446 14240 12452
rect 14370 12200 14426 12209
rect 14370 12135 14426 12144
rect 14186 11656 14242 11665
rect 14186 11591 14242 11600
rect 9272 11452 9568 11472
rect 9328 11450 9352 11452
rect 9408 11450 9432 11452
rect 9488 11450 9512 11452
rect 9350 11398 9352 11450
rect 9414 11398 9426 11450
rect 9488 11398 9490 11450
rect 9328 11396 9352 11398
rect 9408 11396 9432 11398
rect 9488 11396 9512 11398
rect 9272 11376 9568 11396
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5908 11076 5960 11082
rect 5908 11018 5960 11024
rect 1272 10908 1568 10928
rect 1328 10906 1352 10908
rect 1408 10906 1432 10908
rect 1488 10906 1512 10908
rect 1350 10854 1352 10906
rect 1414 10854 1426 10906
rect 1488 10854 1490 10906
rect 1328 10852 1352 10854
rect 1408 10852 1432 10854
rect 1488 10852 1512 10854
rect 1272 10832 1568 10852
rect 4472 10908 4768 10928
rect 4528 10906 4552 10908
rect 4608 10906 4632 10908
rect 4688 10906 4712 10908
rect 4550 10854 4552 10906
rect 4614 10854 4626 10906
rect 4688 10854 4690 10906
rect 4528 10852 4552 10854
rect 4608 10852 4632 10854
rect 4688 10852 4712 10854
rect 4472 10832 4768 10852
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 2872 10364 3168 10384
rect 2928 10362 2952 10364
rect 3008 10362 3032 10364
rect 3088 10362 3112 10364
rect 2950 10310 2952 10362
rect 3014 10310 3026 10362
rect 3088 10310 3090 10362
rect 2928 10308 2952 10310
rect 3008 10308 3032 10310
rect 3088 10308 3112 10310
rect 2872 10288 3168 10308
rect 5368 10130 5396 10406
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 1272 9820 1568 9840
rect 1328 9818 1352 9820
rect 1408 9818 1432 9820
rect 1488 9818 1512 9820
rect 1350 9766 1352 9818
rect 1414 9766 1426 9818
rect 1488 9766 1490 9818
rect 1328 9764 1352 9766
rect 1408 9764 1432 9766
rect 1488 9764 1512 9766
rect 1272 9744 1568 9764
rect 4472 9820 4768 9840
rect 4528 9818 4552 9820
rect 4608 9818 4632 9820
rect 4688 9818 4712 9820
rect 4550 9766 4552 9818
rect 4614 9766 4626 9818
rect 4688 9766 4690 9818
rect 4528 9764 4552 9766
rect 4608 9764 4632 9766
rect 4688 9764 4712 9766
rect 4472 9744 4768 9764
rect 5368 9722 5396 10066
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 2872 9276 3168 9296
rect 2928 9274 2952 9276
rect 3008 9274 3032 9276
rect 3088 9274 3112 9276
rect 2950 9222 2952 9274
rect 3014 9222 3026 9274
rect 3088 9222 3090 9274
rect 2928 9220 2952 9222
rect 3008 9220 3032 9222
rect 3088 9220 3112 9222
rect 2872 9200 3168 9220
rect 1272 8732 1568 8752
rect 1328 8730 1352 8732
rect 1408 8730 1432 8732
rect 1488 8730 1512 8732
rect 1350 8678 1352 8730
rect 1414 8678 1426 8730
rect 1488 8678 1490 8730
rect 1328 8676 1352 8678
rect 1408 8676 1432 8678
rect 1488 8676 1512 8678
rect 1272 8656 1568 8676
rect 4356 8430 4384 9658
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5540 9512 5592 9518
rect 5736 9489 5764 11018
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5828 9722 5856 10542
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5540 9454 5592 9460
rect 5722 9480 5778 9489
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4472 8732 4768 8752
rect 4528 8730 4552 8732
rect 4608 8730 4632 8732
rect 4688 8730 4712 8732
rect 4550 8678 4552 8730
rect 4614 8678 4626 8730
rect 4688 8678 4690 8730
rect 4528 8676 4552 8678
rect 4608 8676 4632 8678
rect 4688 8676 4712 8678
rect 4472 8656 4768 8676
rect 4816 8514 4844 9114
rect 4724 8486 4844 8514
rect 4724 8430 4752 8486
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 2872 8188 3168 8208
rect 2928 8186 2952 8188
rect 3008 8186 3032 8188
rect 3088 8186 3112 8188
rect 2950 8134 2952 8186
rect 3014 8134 3026 8186
rect 3088 8134 3090 8186
rect 2928 8132 2952 8134
rect 3008 8132 3032 8134
rect 3088 8132 3112 8134
rect 2872 8112 3168 8132
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 1272 7644 1568 7664
rect 1328 7642 1352 7644
rect 1408 7642 1432 7644
rect 1488 7642 1512 7644
rect 1350 7590 1352 7642
rect 1414 7590 1426 7642
rect 1488 7590 1490 7642
rect 1328 7588 1352 7590
rect 1408 7588 1432 7590
rect 1488 7588 1512 7590
rect 1272 7568 1568 7588
rect 2872 7100 3168 7120
rect 2928 7098 2952 7100
rect 3008 7098 3032 7100
rect 3088 7098 3112 7100
rect 2950 7046 2952 7098
rect 3014 7046 3026 7098
rect 3088 7046 3090 7098
rect 2928 7044 2952 7046
rect 3008 7044 3032 7046
rect 3088 7044 3112 7046
rect 2872 7024 3168 7044
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 1272 6556 1568 6576
rect 1328 6554 1352 6556
rect 1408 6554 1432 6556
rect 1488 6554 1512 6556
rect 1350 6502 1352 6554
rect 1414 6502 1426 6554
rect 1488 6502 1490 6554
rect 1328 6500 1352 6502
rect 1408 6500 1432 6502
rect 1488 6500 1512 6502
rect 1272 6480 1568 6500
rect 3436 6458 3464 6598
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 2872 6012 3168 6032
rect 2928 6010 2952 6012
rect 3008 6010 3032 6012
rect 3088 6010 3112 6012
rect 2950 5958 2952 6010
rect 3014 5958 3026 6010
rect 3088 5958 3090 6010
rect 2928 5956 2952 5958
rect 3008 5956 3032 5958
rect 3088 5956 3112 5958
rect 2872 5936 3168 5956
rect 3804 5778 3832 7890
rect 4172 7342 4200 8366
rect 4988 8356 5040 8362
rect 4988 8298 5040 8304
rect 4344 7744 4396 7750
rect 4264 7692 4344 7698
rect 4264 7686 4396 7692
rect 4264 7670 4384 7686
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4080 6322 4108 6802
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4172 6254 4200 6666
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 1272 5468 1568 5488
rect 1328 5466 1352 5468
rect 1408 5466 1432 5468
rect 1488 5466 1512 5468
rect 1350 5414 1352 5466
rect 1414 5414 1426 5466
rect 1488 5414 1490 5466
rect 1328 5412 1352 5414
rect 1408 5412 1432 5414
rect 1488 5412 1512 5414
rect 1272 5392 1568 5412
rect 4080 5030 4108 5578
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 2872 4924 3168 4944
rect 2928 4922 2952 4924
rect 3008 4922 3032 4924
rect 3088 4922 3112 4924
rect 2950 4870 2952 4922
rect 3014 4870 3026 4922
rect 3088 4870 3090 4922
rect 2928 4868 2952 4870
rect 3008 4868 3032 4870
rect 3088 4868 3112 4870
rect 2872 4848 3168 4868
rect 4172 4826 4200 6190
rect 4264 5166 4292 7670
rect 4472 7644 4768 7664
rect 4528 7642 4552 7644
rect 4608 7642 4632 7644
rect 4688 7642 4712 7644
rect 4550 7590 4552 7642
rect 4614 7590 4626 7642
rect 4688 7590 4690 7642
rect 4528 7588 4552 7590
rect 4608 7588 4632 7590
rect 4688 7588 4712 7590
rect 4472 7568 4768 7588
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4356 6798 4384 7278
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4356 5710 4384 6734
rect 4472 6556 4768 6576
rect 4528 6554 4552 6556
rect 4608 6554 4632 6556
rect 4688 6554 4712 6556
rect 4550 6502 4552 6554
rect 4614 6502 4626 6554
rect 4688 6502 4690 6554
rect 4528 6500 4552 6502
rect 4608 6500 4632 6502
rect 4688 6500 4712 6502
rect 4472 6480 4768 6500
rect 4528 6248 4580 6254
rect 4526 6216 4528 6225
rect 4580 6216 4582 6225
rect 4526 6151 4582 6160
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 4896 6180 4948 6186
rect 4896 6122 4948 6128
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4816 5574 4844 6122
rect 4908 5914 4936 6122
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4356 5370 4384 5510
rect 4472 5468 4768 5488
rect 4528 5466 4552 5468
rect 4608 5466 4632 5468
rect 4688 5466 4712 5468
rect 4550 5414 4552 5466
rect 4614 5414 4626 5466
rect 4688 5414 4690 5466
rect 4528 5412 4552 5414
rect 4608 5412 4632 5414
rect 4688 5412 4712 5414
rect 4472 5392 4768 5412
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4816 5250 4844 5510
rect 4724 5234 4844 5250
rect 4712 5228 4844 5234
rect 4764 5222 4844 5228
rect 4712 5170 4764 5176
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4356 4690 4384 4966
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4356 4146 4384 4626
rect 4472 4380 4768 4400
rect 4528 4378 4552 4380
rect 4608 4378 4632 4380
rect 4688 4378 4712 4380
rect 4550 4326 4552 4378
rect 4614 4326 4626 4378
rect 4688 4326 4690 4378
rect 4528 4324 4552 4326
rect 4608 4324 4632 4326
rect 4688 4324 4712 4326
rect 4472 4304 4768 4324
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4356 3602 4384 4082
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4356 3194 4384 3538
rect 5000 3534 5028 8298
rect 5092 7818 5120 9454
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 5092 4146 5120 7754
rect 5184 7750 5212 8978
rect 5276 8362 5304 9318
rect 5552 9178 5580 9454
rect 5722 9415 5778 9424
rect 5920 9178 5948 11018
rect 6012 10810 6040 11154
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6012 10130 6040 10746
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6072 10364 6368 10384
rect 6128 10362 6152 10364
rect 6208 10362 6232 10364
rect 6288 10362 6312 10364
rect 6150 10310 6152 10362
rect 6214 10310 6226 10362
rect 6288 10310 6290 10362
rect 6128 10308 6152 10310
rect 6208 10308 6232 10310
rect 6288 10308 6312 10310
rect 6072 10288 6368 10308
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6656 10062 6684 10474
rect 6932 10198 6960 11086
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7116 10674 7144 11018
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 7672 10908 7968 10928
rect 7728 10906 7752 10908
rect 7808 10906 7832 10908
rect 7888 10906 7912 10908
rect 7750 10854 7752 10906
rect 7814 10854 7826 10906
rect 7888 10854 7890 10906
rect 7728 10852 7752 10854
rect 7808 10852 7832 10854
rect 7888 10852 7912 10854
rect 7672 10832 7968 10852
rect 8220 10810 8248 10950
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 7208 10266 7236 10474
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 6736 10192 6788 10198
rect 6920 10192 6972 10198
rect 6788 10140 6868 10146
rect 6736 10134 6868 10140
rect 6920 10134 6972 10140
rect 6748 10118 6868 10134
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6472 9382 6500 9862
rect 6564 9722 6592 9862
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6072 9276 6368 9296
rect 6128 9274 6152 9276
rect 6208 9274 6232 9276
rect 6288 9274 6312 9276
rect 6150 9222 6152 9274
rect 6214 9222 6226 9274
rect 6288 9222 6290 9274
rect 6128 9220 6152 9222
rect 6208 9220 6232 9222
rect 6288 9220 6312 9222
rect 6072 9200 6368 9220
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8634 5396 8774
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5552 7954 5580 9114
rect 6460 9104 6512 9110
rect 6458 9072 6460 9081
rect 6512 9072 6514 9081
rect 6368 9036 6420 9042
rect 6458 9007 6514 9016
rect 6368 8978 6420 8984
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6380 8922 6408 8978
rect 6564 8922 6592 9658
rect 6656 9518 6684 9998
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 5908 8832 5960 8838
rect 6012 8809 6040 8910
rect 6380 8894 6592 8922
rect 6642 8936 6698 8945
rect 6642 8871 6698 8880
rect 5908 8774 5960 8780
rect 5998 8800 6054 8809
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5920 7886 5948 8774
rect 5998 8735 6054 8744
rect 6550 8528 6606 8537
rect 6460 8492 6512 8498
rect 6550 8463 6606 8472
rect 6460 8434 6512 8440
rect 6072 8188 6368 8208
rect 6128 8186 6152 8188
rect 6208 8186 6232 8188
rect 6288 8186 6312 8188
rect 6150 8134 6152 8186
rect 6214 8134 6226 8186
rect 6288 8134 6290 8186
rect 6128 8132 6152 8134
rect 6208 8132 6232 8134
rect 6288 8132 6312 8134
rect 6072 8112 6368 8132
rect 6472 8022 6500 8434
rect 6564 8430 6592 8463
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 5184 6662 5212 7210
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5552 6118 5580 7754
rect 5920 6866 5948 7822
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 6012 6798 6040 7346
rect 6564 7274 6592 8366
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 6072 7100 6368 7120
rect 6128 7098 6152 7100
rect 6208 7098 6232 7100
rect 6288 7098 6312 7100
rect 6150 7046 6152 7098
rect 6214 7046 6226 7098
rect 6288 7046 6290 7098
rect 6128 7044 6152 7046
rect 6208 7044 6232 7046
rect 6288 7044 6312 7046
rect 6072 7024 6368 7044
rect 6564 7002 6592 7210
rect 6552 6996 6604 7002
rect 6472 6956 6552 6984
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5828 6322 5856 6666
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 6012 6322 6040 6598
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5828 5794 5856 6258
rect 5828 5778 5948 5794
rect 5828 5772 5960 5778
rect 5828 5766 5908 5772
rect 5908 5714 5960 5720
rect 6012 5710 6040 6258
rect 6368 6248 6420 6254
rect 6366 6216 6368 6225
rect 6472 6236 6500 6956
rect 6552 6938 6604 6944
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6420 6216 6500 6236
rect 6422 6208 6500 6216
rect 6366 6151 6422 6160
rect 6072 6012 6368 6032
rect 6128 6010 6152 6012
rect 6208 6010 6232 6012
rect 6288 6010 6312 6012
rect 6150 5958 6152 6010
rect 6214 5958 6226 6010
rect 6288 5958 6290 6010
rect 6128 5956 6152 5958
rect 6208 5956 6232 5958
rect 6288 5956 6312 5958
rect 6072 5936 6368 5956
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5736 4554 5764 5238
rect 6288 5166 6316 5714
rect 6472 5710 6500 6208
rect 6564 5846 6592 6598
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 6472 5098 6500 5510
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6072 4924 6368 4944
rect 6128 4922 6152 4924
rect 6208 4922 6232 4924
rect 6288 4922 6312 4924
rect 6150 4870 6152 4922
rect 6214 4870 6226 4922
rect 6288 4870 6290 4922
rect 6128 4868 6152 4870
rect 6208 4868 6232 4870
rect 6288 4868 6312 4870
rect 6072 4848 6368 4868
rect 6564 4758 6592 4966
rect 6552 4752 6604 4758
rect 6552 4694 6604 4700
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4472 3292 4768 3312
rect 4528 3290 4552 3292
rect 4608 3290 4632 3292
rect 4688 3290 4712 3292
rect 4550 3238 4552 3290
rect 4614 3238 4626 3290
rect 4688 3238 4690 3290
rect 4528 3236 4552 3238
rect 4608 3236 4632 3238
rect 4688 3236 4712 3238
rect 4472 3216 4768 3236
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4434 2952 4490 2961
rect 5092 2922 5120 4082
rect 5736 2922 5764 4490
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5828 3942 5856 4082
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5828 3058 5856 3878
rect 5920 3670 5948 3878
rect 6012 3738 6040 4422
rect 6196 4078 6224 4626
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6288 4010 6316 4422
rect 6656 4162 6684 8871
rect 6748 8362 6776 9930
rect 6840 8945 6868 10118
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7194 9480 7250 9489
rect 7012 9444 7064 9450
rect 7194 9415 7250 9424
rect 7012 9386 7064 9392
rect 6826 8936 6882 8945
rect 6826 8871 6882 8880
rect 6840 8498 6960 8514
rect 6840 8492 6972 8498
rect 6840 8486 6920 8492
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6840 8242 6868 8486
rect 6920 8434 6972 8440
rect 6748 8214 6868 8242
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6748 6934 6776 8214
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6748 6322 6776 6870
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6932 6186 6960 8230
rect 7024 8022 7052 9386
rect 7208 9042 7236 9415
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7300 8537 7328 9998
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 8974 7512 9862
rect 7576 9674 7604 10066
rect 8220 10062 8248 10406
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 7672 9820 7968 9840
rect 7728 9818 7752 9820
rect 7808 9818 7832 9820
rect 7888 9818 7912 9820
rect 7750 9766 7752 9818
rect 7814 9766 7826 9818
rect 7888 9766 7890 9818
rect 7728 9764 7752 9766
rect 7808 9764 7832 9766
rect 7888 9764 7912 9766
rect 7672 9744 7968 9764
rect 8024 9716 8076 9722
rect 7576 9646 7788 9674
rect 8024 9658 8076 9664
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7654 9344 7710 9353
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7484 8809 7512 8910
rect 7470 8800 7526 8809
rect 7470 8735 7526 8744
rect 7286 8528 7342 8537
rect 7286 8463 7342 8472
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6748 4622 6776 5578
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6564 4134 6684 4162
rect 6564 4078 6592 4134
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6072 3836 6368 3856
rect 6128 3834 6152 3836
rect 6208 3834 6232 3836
rect 6288 3834 6312 3836
rect 6150 3782 6152 3834
rect 6214 3782 6226 3834
rect 6288 3782 6290 3834
rect 6128 3780 6152 3782
rect 6208 3780 6232 3782
rect 6288 3780 6312 3782
rect 6072 3760 6368 3780
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 6472 3534 6500 3946
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6564 3670 6592 3878
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6184 3528 6236 3534
rect 6104 3488 6184 3516
rect 6104 3058 6132 3488
rect 6184 3470 6236 3476
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6656 3210 6684 4134
rect 6748 3942 6776 4558
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6196 3182 6684 3210
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6196 2990 6224 3182
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 4434 2887 4490 2896
rect 5080 2916 5132 2922
rect 4448 2650 4476 2887
rect 5080 2858 5132 2864
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 6012 2514 6040 2926
rect 6644 2848 6696 2854
rect 6550 2816 6606 2825
rect 6072 2748 6368 2768
rect 6644 2790 6696 2796
rect 6550 2751 6606 2760
rect 6128 2746 6152 2748
rect 6208 2746 6232 2748
rect 6288 2746 6312 2748
rect 6150 2694 6152 2746
rect 6214 2694 6226 2746
rect 6288 2694 6290 2746
rect 6128 2692 6152 2694
rect 6208 2692 6232 2694
rect 6288 2692 6312 2694
rect 6072 2672 6368 2692
rect 6564 2650 6592 2751
rect 6656 2650 6684 2790
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6748 2514 6776 3878
rect 6932 3194 6960 4558
rect 7024 4010 7052 5510
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7116 4622 7144 5034
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7208 4434 7236 7686
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7300 7426 7328 7482
rect 7576 7426 7604 9318
rect 7654 9279 7710 9288
rect 7668 9110 7696 9279
rect 7760 9217 7788 9646
rect 8036 9330 8064 9658
rect 8220 9586 8248 9998
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 7852 9302 8064 9330
rect 7746 9208 7802 9217
rect 7746 9143 7802 9152
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7760 9042 7788 9143
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7852 8922 7880 9302
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 7852 8894 8064 8922
rect 7672 8732 7968 8752
rect 7728 8730 7752 8732
rect 7808 8730 7832 8732
rect 7888 8730 7912 8732
rect 7750 8678 7752 8730
rect 7814 8678 7826 8730
rect 7888 8678 7890 8730
rect 7728 8676 7752 8678
rect 7808 8676 7832 8678
rect 7888 8676 7912 8678
rect 7672 8656 7968 8676
rect 8036 8090 8064 8894
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7672 7644 7968 7664
rect 7728 7642 7752 7644
rect 7808 7642 7832 7644
rect 7888 7642 7912 7644
rect 7750 7590 7752 7642
rect 7814 7590 7826 7642
rect 7888 7590 7890 7642
rect 7728 7588 7752 7590
rect 7808 7588 7832 7590
rect 7888 7588 7912 7590
rect 7672 7568 7968 7588
rect 7300 7398 7604 7426
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7392 5846 7420 7142
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 4758 7328 5510
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7116 4406 7236 4434
rect 7116 4282 7144 4406
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 7484 3505 7512 6938
rect 7576 6798 7604 7398
rect 8036 7002 8064 7822
rect 8128 7750 8156 9046
rect 8206 8936 8262 8945
rect 8206 8871 8262 8880
rect 8220 8566 8248 8871
rect 8312 8634 8340 9386
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7672 6556 7968 6576
rect 7728 6554 7752 6556
rect 7808 6554 7832 6556
rect 7888 6554 7912 6556
rect 7750 6502 7752 6554
rect 7814 6502 7826 6554
rect 7888 6502 7890 6554
rect 7728 6500 7752 6502
rect 7808 6500 7832 6502
rect 7888 6500 7912 6502
rect 7672 6480 7968 6500
rect 8128 6186 8156 7278
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 8128 5914 8156 6122
rect 8220 6118 8248 7822
rect 8404 7290 8432 10474
rect 8482 9072 8538 9081
rect 8482 9007 8538 9016
rect 8312 7262 8432 7290
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8024 5704 8076 5710
rect 8312 5658 8340 7262
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8404 6934 8432 7142
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8076 5652 8340 5658
rect 8024 5646 8340 5652
rect 8036 5630 8340 5646
rect 7672 5468 7968 5488
rect 7728 5466 7752 5468
rect 7808 5466 7832 5468
rect 7888 5466 7912 5468
rect 7750 5414 7752 5466
rect 7814 5414 7826 5466
rect 7888 5414 7890 5466
rect 7728 5412 7752 5414
rect 7808 5412 7832 5414
rect 7888 5412 7912 5414
rect 7672 5392 7968 5412
rect 8312 5234 8340 5630
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 7672 4380 7968 4400
rect 7728 4378 7752 4380
rect 7808 4378 7832 4380
rect 7888 4378 7912 4380
rect 7750 4326 7752 4378
rect 7814 4326 7826 4378
rect 7888 4326 7890 4378
rect 7728 4324 7752 4326
rect 7808 4324 7832 4326
rect 7888 4324 7912 4326
rect 7672 4304 7968 4324
rect 8496 3738 8524 9007
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8430 8616 8774
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8772 8022 8800 11222
rect 14200 11218 14228 11591
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8864 10198 8892 10950
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8956 10062 8984 10542
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8956 9586 8984 9998
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 9048 9518 9076 11018
rect 9140 10606 9168 11154
rect 14292 11121 14320 11494
rect 14278 11112 14334 11121
rect 14188 11076 14240 11082
rect 14278 11047 14334 11056
rect 14188 11018 14240 11024
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9272 10364 9568 10384
rect 9328 10362 9352 10364
rect 9408 10362 9432 10364
rect 9488 10362 9512 10364
rect 9350 10310 9352 10362
rect 9414 10310 9426 10362
rect 9488 10310 9490 10362
rect 9328 10308 9352 10310
rect 9408 10308 9432 10310
rect 9488 10308 9512 10310
rect 9272 10288 9568 10308
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9126 9344 9182 9353
rect 9048 9217 9076 9318
rect 9126 9279 9182 9288
rect 9034 9208 9090 9217
rect 9034 9143 9090 9152
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 9140 7546 9168 9279
rect 9272 9276 9568 9296
rect 9328 9274 9352 9276
rect 9408 9274 9432 9276
rect 9488 9274 9512 9276
rect 9350 9222 9352 9274
rect 9414 9222 9426 9274
rect 9488 9222 9490 9274
rect 9328 9220 9352 9222
rect 9408 9220 9432 9222
rect 9488 9220 9512 9222
rect 9272 9200 9568 9220
rect 9600 9110 9628 10406
rect 14200 10169 14228 11018
rect 14384 10742 14412 12135
rect 14372 10736 14424 10742
rect 14278 10704 14334 10713
rect 14372 10678 14424 10684
rect 14278 10639 14334 10648
rect 14186 10160 14242 10169
rect 14186 10095 14242 10104
rect 14292 9926 14320 10639
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14186 9616 14242 9625
rect 14186 9551 14188 9560
rect 14240 9551 14242 9560
rect 14188 9522 14240 9528
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14186 9208 14242 9217
rect 14186 9143 14188 9152
rect 14240 9143 14242 9152
rect 14188 9114 14240 9120
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 14292 8673 14320 9386
rect 14278 8664 14334 8673
rect 14278 8599 14334 8608
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 9272 8188 9568 8208
rect 9328 8186 9352 8188
rect 9408 8186 9432 8188
rect 9488 8186 9512 8188
rect 9350 8134 9352 8186
rect 9414 8134 9426 8186
rect 9488 8134 9490 8186
rect 9328 8132 9352 8134
rect 9408 8132 9432 8134
rect 9488 8132 9512 8134
rect 9272 8112 9568 8132
rect 14200 8129 14228 8502
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14186 8120 14242 8129
rect 14186 8055 14242 8064
rect 14004 7812 14056 7818
rect 14004 7754 14056 7760
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8956 6866 8984 7142
rect 9048 6866 9076 7278
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8680 4146 8708 5102
rect 8772 4758 8800 6598
rect 8956 6458 8984 6802
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9140 6338 9168 7278
rect 9272 7100 9568 7120
rect 9328 7098 9352 7100
rect 9408 7098 9432 7100
rect 9488 7098 9512 7100
rect 9350 7046 9352 7098
rect 9414 7046 9426 7098
rect 9488 7046 9490 7098
rect 9328 7044 9352 7046
rect 9408 7044 9432 7046
rect 9488 7044 9512 7046
rect 9272 7024 9568 7044
rect 8956 6310 9168 6338
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8760 4752 8812 4758
rect 8760 4694 8812 4700
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8576 3528 8628 3534
rect 7470 3496 7526 3505
rect 8576 3470 8628 3476
rect 7470 3431 7526 3440
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7024 3074 7052 3334
rect 7672 3292 7968 3312
rect 7728 3290 7752 3292
rect 7808 3290 7832 3292
rect 7888 3290 7912 3292
rect 7750 3238 7752 3290
rect 7814 3238 7826 3290
rect 7888 3238 7890 3290
rect 7728 3236 7752 3238
rect 7808 3236 7832 3238
rect 7888 3236 7912 3238
rect 7672 3216 7968 3236
rect 8588 3194 8616 3470
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 6932 3046 7052 3074
rect 7104 3052 7156 3058
rect 6932 2582 6960 3046
rect 7104 2994 7156 3000
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 4472 2204 4768 2224
rect 4528 2202 4552 2204
rect 4608 2202 4632 2204
rect 4688 2202 4712 2204
rect 4550 2150 4552 2202
rect 4614 2150 4626 2202
rect 4688 2150 4690 2202
rect 4528 2148 4552 2150
rect 4608 2148 4632 2150
rect 4688 2148 4712 2150
rect 4472 2128 4768 2148
rect 4908 1902 4936 2450
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 5000 2038 5028 2246
rect 4988 2032 5040 2038
rect 4988 1974 5040 1980
rect 4896 1896 4948 1902
rect 4896 1838 4948 1844
rect 5276 1834 5304 2246
rect 5644 2106 5672 2450
rect 6644 2372 6696 2378
rect 6644 2314 6696 2320
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 5264 1828 5316 1834
rect 5264 1770 5316 1776
rect 6656 66 6684 2314
rect 7024 2310 7052 2858
rect 7116 2825 7144 2994
rect 7102 2816 7158 2825
rect 7102 2751 7158 2760
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7672 2204 7968 2224
rect 7728 2202 7752 2204
rect 7808 2202 7832 2204
rect 7888 2202 7912 2204
rect 7750 2150 7752 2202
rect 7814 2150 7826 2202
rect 7888 2150 7890 2202
rect 7728 2148 7752 2150
rect 7808 2148 7832 2150
rect 7888 2148 7912 2150
rect 7672 2128 7968 2148
rect 8680 2106 8708 4082
rect 8864 4078 8892 4762
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8772 2650 8800 3878
rect 8956 3754 8984 6310
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 14016 6202 14044 7754
rect 14292 7721 14320 8298
rect 14278 7712 14334 7721
rect 14278 7647 14334 7656
rect 14188 7268 14240 7274
rect 14188 7210 14240 7216
rect 14200 7177 14228 7210
rect 14186 7168 14242 7177
rect 14186 7103 14242 7112
rect 14186 6624 14242 6633
rect 14186 6559 14242 6568
rect 14200 6458 14228 6559
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14186 6216 14242 6225
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 9048 5846 9076 6054
rect 9036 5840 9088 5846
rect 9036 5782 9088 5788
rect 9140 5574 9168 6190
rect 9272 6012 9568 6032
rect 9328 6010 9352 6012
rect 9408 6010 9432 6012
rect 9488 6010 9512 6012
rect 9350 5958 9352 6010
rect 9414 5958 9426 6010
rect 9488 5958 9490 6010
rect 9328 5956 9352 5958
rect 9408 5956 9432 5958
rect 9488 5956 9512 5958
rect 9272 5936 9568 5956
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8864 3726 8984 3754
rect 8864 3466 8892 3726
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8956 2990 8984 3538
rect 8944 2984 8996 2990
rect 8942 2952 8944 2961
rect 8996 2952 8998 2961
rect 8942 2887 8998 2896
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 9048 2582 9076 4558
rect 9140 4146 9168 5510
rect 9272 4924 9568 4944
rect 9328 4922 9352 4924
rect 9408 4922 9432 4924
rect 9488 4922 9512 4924
rect 9350 4870 9352 4922
rect 9414 4870 9426 4922
rect 9488 4870 9490 4922
rect 9328 4868 9352 4870
rect 9408 4868 9432 4870
rect 9488 4868 9512 4870
rect 9272 4848 9568 4868
rect 9600 4826 9628 6190
rect 14016 6174 14186 6202
rect 14186 6151 14242 6160
rect 14188 5704 14240 5710
rect 14186 5672 14188 5681
rect 14240 5672 14242 5681
rect 14186 5607 14242 5616
rect 14292 5137 14320 6258
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14278 5128 14334 5137
rect 14188 5092 14240 5098
rect 14278 5063 14334 5072
rect 14188 5034 14240 5040
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 14200 4185 14228 5034
rect 14384 4729 14412 6122
rect 14370 4720 14426 4729
rect 14370 4655 14426 4664
rect 14186 4176 14242 4185
rect 9128 4140 9180 4146
rect 14186 4111 14242 4120
rect 9128 4082 9180 4088
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 3058 9168 3878
rect 9272 3836 9568 3856
rect 9328 3834 9352 3836
rect 9408 3834 9432 3836
rect 9488 3834 9512 3836
rect 9350 3782 9352 3834
rect 9414 3782 9426 3834
rect 9488 3782 9490 3834
rect 9328 3780 9352 3782
rect 9408 3780 9432 3782
rect 9488 3780 9512 3782
rect 9272 3760 9568 3780
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9272 2748 9568 2768
rect 9328 2746 9352 2748
rect 9408 2746 9432 2748
rect 9488 2746 9512 2748
rect 9350 2694 9352 2746
rect 9414 2694 9426 2746
rect 9488 2694 9490 2746
rect 9328 2692 9352 2694
rect 9408 2692 9432 2694
rect 9488 2692 9512 2694
rect 9272 2672 9568 2692
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 9600 1834 9628 3402
rect 14200 3233 14228 3946
rect 14280 3664 14332 3670
rect 14278 3632 14280 3641
rect 14332 3632 14334 3641
rect 14278 3567 14334 3576
rect 14186 3224 14242 3233
rect 14186 3159 14242 3168
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 14200 2689 14228 2858
rect 14186 2680 14242 2689
rect 14186 2615 14242 2624
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 14096 2032 14148 2038
rect 14096 1974 14148 1980
rect 9588 1828 9640 1834
rect 9588 1770 9640 1776
rect 14108 1737 14136 1974
rect 14094 1728 14150 1737
rect 14094 1663 14150 1672
rect 14200 1193 14228 2314
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 14278 2136 14334 2145
rect 14278 2071 14334 2080
rect 14292 1902 14320 2071
rect 14280 1896 14332 1902
rect 14280 1838 14332 1844
rect 14186 1184 14242 1193
rect 14186 1119 14242 1128
rect 14384 649 14412 2246
rect 14370 640 14426 649
rect 14370 575 14426 584
rect 14186 232 14242 241
rect 14186 167 14242 176
rect 14200 66 14228 167
rect 6644 60 6696 66
rect 6644 2 6696 8
rect 14188 60 14240 66
rect 14188 2 14240 8
<< via2 >>
rect 14278 13640 14334 13696
rect 14186 13096 14242 13152
rect 2872 11450 2928 11452
rect 2952 11450 3008 11452
rect 3032 11450 3088 11452
rect 3112 11450 3168 11452
rect 2872 11398 2898 11450
rect 2898 11398 2928 11450
rect 2952 11398 2962 11450
rect 2962 11398 3008 11450
rect 3032 11398 3078 11450
rect 3078 11398 3088 11450
rect 3112 11398 3142 11450
rect 3142 11398 3168 11450
rect 2872 11396 2928 11398
rect 2952 11396 3008 11398
rect 3032 11396 3088 11398
rect 3112 11396 3168 11398
rect 6072 11450 6128 11452
rect 6152 11450 6208 11452
rect 6232 11450 6288 11452
rect 6312 11450 6368 11452
rect 6072 11398 6098 11450
rect 6098 11398 6128 11450
rect 6152 11398 6162 11450
rect 6162 11398 6208 11450
rect 6232 11398 6278 11450
rect 6278 11398 6288 11450
rect 6312 11398 6342 11450
rect 6342 11398 6368 11450
rect 6072 11396 6128 11398
rect 6152 11396 6208 11398
rect 6232 11396 6288 11398
rect 6312 11396 6368 11398
rect 14370 12588 14372 12608
rect 14372 12588 14424 12608
rect 14424 12588 14426 12608
rect 14370 12552 14426 12588
rect 14370 12144 14426 12200
rect 14186 11600 14242 11656
rect 9272 11450 9328 11452
rect 9352 11450 9408 11452
rect 9432 11450 9488 11452
rect 9512 11450 9568 11452
rect 9272 11398 9298 11450
rect 9298 11398 9328 11450
rect 9352 11398 9362 11450
rect 9362 11398 9408 11450
rect 9432 11398 9478 11450
rect 9478 11398 9488 11450
rect 9512 11398 9542 11450
rect 9542 11398 9568 11450
rect 9272 11396 9328 11398
rect 9352 11396 9408 11398
rect 9432 11396 9488 11398
rect 9512 11396 9568 11398
rect 1272 10906 1328 10908
rect 1352 10906 1408 10908
rect 1432 10906 1488 10908
rect 1512 10906 1568 10908
rect 1272 10854 1298 10906
rect 1298 10854 1328 10906
rect 1352 10854 1362 10906
rect 1362 10854 1408 10906
rect 1432 10854 1478 10906
rect 1478 10854 1488 10906
rect 1512 10854 1542 10906
rect 1542 10854 1568 10906
rect 1272 10852 1328 10854
rect 1352 10852 1408 10854
rect 1432 10852 1488 10854
rect 1512 10852 1568 10854
rect 4472 10906 4528 10908
rect 4552 10906 4608 10908
rect 4632 10906 4688 10908
rect 4712 10906 4768 10908
rect 4472 10854 4498 10906
rect 4498 10854 4528 10906
rect 4552 10854 4562 10906
rect 4562 10854 4608 10906
rect 4632 10854 4678 10906
rect 4678 10854 4688 10906
rect 4712 10854 4742 10906
rect 4742 10854 4768 10906
rect 4472 10852 4528 10854
rect 4552 10852 4608 10854
rect 4632 10852 4688 10854
rect 4712 10852 4768 10854
rect 2872 10362 2928 10364
rect 2952 10362 3008 10364
rect 3032 10362 3088 10364
rect 3112 10362 3168 10364
rect 2872 10310 2898 10362
rect 2898 10310 2928 10362
rect 2952 10310 2962 10362
rect 2962 10310 3008 10362
rect 3032 10310 3078 10362
rect 3078 10310 3088 10362
rect 3112 10310 3142 10362
rect 3142 10310 3168 10362
rect 2872 10308 2928 10310
rect 2952 10308 3008 10310
rect 3032 10308 3088 10310
rect 3112 10308 3168 10310
rect 1272 9818 1328 9820
rect 1352 9818 1408 9820
rect 1432 9818 1488 9820
rect 1512 9818 1568 9820
rect 1272 9766 1298 9818
rect 1298 9766 1328 9818
rect 1352 9766 1362 9818
rect 1362 9766 1408 9818
rect 1432 9766 1478 9818
rect 1478 9766 1488 9818
rect 1512 9766 1542 9818
rect 1542 9766 1568 9818
rect 1272 9764 1328 9766
rect 1352 9764 1408 9766
rect 1432 9764 1488 9766
rect 1512 9764 1568 9766
rect 4472 9818 4528 9820
rect 4552 9818 4608 9820
rect 4632 9818 4688 9820
rect 4712 9818 4768 9820
rect 4472 9766 4498 9818
rect 4498 9766 4528 9818
rect 4552 9766 4562 9818
rect 4562 9766 4608 9818
rect 4632 9766 4678 9818
rect 4678 9766 4688 9818
rect 4712 9766 4742 9818
rect 4742 9766 4768 9818
rect 4472 9764 4528 9766
rect 4552 9764 4608 9766
rect 4632 9764 4688 9766
rect 4712 9764 4768 9766
rect 2872 9274 2928 9276
rect 2952 9274 3008 9276
rect 3032 9274 3088 9276
rect 3112 9274 3168 9276
rect 2872 9222 2898 9274
rect 2898 9222 2928 9274
rect 2952 9222 2962 9274
rect 2962 9222 3008 9274
rect 3032 9222 3078 9274
rect 3078 9222 3088 9274
rect 3112 9222 3142 9274
rect 3142 9222 3168 9274
rect 2872 9220 2928 9222
rect 2952 9220 3008 9222
rect 3032 9220 3088 9222
rect 3112 9220 3168 9222
rect 1272 8730 1328 8732
rect 1352 8730 1408 8732
rect 1432 8730 1488 8732
rect 1512 8730 1568 8732
rect 1272 8678 1298 8730
rect 1298 8678 1328 8730
rect 1352 8678 1362 8730
rect 1362 8678 1408 8730
rect 1432 8678 1478 8730
rect 1478 8678 1488 8730
rect 1512 8678 1542 8730
rect 1542 8678 1568 8730
rect 1272 8676 1328 8678
rect 1352 8676 1408 8678
rect 1432 8676 1488 8678
rect 1512 8676 1568 8678
rect 4472 8730 4528 8732
rect 4552 8730 4608 8732
rect 4632 8730 4688 8732
rect 4712 8730 4768 8732
rect 4472 8678 4498 8730
rect 4498 8678 4528 8730
rect 4552 8678 4562 8730
rect 4562 8678 4608 8730
rect 4632 8678 4678 8730
rect 4678 8678 4688 8730
rect 4712 8678 4742 8730
rect 4742 8678 4768 8730
rect 4472 8676 4528 8678
rect 4552 8676 4608 8678
rect 4632 8676 4688 8678
rect 4712 8676 4768 8678
rect 2872 8186 2928 8188
rect 2952 8186 3008 8188
rect 3032 8186 3088 8188
rect 3112 8186 3168 8188
rect 2872 8134 2898 8186
rect 2898 8134 2928 8186
rect 2952 8134 2962 8186
rect 2962 8134 3008 8186
rect 3032 8134 3078 8186
rect 3078 8134 3088 8186
rect 3112 8134 3142 8186
rect 3142 8134 3168 8186
rect 2872 8132 2928 8134
rect 2952 8132 3008 8134
rect 3032 8132 3088 8134
rect 3112 8132 3168 8134
rect 1272 7642 1328 7644
rect 1352 7642 1408 7644
rect 1432 7642 1488 7644
rect 1512 7642 1568 7644
rect 1272 7590 1298 7642
rect 1298 7590 1328 7642
rect 1352 7590 1362 7642
rect 1362 7590 1408 7642
rect 1432 7590 1478 7642
rect 1478 7590 1488 7642
rect 1512 7590 1542 7642
rect 1542 7590 1568 7642
rect 1272 7588 1328 7590
rect 1352 7588 1408 7590
rect 1432 7588 1488 7590
rect 1512 7588 1568 7590
rect 2872 7098 2928 7100
rect 2952 7098 3008 7100
rect 3032 7098 3088 7100
rect 3112 7098 3168 7100
rect 2872 7046 2898 7098
rect 2898 7046 2928 7098
rect 2952 7046 2962 7098
rect 2962 7046 3008 7098
rect 3032 7046 3078 7098
rect 3078 7046 3088 7098
rect 3112 7046 3142 7098
rect 3142 7046 3168 7098
rect 2872 7044 2928 7046
rect 2952 7044 3008 7046
rect 3032 7044 3088 7046
rect 3112 7044 3168 7046
rect 1272 6554 1328 6556
rect 1352 6554 1408 6556
rect 1432 6554 1488 6556
rect 1512 6554 1568 6556
rect 1272 6502 1298 6554
rect 1298 6502 1328 6554
rect 1352 6502 1362 6554
rect 1362 6502 1408 6554
rect 1432 6502 1478 6554
rect 1478 6502 1488 6554
rect 1512 6502 1542 6554
rect 1542 6502 1568 6554
rect 1272 6500 1328 6502
rect 1352 6500 1408 6502
rect 1432 6500 1488 6502
rect 1512 6500 1568 6502
rect 2872 6010 2928 6012
rect 2952 6010 3008 6012
rect 3032 6010 3088 6012
rect 3112 6010 3168 6012
rect 2872 5958 2898 6010
rect 2898 5958 2928 6010
rect 2952 5958 2962 6010
rect 2962 5958 3008 6010
rect 3032 5958 3078 6010
rect 3078 5958 3088 6010
rect 3112 5958 3142 6010
rect 3142 5958 3168 6010
rect 2872 5956 2928 5958
rect 2952 5956 3008 5958
rect 3032 5956 3088 5958
rect 3112 5956 3168 5958
rect 1272 5466 1328 5468
rect 1352 5466 1408 5468
rect 1432 5466 1488 5468
rect 1512 5466 1568 5468
rect 1272 5414 1298 5466
rect 1298 5414 1328 5466
rect 1352 5414 1362 5466
rect 1362 5414 1408 5466
rect 1432 5414 1478 5466
rect 1478 5414 1488 5466
rect 1512 5414 1542 5466
rect 1542 5414 1568 5466
rect 1272 5412 1328 5414
rect 1352 5412 1408 5414
rect 1432 5412 1488 5414
rect 1512 5412 1568 5414
rect 2872 4922 2928 4924
rect 2952 4922 3008 4924
rect 3032 4922 3088 4924
rect 3112 4922 3168 4924
rect 2872 4870 2898 4922
rect 2898 4870 2928 4922
rect 2952 4870 2962 4922
rect 2962 4870 3008 4922
rect 3032 4870 3078 4922
rect 3078 4870 3088 4922
rect 3112 4870 3142 4922
rect 3142 4870 3168 4922
rect 2872 4868 2928 4870
rect 2952 4868 3008 4870
rect 3032 4868 3088 4870
rect 3112 4868 3168 4870
rect 4472 7642 4528 7644
rect 4552 7642 4608 7644
rect 4632 7642 4688 7644
rect 4712 7642 4768 7644
rect 4472 7590 4498 7642
rect 4498 7590 4528 7642
rect 4552 7590 4562 7642
rect 4562 7590 4608 7642
rect 4632 7590 4678 7642
rect 4678 7590 4688 7642
rect 4712 7590 4742 7642
rect 4742 7590 4768 7642
rect 4472 7588 4528 7590
rect 4552 7588 4608 7590
rect 4632 7588 4688 7590
rect 4712 7588 4768 7590
rect 4472 6554 4528 6556
rect 4552 6554 4608 6556
rect 4632 6554 4688 6556
rect 4712 6554 4768 6556
rect 4472 6502 4498 6554
rect 4498 6502 4528 6554
rect 4552 6502 4562 6554
rect 4562 6502 4608 6554
rect 4632 6502 4678 6554
rect 4678 6502 4688 6554
rect 4712 6502 4742 6554
rect 4742 6502 4768 6554
rect 4472 6500 4528 6502
rect 4552 6500 4608 6502
rect 4632 6500 4688 6502
rect 4712 6500 4768 6502
rect 4526 6196 4528 6216
rect 4528 6196 4580 6216
rect 4580 6196 4582 6216
rect 4526 6160 4582 6196
rect 4472 5466 4528 5468
rect 4552 5466 4608 5468
rect 4632 5466 4688 5468
rect 4712 5466 4768 5468
rect 4472 5414 4498 5466
rect 4498 5414 4528 5466
rect 4552 5414 4562 5466
rect 4562 5414 4608 5466
rect 4632 5414 4678 5466
rect 4678 5414 4688 5466
rect 4712 5414 4742 5466
rect 4742 5414 4768 5466
rect 4472 5412 4528 5414
rect 4552 5412 4608 5414
rect 4632 5412 4688 5414
rect 4712 5412 4768 5414
rect 4472 4378 4528 4380
rect 4552 4378 4608 4380
rect 4632 4378 4688 4380
rect 4712 4378 4768 4380
rect 4472 4326 4498 4378
rect 4498 4326 4528 4378
rect 4552 4326 4562 4378
rect 4562 4326 4608 4378
rect 4632 4326 4678 4378
rect 4678 4326 4688 4378
rect 4712 4326 4742 4378
rect 4742 4326 4768 4378
rect 4472 4324 4528 4326
rect 4552 4324 4608 4326
rect 4632 4324 4688 4326
rect 4712 4324 4768 4326
rect 5722 9424 5778 9480
rect 6072 10362 6128 10364
rect 6152 10362 6208 10364
rect 6232 10362 6288 10364
rect 6312 10362 6368 10364
rect 6072 10310 6098 10362
rect 6098 10310 6128 10362
rect 6152 10310 6162 10362
rect 6162 10310 6208 10362
rect 6232 10310 6278 10362
rect 6278 10310 6288 10362
rect 6312 10310 6342 10362
rect 6342 10310 6368 10362
rect 6072 10308 6128 10310
rect 6152 10308 6208 10310
rect 6232 10308 6288 10310
rect 6312 10308 6368 10310
rect 7672 10906 7728 10908
rect 7752 10906 7808 10908
rect 7832 10906 7888 10908
rect 7912 10906 7968 10908
rect 7672 10854 7698 10906
rect 7698 10854 7728 10906
rect 7752 10854 7762 10906
rect 7762 10854 7808 10906
rect 7832 10854 7878 10906
rect 7878 10854 7888 10906
rect 7912 10854 7942 10906
rect 7942 10854 7968 10906
rect 7672 10852 7728 10854
rect 7752 10852 7808 10854
rect 7832 10852 7888 10854
rect 7912 10852 7968 10854
rect 6072 9274 6128 9276
rect 6152 9274 6208 9276
rect 6232 9274 6288 9276
rect 6312 9274 6368 9276
rect 6072 9222 6098 9274
rect 6098 9222 6128 9274
rect 6152 9222 6162 9274
rect 6162 9222 6208 9274
rect 6232 9222 6278 9274
rect 6278 9222 6288 9274
rect 6312 9222 6342 9274
rect 6342 9222 6368 9274
rect 6072 9220 6128 9222
rect 6152 9220 6208 9222
rect 6232 9220 6288 9222
rect 6312 9220 6368 9222
rect 6458 9052 6460 9072
rect 6460 9052 6512 9072
rect 6512 9052 6514 9072
rect 6458 9016 6514 9052
rect 6642 8880 6698 8936
rect 5998 8744 6054 8800
rect 6550 8472 6606 8528
rect 6072 8186 6128 8188
rect 6152 8186 6208 8188
rect 6232 8186 6288 8188
rect 6312 8186 6368 8188
rect 6072 8134 6098 8186
rect 6098 8134 6128 8186
rect 6152 8134 6162 8186
rect 6162 8134 6208 8186
rect 6232 8134 6278 8186
rect 6278 8134 6288 8186
rect 6312 8134 6342 8186
rect 6342 8134 6368 8186
rect 6072 8132 6128 8134
rect 6152 8132 6208 8134
rect 6232 8132 6288 8134
rect 6312 8132 6368 8134
rect 6072 7098 6128 7100
rect 6152 7098 6208 7100
rect 6232 7098 6288 7100
rect 6312 7098 6368 7100
rect 6072 7046 6098 7098
rect 6098 7046 6128 7098
rect 6152 7046 6162 7098
rect 6162 7046 6208 7098
rect 6232 7046 6278 7098
rect 6278 7046 6288 7098
rect 6312 7046 6342 7098
rect 6342 7046 6368 7098
rect 6072 7044 6128 7046
rect 6152 7044 6208 7046
rect 6232 7044 6288 7046
rect 6312 7044 6368 7046
rect 6366 6196 6368 6216
rect 6368 6196 6420 6216
rect 6420 6196 6422 6216
rect 6366 6160 6422 6196
rect 6072 6010 6128 6012
rect 6152 6010 6208 6012
rect 6232 6010 6288 6012
rect 6312 6010 6368 6012
rect 6072 5958 6098 6010
rect 6098 5958 6128 6010
rect 6152 5958 6162 6010
rect 6162 5958 6208 6010
rect 6232 5958 6278 6010
rect 6278 5958 6288 6010
rect 6312 5958 6342 6010
rect 6342 5958 6368 6010
rect 6072 5956 6128 5958
rect 6152 5956 6208 5958
rect 6232 5956 6288 5958
rect 6312 5956 6368 5958
rect 6072 4922 6128 4924
rect 6152 4922 6208 4924
rect 6232 4922 6288 4924
rect 6312 4922 6368 4924
rect 6072 4870 6098 4922
rect 6098 4870 6128 4922
rect 6152 4870 6162 4922
rect 6162 4870 6208 4922
rect 6232 4870 6278 4922
rect 6278 4870 6288 4922
rect 6312 4870 6342 4922
rect 6342 4870 6368 4922
rect 6072 4868 6128 4870
rect 6152 4868 6208 4870
rect 6232 4868 6288 4870
rect 6312 4868 6368 4870
rect 4472 3290 4528 3292
rect 4552 3290 4608 3292
rect 4632 3290 4688 3292
rect 4712 3290 4768 3292
rect 4472 3238 4498 3290
rect 4498 3238 4528 3290
rect 4552 3238 4562 3290
rect 4562 3238 4608 3290
rect 4632 3238 4678 3290
rect 4678 3238 4688 3290
rect 4712 3238 4742 3290
rect 4742 3238 4768 3290
rect 4472 3236 4528 3238
rect 4552 3236 4608 3238
rect 4632 3236 4688 3238
rect 4712 3236 4768 3238
rect 4434 2896 4490 2952
rect 7194 9424 7250 9480
rect 6826 8880 6882 8936
rect 7672 9818 7728 9820
rect 7752 9818 7808 9820
rect 7832 9818 7888 9820
rect 7912 9818 7968 9820
rect 7672 9766 7698 9818
rect 7698 9766 7728 9818
rect 7752 9766 7762 9818
rect 7762 9766 7808 9818
rect 7832 9766 7878 9818
rect 7878 9766 7888 9818
rect 7912 9766 7942 9818
rect 7942 9766 7968 9818
rect 7672 9764 7728 9766
rect 7752 9764 7808 9766
rect 7832 9764 7888 9766
rect 7912 9764 7968 9766
rect 7470 8744 7526 8800
rect 7286 8472 7342 8528
rect 6072 3834 6128 3836
rect 6152 3834 6208 3836
rect 6232 3834 6288 3836
rect 6312 3834 6368 3836
rect 6072 3782 6098 3834
rect 6098 3782 6128 3834
rect 6152 3782 6162 3834
rect 6162 3782 6208 3834
rect 6232 3782 6278 3834
rect 6278 3782 6288 3834
rect 6312 3782 6342 3834
rect 6342 3782 6368 3834
rect 6072 3780 6128 3782
rect 6152 3780 6208 3782
rect 6232 3780 6288 3782
rect 6312 3780 6368 3782
rect 6550 2760 6606 2816
rect 6072 2746 6128 2748
rect 6152 2746 6208 2748
rect 6232 2746 6288 2748
rect 6312 2746 6368 2748
rect 6072 2694 6098 2746
rect 6098 2694 6128 2746
rect 6152 2694 6162 2746
rect 6162 2694 6208 2746
rect 6232 2694 6278 2746
rect 6278 2694 6288 2746
rect 6312 2694 6342 2746
rect 6342 2694 6368 2746
rect 6072 2692 6128 2694
rect 6152 2692 6208 2694
rect 6232 2692 6288 2694
rect 6312 2692 6368 2694
rect 7654 9288 7710 9344
rect 7746 9152 7802 9208
rect 7672 8730 7728 8732
rect 7752 8730 7808 8732
rect 7832 8730 7888 8732
rect 7912 8730 7968 8732
rect 7672 8678 7698 8730
rect 7698 8678 7728 8730
rect 7752 8678 7762 8730
rect 7762 8678 7808 8730
rect 7832 8678 7878 8730
rect 7878 8678 7888 8730
rect 7912 8678 7942 8730
rect 7942 8678 7968 8730
rect 7672 8676 7728 8678
rect 7752 8676 7808 8678
rect 7832 8676 7888 8678
rect 7912 8676 7968 8678
rect 7672 7642 7728 7644
rect 7752 7642 7808 7644
rect 7832 7642 7888 7644
rect 7912 7642 7968 7644
rect 7672 7590 7698 7642
rect 7698 7590 7728 7642
rect 7752 7590 7762 7642
rect 7762 7590 7808 7642
rect 7832 7590 7878 7642
rect 7878 7590 7888 7642
rect 7912 7590 7942 7642
rect 7942 7590 7968 7642
rect 7672 7588 7728 7590
rect 7752 7588 7808 7590
rect 7832 7588 7888 7590
rect 7912 7588 7968 7590
rect 8206 8880 8262 8936
rect 7672 6554 7728 6556
rect 7752 6554 7808 6556
rect 7832 6554 7888 6556
rect 7912 6554 7968 6556
rect 7672 6502 7698 6554
rect 7698 6502 7728 6554
rect 7752 6502 7762 6554
rect 7762 6502 7808 6554
rect 7832 6502 7878 6554
rect 7878 6502 7888 6554
rect 7912 6502 7942 6554
rect 7942 6502 7968 6554
rect 7672 6500 7728 6502
rect 7752 6500 7808 6502
rect 7832 6500 7888 6502
rect 7912 6500 7968 6502
rect 8482 9016 8538 9072
rect 7672 5466 7728 5468
rect 7752 5466 7808 5468
rect 7832 5466 7888 5468
rect 7912 5466 7968 5468
rect 7672 5414 7698 5466
rect 7698 5414 7728 5466
rect 7752 5414 7762 5466
rect 7762 5414 7808 5466
rect 7832 5414 7878 5466
rect 7878 5414 7888 5466
rect 7912 5414 7942 5466
rect 7942 5414 7968 5466
rect 7672 5412 7728 5414
rect 7752 5412 7808 5414
rect 7832 5412 7888 5414
rect 7912 5412 7968 5414
rect 7672 4378 7728 4380
rect 7752 4378 7808 4380
rect 7832 4378 7888 4380
rect 7912 4378 7968 4380
rect 7672 4326 7698 4378
rect 7698 4326 7728 4378
rect 7752 4326 7762 4378
rect 7762 4326 7808 4378
rect 7832 4326 7878 4378
rect 7878 4326 7888 4378
rect 7912 4326 7942 4378
rect 7942 4326 7968 4378
rect 7672 4324 7728 4326
rect 7752 4324 7808 4326
rect 7832 4324 7888 4326
rect 7912 4324 7968 4326
rect 14278 11056 14334 11112
rect 9272 10362 9328 10364
rect 9352 10362 9408 10364
rect 9432 10362 9488 10364
rect 9512 10362 9568 10364
rect 9272 10310 9298 10362
rect 9298 10310 9328 10362
rect 9352 10310 9362 10362
rect 9362 10310 9408 10362
rect 9432 10310 9478 10362
rect 9478 10310 9488 10362
rect 9512 10310 9542 10362
rect 9542 10310 9568 10362
rect 9272 10308 9328 10310
rect 9352 10308 9408 10310
rect 9432 10308 9488 10310
rect 9512 10308 9568 10310
rect 9126 9288 9182 9344
rect 9034 9152 9090 9208
rect 9272 9274 9328 9276
rect 9352 9274 9408 9276
rect 9432 9274 9488 9276
rect 9512 9274 9568 9276
rect 9272 9222 9298 9274
rect 9298 9222 9328 9274
rect 9352 9222 9362 9274
rect 9362 9222 9408 9274
rect 9432 9222 9478 9274
rect 9478 9222 9488 9274
rect 9512 9222 9542 9274
rect 9542 9222 9568 9274
rect 9272 9220 9328 9222
rect 9352 9220 9408 9222
rect 9432 9220 9488 9222
rect 9512 9220 9568 9222
rect 14278 10648 14334 10704
rect 14186 10104 14242 10160
rect 14186 9580 14242 9616
rect 14186 9560 14188 9580
rect 14188 9560 14240 9580
rect 14240 9560 14242 9580
rect 14186 9172 14242 9208
rect 14186 9152 14188 9172
rect 14188 9152 14240 9172
rect 14240 9152 14242 9172
rect 14278 8608 14334 8664
rect 9272 8186 9328 8188
rect 9352 8186 9408 8188
rect 9432 8186 9488 8188
rect 9512 8186 9568 8188
rect 9272 8134 9298 8186
rect 9298 8134 9328 8186
rect 9352 8134 9362 8186
rect 9362 8134 9408 8186
rect 9432 8134 9478 8186
rect 9478 8134 9488 8186
rect 9512 8134 9542 8186
rect 9542 8134 9568 8186
rect 9272 8132 9328 8134
rect 9352 8132 9408 8134
rect 9432 8132 9488 8134
rect 9512 8132 9568 8134
rect 14186 8064 14242 8120
rect 9272 7098 9328 7100
rect 9352 7098 9408 7100
rect 9432 7098 9488 7100
rect 9512 7098 9568 7100
rect 9272 7046 9298 7098
rect 9298 7046 9328 7098
rect 9352 7046 9362 7098
rect 9362 7046 9408 7098
rect 9432 7046 9478 7098
rect 9478 7046 9488 7098
rect 9512 7046 9542 7098
rect 9542 7046 9568 7098
rect 9272 7044 9328 7046
rect 9352 7044 9408 7046
rect 9432 7044 9488 7046
rect 9512 7044 9568 7046
rect 7470 3440 7526 3496
rect 7672 3290 7728 3292
rect 7752 3290 7808 3292
rect 7832 3290 7888 3292
rect 7912 3290 7968 3292
rect 7672 3238 7698 3290
rect 7698 3238 7728 3290
rect 7752 3238 7762 3290
rect 7762 3238 7808 3290
rect 7832 3238 7878 3290
rect 7878 3238 7888 3290
rect 7912 3238 7942 3290
rect 7942 3238 7968 3290
rect 7672 3236 7728 3238
rect 7752 3236 7808 3238
rect 7832 3236 7888 3238
rect 7912 3236 7968 3238
rect 4472 2202 4528 2204
rect 4552 2202 4608 2204
rect 4632 2202 4688 2204
rect 4712 2202 4768 2204
rect 4472 2150 4498 2202
rect 4498 2150 4528 2202
rect 4552 2150 4562 2202
rect 4562 2150 4608 2202
rect 4632 2150 4678 2202
rect 4678 2150 4688 2202
rect 4712 2150 4742 2202
rect 4742 2150 4768 2202
rect 4472 2148 4528 2150
rect 4552 2148 4608 2150
rect 4632 2148 4688 2150
rect 4712 2148 4768 2150
rect 7102 2760 7158 2816
rect 7672 2202 7728 2204
rect 7752 2202 7808 2204
rect 7832 2202 7888 2204
rect 7912 2202 7968 2204
rect 7672 2150 7698 2202
rect 7698 2150 7728 2202
rect 7752 2150 7762 2202
rect 7762 2150 7808 2202
rect 7832 2150 7878 2202
rect 7878 2150 7888 2202
rect 7912 2150 7942 2202
rect 7942 2150 7968 2202
rect 7672 2148 7728 2150
rect 7752 2148 7808 2150
rect 7832 2148 7888 2150
rect 7912 2148 7968 2150
rect 14278 7656 14334 7712
rect 14186 7112 14242 7168
rect 14186 6568 14242 6624
rect 9272 6010 9328 6012
rect 9352 6010 9408 6012
rect 9432 6010 9488 6012
rect 9512 6010 9568 6012
rect 9272 5958 9298 6010
rect 9298 5958 9328 6010
rect 9352 5958 9362 6010
rect 9362 5958 9408 6010
rect 9432 5958 9478 6010
rect 9478 5958 9488 6010
rect 9512 5958 9542 6010
rect 9542 5958 9568 6010
rect 9272 5956 9328 5958
rect 9352 5956 9408 5958
rect 9432 5956 9488 5958
rect 9512 5956 9568 5958
rect 8942 2932 8944 2952
rect 8944 2932 8996 2952
rect 8996 2932 8998 2952
rect 8942 2896 8998 2932
rect 9272 4922 9328 4924
rect 9352 4922 9408 4924
rect 9432 4922 9488 4924
rect 9512 4922 9568 4924
rect 9272 4870 9298 4922
rect 9298 4870 9328 4922
rect 9352 4870 9362 4922
rect 9362 4870 9408 4922
rect 9432 4870 9478 4922
rect 9478 4870 9488 4922
rect 9512 4870 9542 4922
rect 9542 4870 9568 4922
rect 9272 4868 9328 4870
rect 9352 4868 9408 4870
rect 9432 4868 9488 4870
rect 9512 4868 9568 4870
rect 14186 6160 14242 6216
rect 14186 5652 14188 5672
rect 14188 5652 14240 5672
rect 14240 5652 14242 5672
rect 14186 5616 14242 5652
rect 14278 5072 14334 5128
rect 14370 4664 14426 4720
rect 14186 4120 14242 4176
rect 9272 3834 9328 3836
rect 9352 3834 9408 3836
rect 9432 3834 9488 3836
rect 9512 3834 9568 3836
rect 9272 3782 9298 3834
rect 9298 3782 9328 3834
rect 9352 3782 9362 3834
rect 9362 3782 9408 3834
rect 9432 3782 9478 3834
rect 9478 3782 9488 3834
rect 9512 3782 9542 3834
rect 9542 3782 9568 3834
rect 9272 3780 9328 3782
rect 9352 3780 9408 3782
rect 9432 3780 9488 3782
rect 9512 3780 9568 3782
rect 9272 2746 9328 2748
rect 9352 2746 9408 2748
rect 9432 2746 9488 2748
rect 9512 2746 9568 2748
rect 9272 2694 9298 2746
rect 9298 2694 9328 2746
rect 9352 2694 9362 2746
rect 9362 2694 9408 2746
rect 9432 2694 9478 2746
rect 9478 2694 9488 2746
rect 9512 2694 9542 2746
rect 9542 2694 9568 2746
rect 9272 2692 9328 2694
rect 9352 2692 9408 2694
rect 9432 2692 9488 2694
rect 9512 2692 9568 2694
rect 14278 3612 14280 3632
rect 14280 3612 14332 3632
rect 14332 3612 14334 3632
rect 14278 3576 14334 3612
rect 14186 3168 14242 3224
rect 14186 2624 14242 2680
rect 14094 1672 14150 1728
rect 14278 2080 14334 2136
rect 14186 1128 14242 1184
rect 14370 584 14426 640
rect 14186 176 14242 232
<< metal3 >>
rect 14000 13696 34000 13728
rect 14000 13640 14278 13696
rect 14334 13640 34000 13696
rect 14000 13608 34000 13640
rect 14000 13152 34000 13184
rect 14000 13096 14186 13152
rect 14242 13096 34000 13152
rect 14000 13064 34000 13096
rect 14000 12608 34000 12640
rect 14000 12552 14370 12608
rect 14426 12552 34000 12608
rect 14000 12520 34000 12552
rect 14000 12200 34000 12232
rect 14000 12144 14370 12200
rect 14426 12144 34000 12200
rect 14000 12112 34000 12144
rect 14000 11656 34000 11688
rect 14000 11600 14186 11656
rect 14242 11600 34000 11656
rect 14000 11568 34000 11600
rect 2860 11456 3180 11457
rect 2860 11392 2868 11456
rect 2932 11392 2948 11456
rect 3012 11392 3028 11456
rect 3092 11392 3108 11456
rect 3172 11392 3180 11456
rect 2860 11391 3180 11392
rect 6060 11456 6380 11457
rect 6060 11392 6068 11456
rect 6132 11392 6148 11456
rect 6212 11392 6228 11456
rect 6292 11392 6308 11456
rect 6372 11392 6380 11456
rect 6060 11391 6380 11392
rect 9260 11456 9580 11457
rect 9260 11392 9268 11456
rect 9332 11392 9348 11456
rect 9412 11392 9428 11456
rect 9492 11392 9508 11456
rect 9572 11392 9580 11456
rect 9260 11391 9580 11392
rect 14000 11112 34000 11144
rect 14000 11056 14278 11112
rect 14334 11056 34000 11112
rect 14000 11024 34000 11056
rect 1260 10912 1580 10913
rect 1260 10848 1268 10912
rect 1332 10848 1348 10912
rect 1412 10848 1428 10912
rect 1492 10848 1508 10912
rect 1572 10848 1580 10912
rect 1260 10847 1580 10848
rect 4460 10912 4780 10913
rect 4460 10848 4468 10912
rect 4532 10848 4548 10912
rect 4612 10848 4628 10912
rect 4692 10848 4708 10912
rect 4772 10848 4780 10912
rect 4460 10847 4780 10848
rect 7660 10912 7980 10913
rect 7660 10848 7668 10912
rect 7732 10848 7748 10912
rect 7812 10848 7828 10912
rect 7892 10848 7908 10912
rect 7972 10848 7980 10912
rect 7660 10847 7980 10848
rect 14000 10704 34000 10736
rect 14000 10648 14278 10704
rect 14334 10648 34000 10704
rect 14000 10616 34000 10648
rect 2860 10368 3180 10369
rect 2860 10304 2868 10368
rect 2932 10304 2948 10368
rect 3012 10304 3028 10368
rect 3092 10304 3108 10368
rect 3172 10304 3180 10368
rect 2860 10303 3180 10304
rect 6060 10368 6380 10369
rect 6060 10304 6068 10368
rect 6132 10304 6148 10368
rect 6212 10304 6228 10368
rect 6292 10304 6308 10368
rect 6372 10304 6380 10368
rect 6060 10303 6380 10304
rect 9260 10368 9580 10369
rect 9260 10304 9268 10368
rect 9332 10304 9348 10368
rect 9412 10304 9428 10368
rect 9492 10304 9508 10368
rect 9572 10304 9580 10368
rect 9260 10303 9580 10304
rect 14000 10160 34000 10192
rect 14000 10104 14186 10160
rect 14242 10104 34000 10160
rect 14000 10072 34000 10104
rect 1260 9824 1580 9825
rect 1260 9760 1268 9824
rect 1332 9760 1348 9824
rect 1412 9760 1428 9824
rect 1492 9760 1508 9824
rect 1572 9760 1580 9824
rect 1260 9759 1580 9760
rect 4460 9824 4780 9825
rect 4460 9760 4468 9824
rect 4532 9760 4548 9824
rect 4612 9760 4628 9824
rect 4692 9760 4708 9824
rect 4772 9760 4780 9824
rect 4460 9759 4780 9760
rect 7660 9824 7980 9825
rect 7660 9760 7668 9824
rect 7732 9760 7748 9824
rect 7812 9760 7828 9824
rect 7892 9760 7908 9824
rect 7972 9760 7980 9824
rect 7660 9759 7980 9760
rect 14000 9616 34000 9648
rect 14000 9560 14186 9616
rect 14242 9560 34000 9616
rect 14000 9528 34000 9560
rect 5717 9482 5783 9485
rect 7189 9482 7255 9485
rect 5717 9480 7255 9482
rect 5717 9424 5722 9480
rect 5778 9424 7194 9480
rect 7250 9424 7255 9480
rect 5717 9422 7255 9424
rect 5717 9419 5783 9422
rect 7189 9419 7255 9422
rect 7649 9346 7715 9349
rect 9121 9346 9187 9349
rect 7649 9344 9187 9346
rect 7649 9288 7654 9344
rect 7710 9288 9126 9344
rect 9182 9288 9187 9344
rect 7649 9286 9187 9288
rect 7649 9283 7715 9286
rect 9121 9283 9187 9286
rect 2860 9280 3180 9281
rect 2860 9216 2868 9280
rect 2932 9216 2948 9280
rect 3012 9216 3028 9280
rect 3092 9216 3108 9280
rect 3172 9216 3180 9280
rect 2860 9215 3180 9216
rect 6060 9280 6380 9281
rect 6060 9216 6068 9280
rect 6132 9216 6148 9280
rect 6212 9216 6228 9280
rect 6292 9216 6308 9280
rect 6372 9216 6380 9280
rect 6060 9215 6380 9216
rect 9260 9280 9580 9281
rect 9260 9216 9268 9280
rect 9332 9216 9348 9280
rect 9412 9216 9428 9280
rect 9492 9216 9508 9280
rect 9572 9216 9580 9280
rect 9260 9215 9580 9216
rect 7741 9210 7807 9213
rect 9029 9210 9095 9213
rect 7741 9208 9095 9210
rect 7741 9152 7746 9208
rect 7802 9152 9034 9208
rect 9090 9152 9095 9208
rect 7741 9150 9095 9152
rect 7741 9147 7807 9150
rect 9029 9147 9095 9150
rect 14000 9208 34000 9240
rect 14000 9152 14186 9208
rect 14242 9152 34000 9208
rect 14000 9120 34000 9152
rect 6453 9074 6519 9077
rect 8477 9074 8543 9077
rect 6453 9072 8543 9074
rect 6453 9016 6458 9072
rect 6514 9016 8482 9072
rect 8538 9016 8543 9072
rect 6453 9014 8543 9016
rect 6453 9011 6519 9014
rect 8477 9011 8543 9014
rect 6637 8938 6703 8941
rect 6821 8938 6887 8941
rect 8201 8938 8267 8941
rect 6637 8936 8267 8938
rect 6637 8880 6642 8936
rect 6698 8880 6826 8936
rect 6882 8880 8206 8936
rect 8262 8880 8267 8936
rect 6637 8878 8267 8880
rect 6637 8875 6703 8878
rect 6821 8875 6887 8878
rect 8201 8875 8267 8878
rect 5993 8802 6059 8805
rect 7465 8802 7531 8805
rect 5993 8800 7531 8802
rect 5993 8744 5998 8800
rect 6054 8744 7470 8800
rect 7526 8744 7531 8800
rect 5993 8742 7531 8744
rect 5993 8739 6059 8742
rect 7465 8739 7531 8742
rect 1260 8736 1580 8737
rect 1260 8672 1268 8736
rect 1332 8672 1348 8736
rect 1412 8672 1428 8736
rect 1492 8672 1508 8736
rect 1572 8672 1580 8736
rect 1260 8671 1580 8672
rect 4460 8736 4780 8737
rect 4460 8672 4468 8736
rect 4532 8672 4548 8736
rect 4612 8672 4628 8736
rect 4692 8672 4708 8736
rect 4772 8672 4780 8736
rect 4460 8671 4780 8672
rect 7660 8736 7980 8737
rect 7660 8672 7668 8736
rect 7732 8672 7748 8736
rect 7812 8672 7828 8736
rect 7892 8672 7908 8736
rect 7972 8672 7980 8736
rect 7660 8671 7980 8672
rect 14000 8664 34000 8696
rect 14000 8608 14278 8664
rect 14334 8608 34000 8664
rect 14000 8576 34000 8608
rect 6545 8530 6611 8533
rect 7281 8530 7347 8533
rect 6545 8528 7347 8530
rect 6545 8472 6550 8528
rect 6606 8472 7286 8528
rect 7342 8472 7347 8528
rect 6545 8470 7347 8472
rect 6545 8467 6611 8470
rect 7281 8467 7347 8470
rect 2860 8192 3180 8193
rect 2860 8128 2868 8192
rect 2932 8128 2948 8192
rect 3012 8128 3028 8192
rect 3092 8128 3108 8192
rect 3172 8128 3180 8192
rect 2860 8127 3180 8128
rect 6060 8192 6380 8193
rect 6060 8128 6068 8192
rect 6132 8128 6148 8192
rect 6212 8128 6228 8192
rect 6292 8128 6308 8192
rect 6372 8128 6380 8192
rect 6060 8127 6380 8128
rect 9260 8192 9580 8193
rect 9260 8128 9268 8192
rect 9332 8128 9348 8192
rect 9412 8128 9428 8192
rect 9492 8128 9508 8192
rect 9572 8128 9580 8192
rect 9260 8127 9580 8128
rect 14000 8120 34000 8152
rect 14000 8064 14186 8120
rect 14242 8064 34000 8120
rect 14000 8032 34000 8064
rect 14000 7712 34000 7744
rect 14000 7656 14278 7712
rect 14334 7656 34000 7712
rect 1260 7648 1580 7649
rect 1260 7584 1268 7648
rect 1332 7584 1348 7648
rect 1412 7584 1428 7648
rect 1492 7584 1508 7648
rect 1572 7584 1580 7648
rect 1260 7583 1580 7584
rect 4460 7648 4780 7649
rect 4460 7584 4468 7648
rect 4532 7584 4548 7648
rect 4612 7584 4628 7648
rect 4692 7584 4708 7648
rect 4772 7584 4780 7648
rect 4460 7583 4780 7584
rect 7660 7648 7980 7649
rect 7660 7584 7668 7648
rect 7732 7584 7748 7648
rect 7812 7584 7828 7648
rect 7892 7584 7908 7648
rect 7972 7584 7980 7648
rect 14000 7624 34000 7656
rect 7660 7583 7980 7584
rect 14000 7168 34000 7200
rect 14000 7112 14186 7168
rect 14242 7112 34000 7168
rect 2860 7104 3180 7105
rect 2860 7040 2868 7104
rect 2932 7040 2948 7104
rect 3012 7040 3028 7104
rect 3092 7040 3108 7104
rect 3172 7040 3180 7104
rect 2860 7039 3180 7040
rect 6060 7104 6380 7105
rect 6060 7040 6068 7104
rect 6132 7040 6148 7104
rect 6212 7040 6228 7104
rect 6292 7040 6308 7104
rect 6372 7040 6380 7104
rect 6060 7039 6380 7040
rect 9260 7104 9580 7105
rect 9260 7040 9268 7104
rect 9332 7040 9348 7104
rect 9412 7040 9428 7104
rect 9492 7040 9508 7104
rect 9572 7040 9580 7104
rect 14000 7080 34000 7112
rect 9260 7039 9580 7040
rect 14000 6624 34000 6656
rect 14000 6568 14186 6624
rect 14242 6568 34000 6624
rect 1260 6560 1580 6561
rect 1260 6496 1268 6560
rect 1332 6496 1348 6560
rect 1412 6496 1428 6560
rect 1492 6496 1508 6560
rect 1572 6496 1580 6560
rect 1260 6495 1580 6496
rect 4460 6560 4780 6561
rect 4460 6496 4468 6560
rect 4532 6496 4548 6560
rect 4612 6496 4628 6560
rect 4692 6496 4708 6560
rect 4772 6496 4780 6560
rect 4460 6495 4780 6496
rect 7660 6560 7980 6561
rect 7660 6496 7668 6560
rect 7732 6496 7748 6560
rect 7812 6496 7828 6560
rect 7892 6496 7908 6560
rect 7972 6496 7980 6560
rect 14000 6536 34000 6568
rect 7660 6495 7980 6496
rect 4521 6218 4587 6221
rect 6361 6218 6427 6221
rect 4521 6216 6427 6218
rect 4521 6160 4526 6216
rect 4582 6160 6366 6216
rect 6422 6160 6427 6216
rect 4521 6158 6427 6160
rect 4521 6155 4587 6158
rect 6361 6155 6427 6158
rect 14000 6216 34000 6248
rect 14000 6160 14186 6216
rect 14242 6160 34000 6216
rect 14000 6128 34000 6160
rect 2860 6016 3180 6017
rect 2860 5952 2868 6016
rect 2932 5952 2948 6016
rect 3012 5952 3028 6016
rect 3092 5952 3108 6016
rect 3172 5952 3180 6016
rect 2860 5951 3180 5952
rect 6060 6016 6380 6017
rect 6060 5952 6068 6016
rect 6132 5952 6148 6016
rect 6212 5952 6228 6016
rect 6292 5952 6308 6016
rect 6372 5952 6380 6016
rect 6060 5951 6380 5952
rect 9260 6016 9580 6017
rect 9260 5952 9268 6016
rect 9332 5952 9348 6016
rect 9412 5952 9428 6016
rect 9492 5952 9508 6016
rect 9572 5952 9580 6016
rect 9260 5951 9580 5952
rect 14000 5672 34000 5704
rect 14000 5616 14186 5672
rect 14242 5616 34000 5672
rect 14000 5584 34000 5616
rect 1260 5472 1580 5473
rect 1260 5408 1268 5472
rect 1332 5408 1348 5472
rect 1412 5408 1428 5472
rect 1492 5408 1508 5472
rect 1572 5408 1580 5472
rect 1260 5407 1580 5408
rect 4460 5472 4780 5473
rect 4460 5408 4468 5472
rect 4532 5408 4548 5472
rect 4612 5408 4628 5472
rect 4692 5408 4708 5472
rect 4772 5408 4780 5472
rect 4460 5407 4780 5408
rect 7660 5472 7980 5473
rect 7660 5408 7668 5472
rect 7732 5408 7748 5472
rect 7812 5408 7828 5472
rect 7892 5408 7908 5472
rect 7972 5408 7980 5472
rect 7660 5407 7980 5408
rect 14000 5128 34000 5160
rect 14000 5072 14278 5128
rect 14334 5072 34000 5128
rect 14000 5040 34000 5072
rect 2860 4928 3180 4929
rect 2860 4864 2868 4928
rect 2932 4864 2948 4928
rect 3012 4864 3028 4928
rect 3092 4864 3108 4928
rect 3172 4864 3180 4928
rect 2860 4863 3180 4864
rect 6060 4928 6380 4929
rect 6060 4864 6068 4928
rect 6132 4864 6148 4928
rect 6212 4864 6228 4928
rect 6292 4864 6308 4928
rect 6372 4864 6380 4928
rect 6060 4863 6380 4864
rect 9260 4928 9580 4929
rect 9260 4864 9268 4928
rect 9332 4864 9348 4928
rect 9412 4864 9428 4928
rect 9492 4864 9508 4928
rect 9572 4864 9580 4928
rect 9260 4863 9580 4864
rect 14000 4720 34000 4752
rect 14000 4664 14370 4720
rect 14426 4664 34000 4720
rect 14000 4632 34000 4664
rect 4460 4384 4780 4385
rect 4460 4320 4468 4384
rect 4532 4320 4548 4384
rect 4612 4320 4628 4384
rect 4692 4320 4708 4384
rect 4772 4320 4780 4384
rect 4460 4319 4780 4320
rect 7660 4384 7980 4385
rect 7660 4320 7668 4384
rect 7732 4320 7748 4384
rect 7812 4320 7828 4384
rect 7892 4320 7908 4384
rect 7972 4320 7980 4384
rect 7660 4319 7980 4320
rect 14000 4176 34000 4208
rect 14000 4120 14186 4176
rect 14242 4120 34000 4176
rect 14000 4088 34000 4120
rect 6060 3840 6380 3841
rect 6060 3776 6068 3840
rect 6132 3776 6148 3840
rect 6212 3776 6228 3840
rect 6292 3776 6308 3840
rect 6372 3776 6380 3840
rect 6060 3775 6380 3776
rect 9260 3840 9580 3841
rect 9260 3776 9268 3840
rect 9332 3776 9348 3840
rect 9412 3776 9428 3840
rect 9492 3776 9508 3840
rect 9572 3776 9580 3840
rect 9260 3775 9580 3776
rect 14000 3632 34000 3664
rect 14000 3576 14278 3632
rect 14334 3576 34000 3632
rect 14000 3544 34000 3576
rect 7465 3498 7531 3501
rect 4294 3496 7531 3498
rect 4294 3440 7470 3496
rect 7526 3440 7531 3496
rect 4294 3438 7531 3440
rect 4294 3362 4354 3438
rect 7465 3435 7531 3438
rect 2668 3302 4354 3362
rect 4460 3296 4780 3297
rect 4460 3232 4468 3296
rect 4532 3232 4548 3296
rect 4612 3232 4628 3296
rect 4692 3232 4708 3296
rect 4772 3232 4780 3296
rect 4460 3231 4780 3232
rect 7660 3296 7980 3297
rect 7660 3232 7668 3296
rect 7732 3232 7748 3296
rect 7812 3232 7828 3296
rect 7892 3232 7908 3296
rect 7972 3232 7980 3296
rect 7660 3231 7980 3232
rect 14000 3224 34000 3256
rect 14000 3168 14186 3224
rect 14242 3168 34000 3224
rect 14000 3136 34000 3168
rect 4429 2954 4495 2957
rect 8937 2954 9003 2957
rect 4429 2952 9003 2954
rect 4429 2896 4434 2952
rect 4490 2896 8942 2952
rect 8998 2896 9003 2952
rect 4429 2894 9003 2896
rect 4429 2891 4495 2894
rect 8937 2891 9003 2894
rect 6545 2818 6611 2821
rect 7097 2818 7163 2821
rect 6545 2816 7163 2818
rect 6545 2760 6550 2816
rect 6606 2760 7102 2816
rect 7158 2760 7163 2816
rect 6545 2758 7163 2760
rect 6545 2755 6611 2758
rect 7097 2755 7163 2758
rect 6060 2752 6380 2753
rect 6060 2688 6068 2752
rect 6132 2688 6148 2752
rect 6212 2688 6228 2752
rect 6292 2688 6308 2752
rect 6372 2688 6380 2752
rect 6060 2687 6380 2688
rect 9260 2752 9580 2753
rect 9260 2688 9268 2752
rect 9332 2688 9348 2752
rect 9412 2688 9428 2752
rect 9492 2688 9508 2752
rect 9572 2688 9580 2752
rect 9260 2687 9580 2688
rect 14000 2680 34000 2712
rect 14000 2624 14186 2680
rect 14242 2624 34000 2680
rect 14000 2592 34000 2624
rect 4460 2208 4780 2209
rect 4460 2144 4468 2208
rect 4532 2144 4548 2208
rect 4612 2144 4628 2208
rect 4692 2144 4708 2208
rect 4772 2144 4780 2208
rect 4460 2143 4780 2144
rect 7660 2208 7980 2209
rect 7660 2144 7668 2208
rect 7732 2144 7748 2208
rect 7812 2144 7828 2208
rect 7892 2144 7908 2208
rect 7972 2144 7980 2208
rect 7660 2143 7980 2144
rect 14000 2136 34000 2168
rect 14000 2080 14278 2136
rect 14334 2080 34000 2136
rect 14000 2048 34000 2080
rect 14000 1728 34000 1760
rect 14000 1672 14094 1728
rect 14150 1672 34000 1728
rect 14000 1640 34000 1672
rect 14000 1184 34000 1216
rect 14000 1128 14186 1184
rect 14242 1128 34000 1184
rect 14000 1096 34000 1128
rect 14000 640 34000 672
rect 14000 584 14370 640
rect 14426 584 34000 640
rect 14000 552 34000 584
rect 14000 232 34000 264
rect 14000 176 14186 232
rect 14242 176 34000 232
rect 14000 144 34000 176
<< via3 >>
rect 2868 11452 2932 11456
rect 2868 11396 2872 11452
rect 2872 11396 2928 11452
rect 2928 11396 2932 11452
rect 2868 11392 2932 11396
rect 2948 11452 3012 11456
rect 2948 11396 2952 11452
rect 2952 11396 3008 11452
rect 3008 11396 3012 11452
rect 2948 11392 3012 11396
rect 3028 11452 3092 11456
rect 3028 11396 3032 11452
rect 3032 11396 3088 11452
rect 3088 11396 3092 11452
rect 3028 11392 3092 11396
rect 3108 11452 3172 11456
rect 3108 11396 3112 11452
rect 3112 11396 3168 11452
rect 3168 11396 3172 11452
rect 3108 11392 3172 11396
rect 6068 11452 6132 11456
rect 6068 11396 6072 11452
rect 6072 11396 6128 11452
rect 6128 11396 6132 11452
rect 6068 11392 6132 11396
rect 6148 11452 6212 11456
rect 6148 11396 6152 11452
rect 6152 11396 6208 11452
rect 6208 11396 6212 11452
rect 6148 11392 6212 11396
rect 6228 11452 6292 11456
rect 6228 11396 6232 11452
rect 6232 11396 6288 11452
rect 6288 11396 6292 11452
rect 6228 11392 6292 11396
rect 6308 11452 6372 11456
rect 6308 11396 6312 11452
rect 6312 11396 6368 11452
rect 6368 11396 6372 11452
rect 6308 11392 6372 11396
rect 9268 11452 9332 11456
rect 9268 11396 9272 11452
rect 9272 11396 9328 11452
rect 9328 11396 9332 11452
rect 9268 11392 9332 11396
rect 9348 11452 9412 11456
rect 9348 11396 9352 11452
rect 9352 11396 9408 11452
rect 9408 11396 9412 11452
rect 9348 11392 9412 11396
rect 9428 11452 9492 11456
rect 9428 11396 9432 11452
rect 9432 11396 9488 11452
rect 9488 11396 9492 11452
rect 9428 11392 9492 11396
rect 9508 11452 9572 11456
rect 9508 11396 9512 11452
rect 9512 11396 9568 11452
rect 9568 11396 9572 11452
rect 9508 11392 9572 11396
rect 1268 10908 1332 10912
rect 1268 10852 1272 10908
rect 1272 10852 1328 10908
rect 1328 10852 1332 10908
rect 1268 10848 1332 10852
rect 1348 10908 1412 10912
rect 1348 10852 1352 10908
rect 1352 10852 1408 10908
rect 1408 10852 1412 10908
rect 1348 10848 1412 10852
rect 1428 10908 1492 10912
rect 1428 10852 1432 10908
rect 1432 10852 1488 10908
rect 1488 10852 1492 10908
rect 1428 10848 1492 10852
rect 1508 10908 1572 10912
rect 1508 10852 1512 10908
rect 1512 10852 1568 10908
rect 1568 10852 1572 10908
rect 1508 10848 1572 10852
rect 4468 10908 4532 10912
rect 4468 10852 4472 10908
rect 4472 10852 4528 10908
rect 4528 10852 4532 10908
rect 4468 10848 4532 10852
rect 4548 10908 4612 10912
rect 4548 10852 4552 10908
rect 4552 10852 4608 10908
rect 4608 10852 4612 10908
rect 4548 10848 4612 10852
rect 4628 10908 4692 10912
rect 4628 10852 4632 10908
rect 4632 10852 4688 10908
rect 4688 10852 4692 10908
rect 4628 10848 4692 10852
rect 4708 10908 4772 10912
rect 4708 10852 4712 10908
rect 4712 10852 4768 10908
rect 4768 10852 4772 10908
rect 4708 10848 4772 10852
rect 7668 10908 7732 10912
rect 7668 10852 7672 10908
rect 7672 10852 7728 10908
rect 7728 10852 7732 10908
rect 7668 10848 7732 10852
rect 7748 10908 7812 10912
rect 7748 10852 7752 10908
rect 7752 10852 7808 10908
rect 7808 10852 7812 10908
rect 7748 10848 7812 10852
rect 7828 10908 7892 10912
rect 7828 10852 7832 10908
rect 7832 10852 7888 10908
rect 7888 10852 7892 10908
rect 7828 10848 7892 10852
rect 7908 10908 7972 10912
rect 7908 10852 7912 10908
rect 7912 10852 7968 10908
rect 7968 10852 7972 10908
rect 7908 10848 7972 10852
rect 2868 10364 2932 10368
rect 2868 10308 2872 10364
rect 2872 10308 2928 10364
rect 2928 10308 2932 10364
rect 2868 10304 2932 10308
rect 2948 10364 3012 10368
rect 2948 10308 2952 10364
rect 2952 10308 3008 10364
rect 3008 10308 3012 10364
rect 2948 10304 3012 10308
rect 3028 10364 3092 10368
rect 3028 10308 3032 10364
rect 3032 10308 3088 10364
rect 3088 10308 3092 10364
rect 3028 10304 3092 10308
rect 3108 10364 3172 10368
rect 3108 10308 3112 10364
rect 3112 10308 3168 10364
rect 3168 10308 3172 10364
rect 3108 10304 3172 10308
rect 6068 10364 6132 10368
rect 6068 10308 6072 10364
rect 6072 10308 6128 10364
rect 6128 10308 6132 10364
rect 6068 10304 6132 10308
rect 6148 10364 6212 10368
rect 6148 10308 6152 10364
rect 6152 10308 6208 10364
rect 6208 10308 6212 10364
rect 6148 10304 6212 10308
rect 6228 10364 6292 10368
rect 6228 10308 6232 10364
rect 6232 10308 6288 10364
rect 6288 10308 6292 10364
rect 6228 10304 6292 10308
rect 6308 10364 6372 10368
rect 6308 10308 6312 10364
rect 6312 10308 6368 10364
rect 6368 10308 6372 10364
rect 6308 10304 6372 10308
rect 9268 10364 9332 10368
rect 9268 10308 9272 10364
rect 9272 10308 9328 10364
rect 9328 10308 9332 10364
rect 9268 10304 9332 10308
rect 9348 10364 9412 10368
rect 9348 10308 9352 10364
rect 9352 10308 9408 10364
rect 9408 10308 9412 10364
rect 9348 10304 9412 10308
rect 9428 10364 9492 10368
rect 9428 10308 9432 10364
rect 9432 10308 9488 10364
rect 9488 10308 9492 10364
rect 9428 10304 9492 10308
rect 9508 10364 9572 10368
rect 9508 10308 9512 10364
rect 9512 10308 9568 10364
rect 9568 10308 9572 10364
rect 9508 10304 9572 10308
rect 1268 9820 1332 9824
rect 1268 9764 1272 9820
rect 1272 9764 1328 9820
rect 1328 9764 1332 9820
rect 1268 9760 1332 9764
rect 1348 9820 1412 9824
rect 1348 9764 1352 9820
rect 1352 9764 1408 9820
rect 1408 9764 1412 9820
rect 1348 9760 1412 9764
rect 1428 9820 1492 9824
rect 1428 9764 1432 9820
rect 1432 9764 1488 9820
rect 1488 9764 1492 9820
rect 1428 9760 1492 9764
rect 1508 9820 1572 9824
rect 1508 9764 1512 9820
rect 1512 9764 1568 9820
rect 1568 9764 1572 9820
rect 1508 9760 1572 9764
rect 4468 9820 4532 9824
rect 4468 9764 4472 9820
rect 4472 9764 4528 9820
rect 4528 9764 4532 9820
rect 4468 9760 4532 9764
rect 4548 9820 4612 9824
rect 4548 9764 4552 9820
rect 4552 9764 4608 9820
rect 4608 9764 4612 9820
rect 4548 9760 4612 9764
rect 4628 9820 4692 9824
rect 4628 9764 4632 9820
rect 4632 9764 4688 9820
rect 4688 9764 4692 9820
rect 4628 9760 4692 9764
rect 4708 9820 4772 9824
rect 4708 9764 4712 9820
rect 4712 9764 4768 9820
rect 4768 9764 4772 9820
rect 4708 9760 4772 9764
rect 7668 9820 7732 9824
rect 7668 9764 7672 9820
rect 7672 9764 7728 9820
rect 7728 9764 7732 9820
rect 7668 9760 7732 9764
rect 7748 9820 7812 9824
rect 7748 9764 7752 9820
rect 7752 9764 7808 9820
rect 7808 9764 7812 9820
rect 7748 9760 7812 9764
rect 7828 9820 7892 9824
rect 7828 9764 7832 9820
rect 7832 9764 7888 9820
rect 7888 9764 7892 9820
rect 7828 9760 7892 9764
rect 7908 9820 7972 9824
rect 7908 9764 7912 9820
rect 7912 9764 7968 9820
rect 7968 9764 7972 9820
rect 7908 9760 7972 9764
rect 2868 9276 2932 9280
rect 2868 9220 2872 9276
rect 2872 9220 2928 9276
rect 2928 9220 2932 9276
rect 2868 9216 2932 9220
rect 2948 9276 3012 9280
rect 2948 9220 2952 9276
rect 2952 9220 3008 9276
rect 3008 9220 3012 9276
rect 2948 9216 3012 9220
rect 3028 9276 3092 9280
rect 3028 9220 3032 9276
rect 3032 9220 3088 9276
rect 3088 9220 3092 9276
rect 3028 9216 3092 9220
rect 3108 9276 3172 9280
rect 3108 9220 3112 9276
rect 3112 9220 3168 9276
rect 3168 9220 3172 9276
rect 3108 9216 3172 9220
rect 6068 9276 6132 9280
rect 6068 9220 6072 9276
rect 6072 9220 6128 9276
rect 6128 9220 6132 9276
rect 6068 9216 6132 9220
rect 6148 9276 6212 9280
rect 6148 9220 6152 9276
rect 6152 9220 6208 9276
rect 6208 9220 6212 9276
rect 6148 9216 6212 9220
rect 6228 9276 6292 9280
rect 6228 9220 6232 9276
rect 6232 9220 6288 9276
rect 6288 9220 6292 9276
rect 6228 9216 6292 9220
rect 6308 9276 6372 9280
rect 6308 9220 6312 9276
rect 6312 9220 6368 9276
rect 6368 9220 6372 9276
rect 6308 9216 6372 9220
rect 9268 9276 9332 9280
rect 9268 9220 9272 9276
rect 9272 9220 9328 9276
rect 9328 9220 9332 9276
rect 9268 9216 9332 9220
rect 9348 9276 9412 9280
rect 9348 9220 9352 9276
rect 9352 9220 9408 9276
rect 9408 9220 9412 9276
rect 9348 9216 9412 9220
rect 9428 9276 9492 9280
rect 9428 9220 9432 9276
rect 9432 9220 9488 9276
rect 9488 9220 9492 9276
rect 9428 9216 9492 9220
rect 9508 9276 9572 9280
rect 9508 9220 9512 9276
rect 9512 9220 9568 9276
rect 9568 9220 9572 9276
rect 9508 9216 9572 9220
rect 1268 8732 1332 8736
rect 1268 8676 1272 8732
rect 1272 8676 1328 8732
rect 1328 8676 1332 8732
rect 1268 8672 1332 8676
rect 1348 8732 1412 8736
rect 1348 8676 1352 8732
rect 1352 8676 1408 8732
rect 1408 8676 1412 8732
rect 1348 8672 1412 8676
rect 1428 8732 1492 8736
rect 1428 8676 1432 8732
rect 1432 8676 1488 8732
rect 1488 8676 1492 8732
rect 1428 8672 1492 8676
rect 1508 8732 1572 8736
rect 1508 8676 1512 8732
rect 1512 8676 1568 8732
rect 1568 8676 1572 8732
rect 1508 8672 1572 8676
rect 4468 8732 4532 8736
rect 4468 8676 4472 8732
rect 4472 8676 4528 8732
rect 4528 8676 4532 8732
rect 4468 8672 4532 8676
rect 4548 8732 4612 8736
rect 4548 8676 4552 8732
rect 4552 8676 4608 8732
rect 4608 8676 4612 8732
rect 4548 8672 4612 8676
rect 4628 8732 4692 8736
rect 4628 8676 4632 8732
rect 4632 8676 4688 8732
rect 4688 8676 4692 8732
rect 4628 8672 4692 8676
rect 4708 8732 4772 8736
rect 4708 8676 4712 8732
rect 4712 8676 4768 8732
rect 4768 8676 4772 8732
rect 4708 8672 4772 8676
rect 7668 8732 7732 8736
rect 7668 8676 7672 8732
rect 7672 8676 7728 8732
rect 7728 8676 7732 8732
rect 7668 8672 7732 8676
rect 7748 8732 7812 8736
rect 7748 8676 7752 8732
rect 7752 8676 7808 8732
rect 7808 8676 7812 8732
rect 7748 8672 7812 8676
rect 7828 8732 7892 8736
rect 7828 8676 7832 8732
rect 7832 8676 7888 8732
rect 7888 8676 7892 8732
rect 7828 8672 7892 8676
rect 7908 8732 7972 8736
rect 7908 8676 7912 8732
rect 7912 8676 7968 8732
rect 7968 8676 7972 8732
rect 7908 8672 7972 8676
rect 2868 8188 2932 8192
rect 2868 8132 2872 8188
rect 2872 8132 2928 8188
rect 2928 8132 2932 8188
rect 2868 8128 2932 8132
rect 2948 8188 3012 8192
rect 2948 8132 2952 8188
rect 2952 8132 3008 8188
rect 3008 8132 3012 8188
rect 2948 8128 3012 8132
rect 3028 8188 3092 8192
rect 3028 8132 3032 8188
rect 3032 8132 3088 8188
rect 3088 8132 3092 8188
rect 3028 8128 3092 8132
rect 3108 8188 3172 8192
rect 3108 8132 3112 8188
rect 3112 8132 3168 8188
rect 3168 8132 3172 8188
rect 3108 8128 3172 8132
rect 6068 8188 6132 8192
rect 6068 8132 6072 8188
rect 6072 8132 6128 8188
rect 6128 8132 6132 8188
rect 6068 8128 6132 8132
rect 6148 8188 6212 8192
rect 6148 8132 6152 8188
rect 6152 8132 6208 8188
rect 6208 8132 6212 8188
rect 6148 8128 6212 8132
rect 6228 8188 6292 8192
rect 6228 8132 6232 8188
rect 6232 8132 6288 8188
rect 6288 8132 6292 8188
rect 6228 8128 6292 8132
rect 6308 8188 6372 8192
rect 6308 8132 6312 8188
rect 6312 8132 6368 8188
rect 6368 8132 6372 8188
rect 6308 8128 6372 8132
rect 9268 8188 9332 8192
rect 9268 8132 9272 8188
rect 9272 8132 9328 8188
rect 9328 8132 9332 8188
rect 9268 8128 9332 8132
rect 9348 8188 9412 8192
rect 9348 8132 9352 8188
rect 9352 8132 9408 8188
rect 9408 8132 9412 8188
rect 9348 8128 9412 8132
rect 9428 8188 9492 8192
rect 9428 8132 9432 8188
rect 9432 8132 9488 8188
rect 9488 8132 9492 8188
rect 9428 8128 9492 8132
rect 9508 8188 9572 8192
rect 9508 8132 9512 8188
rect 9512 8132 9568 8188
rect 9568 8132 9572 8188
rect 9508 8128 9572 8132
rect 1268 7644 1332 7648
rect 1268 7588 1272 7644
rect 1272 7588 1328 7644
rect 1328 7588 1332 7644
rect 1268 7584 1332 7588
rect 1348 7644 1412 7648
rect 1348 7588 1352 7644
rect 1352 7588 1408 7644
rect 1408 7588 1412 7644
rect 1348 7584 1412 7588
rect 1428 7644 1492 7648
rect 1428 7588 1432 7644
rect 1432 7588 1488 7644
rect 1488 7588 1492 7644
rect 1428 7584 1492 7588
rect 1508 7644 1572 7648
rect 1508 7588 1512 7644
rect 1512 7588 1568 7644
rect 1568 7588 1572 7644
rect 1508 7584 1572 7588
rect 4468 7644 4532 7648
rect 4468 7588 4472 7644
rect 4472 7588 4528 7644
rect 4528 7588 4532 7644
rect 4468 7584 4532 7588
rect 4548 7644 4612 7648
rect 4548 7588 4552 7644
rect 4552 7588 4608 7644
rect 4608 7588 4612 7644
rect 4548 7584 4612 7588
rect 4628 7644 4692 7648
rect 4628 7588 4632 7644
rect 4632 7588 4688 7644
rect 4688 7588 4692 7644
rect 4628 7584 4692 7588
rect 4708 7644 4772 7648
rect 4708 7588 4712 7644
rect 4712 7588 4768 7644
rect 4768 7588 4772 7644
rect 4708 7584 4772 7588
rect 7668 7644 7732 7648
rect 7668 7588 7672 7644
rect 7672 7588 7728 7644
rect 7728 7588 7732 7644
rect 7668 7584 7732 7588
rect 7748 7644 7812 7648
rect 7748 7588 7752 7644
rect 7752 7588 7808 7644
rect 7808 7588 7812 7644
rect 7748 7584 7812 7588
rect 7828 7644 7892 7648
rect 7828 7588 7832 7644
rect 7832 7588 7888 7644
rect 7888 7588 7892 7644
rect 7828 7584 7892 7588
rect 7908 7644 7972 7648
rect 7908 7588 7912 7644
rect 7912 7588 7968 7644
rect 7968 7588 7972 7644
rect 7908 7584 7972 7588
rect 2868 7100 2932 7104
rect 2868 7044 2872 7100
rect 2872 7044 2928 7100
rect 2928 7044 2932 7100
rect 2868 7040 2932 7044
rect 2948 7100 3012 7104
rect 2948 7044 2952 7100
rect 2952 7044 3008 7100
rect 3008 7044 3012 7100
rect 2948 7040 3012 7044
rect 3028 7100 3092 7104
rect 3028 7044 3032 7100
rect 3032 7044 3088 7100
rect 3088 7044 3092 7100
rect 3028 7040 3092 7044
rect 3108 7100 3172 7104
rect 3108 7044 3112 7100
rect 3112 7044 3168 7100
rect 3168 7044 3172 7100
rect 3108 7040 3172 7044
rect 6068 7100 6132 7104
rect 6068 7044 6072 7100
rect 6072 7044 6128 7100
rect 6128 7044 6132 7100
rect 6068 7040 6132 7044
rect 6148 7100 6212 7104
rect 6148 7044 6152 7100
rect 6152 7044 6208 7100
rect 6208 7044 6212 7100
rect 6148 7040 6212 7044
rect 6228 7100 6292 7104
rect 6228 7044 6232 7100
rect 6232 7044 6288 7100
rect 6288 7044 6292 7100
rect 6228 7040 6292 7044
rect 6308 7100 6372 7104
rect 6308 7044 6312 7100
rect 6312 7044 6368 7100
rect 6368 7044 6372 7100
rect 6308 7040 6372 7044
rect 9268 7100 9332 7104
rect 9268 7044 9272 7100
rect 9272 7044 9328 7100
rect 9328 7044 9332 7100
rect 9268 7040 9332 7044
rect 9348 7100 9412 7104
rect 9348 7044 9352 7100
rect 9352 7044 9408 7100
rect 9408 7044 9412 7100
rect 9348 7040 9412 7044
rect 9428 7100 9492 7104
rect 9428 7044 9432 7100
rect 9432 7044 9488 7100
rect 9488 7044 9492 7100
rect 9428 7040 9492 7044
rect 9508 7100 9572 7104
rect 9508 7044 9512 7100
rect 9512 7044 9568 7100
rect 9568 7044 9572 7100
rect 9508 7040 9572 7044
rect 1268 6556 1332 6560
rect 1268 6500 1272 6556
rect 1272 6500 1328 6556
rect 1328 6500 1332 6556
rect 1268 6496 1332 6500
rect 1348 6556 1412 6560
rect 1348 6500 1352 6556
rect 1352 6500 1408 6556
rect 1408 6500 1412 6556
rect 1348 6496 1412 6500
rect 1428 6556 1492 6560
rect 1428 6500 1432 6556
rect 1432 6500 1488 6556
rect 1488 6500 1492 6556
rect 1428 6496 1492 6500
rect 1508 6556 1572 6560
rect 1508 6500 1512 6556
rect 1512 6500 1568 6556
rect 1568 6500 1572 6556
rect 1508 6496 1572 6500
rect 4468 6556 4532 6560
rect 4468 6500 4472 6556
rect 4472 6500 4528 6556
rect 4528 6500 4532 6556
rect 4468 6496 4532 6500
rect 4548 6556 4612 6560
rect 4548 6500 4552 6556
rect 4552 6500 4608 6556
rect 4608 6500 4612 6556
rect 4548 6496 4612 6500
rect 4628 6556 4692 6560
rect 4628 6500 4632 6556
rect 4632 6500 4688 6556
rect 4688 6500 4692 6556
rect 4628 6496 4692 6500
rect 4708 6556 4772 6560
rect 4708 6500 4712 6556
rect 4712 6500 4768 6556
rect 4768 6500 4772 6556
rect 4708 6496 4772 6500
rect 7668 6556 7732 6560
rect 7668 6500 7672 6556
rect 7672 6500 7728 6556
rect 7728 6500 7732 6556
rect 7668 6496 7732 6500
rect 7748 6556 7812 6560
rect 7748 6500 7752 6556
rect 7752 6500 7808 6556
rect 7808 6500 7812 6556
rect 7748 6496 7812 6500
rect 7828 6556 7892 6560
rect 7828 6500 7832 6556
rect 7832 6500 7888 6556
rect 7888 6500 7892 6556
rect 7828 6496 7892 6500
rect 7908 6556 7972 6560
rect 7908 6500 7912 6556
rect 7912 6500 7968 6556
rect 7968 6500 7972 6556
rect 7908 6496 7972 6500
rect 2868 6012 2932 6016
rect 2868 5956 2872 6012
rect 2872 5956 2928 6012
rect 2928 5956 2932 6012
rect 2868 5952 2932 5956
rect 2948 6012 3012 6016
rect 2948 5956 2952 6012
rect 2952 5956 3008 6012
rect 3008 5956 3012 6012
rect 2948 5952 3012 5956
rect 3028 6012 3092 6016
rect 3028 5956 3032 6012
rect 3032 5956 3088 6012
rect 3088 5956 3092 6012
rect 3028 5952 3092 5956
rect 3108 6012 3172 6016
rect 3108 5956 3112 6012
rect 3112 5956 3168 6012
rect 3168 5956 3172 6012
rect 3108 5952 3172 5956
rect 6068 6012 6132 6016
rect 6068 5956 6072 6012
rect 6072 5956 6128 6012
rect 6128 5956 6132 6012
rect 6068 5952 6132 5956
rect 6148 6012 6212 6016
rect 6148 5956 6152 6012
rect 6152 5956 6208 6012
rect 6208 5956 6212 6012
rect 6148 5952 6212 5956
rect 6228 6012 6292 6016
rect 6228 5956 6232 6012
rect 6232 5956 6288 6012
rect 6288 5956 6292 6012
rect 6228 5952 6292 5956
rect 6308 6012 6372 6016
rect 6308 5956 6312 6012
rect 6312 5956 6368 6012
rect 6368 5956 6372 6012
rect 6308 5952 6372 5956
rect 9268 6012 9332 6016
rect 9268 5956 9272 6012
rect 9272 5956 9328 6012
rect 9328 5956 9332 6012
rect 9268 5952 9332 5956
rect 9348 6012 9412 6016
rect 9348 5956 9352 6012
rect 9352 5956 9408 6012
rect 9408 5956 9412 6012
rect 9348 5952 9412 5956
rect 9428 6012 9492 6016
rect 9428 5956 9432 6012
rect 9432 5956 9488 6012
rect 9488 5956 9492 6012
rect 9428 5952 9492 5956
rect 9508 6012 9572 6016
rect 9508 5956 9512 6012
rect 9512 5956 9568 6012
rect 9568 5956 9572 6012
rect 9508 5952 9572 5956
rect 1268 5468 1332 5472
rect 1268 5412 1272 5468
rect 1272 5412 1328 5468
rect 1328 5412 1332 5468
rect 1268 5408 1332 5412
rect 1348 5468 1412 5472
rect 1348 5412 1352 5468
rect 1352 5412 1408 5468
rect 1408 5412 1412 5468
rect 1348 5408 1412 5412
rect 1428 5468 1492 5472
rect 1428 5412 1432 5468
rect 1432 5412 1488 5468
rect 1488 5412 1492 5468
rect 1428 5408 1492 5412
rect 1508 5468 1572 5472
rect 1508 5412 1512 5468
rect 1512 5412 1568 5468
rect 1568 5412 1572 5468
rect 1508 5408 1572 5412
rect 4468 5468 4532 5472
rect 4468 5412 4472 5468
rect 4472 5412 4528 5468
rect 4528 5412 4532 5468
rect 4468 5408 4532 5412
rect 4548 5468 4612 5472
rect 4548 5412 4552 5468
rect 4552 5412 4608 5468
rect 4608 5412 4612 5468
rect 4548 5408 4612 5412
rect 4628 5468 4692 5472
rect 4628 5412 4632 5468
rect 4632 5412 4688 5468
rect 4688 5412 4692 5468
rect 4628 5408 4692 5412
rect 4708 5468 4772 5472
rect 4708 5412 4712 5468
rect 4712 5412 4768 5468
rect 4768 5412 4772 5468
rect 4708 5408 4772 5412
rect 7668 5468 7732 5472
rect 7668 5412 7672 5468
rect 7672 5412 7728 5468
rect 7728 5412 7732 5468
rect 7668 5408 7732 5412
rect 7748 5468 7812 5472
rect 7748 5412 7752 5468
rect 7752 5412 7808 5468
rect 7808 5412 7812 5468
rect 7748 5408 7812 5412
rect 7828 5468 7892 5472
rect 7828 5412 7832 5468
rect 7832 5412 7888 5468
rect 7888 5412 7892 5468
rect 7828 5408 7892 5412
rect 7908 5468 7972 5472
rect 7908 5412 7912 5468
rect 7912 5412 7968 5468
rect 7968 5412 7972 5468
rect 7908 5408 7972 5412
rect 2868 4924 2932 4928
rect 2868 4868 2872 4924
rect 2872 4868 2928 4924
rect 2928 4868 2932 4924
rect 2868 4864 2932 4868
rect 2948 4924 3012 4928
rect 2948 4868 2952 4924
rect 2952 4868 3008 4924
rect 3008 4868 3012 4924
rect 2948 4864 3012 4868
rect 3028 4924 3092 4928
rect 3028 4868 3032 4924
rect 3032 4868 3088 4924
rect 3088 4868 3092 4924
rect 3028 4864 3092 4868
rect 3108 4924 3172 4928
rect 3108 4868 3112 4924
rect 3112 4868 3168 4924
rect 3168 4868 3172 4924
rect 3108 4864 3172 4868
rect 6068 4924 6132 4928
rect 6068 4868 6072 4924
rect 6072 4868 6128 4924
rect 6128 4868 6132 4924
rect 6068 4864 6132 4868
rect 6148 4924 6212 4928
rect 6148 4868 6152 4924
rect 6152 4868 6208 4924
rect 6208 4868 6212 4924
rect 6148 4864 6212 4868
rect 6228 4924 6292 4928
rect 6228 4868 6232 4924
rect 6232 4868 6288 4924
rect 6288 4868 6292 4924
rect 6228 4864 6292 4868
rect 6308 4924 6372 4928
rect 6308 4868 6312 4924
rect 6312 4868 6368 4924
rect 6368 4868 6372 4924
rect 6308 4864 6372 4868
rect 9268 4924 9332 4928
rect 9268 4868 9272 4924
rect 9272 4868 9328 4924
rect 9328 4868 9332 4924
rect 9268 4864 9332 4868
rect 9348 4924 9412 4928
rect 9348 4868 9352 4924
rect 9352 4868 9408 4924
rect 9408 4868 9412 4924
rect 9348 4864 9412 4868
rect 9428 4924 9492 4928
rect 9428 4868 9432 4924
rect 9432 4868 9488 4924
rect 9488 4868 9492 4924
rect 9428 4864 9492 4868
rect 9508 4924 9572 4928
rect 9508 4868 9512 4924
rect 9512 4868 9568 4924
rect 9568 4868 9572 4924
rect 9508 4864 9572 4868
rect 4468 4380 4532 4384
rect 4468 4324 4472 4380
rect 4472 4324 4528 4380
rect 4528 4324 4532 4380
rect 4468 4320 4532 4324
rect 4548 4380 4612 4384
rect 4548 4324 4552 4380
rect 4552 4324 4608 4380
rect 4608 4324 4612 4380
rect 4548 4320 4612 4324
rect 4628 4380 4692 4384
rect 4628 4324 4632 4380
rect 4632 4324 4688 4380
rect 4688 4324 4692 4380
rect 4628 4320 4692 4324
rect 4708 4380 4772 4384
rect 4708 4324 4712 4380
rect 4712 4324 4768 4380
rect 4768 4324 4772 4380
rect 4708 4320 4772 4324
rect 7668 4380 7732 4384
rect 7668 4324 7672 4380
rect 7672 4324 7728 4380
rect 7728 4324 7732 4380
rect 7668 4320 7732 4324
rect 7748 4380 7812 4384
rect 7748 4324 7752 4380
rect 7752 4324 7808 4380
rect 7808 4324 7812 4380
rect 7748 4320 7812 4324
rect 7828 4380 7892 4384
rect 7828 4324 7832 4380
rect 7832 4324 7888 4380
rect 7888 4324 7892 4380
rect 7828 4320 7892 4324
rect 7908 4380 7972 4384
rect 7908 4324 7912 4380
rect 7912 4324 7968 4380
rect 7968 4324 7972 4380
rect 7908 4320 7972 4324
rect 6068 3836 6132 3840
rect 6068 3780 6072 3836
rect 6072 3780 6128 3836
rect 6128 3780 6132 3836
rect 6068 3776 6132 3780
rect 6148 3836 6212 3840
rect 6148 3780 6152 3836
rect 6152 3780 6208 3836
rect 6208 3780 6212 3836
rect 6148 3776 6212 3780
rect 6228 3836 6292 3840
rect 6228 3780 6232 3836
rect 6232 3780 6288 3836
rect 6288 3780 6292 3836
rect 6228 3776 6292 3780
rect 6308 3836 6372 3840
rect 6308 3780 6312 3836
rect 6312 3780 6368 3836
rect 6368 3780 6372 3836
rect 6308 3776 6372 3780
rect 9268 3836 9332 3840
rect 9268 3780 9272 3836
rect 9272 3780 9328 3836
rect 9328 3780 9332 3836
rect 9268 3776 9332 3780
rect 9348 3836 9412 3840
rect 9348 3780 9352 3836
rect 9352 3780 9408 3836
rect 9408 3780 9412 3836
rect 9348 3776 9412 3780
rect 9428 3836 9492 3840
rect 9428 3780 9432 3836
rect 9432 3780 9488 3836
rect 9488 3780 9492 3836
rect 9428 3776 9492 3780
rect 9508 3836 9572 3840
rect 9508 3780 9512 3836
rect 9512 3780 9568 3836
rect 9568 3780 9572 3836
rect 9508 3776 9572 3780
rect 4468 3292 4532 3296
rect 4468 3236 4472 3292
rect 4472 3236 4528 3292
rect 4528 3236 4532 3292
rect 4468 3232 4532 3236
rect 4548 3292 4612 3296
rect 4548 3236 4552 3292
rect 4552 3236 4608 3292
rect 4608 3236 4612 3292
rect 4548 3232 4612 3236
rect 4628 3292 4692 3296
rect 4628 3236 4632 3292
rect 4632 3236 4688 3292
rect 4688 3236 4692 3292
rect 4628 3232 4692 3236
rect 4708 3292 4772 3296
rect 4708 3236 4712 3292
rect 4712 3236 4768 3292
rect 4768 3236 4772 3292
rect 4708 3232 4772 3236
rect 7668 3292 7732 3296
rect 7668 3236 7672 3292
rect 7672 3236 7728 3292
rect 7728 3236 7732 3292
rect 7668 3232 7732 3236
rect 7748 3292 7812 3296
rect 7748 3236 7752 3292
rect 7752 3236 7808 3292
rect 7808 3236 7812 3292
rect 7748 3232 7812 3236
rect 7828 3292 7892 3296
rect 7828 3236 7832 3292
rect 7832 3236 7888 3292
rect 7888 3236 7892 3292
rect 7828 3232 7892 3236
rect 7908 3292 7972 3296
rect 7908 3236 7912 3292
rect 7912 3236 7968 3292
rect 7968 3236 7972 3292
rect 7908 3232 7972 3236
rect 6068 2748 6132 2752
rect 6068 2692 6072 2748
rect 6072 2692 6128 2748
rect 6128 2692 6132 2748
rect 6068 2688 6132 2692
rect 6148 2748 6212 2752
rect 6148 2692 6152 2748
rect 6152 2692 6208 2748
rect 6208 2692 6212 2748
rect 6148 2688 6212 2692
rect 6228 2748 6292 2752
rect 6228 2692 6232 2748
rect 6232 2692 6288 2748
rect 6288 2692 6292 2748
rect 6228 2688 6292 2692
rect 6308 2748 6372 2752
rect 6308 2692 6312 2748
rect 6312 2692 6368 2748
rect 6368 2692 6372 2748
rect 6308 2688 6372 2692
rect 9268 2748 9332 2752
rect 9268 2692 9272 2748
rect 9272 2692 9328 2748
rect 9328 2692 9332 2748
rect 9268 2688 9332 2692
rect 9348 2748 9412 2752
rect 9348 2692 9352 2748
rect 9352 2692 9408 2748
rect 9408 2692 9412 2748
rect 9348 2688 9412 2692
rect 9428 2748 9492 2752
rect 9428 2692 9432 2748
rect 9432 2692 9488 2748
rect 9488 2692 9492 2748
rect 9428 2688 9492 2692
rect 9508 2748 9572 2752
rect 9508 2692 9512 2748
rect 9512 2692 9568 2748
rect 9568 2692 9572 2748
rect 9508 2688 9572 2692
rect 4468 2204 4532 2208
rect 4468 2148 4472 2204
rect 4472 2148 4528 2204
rect 4528 2148 4532 2204
rect 4468 2144 4532 2148
rect 4548 2204 4612 2208
rect 4548 2148 4552 2204
rect 4552 2148 4608 2204
rect 4608 2148 4612 2204
rect 4548 2144 4612 2148
rect 4628 2204 4692 2208
rect 4628 2148 4632 2204
rect 4632 2148 4688 2204
rect 4688 2148 4692 2204
rect 4628 2144 4692 2148
rect 4708 2204 4772 2208
rect 4708 2148 4712 2204
rect 4712 2148 4768 2204
rect 4768 2148 4772 2204
rect 4708 2144 4772 2148
rect 7668 2204 7732 2208
rect 7668 2148 7672 2204
rect 7672 2148 7728 2204
rect 7728 2148 7732 2204
rect 7668 2144 7732 2148
rect 7748 2204 7812 2208
rect 7748 2148 7752 2204
rect 7752 2148 7808 2204
rect 7808 2148 7812 2204
rect 7748 2144 7812 2148
rect 7828 2204 7892 2208
rect 7828 2148 7832 2204
rect 7832 2148 7888 2204
rect 7888 2148 7892 2204
rect 7828 2144 7892 2148
rect 7908 2204 7972 2208
rect 7908 2148 7912 2204
rect 7912 2148 7968 2204
rect 7968 2148 7972 2204
rect 7908 2144 7972 2148
<< metal4 >>
rect -1620 13922 -1300 13964
rect -1620 13686 -1578 13922
rect -1342 13686 -1300 13922
rect -1620 8494 -1300 13686
rect -1620 8258 -1578 8494
rect -1342 8258 -1300 8494
rect -1620 5294 -1300 8258
rect -1620 5058 -1578 5294
rect -1342 5058 -1300 5294
rect -1620 -86 -1300 5058
rect -960 13262 -640 13304
rect -960 13026 -918 13262
rect -682 13026 -640 13262
rect -960 10094 -640 13026
rect 2160 13262 2480 13964
rect 2160 13026 2202 13262
rect 2438 13026 2480 13262
rect -960 9858 -918 10094
rect -682 9858 -640 10094
rect -960 6894 -640 9858
rect -960 6658 -918 6894
rect -682 6658 -640 6894
rect -960 3694 -640 6658
rect -960 3458 -918 3694
rect -682 3458 -640 3694
rect -960 574 -640 3458
rect -300 12602 20 12644
rect -300 12366 -258 12602
rect -22 12366 20 12602
rect -300 10794 20 12366
rect -300 10558 -258 10794
rect -22 10558 20 10794
rect -300 7594 20 10558
rect -300 7358 -258 7594
rect -22 7358 20 7594
rect -300 4394 20 7358
rect -300 4158 -258 4394
rect -22 4158 20 4394
rect -300 1234 20 4158
rect 360 11942 680 11984
rect 360 11706 402 11942
rect 638 11706 680 11942
rect 360 9194 680 11706
rect 360 8958 402 9194
rect 638 8958 680 9194
rect 360 5994 680 8958
rect 360 5758 402 5994
rect 638 5758 680 5994
rect 360 2794 680 5758
rect 1260 11942 1580 12644
rect 1260 11706 1302 11942
rect 1538 11706 1580 11942
rect 1260 10912 1580 11706
rect 1260 10848 1268 10912
rect 1332 10848 1348 10912
rect 1412 10848 1428 10912
rect 1492 10848 1508 10912
rect 1572 10848 1580 10912
rect 1260 9824 1580 10848
rect 1260 9760 1268 9824
rect 1332 9760 1348 9824
rect 1412 9760 1428 9824
rect 1492 9760 1508 9824
rect 1572 9760 1580 9824
rect 1260 9194 1580 9760
rect 1260 8958 1302 9194
rect 1538 8958 1580 9194
rect 1260 8736 1580 8958
rect 1260 8672 1268 8736
rect 1332 8672 1348 8736
rect 1412 8672 1428 8736
rect 1492 8672 1508 8736
rect 1572 8672 1580 8736
rect 1260 7648 1580 8672
rect 1260 7584 1268 7648
rect 1332 7584 1348 7648
rect 1412 7584 1428 7648
rect 1492 7584 1508 7648
rect 1572 7584 1580 7648
rect 1260 6560 1580 7584
rect 1260 6496 1268 6560
rect 1332 6496 1348 6560
rect 1412 6496 1428 6560
rect 1492 6496 1508 6560
rect 1572 6496 1580 6560
rect 1260 5994 1580 6496
rect 1260 5758 1302 5994
rect 1538 5758 1580 5994
rect 1260 5472 1580 5758
rect 1260 5408 1268 5472
rect 1332 5408 1348 5472
rect 1412 5408 1428 5472
rect 1492 5408 1508 5472
rect 1572 5408 1580 5472
rect 1260 4432 1580 5408
rect 2160 10094 2480 13026
rect 3760 13922 4080 13964
rect 3760 13686 3802 13922
rect 4038 13686 4080 13922
rect 2160 9858 2202 10094
rect 2438 9858 2480 10094
rect 2160 6894 2480 9858
rect 2160 6658 2202 6894
rect 2438 6658 2480 6894
rect 2160 4480 2480 6658
rect 2860 12602 3180 12644
rect 2860 12366 2902 12602
rect 3138 12366 3180 12602
rect 2860 11456 3180 12366
rect 2860 11392 2868 11456
rect 2932 11392 2948 11456
rect 3012 11392 3028 11456
rect 3092 11392 3108 11456
rect 3172 11392 3180 11456
rect 2860 10794 3180 11392
rect 2860 10558 2902 10794
rect 3138 10558 3180 10794
rect 2860 10368 3180 10558
rect 2860 10304 2868 10368
rect 2932 10304 2948 10368
rect 3012 10304 3028 10368
rect 3092 10304 3108 10368
rect 3172 10304 3180 10368
rect 2860 9280 3180 10304
rect 2860 9216 2868 9280
rect 2932 9216 2948 9280
rect 3012 9216 3028 9280
rect 3092 9216 3108 9280
rect 3172 9216 3180 9280
rect 2860 8192 3180 9216
rect 2860 8128 2868 8192
rect 2932 8128 2948 8192
rect 3012 8128 3028 8192
rect 3092 8128 3108 8192
rect 3172 8128 3180 8192
rect 2860 7594 3180 8128
rect 2860 7358 2902 7594
rect 3138 7358 3180 7594
rect 2860 7104 3180 7358
rect 2860 7040 2868 7104
rect 2932 7040 2948 7104
rect 3012 7040 3028 7104
rect 3092 7040 3108 7104
rect 3172 7040 3180 7104
rect 2860 6016 3180 7040
rect 2860 5952 2868 6016
rect 2932 5952 2948 6016
rect 3012 5952 3028 6016
rect 3092 5952 3108 6016
rect 3172 5952 3180 6016
rect 2860 4928 3180 5952
rect 2860 4864 2868 4928
rect 2932 4864 2948 4928
rect 3012 4864 3028 4928
rect 3092 4864 3108 4928
rect 3172 4864 3180 4928
rect 2860 4432 3180 4864
rect 3760 8494 4080 13686
rect 5360 13262 5680 13964
rect 5360 13026 5402 13262
rect 5638 13026 5680 13262
rect 3760 8258 3802 8494
rect 4038 8258 4080 8494
rect 3760 5294 4080 8258
rect 3760 5058 3802 5294
rect 4038 5058 4080 5294
rect 360 2558 402 2794
rect 638 2558 680 2794
rect 360 1894 680 2558
rect 360 1658 402 1894
rect 638 1658 680 1894
rect 360 1616 680 1658
rect 1260 1894 1580 2128
rect 1260 1658 1302 1894
rect 1538 1658 1580 1894
rect -300 998 -258 1234
rect -22 998 20 1234
rect -300 956 20 998
rect 1260 956 1580 1658
rect -960 338 -918 574
rect -682 338 -640 574
rect -960 296 -640 338
rect 2160 574 2480 2080
rect 2860 1234 3180 2128
rect 2860 998 2902 1234
rect 3138 998 3180 1234
rect 2860 956 3180 998
rect 2160 338 2202 574
rect 2438 338 2480 574
rect -1620 -322 -1578 -86
rect -1342 -322 -1300 -86
rect -1620 -364 -1300 -322
rect 2160 -364 2480 338
rect 3760 -86 4080 5058
rect 4460 11942 4780 12644
rect 4460 11706 4502 11942
rect 4738 11706 4780 11942
rect 4460 10912 4780 11706
rect 4460 10848 4468 10912
rect 4532 10848 4548 10912
rect 4612 10848 4628 10912
rect 4692 10848 4708 10912
rect 4772 10848 4780 10912
rect 4460 9824 4780 10848
rect 4460 9760 4468 9824
rect 4532 9760 4548 9824
rect 4612 9760 4628 9824
rect 4692 9760 4708 9824
rect 4772 9760 4780 9824
rect 4460 9194 4780 9760
rect 4460 8958 4502 9194
rect 4738 8958 4780 9194
rect 4460 8736 4780 8958
rect 4460 8672 4468 8736
rect 4532 8672 4548 8736
rect 4612 8672 4628 8736
rect 4692 8672 4708 8736
rect 4772 8672 4780 8736
rect 4460 7648 4780 8672
rect 4460 7584 4468 7648
rect 4532 7584 4548 7648
rect 4612 7584 4628 7648
rect 4692 7584 4708 7648
rect 4772 7584 4780 7648
rect 4460 6560 4780 7584
rect 4460 6496 4468 6560
rect 4532 6496 4548 6560
rect 4612 6496 4628 6560
rect 4692 6496 4708 6560
rect 4772 6496 4780 6560
rect 4460 5994 4780 6496
rect 4460 5758 4502 5994
rect 4738 5758 4780 5994
rect 4460 5472 4780 5758
rect 4460 5408 4468 5472
rect 4532 5408 4548 5472
rect 4612 5408 4628 5472
rect 4692 5408 4708 5472
rect 4772 5408 4780 5472
rect 4460 4384 4780 5408
rect 4460 4320 4468 4384
rect 4532 4320 4548 4384
rect 4612 4320 4628 4384
rect 4692 4320 4708 4384
rect 4772 4320 4780 4384
rect 4460 3296 4780 4320
rect 4460 3232 4468 3296
rect 4532 3232 4548 3296
rect 4612 3232 4628 3296
rect 4692 3232 4708 3296
rect 4772 3232 4780 3296
rect 4460 2794 4780 3232
rect 4460 2558 4502 2794
rect 4738 2558 4780 2794
rect 4460 2208 4780 2558
rect 4460 2144 4468 2208
rect 4532 2144 4548 2208
rect 4612 2144 4628 2208
rect 4692 2144 4708 2208
rect 4772 2144 4780 2208
rect 4460 1894 4780 2144
rect 4460 1658 4502 1894
rect 4738 1658 4780 1894
rect 4460 956 4780 1658
rect 5360 10094 5680 13026
rect 6960 13922 7280 13964
rect 6960 13686 7002 13922
rect 7238 13686 7280 13922
rect 5360 9858 5402 10094
rect 5638 9858 5680 10094
rect 5360 6894 5680 9858
rect 5360 6658 5402 6894
rect 5638 6658 5680 6894
rect 5360 3694 5680 6658
rect 5360 3458 5402 3694
rect 5638 3458 5680 3694
rect 3760 -322 3802 -86
rect 4038 -322 4080 -86
rect 3760 -364 4080 -322
rect 5360 574 5680 3458
rect 6060 12602 6380 12644
rect 6060 12366 6102 12602
rect 6338 12366 6380 12602
rect 6060 11456 6380 12366
rect 6060 11392 6068 11456
rect 6132 11392 6148 11456
rect 6212 11392 6228 11456
rect 6292 11392 6308 11456
rect 6372 11392 6380 11456
rect 6060 10794 6380 11392
rect 6060 10558 6102 10794
rect 6338 10558 6380 10794
rect 6060 10368 6380 10558
rect 6060 10304 6068 10368
rect 6132 10304 6148 10368
rect 6212 10304 6228 10368
rect 6292 10304 6308 10368
rect 6372 10304 6380 10368
rect 6060 9280 6380 10304
rect 6060 9216 6068 9280
rect 6132 9216 6148 9280
rect 6212 9216 6228 9280
rect 6292 9216 6308 9280
rect 6372 9216 6380 9280
rect 6060 8192 6380 9216
rect 6060 8128 6068 8192
rect 6132 8128 6148 8192
rect 6212 8128 6228 8192
rect 6292 8128 6308 8192
rect 6372 8128 6380 8192
rect 6060 7594 6380 8128
rect 6060 7358 6102 7594
rect 6338 7358 6380 7594
rect 6060 7104 6380 7358
rect 6060 7040 6068 7104
rect 6132 7040 6148 7104
rect 6212 7040 6228 7104
rect 6292 7040 6308 7104
rect 6372 7040 6380 7104
rect 6060 6016 6380 7040
rect 6060 5952 6068 6016
rect 6132 5952 6148 6016
rect 6212 5952 6228 6016
rect 6292 5952 6308 6016
rect 6372 5952 6380 6016
rect 6060 4928 6380 5952
rect 6060 4864 6068 4928
rect 6132 4864 6148 4928
rect 6212 4864 6228 4928
rect 6292 4864 6308 4928
rect 6372 4864 6380 4928
rect 6060 4394 6380 4864
rect 6060 4158 6102 4394
rect 6338 4158 6380 4394
rect 6060 3840 6380 4158
rect 6060 3776 6068 3840
rect 6132 3776 6148 3840
rect 6212 3776 6228 3840
rect 6292 3776 6308 3840
rect 6372 3776 6380 3840
rect 6060 2752 6380 3776
rect 6060 2688 6068 2752
rect 6132 2688 6148 2752
rect 6212 2688 6228 2752
rect 6292 2688 6308 2752
rect 6372 2688 6380 2752
rect 6060 1234 6380 2688
rect 6060 998 6102 1234
rect 6338 998 6380 1234
rect 6060 956 6380 998
rect 6960 8494 7280 13686
rect 8560 13262 8880 13964
rect 12064 13922 12384 13964
rect 12064 13686 12106 13922
rect 12342 13686 12384 13922
rect 8560 13026 8602 13262
rect 8838 13026 8880 13262
rect 6960 8258 7002 8494
rect 7238 8258 7280 8494
rect 6960 5294 7280 8258
rect 6960 5058 7002 5294
rect 7238 5058 7280 5294
rect 5360 338 5402 574
rect 5638 338 5680 574
rect 5360 -364 5680 338
rect 6960 -86 7280 5058
rect 7660 11942 7980 12644
rect 7660 11706 7702 11942
rect 7938 11706 7980 11942
rect 7660 10912 7980 11706
rect 7660 10848 7668 10912
rect 7732 10848 7748 10912
rect 7812 10848 7828 10912
rect 7892 10848 7908 10912
rect 7972 10848 7980 10912
rect 7660 9824 7980 10848
rect 7660 9760 7668 9824
rect 7732 9760 7748 9824
rect 7812 9760 7828 9824
rect 7892 9760 7908 9824
rect 7972 9760 7980 9824
rect 7660 9194 7980 9760
rect 7660 8958 7702 9194
rect 7938 8958 7980 9194
rect 7660 8736 7980 8958
rect 7660 8672 7668 8736
rect 7732 8672 7748 8736
rect 7812 8672 7828 8736
rect 7892 8672 7908 8736
rect 7972 8672 7980 8736
rect 7660 7648 7980 8672
rect 7660 7584 7668 7648
rect 7732 7584 7748 7648
rect 7812 7584 7828 7648
rect 7892 7584 7908 7648
rect 7972 7584 7980 7648
rect 7660 6560 7980 7584
rect 7660 6496 7668 6560
rect 7732 6496 7748 6560
rect 7812 6496 7828 6560
rect 7892 6496 7908 6560
rect 7972 6496 7980 6560
rect 7660 5994 7980 6496
rect 7660 5758 7702 5994
rect 7938 5758 7980 5994
rect 7660 5472 7980 5758
rect 7660 5408 7668 5472
rect 7732 5408 7748 5472
rect 7812 5408 7828 5472
rect 7892 5408 7908 5472
rect 7972 5408 7980 5472
rect 7660 4384 7980 5408
rect 7660 4320 7668 4384
rect 7732 4320 7748 4384
rect 7812 4320 7828 4384
rect 7892 4320 7908 4384
rect 7972 4320 7980 4384
rect 7660 3296 7980 4320
rect 7660 3232 7668 3296
rect 7732 3232 7748 3296
rect 7812 3232 7828 3296
rect 7892 3232 7908 3296
rect 7972 3232 7980 3296
rect 7660 2794 7980 3232
rect 7660 2558 7702 2794
rect 7938 2558 7980 2794
rect 7660 2208 7980 2558
rect 7660 2144 7668 2208
rect 7732 2144 7748 2208
rect 7812 2144 7828 2208
rect 7892 2144 7908 2208
rect 7972 2144 7980 2208
rect 7660 1894 7980 2144
rect 7660 1658 7702 1894
rect 7938 1658 7980 1894
rect 7660 956 7980 1658
rect 8560 10094 8880 13026
rect 11404 13262 11724 13304
rect 11404 13026 11446 13262
rect 11682 13026 11724 13262
rect 8560 9858 8602 10094
rect 8838 9858 8880 10094
rect 8560 6894 8880 9858
rect 8560 6658 8602 6894
rect 8838 6658 8880 6894
rect 8560 3694 8880 6658
rect 8560 3458 8602 3694
rect 8838 3458 8880 3694
rect 6960 -322 7002 -86
rect 7238 -322 7280 -86
rect 6960 -364 7280 -322
rect 8560 574 8880 3458
rect 9260 12602 9580 12644
rect 9260 12366 9302 12602
rect 9538 12366 9580 12602
rect 9260 11456 9580 12366
rect 10744 12602 11064 12644
rect 10744 12366 10786 12602
rect 11022 12366 11064 12602
rect 9260 11392 9268 11456
rect 9332 11392 9348 11456
rect 9412 11392 9428 11456
rect 9492 11392 9508 11456
rect 9572 11392 9580 11456
rect 9260 10794 9580 11392
rect 9260 10558 9302 10794
rect 9538 10558 9580 10794
rect 9260 10368 9580 10558
rect 9260 10304 9268 10368
rect 9332 10304 9348 10368
rect 9412 10304 9428 10368
rect 9492 10304 9508 10368
rect 9572 10304 9580 10368
rect 9260 9280 9580 10304
rect 9260 9216 9268 9280
rect 9332 9216 9348 9280
rect 9412 9216 9428 9280
rect 9492 9216 9508 9280
rect 9572 9216 9580 9280
rect 9260 8192 9580 9216
rect 9260 8128 9268 8192
rect 9332 8128 9348 8192
rect 9412 8128 9428 8192
rect 9492 8128 9508 8192
rect 9572 8128 9580 8192
rect 9260 7594 9580 8128
rect 9260 7358 9302 7594
rect 9538 7358 9580 7594
rect 9260 7104 9580 7358
rect 9260 7040 9268 7104
rect 9332 7040 9348 7104
rect 9412 7040 9428 7104
rect 9492 7040 9508 7104
rect 9572 7040 9580 7104
rect 9260 6016 9580 7040
rect 9260 5952 9268 6016
rect 9332 5952 9348 6016
rect 9412 5952 9428 6016
rect 9492 5952 9508 6016
rect 9572 5952 9580 6016
rect 9260 4928 9580 5952
rect 9260 4864 9268 4928
rect 9332 4864 9348 4928
rect 9412 4864 9428 4928
rect 9492 4864 9508 4928
rect 9572 4864 9580 4928
rect 9260 4394 9580 4864
rect 9260 4158 9302 4394
rect 9538 4158 9580 4394
rect 9260 3840 9580 4158
rect 9260 3776 9268 3840
rect 9332 3776 9348 3840
rect 9412 3776 9428 3840
rect 9492 3776 9508 3840
rect 9572 3776 9580 3840
rect 9260 2752 9580 3776
rect 9260 2688 9268 2752
rect 9332 2688 9348 2752
rect 9412 2688 9428 2752
rect 9492 2688 9508 2752
rect 9572 2688 9580 2752
rect 9260 1234 9580 2688
rect 10084 11942 10404 11984
rect 10084 11706 10126 11942
rect 10362 11706 10404 11942
rect 10084 9194 10404 11706
rect 10084 8958 10126 9194
rect 10362 8958 10404 9194
rect 10084 5994 10404 8958
rect 10084 5758 10126 5994
rect 10362 5758 10404 5994
rect 10084 2794 10404 5758
rect 10084 2558 10126 2794
rect 10362 2558 10404 2794
rect 10084 1894 10404 2558
rect 10084 1658 10126 1894
rect 10362 1658 10404 1894
rect 10084 1616 10404 1658
rect 10744 10794 11064 12366
rect 10744 10558 10786 10794
rect 11022 10558 11064 10794
rect 10744 7594 11064 10558
rect 10744 7358 10786 7594
rect 11022 7358 11064 7594
rect 10744 4394 11064 7358
rect 10744 4158 10786 4394
rect 11022 4158 11064 4394
rect 9260 998 9302 1234
rect 9538 998 9580 1234
rect 9260 956 9580 998
rect 10744 1234 11064 4158
rect 10744 998 10786 1234
rect 11022 998 11064 1234
rect 10744 956 11064 998
rect 11404 10094 11724 13026
rect 11404 9858 11446 10094
rect 11682 9858 11724 10094
rect 11404 6894 11724 9858
rect 11404 6658 11446 6894
rect 11682 6658 11724 6894
rect 11404 3694 11724 6658
rect 11404 3458 11446 3694
rect 11682 3458 11724 3694
rect 8560 338 8602 574
rect 8838 338 8880 574
rect 8560 -364 8880 338
rect 11404 574 11724 3458
rect 11404 338 11446 574
rect 11682 338 11724 574
rect 11404 296 11724 338
rect 12064 8494 12384 13686
rect 12064 8258 12106 8494
rect 12342 8258 12384 8494
rect 12064 5294 12384 8258
rect 12064 5058 12106 5294
rect 12342 5058 12384 5294
rect 12064 -86 12384 5058
rect 12064 -322 12106 -86
rect 12342 -322 12384 -86
rect 12064 -364 12384 -322
<< via4 >>
rect -1578 13686 -1342 13922
rect -1578 8258 -1342 8494
rect -1578 5058 -1342 5294
rect -918 13026 -682 13262
rect 2202 13026 2438 13262
rect -918 9858 -682 10094
rect -918 6658 -682 6894
rect -918 3458 -682 3694
rect -258 12366 -22 12602
rect -258 10558 -22 10794
rect -258 7358 -22 7594
rect -258 4158 -22 4394
rect 402 11706 638 11942
rect 402 8958 638 9194
rect 402 5758 638 5994
rect 1302 11706 1538 11942
rect 1302 8958 1538 9194
rect 1302 5758 1538 5994
rect 3802 13686 4038 13922
rect 2202 9858 2438 10094
rect 2202 6658 2438 6894
rect 2902 12366 3138 12602
rect 2902 10558 3138 10794
rect 2902 7358 3138 7594
rect 5402 13026 5638 13262
rect 3802 8258 4038 8494
rect 3802 5058 4038 5294
rect 402 2558 638 2794
rect 402 1658 638 1894
rect 1302 1658 1538 1894
rect -258 998 -22 1234
rect -918 338 -682 574
rect 2902 998 3138 1234
rect 2202 338 2438 574
rect -1578 -322 -1342 -86
rect 4502 11706 4738 11942
rect 4502 8958 4738 9194
rect 4502 5758 4738 5994
rect 4502 2558 4738 2794
rect 4502 1658 4738 1894
rect 7002 13686 7238 13922
rect 5402 9858 5638 10094
rect 5402 6658 5638 6894
rect 5402 3458 5638 3694
rect 3802 -322 4038 -86
rect 6102 12366 6338 12602
rect 6102 10558 6338 10794
rect 6102 7358 6338 7594
rect 6102 4158 6338 4394
rect 6102 998 6338 1234
rect 12106 13686 12342 13922
rect 8602 13026 8838 13262
rect 7002 8258 7238 8494
rect 7002 5058 7238 5294
rect 5402 338 5638 574
rect 7702 11706 7938 11942
rect 7702 8958 7938 9194
rect 7702 5758 7938 5994
rect 7702 2558 7938 2794
rect 7702 1658 7938 1894
rect 11446 13026 11682 13262
rect 8602 9858 8838 10094
rect 8602 6658 8838 6894
rect 8602 3458 8838 3694
rect 7002 -322 7238 -86
rect 9302 12366 9538 12602
rect 10786 12366 11022 12602
rect 9302 10558 9538 10794
rect 9302 7358 9538 7594
rect 9302 4158 9538 4394
rect 10126 11706 10362 11942
rect 10126 8958 10362 9194
rect 10126 5758 10362 5994
rect 10126 2558 10362 2794
rect 10126 1658 10362 1894
rect 10786 10558 11022 10794
rect 10786 7358 11022 7594
rect 10786 4158 11022 4394
rect 9302 998 9538 1234
rect 10786 998 11022 1234
rect 11446 9858 11682 10094
rect 11446 6658 11682 6894
rect 11446 3458 11682 3694
rect 8602 338 8838 574
rect 11446 338 11682 574
rect 12106 8258 12342 8494
rect 12106 5058 12342 5294
rect 12106 -322 12342 -86
<< metal5 >>
rect -1620 13922 12384 13964
rect -1620 13686 -1578 13922
rect -1342 13686 3802 13922
rect 4038 13686 7002 13922
rect 7238 13686 12106 13922
rect 12342 13686 12384 13922
rect -1620 13644 12384 13686
rect -960 13262 11724 13304
rect -960 13026 -918 13262
rect -682 13026 2202 13262
rect 2438 13026 5402 13262
rect 5638 13026 8602 13262
rect 8838 13026 11446 13262
rect 11682 13026 11724 13262
rect -960 12984 11724 13026
rect -300 12602 11064 12644
rect -300 12366 -258 12602
rect -22 12366 2902 12602
rect 3138 12366 6102 12602
rect 6338 12366 9302 12602
rect 9538 12366 10786 12602
rect 11022 12366 11064 12602
rect -300 12324 11064 12366
rect 360 11942 10404 11984
rect 360 11706 402 11942
rect 638 11706 1302 11942
rect 1538 11706 4502 11942
rect 4738 11706 7702 11942
rect 7938 11706 10126 11942
rect 10362 11706 10404 11942
rect 360 11664 10404 11706
rect -300 10794 11064 10836
rect -300 10558 -258 10794
rect -22 10558 2902 10794
rect 3138 10558 6102 10794
rect 6338 10558 9302 10794
rect 9538 10558 10786 10794
rect 11022 10558 11064 10794
rect -300 10516 11064 10558
rect -1620 10094 12384 10136
rect -1620 9858 -918 10094
rect -682 9858 2202 10094
rect 2438 9858 5402 10094
rect 5638 9858 8602 10094
rect 8838 9858 11446 10094
rect 11682 9858 12384 10094
rect -1620 9816 12384 9858
rect -300 9194 11064 9236
rect -300 8958 402 9194
rect 638 8958 1302 9194
rect 1538 8958 4502 9194
rect 4738 8958 7702 9194
rect 7938 8958 10126 9194
rect 10362 8958 11064 9194
rect -300 8916 11064 8958
rect -1620 8494 12384 8536
rect -1620 8258 -1578 8494
rect -1342 8258 3802 8494
rect 4038 8258 7002 8494
rect 7238 8258 12106 8494
rect 12342 8258 12384 8494
rect -1620 8216 12384 8258
rect -300 7594 11064 7636
rect -300 7358 -258 7594
rect -22 7358 2902 7594
rect 3138 7358 6102 7594
rect 6338 7358 9302 7594
rect 9538 7358 10786 7594
rect 11022 7358 11064 7594
rect -300 7316 11064 7358
rect -1620 6894 12384 6936
rect -1620 6658 -918 6894
rect -682 6658 2202 6894
rect 2438 6658 5402 6894
rect 5638 6658 8602 6894
rect 8838 6658 11446 6894
rect 11682 6658 12384 6894
rect -1620 6616 12384 6658
rect -300 5994 11064 6036
rect -300 5758 402 5994
rect 638 5758 1302 5994
rect 1538 5758 4502 5994
rect 4738 5758 7702 5994
rect 7938 5758 10126 5994
rect 10362 5758 11064 5994
rect -300 5716 11064 5758
rect -1620 5294 12384 5336
rect -1620 5058 -1578 5294
rect -1342 5058 3802 5294
rect 4038 5058 7002 5294
rect 7238 5058 12106 5294
rect 12342 5058 12384 5294
rect -1620 5016 12384 5058
rect -300 4394 11064 4436
rect -300 4158 -258 4394
rect -22 4158 6102 4394
rect 6338 4158 9302 4394
rect 9538 4158 10786 4394
rect 11022 4158 11064 4394
rect -300 4116 11064 4158
rect -1620 3694 12384 3736
rect -1620 3458 -918 3694
rect -682 3458 5402 3694
rect 5638 3458 8602 3694
rect 8838 3458 11446 3694
rect 11682 3458 12384 3694
rect -1620 3416 12384 3458
rect -300 2794 11064 2836
rect -300 2558 402 2794
rect 638 2558 4502 2794
rect 4738 2558 7702 2794
rect 7938 2558 10126 2794
rect 10362 2558 11064 2794
rect -300 2516 11064 2558
rect 360 1894 10404 1936
rect 360 1658 402 1894
rect 638 1658 1302 1894
rect 1538 1658 4502 1894
rect 4738 1658 7702 1894
rect 7938 1658 10126 1894
rect 10362 1658 10404 1894
rect 360 1616 10404 1658
rect -300 1234 11064 1276
rect -300 998 -258 1234
rect -22 998 2902 1234
rect 3138 998 6102 1234
rect 6338 998 9302 1234
rect 9538 998 10786 1234
rect 11022 998 11064 1234
rect -300 956 11064 998
rect -960 574 11724 616
rect -960 338 -918 574
rect -682 338 2202 574
rect 2438 338 5402 574
rect 5638 338 8602 574
rect 8838 338 11446 574
rect 11682 338 11724 574
rect -960 296 11724 338
rect -1620 -86 12384 -44
rect -1620 -322 -1578 -86
rect -1342 -322 3802 -86
rect 4038 -322 7002 -86
rect 7238 -322 12106 -86
rect 12342 -322 12384 -86
rect -1620 -364 12384 -322
use gpio_logic_high  gpio_logic_high
timestamp 1621458646
transform 1 0 1196 0 1 2480
box -38 -48 1602 1136
use sky130_fd_sc_hd__decap_8  FILLER_2_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 3496 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 3496 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28
timestamp 1618914159
transform 1 0 3496 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 3220 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1618914159
transform 1 0 3220 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1618914159
transform 1 0 3220 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 4232 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36
timestamp 1618914159
transform 1 0 4232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 4416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 5060 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 4048 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _104_
timestamp 1618914159
transform 1 0 4324 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1618914159
transform 1 0 5980 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 6348 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 5888 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34
timestamp 1618914159
transform 1 0 5888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 5336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 5612 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _057_
timestamp 1618914159
transform 1 0 6072 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp 1618914159
transform 1 0 5980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _096_
timestamp 1618914159
transform 1 0 6716 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _095_
timestamp 1618914159
transform 1 0 6164 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _094_
timestamp 1618914159
transform 1 0 6256 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_2_77
timestamp 1618914159
transform 1 0 8004 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1618914159
transform 1 0 8096 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output12
timestamp 1618914159
transform 1 0 8096 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1618914159
transform 1 0 8188 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_84
timestamp 1618914159
transform 1 0 8648 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output9
timestamp 1618914159
transform 1 0 8832 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output8
timestamp 1618914159
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1618914159
transform 1 0 8556 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1618914159
transform 1 0 8464 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 8556 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _080_
timestamp 1618914159
transform 1 0 8556 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_92
timestamp 1618914159
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1618914159
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1618914159
transform -1 0 9844 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1618914159
transform -1 0 9844 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1618914159
transform -1 0 9844 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _103_
timestamp 1618914159
transform 1 0 4324 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _107_
timestamp 1618914159
transform 1 0 4048 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1618914159
transform 1 0 3220 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1618914159
transform 1 0 3220 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_28
timestamp 1618914159
transform 1 0 3496 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_28
timestamp 1618914159
transform 1 0 3496 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1618914159
transform 1 0 4232 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _042_
timestamp 1618914159
transform 1 0 6164 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _045_
timestamp 1618914159
transform 1 0 5980 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp 1618914159
transform 1 0 6348 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 6624 0 1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 6532 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1618914159
transform 1 0 5888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_58
timestamp 1618914159
transform 1 0 6256 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_60
timestamp 1618914159
transform 1 0 6440 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__nand2b_1  _073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 8740 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__ebufn_2  _083_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 8556 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1618914159
transform -1 0 9844 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1618914159
transform -1 0 9844 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1618914159
transform 1 0 8464 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output11
timestamp 1618914159
transform 1 0 9200 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_92
timestamp 1618914159
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1618914159
transform 1 0 920 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1618914159
transform 1 0 920 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 1196 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1618914159
transform 1 0 2300 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1618914159
transform 1 0 1196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1618914159
transform 1 0 2300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _063_
timestamp 1618914159
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _076_
timestamp 1618914159
transform 1 0 3772 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _101_
timestamp 1618914159
transform 1 0 4324 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _102_
timestamp 1618914159
transform 1 0 4324 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1618914159
transform 1 0 3588 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_serial_clock
timestamp 1618914159
transform 1 0 4048 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_27
timestamp 1618914159
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 3680 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1618914159
transform 1 0 3404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1618914159
transform 1 0 6164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1618914159
transform 1 0 6164 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1618914159
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _048_
timestamp 1618914159
transform 1 0 6256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _047_
timestamp 1618914159
transform 1 0 6348 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_61
timestamp 1618914159
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1618914159
transform 1 0 6624 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output16
timestamp 1618914159
transform 1 0 7268 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _061_
timestamp 1618914159
transform 1 0 6716 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp 1618914159
transform 1 0 6992 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _109_
timestamp 1618914159
transform 1 0 6808 0 1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _093_
timestamp 1618914159
transform 1 0 7636 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1618914159
transform -1 0 9844 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1618914159
transform -1 0 9844 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1618914159
transform 1 0 8924 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output13
timestamp 1618914159
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_88
timestamp 1618914159
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1618914159
transform 1 0 920 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1618914159
transform 1 0 920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1618914159
transform 1 0 1196 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1618914159
transform 1 0 2300 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1618914159
transform 1 0 1196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_15
timestamp 1618914159
transform 1 0 2300 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_23
timestamp 1618914159
transform 1 0 3036 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_30
timestamp 1618914159
transform 1 0 3680 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_27
timestamp 1618914159
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1618914159
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1618914159
transform 1 0 3496 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1618914159
transform 1 0 3588 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _051_
timestamp 1618914159
transform 1 0 3772 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _050_
timestamp 1618914159
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 1618914159
transform 1 0 4232 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _100_
timestamp 1618914159
transform 1 0 4324 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _089_
timestamp 1618914159
transform 1 0 4508 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _046_
timestamp 1618914159
transform 1 0 6256 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _049_
timestamp 1618914159
transform 1 0 6532 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _088_
timestamp 1618914159
transform 1 0 6348 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _090_
timestamp 1618914159
transform 1 0 6992 0 -1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1618914159
transform 1 0 6164 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_64
timestamp 1618914159
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp 1618914159
transform 1 0 8188 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _059_
timestamp 1618914159
transform 1 0 8924 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _070_
timestamp 1618914159
transform 1 0 8924 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1618914159
transform -1 0 9844 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1618914159
transform -1 0 9844 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1618914159
transform 1 0 8832 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output14
timestamp 1618914159
transform 1 0 9200 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output15
timestamp 1618914159
transform 1 0 8464 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_92
timestamp 1618914159
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1618914159
transform 1 0 920 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1618914159
transform 1 0 920 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1618914159
transform 1 0 1196 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1618914159
transform 1 0 2300 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1618914159
transform 1 0 1196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1618914159
transform 1 0 2300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp 1618914159
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_27
timestamp 1618914159
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_34
timestamp 1618914159
transform 1 0 4048 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1618914159
transform 1 0 3680 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 1618914159
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1618914159
transform 1 0 3588 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _068_
timestamp 1618914159
transform 1 0 4140 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _041_
timestamp 1618914159
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 4324 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _099_
timestamp 1618914159
transform 1 0 4416 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _085_
timestamp 1618914159
transform 1 0 6348 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _106_
timestamp 1618914159
transform 1 0 6256 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1618914159
transform 1 0 6164 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_58
timestamp 1618914159
transform 1 0 6256 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output18
timestamp 1618914159
transform 1 0 8464 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_4  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 8096 0 -1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp 1618914159
transform 1 0 8188 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1618914159
transform 1 0 9108 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_92
timestamp 1618914159
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output17
timestamp 1618914159
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1618914159
transform 1 0 8832 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1618914159
transform -1 0 9844 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1618914159
transform -1 0 9844 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 8924 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1618914159
transform 1 0 920 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1618914159
transform 1 0 920 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1618914159
transform 1 0 920 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1618914159
transform 1 0 1196 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1618914159
transform 1 0 2300 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1618914159
transform 1 0 1196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1618914159
transform 1 0 2300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1618914159
transform 1 0 1196 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1618914159
transform 1 0 2300 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_30
timestamp 1618914159
transform 1 0 3680 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1618914159
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_30
timestamp 1618914159
transform 1 0 3680 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_27
timestamp 1618914159
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1618914159
transform 1 0 3588 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1618914159
transform 1 0 3588 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_38
timestamp 1618914159
transform 1 0 4416 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_39
timestamp 1618914159
transform 1 0 4508 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_serial_clock
timestamp 1618914159
transform 1 0 5060 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _065_
timestamp 1618914159
transform 1 0 4416 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _064_
timestamp 1618914159
transform 1 0 4692 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _044_
timestamp 1618914159
transform 1 0 4968 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _043_
timestamp 1618914159
transform 1 0 5244 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1618914159
transform 1 0 3404 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _105_
timestamp 1618914159
transform 1 0 4692 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1618914159
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1618914159
transform -1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform -1 0 6624 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1618914159
transform 1 0 6164 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _082_
timestamp 1618914159
transform 1 0 5336 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _040_
timestamp 1618914159
transform 1 0 6256 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output22
timestamp 1618914159
transform 1 0 6532 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _079_
timestamp 1618914159
transform 1 0 6900 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _098_
timestamp 1618914159
transform 1 0 6624 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _086_
timestamp 1618914159
transform 1 0 6532 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_11_81
timestamp 1618914159
transform 1 0 8372 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output21
timestamp 1618914159
transform 1 0 8464 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output20
timestamp 1618914159
transform 1 0 8464 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output19
timestamp 1618914159
transform 1 0 9200 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1618914159
transform 1 0 8832 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1618914159
transform 1 0 8832 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1618914159
transform -1 0 9844 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1618914159
transform -1 0 9844 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1618914159
transform -1 0 9844 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_2  _075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 8924 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _052_
timestamp 1618914159
transform 1 0 8924 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _087_
timestamp 1618914159
transform 1 0 7728 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1618914159
transform 1 0 920 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1618914159
transform 1 0 920 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1618914159
transform 1 0 1196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1618914159
transform 1 0 2300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1618914159
transform 1 0 1196 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1618914159
transform 1 0 2300 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1618914159
transform 1 0 3588 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_27
timestamp 1618914159
transform 1 0 3404 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_39
timestamp 1618914159
transform 1 0 4508 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_47
timestamp 1618914159
transform 1 0 5244 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_27
timestamp 1618914159
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_30
timestamp 1618914159
transform 1 0 3680 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_42
timestamp 1618914159
transform 1 0 4784 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_56
timestamp 1618914159
transform 1 0 6072 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_50
timestamp 1618914159
transform 1 0 5520 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1618914159
transform 1 0 6256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1618914159
transform 1 0 5796 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1618914159
transform 1 0 6164 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _067_
timestamp 1618914159
transform 1 0 5336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp 1618914159
transform 1 0 5612 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _053_
timestamp 1618914159
transform 1 0 5888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _039_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 6992 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _097_
timestamp 1618914159
transform 1 0 6440 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _084_
timestamp 1618914159
transform 1 0 7452 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp 1618914159
transform 1 0 9292 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618914159
transform 1 0 8924 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1618914159
transform -1 0 9844 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1618914159
transform -1 0 9844 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1618914159
transform 1 0 8832 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output25
timestamp 1618914159
transform 1 0 8464 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_92
timestamp 1618914159
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_80
timestamp 1618914159
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1618914159
transform 1 0 920 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1618914159
transform 1 0 1196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1618914159
transform 1 0 2300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1618914159
transform 1 0 3588 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1618914159
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1618914159
transform 1 0 3680 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_42
timestamp 1618914159
transform 1 0 4784 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_48
timestamp 1618914159
transform 1 0 5336 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  output24
timestamp 1618914159
transform 1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1618914159
transform 1 0 5704 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _077_
timestamp 1618914159
transform 1 0 5980 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1618914159
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1618914159
transform 1 0 6348 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1618914159
transform 1 0 6256 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_64
timestamp 1618914159
transform 1 0 6808 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output26
timestamp 1618914159
transform 1 0 6900 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1618914159
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1618914159
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _069_
timestamp 1618914159
transform 1 0 8648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1618914159
transform -1 0 9844 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1618914159
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1618914159
transform 1 0 7636 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output23
timestamp 1618914159
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1618914159
transform 1 0 7912 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_88
timestamp 1618914159
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
<< labels >>
rlabel metal3 s 14000 1096 34000 1216 6 mgmt_gpio_in
port 0 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 1 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 2 nsew signal input
rlabel metal3 s 14000 552 34000 672 6 one
port 3 nsew signal tristate
rlabel metal3 s 14000 2592 34000 2712 6 pad_gpio_ana_en
port 4 nsew signal tristate
rlabel metal3 s 14000 3136 34000 3256 6 pad_gpio_ana_pol
port 5 nsew signal tristate
rlabel metal3 s 14000 3544 34000 3664 6 pad_gpio_ana_sel
port 6 nsew signal tristate
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[0]
port 7 nsew signal tristate
rlabel metal3 s 14000 4632 34000 4752 6 pad_gpio_dm[1]
port 8 nsew signal tristate
rlabel metal3 s 14000 5040 34000 5160 6 pad_gpio_dm[2]
port 9 nsew signal tristate
rlabel metal3 s 14000 5584 34000 5704 6 pad_gpio_holdover
port 10 nsew signal tristate
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_ib_mode_sel
port 11 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_in
port 12 nsew signal input
rlabel metal3 s 14000 7080 34000 7200 6 pad_gpio_inenb
port 13 nsew signal tristate
rlabel metal3 s 14000 7624 34000 7744 6 pad_gpio_out
port 14 nsew signal tristate
rlabel metal3 s 14000 8032 34000 8152 6 pad_gpio_outenb
port 15 nsew signal tristate
rlabel metal3 s 14000 8576 34000 8696 6 pad_gpio_slow_sel
port 16 nsew signal tristate
rlabel metal3 s 14000 9120 34000 9240 6 pad_gpio_vtrip_sel
port 17 nsew signal tristate
rlabel metal3 s 14000 9528 34000 9648 6 resetn
port 18 nsew signal input
rlabel metal3 s 14000 10072 34000 10192 6 resetn_out
port 19 nsew signal tristate
rlabel metal3 s 14000 10616 34000 10736 6 serial_clock
port 20 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_clock_out
port 21 nsew signal tristate
rlabel metal3 s 14000 11568 34000 11688 6 serial_data_in
port 22 nsew signal input
rlabel metal3 s 14000 12112 34000 12232 6 serial_data_out
port 23 nsew signal tristate
rlabel metal3 s 14000 12520 34000 12640 6 user_gpio_in
port 24 nsew signal tristate
rlabel metal3 s 14000 13064 34000 13184 6 user_gpio_oeb
port 25 nsew signal input
rlabel metal3 s 14000 13608 34000 13728 6 user_gpio_out
port 26 nsew signal input
rlabel metal3 s 14000 144 34000 264 6 zero
port 27 nsew signal tristate
rlabel metal4 s 7660 956 7980 12644 6 vccd
port 28 nsew power bidirectional
rlabel metal4 s 4460 956 4780 12644 6 vccd
port 29 nsew power bidirectional
rlabel metal4 s 1260 4432 1580 12644 6 vccd
port 30 nsew power bidirectional
rlabel metal4 s 10084 1616 10404 11984 6 vccd
port 31 nsew power bidirectional
rlabel metal4 s 360 1616 680 11984 6 vccd
port 32 nsew power bidirectional
rlabel metal4 s 1260 956 1580 2128 6 vccd
port 33 nsew power bidirectional
rlabel metal5 s 360 11664 10404 11984 6 vccd
port 34 nsew power bidirectional
rlabel metal5 s -300 8916 11064 9236 6 vccd
port 35 nsew power bidirectional
rlabel metal5 s -300 5716 11064 6036 6 vccd
port 36 nsew power bidirectional
rlabel metal5 s -300 2516 11064 2836 6 vccd
port 37 nsew power bidirectional
rlabel metal5 s 360 1616 10404 1936 6 vccd
port 38 nsew power bidirectional
rlabel metal4 s 10744 956 11064 12644 6 vssd
port 39 nsew ground bidirectional
rlabel metal4 s 9260 956 9580 12644 6 vssd
port 40 nsew ground bidirectional
rlabel metal4 s 6060 956 6380 12644 6 vssd
port 41 nsew ground bidirectional
rlabel metal4 s 2860 4432 3180 12644 6 vssd
port 42 nsew ground bidirectional
rlabel metal4 s -300 956 20 12644 4 vssd
port 43 nsew ground bidirectional
rlabel metal4 s 2860 956 3180 2128 6 vssd
port 44 nsew ground bidirectional
rlabel metal5 s -300 12324 11064 12644 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s -300 10516 11064 10836 6 vssd
port 46 nsew ground bidirectional
rlabel metal5 s -300 7316 11064 7636 6 vssd
port 47 nsew ground bidirectional
rlabel metal5 s -300 4116 11064 4436 6 vssd
port 48 nsew ground bidirectional
rlabel metal5 s -300 956 11064 1276 6 vssd
port 49 nsew ground bidirectional
rlabel metal4 s 8560 -364 8880 13964 6 vccd1
port 50 nsew power bidirectional
rlabel metal4 s 5360 -364 5680 13964 6 vccd1
port 51 nsew power bidirectional
rlabel metal4 s 2160 4480 2480 13964 6 vccd1
port 52 nsew power bidirectional
rlabel metal4 s 11404 296 11724 13304 6 vccd1
port 53 nsew power bidirectional
rlabel metal4 s -960 296 -640 13304 4 vccd1
port 54 nsew power bidirectional
rlabel metal4 s 2160 -364 2480 2080 6 vccd1
port 55 nsew power bidirectional
rlabel metal5 s -960 12984 11724 13304 6 vccd1
port 56 nsew power bidirectional
rlabel metal5 s -1620 9816 12384 10136 6 vccd1
port 57 nsew power bidirectional
rlabel metal5 s -1620 6616 12384 6936 6 vccd1
port 58 nsew power bidirectional
rlabel metal5 s -1620 3416 12384 3736 6 vccd1
port 59 nsew power bidirectional
rlabel metal5 s -960 296 11724 616 6 vccd1
port 60 nsew power bidirectional
rlabel metal4 s 12064 -364 12384 13964 6 vssd1
port 61 nsew ground bidirectional
rlabel metal4 s 6960 -364 7280 13964 6 vssd1
port 62 nsew ground bidirectional
rlabel metal4 s 3760 -364 4080 13964 6 vssd1
port 63 nsew ground bidirectional
rlabel metal4 s -1620 -364 -1300 13964 4 vssd1
port 64 nsew ground bidirectional
rlabel metal5 s -1620 13644 12384 13964 6 vssd1
port 65 nsew ground bidirectional
rlabel metal5 s -1620 8216 12384 8536 6 vssd1
port 66 nsew ground bidirectional
rlabel metal5 s -1620 5016 12384 5336 6 vssd1
port 67 nsew ground bidirectional
rlabel metal5 s -1620 -364 12384 -44 8 vssd1
port 68 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 34000 14000
<< end >>
