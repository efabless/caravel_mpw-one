magic
tech sky130A
magscale 1 2
timestamp 1603424375
<< metal1 >>
rect 85286 1020000 85338 1020260
rect 133486 1020000 133538 1020260
rect 181486 1020000 181538 1020260
rect 229686 1020000 229738 1020260
rect 277686 1020000 277738 1020260
rect 372886 1020000 372938 1020260
rect 421086 1020000 421138 1020260
rect 469086 1020000 469138 1020260
rect 564286 1020000 564338 1020260
rect 39739 986886 39999 986938
rect 600000 974862 600260 974914
rect 600000 880662 600260 880714
rect 39739 807686 39999 807738
rect 600000 786462 600260 786514
rect 39739 762086 39999 762138
rect 600000 738862 600260 738914
rect 39739 716486 39999 716538
rect 600000 691262 600260 691314
rect 39739 670886 39999 670938
rect 600000 643462 600260 643514
rect 39739 625486 39999 625538
rect 600000 595862 600260 595914
rect 39739 579886 39999 579938
rect 600000 548262 600260 548314
rect 39739 534286 39999 534338
rect 39739 399686 39999 399738
rect 600000 360862 600260 360914
rect 39739 354086 39999 354138
rect 600000 313062 600260 313114
rect 39739 308486 39999 308538
rect 600000 265462 600260 265514
rect 39739 262886 39999 262938
rect 600000 217862 600260 217914
rect 39739 217486 39999 217538
rect 39739 171886 39999 171938
rect 600000 170262 600260 170314
rect 600000 122662 600260 122714
rect 600000 75062 600260 75114
<< metal2 >>
rect 73475 1020000 73521 1020894
rect 73884 1020000 73930 1020894
rect 74026 1020000 74078 1020310
rect 77271 1020000 77323 1021284
rect 78120 1020000 78172 1020540
rect 78498 1020000 78550 1020814
rect 78950 1020000 79002 1020452
rect 79163 1020000 79215 1020668
rect 79892 1020000 79944 1020310
rect 81849 1020000 81901 1021018
rect 82771 1020000 82823 1020108
rect 86167 1020000 86219 1020238
rect 88322 1020000 88374 1020236
rect 121675 1020000 121721 1020894
rect 122084 1020000 122130 1020894
rect 122226 1020000 122278 1020310
rect 125471 1020000 125523 1021284
rect 126320 1020000 126372 1020540
rect 126698 1020000 126750 1020814
rect 127150 1020000 127202 1020452
rect 127363 1020000 127415 1020668
rect 128092 1020000 128144 1020310
rect 130049 1020000 130101 1021018
rect 130971 1020000 131023 1020108
rect 134367 1020000 134419 1020238
rect 136522 1020000 136574 1020236
rect 169675 1020000 169721 1020894
rect 170084 1020000 170130 1020894
rect 170226 1020000 170278 1020310
rect 173471 1020000 173523 1021284
rect 174320 1020000 174372 1020540
rect 174698 1020000 174750 1020814
rect 175150 1020000 175202 1020452
rect 175363 1020000 175415 1020668
rect 176092 1020000 176144 1020310
rect 178049 1020000 178101 1021018
rect 178971 1020000 179023 1020108
rect 182367 1020000 182419 1020238
rect 184522 1020000 184574 1020236
rect 217875 1020000 217921 1020894
rect 218284 1020000 218330 1020894
rect 218426 1020000 218478 1020310
rect 221671 1020000 221723 1021284
rect 222520 1020000 222572 1020540
rect 222898 1020000 222950 1020814
rect 223350 1020000 223402 1020452
rect 223563 1020000 223615 1020668
rect 224292 1020000 224344 1020310
rect 226249 1020000 226301 1021018
rect 227171 1020000 227223 1020108
rect 230567 1020000 230619 1020238
rect 232722 1020000 232774 1020236
rect 265875 1020000 265921 1020894
rect 266284 1020000 266330 1020894
rect 266426 1020000 266478 1020310
rect 269671 1020000 269723 1021284
rect 270520 1020000 270572 1020540
rect 270898 1020000 270950 1020814
rect 271350 1020000 271402 1020452
rect 271563 1020000 271615 1020668
rect 272292 1020000 272344 1020310
rect 274249 1020000 274301 1021018
rect 275171 1020000 275223 1020108
rect 278567 1020000 278619 1020238
rect 280722 1020000 280774 1020236
rect 361075 1020000 361121 1020894
rect 361484 1020000 361530 1020894
rect 361626 1020000 361678 1020310
rect 364871 1020000 364923 1021284
rect 365720 1020000 365772 1020540
rect 366098 1020000 366150 1020814
rect 366550 1020000 366602 1020452
rect 366763 1020000 366815 1020668
rect 367492 1020000 367544 1020310
rect 369449 1020000 369501 1021018
rect 370371 1020000 370423 1020108
rect 373767 1020000 373819 1020238
rect 375922 1020000 375974 1020236
rect 409275 1020000 409321 1020894
rect 409684 1020000 409730 1020894
rect 409826 1020000 409878 1020310
rect 413071 1020000 413123 1021284
rect 413920 1020000 413972 1020540
rect 414298 1020000 414350 1020814
rect 414750 1020000 414802 1020452
rect 414963 1020000 415015 1020668
rect 415692 1020000 415744 1020310
rect 417649 1020000 417701 1021018
rect 418571 1020000 418623 1020108
rect 421967 1020000 422019 1020238
rect 424122 1020000 424174 1020236
rect 457275 1020000 457321 1020894
rect 457684 1020000 457730 1020894
rect 457826 1020000 457878 1020310
rect 461071 1020000 461123 1021284
rect 461920 1020000 461972 1020540
rect 462298 1020000 462350 1020814
rect 462750 1020000 462802 1020452
rect 462963 1020000 463015 1020668
rect 463692 1020000 463744 1020310
rect 465649 1020000 465701 1021018
rect 466571 1020000 466623 1020108
rect 469967 1020000 470019 1020238
rect 472122 1020000 472174 1020236
rect 552475 1020000 552521 1020894
rect 552884 1020000 552930 1020894
rect 553026 1020000 553078 1020310
rect 556271 1020000 556323 1021284
rect 557120 1020000 557172 1020540
rect 557498 1020000 557550 1020814
rect 557950 1020000 558002 1020452
rect 558163 1020000 558215 1020668
rect 558892 1020000 558944 1020310
rect 560849 1020000 560901 1021018
rect 561771 1020000 561823 1020108
rect 565167 1020000 565219 1020238
rect 567322 1020000 567374 1020236
rect 39763 989922 39999 989974
rect 39761 987767 39999 987819
rect 600000 986679 600894 986725
rect 600000 986270 600894 986316
rect 600000 986122 600310 986174
rect 39891 984371 39999 984423
rect 38982 983449 40000 983501
rect 600000 982877 601284 982929
rect 600000 982028 600540 982080
rect 600000 981650 600814 981702
rect 39690 981492 40000 981544
rect 600000 981198 600452 981250
rect 600000 980985 600668 981037
rect 39332 980763 40000 980815
rect 39547 980550 39999 980602
rect 600000 980256 600310 980308
rect 39186 980098 40000 980150
rect 39459 979720 39999 979772
rect 38715 978871 39999 978923
rect 600000 978299 601018 978351
rect 600000 977377 600108 977429
rect 39690 975626 40000 975678
rect 39105 975484 39999 975530
rect 39105 975075 39999 975121
rect 600000 973981 600238 974033
rect 600000 971826 600236 971878
rect 600000 892479 600894 892525
rect 600000 892070 600894 892116
rect 600000 891922 600310 891974
rect 600000 888677 601284 888729
rect 600000 887828 600540 887880
rect 600000 887450 600814 887502
rect 600000 886998 600452 887050
rect 600000 886785 600668 886837
rect 600000 886056 600310 886108
rect 600000 884099 601018 884151
rect 600000 883177 600108 883229
rect 600000 879781 600238 879833
rect 600000 877626 600236 877678
rect 39763 810722 39999 810774
rect 39761 808567 39999 808619
rect 39891 805171 39999 805223
rect 38982 804249 40000 804301
rect 39690 802292 40000 802344
rect 39332 801563 40000 801615
rect 39547 801350 39999 801402
rect 39186 800898 40000 800950
rect 39459 800520 39999 800572
rect 38715 799671 39999 799723
rect 600000 798279 600894 798325
rect 600000 797870 600894 797916
rect 600000 797722 600310 797774
rect 39690 796426 40000 796478
rect 39105 796284 39999 796330
rect 39105 795875 39999 795921
rect 600000 794477 601284 794529
rect 600000 793628 600540 793680
rect 600000 793250 600814 793302
rect 600000 792798 600452 792850
rect 600000 792585 600668 792637
rect 600000 791856 600310 791908
rect 600000 789899 601018 789951
rect 600000 788977 600108 789029
rect 600000 785581 600238 785633
rect 600000 783426 600236 783478
rect 39763 765122 39999 765174
rect 39761 762967 39999 763019
rect 39891 759571 39999 759623
rect 38982 758649 40000 758701
rect 39690 756692 40000 756744
rect 39332 755963 40000 756015
rect 39547 755750 39999 755802
rect 39186 755298 40000 755350
rect 39459 754920 39999 754972
rect 38715 754071 39999 754123
rect 39690 750826 40000 750878
rect 39105 750684 39999 750730
rect 600000 750679 600894 750725
rect 39105 750275 39999 750321
rect 600000 750270 600894 750316
rect 600000 750122 600310 750174
rect 600000 746877 601284 746929
rect 600000 746028 600540 746080
rect 600000 745650 600814 745702
rect 600000 745198 600452 745250
rect 600000 744985 600668 745037
rect 600000 744256 600310 744308
rect 600000 742299 601018 742351
rect 600000 741377 600108 741429
rect 600000 737981 600238 738033
rect 600000 735826 600236 735878
rect 39763 719522 39999 719574
rect 39761 717367 39999 717419
rect 39891 713971 39999 714023
rect 38982 713049 40000 713101
rect 39690 711092 40000 711144
rect 39332 710363 40000 710415
rect 39547 710150 39999 710202
rect 39186 709698 40000 709750
rect 39459 709320 39999 709372
rect 38715 708471 39999 708523
rect 39690 705226 40000 705278
rect 39105 705084 39999 705130
rect 39105 704675 39999 704721
rect 600000 703079 600894 703125
rect 600000 702670 600894 702716
rect 600000 702522 600310 702574
rect 600000 699277 601284 699329
rect 600000 698428 600540 698480
rect 600000 698050 600814 698102
rect 600000 697598 600452 697650
rect 600000 697385 600668 697437
rect 600000 696656 600310 696708
rect 600000 694699 601018 694751
rect 600000 693777 600108 693829
rect 600000 690381 600238 690433
rect 600000 688226 600236 688278
rect 39763 673922 39999 673974
rect 39761 671767 39999 671819
rect 39891 668371 39999 668423
rect 38982 667449 40000 667501
rect 39690 665492 40000 665544
rect 39332 664763 40000 664815
rect 39547 664550 39999 664602
rect 39186 664098 40000 664150
rect 39459 663720 39999 663772
rect 38715 662871 39999 662923
rect 39690 659626 40000 659678
rect 39105 659484 39999 659530
rect 39105 659075 39999 659121
rect 600000 655279 600894 655325
rect 600000 654870 600894 654916
rect 600000 654722 600310 654774
rect 600000 651477 601284 651529
rect 600000 650628 600540 650680
rect 600000 650250 600814 650302
rect 600000 649798 600452 649850
rect 600000 649585 600668 649637
rect 600000 648856 600310 648908
rect 600000 646899 601018 646951
rect 600000 645977 600108 646029
rect 600000 642581 600238 642633
rect 600000 640426 600236 640478
rect 39763 628522 39999 628574
rect 39761 626367 39999 626419
rect 39891 622971 39999 623023
rect 38982 622049 40000 622101
rect 39690 620092 40000 620144
rect 39332 619363 40000 619415
rect 39547 619150 39999 619202
rect 39186 618698 40000 618750
rect 39459 618320 39999 618372
rect 38715 617471 39999 617523
rect 39690 614226 40000 614278
rect 39105 614084 39999 614130
rect 39105 613675 39999 613721
rect 600000 607679 600894 607725
rect 600000 607270 600894 607316
rect 600000 607122 600310 607174
rect 600000 603877 601284 603929
rect 600000 603028 600540 603080
rect 600000 602650 600814 602702
rect 600000 602198 600452 602250
rect 600000 601985 600668 602037
rect 600000 601256 600310 601308
rect 600000 599299 601018 599351
rect 600000 598377 600108 598429
rect 600000 594981 600238 595033
rect 600000 592826 600236 592878
rect 39763 582922 39999 582974
rect 39761 580767 39999 580819
rect 39891 577371 39999 577423
rect 38982 576449 40000 576501
rect 39690 574492 40000 574544
rect 39332 573763 40000 573815
rect 39547 573550 39999 573602
rect 39186 573098 40000 573150
rect 39459 572720 39999 572772
rect 38715 571871 39999 571923
rect 39690 568626 40000 568678
rect 39105 568484 39999 568530
rect 39105 568075 39999 568121
rect 600000 560079 600894 560125
rect 600000 559670 600894 559716
rect 600000 559522 600310 559574
rect 600000 556277 601284 556329
rect 600000 555428 600540 555480
rect 600000 555050 600814 555102
rect 600000 554598 600452 554650
rect 600000 554385 600668 554437
rect 600000 553656 600310 553708
rect 600000 551699 601018 551751
rect 600000 550777 600108 550829
rect 600000 547381 600238 547433
rect 600000 545226 600236 545278
rect 39763 537322 39999 537374
rect 39761 535167 39999 535219
rect 39891 531771 39999 531823
rect 38982 530849 40000 530901
rect 39690 528892 40000 528944
rect 39332 528163 40000 528215
rect 39547 527950 39999 528002
rect 39186 527498 40000 527550
rect 39459 527120 39999 527172
rect 38715 526271 39999 526323
rect 39690 523026 40000 523078
rect 39105 522884 39999 522930
rect 39105 522475 39999 522521
rect 39763 402722 39999 402774
rect 39761 400567 39999 400619
rect 39891 397171 39999 397223
rect 38982 396249 40000 396301
rect 39690 394292 40000 394344
rect 39332 393563 40000 393615
rect 39547 393350 39999 393402
rect 39186 392898 40000 392950
rect 39459 392520 39999 392572
rect 38715 391671 39999 391723
rect 39690 388426 40000 388478
rect 39105 388284 39999 388330
rect 39105 387875 39999 387921
rect 600000 372679 600894 372725
rect 600000 372270 600894 372316
rect 600000 372122 600310 372174
rect 600000 368877 601284 368929
rect 600000 368028 600540 368080
rect 600000 367650 600814 367702
rect 600000 367198 600452 367250
rect 600000 366985 600668 367037
rect 600000 366256 600310 366308
rect 600000 364299 601018 364351
rect 600000 363377 600108 363429
rect 600000 359981 600238 360033
rect 600000 357826 600236 357878
rect 39763 357122 39999 357174
rect 39761 354967 39999 355019
rect 39891 351571 39999 351623
rect 38982 350649 40000 350701
rect 39690 348692 40000 348744
rect 39332 347963 40000 348015
rect 39547 347750 39999 347802
rect 39186 347298 40000 347350
rect 39459 346920 39999 346972
rect 38715 346071 39999 346123
rect 39690 342826 40000 342878
rect 39105 342684 39999 342730
rect 39105 342275 39999 342321
rect 600000 324879 600894 324925
rect 600000 324470 600894 324516
rect 600000 324322 600310 324374
rect 600000 321077 601284 321129
rect 600000 320228 600540 320280
rect 600000 319850 600814 319902
rect 600000 319398 600452 319450
rect 600000 319185 600668 319237
rect 600000 318456 600310 318508
rect 600000 316499 601018 316551
rect 600000 315577 600108 315629
rect 600000 312181 600238 312233
rect 39763 311522 39999 311574
rect 600000 310026 600236 310078
rect 39761 309367 39999 309419
rect 39891 305971 39999 306023
rect 38982 305049 40000 305101
rect 39690 303092 40000 303144
rect 39332 302363 40000 302415
rect 39547 302150 39999 302202
rect 39186 301698 40000 301750
rect 39459 301320 39999 301372
rect 38715 300471 39999 300523
rect 39690 297226 40000 297278
rect 39105 297084 39999 297130
rect 39105 296675 39999 296721
rect 600000 277279 600894 277325
rect 600000 276870 600894 276916
rect 600000 276722 600310 276774
rect 600000 273477 601284 273529
rect 600000 272628 600540 272680
rect 600000 272250 600814 272302
rect 600000 271798 600452 271850
rect 600000 271585 600668 271637
rect 600000 270856 600310 270908
rect 600000 268899 601018 268951
rect 600000 267977 600108 268029
rect 39763 265922 39999 265974
rect 600000 264581 600238 264633
rect 39761 263767 39999 263819
rect 600000 262426 600236 262478
rect 39891 260371 39999 260423
rect 38982 259449 40000 259501
rect 39690 257492 40000 257544
rect 39332 256763 40000 256815
rect 39547 256550 39999 256602
rect 39186 256098 40000 256150
rect 39459 255720 39999 255772
rect 38715 254871 39999 254923
rect 39690 251626 40000 251678
rect 39105 251484 39999 251530
rect 39105 251075 39999 251121
rect 600000 229679 600894 229725
rect 600000 229270 600894 229316
rect 600000 229122 600310 229174
rect 600000 225877 601284 225929
rect 600000 225028 600540 225080
rect 600000 224650 600814 224702
rect 600000 224198 600452 224250
rect 600000 223985 600668 224037
rect 600000 223256 600310 223308
rect 600000 221299 601018 221351
rect 39763 220522 39999 220574
rect 600000 220377 600108 220429
rect 39761 218367 39999 218419
rect 600000 216981 600238 217033
rect 39891 214971 39999 215023
rect 600000 214826 600236 214878
rect 38982 214049 40000 214101
rect 39690 212092 40000 212144
rect 39332 211363 40000 211415
rect 39547 211150 39999 211202
rect 39186 210698 40000 210750
rect 39459 210320 39999 210372
rect 38715 209471 39999 209523
rect 39690 206226 40000 206278
rect 39105 206084 39999 206130
rect 39105 205675 39999 205721
rect 600000 182079 600894 182125
rect 600000 181670 600894 181716
rect 600000 181522 600310 181574
rect 600000 178277 601284 178329
rect 600000 177428 600540 177480
rect 600000 177050 600814 177102
rect 600000 176598 600452 176650
rect 600000 176385 600668 176437
rect 600000 175656 600310 175708
rect 39763 174922 39999 174974
rect 600000 173699 601018 173751
rect 39761 172767 39999 172819
rect 600000 172777 600108 172829
rect 39891 169371 39999 169423
rect 600000 169381 600238 169433
rect 38982 168449 40000 168501
rect 600000 167226 600236 167278
rect 39690 166492 40000 166544
rect 39332 165763 40000 165815
rect 39547 165550 39999 165602
rect 39186 165098 40000 165150
rect 39459 164720 39999 164772
rect 38715 163871 39999 163923
rect 39690 160626 40000 160678
rect 39105 160484 39999 160530
rect 39105 160075 39999 160121
rect 600000 134479 600894 134525
rect 600000 134070 600894 134116
rect 600000 133922 600310 133974
rect 600000 130677 601284 130729
rect 600000 129828 600540 129880
rect 600000 129450 600814 129502
rect 600000 128998 600452 129050
rect 600000 128785 600668 128837
rect 600000 128056 600310 128108
rect 600000 126099 601018 126151
rect 600000 125177 600108 125229
rect 600000 121781 600238 121833
rect 600000 119626 600236 119678
rect 600000 86879 600894 86925
rect 600000 86470 600894 86516
rect 600000 86322 600310 86374
rect 600000 83077 601284 83129
rect 600000 82228 600540 82280
rect 600000 81850 600814 81902
rect 600000 81398 600452 81450
rect 600000 81185 600668 81237
rect 600000 80456 600310 80508
rect 600000 78499 601018 78551
rect 600000 77577 600108 77629
rect 600000 74181 600238 74233
rect 600000 72026 600236 72078
rect 132091 39706 132143 40000
rect 173899 38982 173951 40000
rect 269499 38982 269551 40000
rect 274077 38715 274129 39999
rect 277879 39105 277925 39999
rect 317899 38982 317951 40000
rect 322477 38715 322529 39999
rect 326279 39105 326325 39999
rect 366299 38982 366351 40000
rect 370877 38715 370929 39999
rect 374679 39105 374725 39999
rect 414699 38982 414751 40000
rect 419277 38715 419329 39999
rect 423079 39105 423125 39999
rect 461977 39891 462029 39999
rect 462899 38982 462951 40000
rect 466250 39186 466302 40000
rect 467477 38715 467529 39999
rect 471279 39105 471325 39999
<< metal3 >>
rect 81973 1020000 82039 1027360
rect 88648 1020000 88714 1057912
rect 130173 1020000 130239 1027360
rect 136848 1020000 136914 1057912
rect 178173 1020000 178239 1027360
rect 184848 1020000 184914 1057912
rect 226373 1020000 226439 1027360
rect 233048 1020000 233114 1057912
rect 274373 1020000 274439 1027360
rect 281048 1020000 281114 1057912
rect 369573 1020000 369639 1027360
rect 376248 1020000 376314 1057912
rect 417773 1020000 417839 1027360
rect 424448 1020000 424514 1057912
rect 465773 1020000 465839 1027360
rect 472448 1020000 472514 1057912
rect 560973 1020000 561039 1027360
rect 567648 1020000 567714 1057912
rect 2088 990248 40000 990314
rect 32639 983573 39999 983639
rect 600000 978161 607360 978227
rect 600000 971486 637912 971552
rect 600000 883961 607360 884027
rect 600000 877286 637912 877352
rect 2088 811048 40000 811114
rect 32639 804373 39999 804439
rect 600000 789761 607360 789827
rect 600000 783086 637912 783152
rect 2088 765448 40000 765514
rect 32639 758773 39999 758839
rect 600000 742161 607360 742227
rect 600000 735486 637912 735552
rect 2088 719848 40000 719914
rect 32639 713173 39999 713239
rect 600000 694561 607360 694627
rect 600000 687886 637912 687952
rect 2088 674248 40000 674314
rect 32639 667573 39999 667639
rect 600000 646761 607360 646827
rect 600000 640086 637912 640152
rect 2088 628848 40000 628914
rect 32639 622173 39999 622239
rect 600000 599161 607360 599227
rect 600000 592486 637912 592552
rect 2088 583248 40000 583314
rect 32639 576573 39999 576639
rect 600000 551561 607360 551627
rect 600000 544886 637912 544952
rect 2088 537648 40000 537714
rect 32639 530973 39999 531039
rect 2088 403048 40000 403114
rect 32639 396373 39999 396439
rect 600000 364161 607360 364227
rect 2088 357448 40000 357514
rect 600000 357486 637912 357552
rect 32639 350773 39999 350839
rect 600000 316361 607360 316427
rect 2088 311848 40000 311914
rect 600000 309686 637912 309752
rect 32639 305173 39999 305239
rect 600000 268761 607360 268827
rect 2088 266248 40000 266314
rect 600000 262086 637912 262152
rect 32639 259573 39999 259639
rect 600000 221161 607360 221227
rect 2088 220848 40000 220914
rect 600000 214486 637912 214552
rect 32639 214173 39999 214239
rect 2088 175248 40000 175314
rect 600000 173561 607360 173627
rect 32639 168573 39999 168639
rect 600000 166886 637912 166952
rect 600000 125961 607360 126027
rect 600000 119286 637912 119352
rect 600000 78361 607360 78427
rect 600000 71686 637912 71752
rect 128667 38031 128813 39999
rect 167086 2088 167152 40000
rect 359486 2088 359552 40000
rect 407886 2088 407952 40000
rect 456086 2088 456152 40000
<< metal5 >>
rect 75040 1040912 87560 1053402
rect 123240 1040912 135760 1053402
rect 171240 1040912 183760 1053402
rect 219440 1040912 231960 1053402
rect 267440 1040912 279960 1053402
rect 314620 1040802 327160 1053324
rect 362640 1040912 375160 1053402
rect 410840 1040912 423360 1053402
rect 458840 1040912 471360 1053402
rect 506020 1040802 518560 1053324
rect 554040 1040912 566560 1053402
rect 6598 976640 19088 989160
rect 620912 972640 633402 985160
rect 6086 931663 19572 942991
rect 620428 926609 633914 937937
rect 620912 878440 633402 890960
rect 6675 841820 19197 854360
rect 620802 831840 633324 844380
rect 6598 797440 19088 809960
rect 620912 784240 633402 796760
rect 6598 751840 19088 764360
rect 620912 736640 633402 749160
rect 6598 706240 19088 718760
rect 620912 689040 633402 701560
rect 6598 660640 19088 673160
rect 620912 641240 633402 653760
rect 6598 615240 19088 627760
rect 620912 593640 633402 606160
rect 6598 569640 19088 582160
rect 620912 546040 633402 558560
rect 6598 524040 19088 536560
rect 6675 478420 19197 490960
rect 620428 453409 633914 464737
rect 6086 434463 19572 445791
rect 6598 389440 19088 401960
rect 620912 358640 633402 371160
rect 6598 343840 19088 356360
rect 620912 310840 633402 323360
rect 6598 298240 19088 310760
rect 6598 252640 19088 265160
rect 620912 263240 633402 275760
rect 6598 207240 19088 219760
rect 620912 215640 633402 228160
rect 6598 161640 19088 174160
rect 620912 168040 633402 180560
rect 6675 116020 19197 128560
rect 620912 120440 633402 132960
rect 6086 72063 19572 83391
rect 620912 72840 633402 85360
rect 73440 6675 85980 19197
rect 120840 6675 133380 19197
rect 168240 6598 180760 19088
rect 217209 6086 228537 19572
rect 263840 6598 276360 19088
rect 312240 6598 324760 19088
rect 360640 6598 373160 19088
rect 409040 6598 421560 19088
rect 457240 6598 469760 19088
rect 553040 6675 565580 19197
use sky130_ef_io__corner_pad  mgmt_corner\[0\] /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_118 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_246
timestamp 1603391777
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  mgmt_vssa_hvclamp_pad /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform -1 0 87200 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_119
timestamp 1603391777
transform -1 0 48000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_120
timestamp 1603391777
transform -1 0 52000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_121
timestamp 1603391777
transform -1 0 56000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_122
timestamp 1603391777
transform -1 0 60000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_123
timestamp 1603391777
transform -1 0 64000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_124
timestamp 1603391777
transform -1 0 68000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1603391777
transform -1 0 72000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_126 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform -1 0 72200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_130
timestamp 1603391777
transform -1 0 99200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_129
timestamp 1603391777
transform -1 0 95200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_128
timestamp 1603391777
transform -1 0 91200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_134
timestamp 1603391777
transform -1 0 115200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_133
timestamp 1603391777
transform -1 0 111200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_132
timestamp 1603391777
transform -1 0 107200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1603391777
transform -1 0 103200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_137
timestamp 1603391777
transform -1 0 119600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_136
timestamp 1603391777
transform -1 0 119400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_135
timestamp 1603391777
transform -1 0 119200 0 -1 39593
box 0 0 4000 39593
use sky130_fd_io__top_xres4v2  resetb_pad /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1603391773
transform -1 0 134600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_139
timestamp 1603391777
transform -1 0 138600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_140
timestamp 1603391777
transform -1 0 142600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_141
timestamp 1603391777
transform -1 0 146600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_142
timestamp 1603391777
transform -1 0 150600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_143
timestamp 1603391777
transform -1 0 154600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_144
timestamp 1603391777
transform -1 0 158600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_145
timestamp 1603391777
transform -1 0 162600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_146
timestamp 1603391777
transform -1 0 166600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  clock_pad /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform -1 0 183000 0 -1 39593
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_147
timestamp 1603391777
transform -1 0 166800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_148
timestamp 1603391777
transform -1 0 167000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_150
timestamp 1603391777
transform -1 0 187000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_151
timestamp 1603391777
transform -1 0 191000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_152
timestamp 1603391777
transform -1 0 195000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_153
timestamp 1603391777
transform -1 0 199000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_154
timestamp 1603391777
transform -1 0 203000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_155
timestamp 1603391777
transform -1 0 207000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_pad  mgmt_vssd_lvclmap_pad /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform -1 0 230400 0 -1 39593
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_156
timestamp 1603391777
transform -1 0 211000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_157
timestamp 1603391777
transform -1 0 215000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_158
timestamp 1603391777
transform -1 0 215200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_159
timestamp 1603391777
transform -1 0 215400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_161
timestamp 1603391777
transform -1 0 234400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_162
timestamp 1603391777
transform -1 0 238400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_163
timestamp 1603391777
transform -1 0 242400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_164
timestamp 1603391777
transform -1 0 246400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  flash_csb_pad
timestamp 1603391777
transform -1 0 278600 0 -1 39593
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_165
timestamp 1603391777
transform -1 0 250400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_166
timestamp 1603391777
transform -1 0 254400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_167
timestamp 1603391777
transform -1 0 258400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_168
timestamp 1603391777
transform -1 0 262400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_169
timestamp 1603391777
transform -1 0 262600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_171
timestamp 1603391777
transform -1 0 282600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_172
timestamp 1603391777
transform -1 0 286600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  flash_clk_pad
timestamp 1603391777
transform -1 0 327000 0 -1 39593
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_173
timestamp 1603391777
transform -1 0 290600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_174
timestamp 1603391777
transform -1 0 294600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_175
timestamp 1603391777
transform -1 0 298600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_176
timestamp 1603391777
transform -1 0 302600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_177
timestamp 1603391777
transform -1 0 306600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_178
timestamp 1603391777
transform -1 0 310600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_179
timestamp 1603391777
transform -1 0 310800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_180
timestamp 1603391777
transform -1 0 311000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_185
timestamp 1603391777
transform -1 0 343000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_184
timestamp 1603391777
transform -1 0 339000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_183
timestamp 1603391777
transform -1 0 335000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_182
timestamp 1603391777
transform -1 0 331000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_189
timestamp 1603391777
transform -1 0 359000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_188
timestamp 1603391777
transform -1 0 355000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_187
timestamp 1603391777
transform -1 0 351000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_186
timestamp 1603391777
transform -1 0 347000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_191
timestamp 1603391777
transform -1 0 359400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_190
timestamp 1603391777
transform -1 0 359200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  flash_io0_pad
timestamp 1603391777
transform -1 0 375400 0 -1 39593
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_194
timestamp 1603391777
transform -1 0 383400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_193
timestamp 1603391777
transform -1 0 379400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_198
timestamp 1603391777
transform -1 0 399400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_197
timestamp 1603391777
transform -1 0 395400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_196
timestamp 1603391777
transform -1 0 391400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_195
timestamp 1603391777
transform -1 0 387400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_202
timestamp 1603391777
transform -1 0 407800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_201
timestamp 1603391777
transform -1 0 407600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_200
timestamp 1603391777
transform -1 0 407400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_199
timestamp 1603391777
transform -1 0 403400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  flash_io1_pad
timestamp 1603391777
transform -1 0 423800 0 -1 39593
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_204
timestamp 1603391777
transform -1 0 427800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_205
timestamp 1603391777
transform -1 0 431800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_206
timestamp 1603391777
transform -1 0 435800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_207
timestamp 1603391777
transform -1 0 439800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_208
timestamp 1603391777
transform -1 0 443800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_209
timestamp 1603391777
transform -1 0 447800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_210
timestamp 1603391777
transform -1 0 451800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  gpio_pad
timestamp 1603391777
transform -1 0 472000 0 -1 39593
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_211
timestamp 1603391777
transform -1 0 455800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_212
timestamp 1603391777
transform -1 0 456000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_214
timestamp 1603391777
transform -1 0 476000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_215
timestamp 1603391777
transform -1 0 480000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_216
timestamp 1603391777
transform -1 0 484000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_217
timestamp 1603391777
transform -1 0 488000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_218
timestamp 1603391777
transform -1 0 492000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vssio_hvc_pad  mgmt_vssio_hvclamp_pad\[1\] /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform -1 0 519400 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_219
timestamp 1603391777
transform -1 0 496000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_220
timestamp 1603391777
transform -1 0 500000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_221
timestamp 1603391777
transform -1 0 504000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_222
timestamp 1603391777
transform -1 0 504200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_223
timestamp 1603391777
transform -1 0 504400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_225
timestamp 1603391777
transform -1 0 523400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_226
timestamp 1603391777
transform -1 0 527400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_227
timestamp 1603391777
transform -1 0 531400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_231
timestamp 1603391777
transform -1 0 547400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_230
timestamp 1603391777
transform -1 0 543400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_229
timestamp 1603391777
transform -1 0 539400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_228
timestamp 1603391777
transform -1 0 535400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_234
timestamp 1603391777
transform -1 0 551800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_233
timestamp 1603391777
transform -1 0 551600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_232
timestamp 1603391777
transform -1 0 551400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  mgmt_vdda_hvclamp_pad /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform -1 0 566800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_237
timestamp 1603391777
transform -1 0 574800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_236
timestamp 1603391777
transform -1 0 570800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_242
timestamp 1603391777
transform -1 0 594800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_241
timestamp 1603391777
transform -1 0 590800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_240
timestamp 1603391777
transform -1 0 586800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_239
timestamp 1603391777
transform -1 0 582800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_238
timestamp 1603391777
transform -1 0 578800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_245
timestamp 1603391777
transform -1 0 599200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_244
timestamp 1603391777
transform -1 0 599000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_243
timestamp 1603391777
transform -1 0 598800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_504
timestamp 1603391777
transform 0 1 600407 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1603391777
transform 0 1 599200 -1 0 40000
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_249
timestamp 1603391777
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_248
timestamp 1603391777
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_247
timestamp 1603391777
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_255
timestamp 1603391777
transform 0 -1 39593 1 0 70000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_254
timestamp 1603391777
transform 0 -1 39593 1 0 69800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_253 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform 0 -1 39593 1 0 68800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_252
timestamp 1603391777
transform 0 -1 39593 1 0 64800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_251
timestamp 1603391777
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_250
timestamp 1603391777
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  mgmt_vccd_lvclamp_pad /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform 0 -1 39593 1 0 70200
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_508
timestamp 1603391777
transform 0 1 600407 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_507
timestamp 1603391777
transform 0 1 600407 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1603391777
transform 0 1 600407 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1603391777
transform 0 1 600407 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_515
timestamp 1603391777
transform 0 1 600407 -1 0 71600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_514
timestamp 1603391777
transform 0 1 600407 -1 0 71400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_513
timestamp 1603391777
transform 0 1 600407 -1 0 71200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_512
timestamp 1603391777
transform 0 1 600407 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_511 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform 0 1 600407 -1 0 70000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_510
timestamp 1603391777
transform 0 1 600407 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_509
timestamp 1603391777
transform 0 1 600407 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[0\]
timestamp 1603391777
transform 0 1 600407 -1 0 87600
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_259
timestamp 1603391777
transform 0 -1 39593 1 0 93200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_258
timestamp 1603391777
transform 0 -1 39593 1 0 89200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_257
timestamp 1603391777
transform 0 -1 39593 1 0 85200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_263
timestamp 1603391777
transform 0 -1 39593 1 0 109200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_262
timestamp 1603391777
transform 0 -1 39593 1 0 105200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_261
timestamp 1603391777
transform 0 -1 39593 1 0 101200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_260
timestamp 1603391777
transform 0 -1 39593 1 0 97200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_267
timestamp 1603391777
transform 0 -1 39593 1 0 114600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_266
timestamp 1603391777
transform 0 -1 39593 1 0 114400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_265
timestamp 1603391777
transform 0 -1 39593 1 0 114200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_264
timestamp 1603391777
transform 0 -1 39593 1 0 113200
box 0 0 1000 39593
use sky130_ef_io__vddio_hvc_pad  mgmt_vddio_hvclamp_pad\[0\] /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_ef_io/mag
timestamp 1603391777
transform 0 -1 39593 1 0 114800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_519
timestamp 1603391777
transform 0 1 600407 -1 0 99600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_518
timestamp 1603391777
transform 0 1 600407 -1 0 95600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_517
timestamp 1603391777
transform 0 1 600407 -1 0 91600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_523
timestamp 1603391777
transform 0 1 600407 -1 0 115600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_522
timestamp 1603391777
transform 0 1 600407 -1 0 111600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_521
timestamp 1603391777
transform 0 1 600407 -1 0 107600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_520
timestamp 1603391777
transform 0 1 600407 -1 0 103600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_528
timestamp 1603391777
transform 0 1 600407 -1 0 119200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_527
timestamp 1603391777
transform 0 1 600407 -1 0 119000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_526
timestamp 1603391777
transform 0 1 600407 -1 0 118800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_525
timestamp 1603391777
transform 0 1 600407 -1 0 118600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_524
timestamp 1603391777
transform 0 1 600407 -1 0 117600
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[1\]
timestamp 1603391777
transform 0 1 600407 -1 0 135200
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_271
timestamp 1603391777
transform 0 -1 39593 1 0 137800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_270
timestamp 1603391777
transform 0 -1 39593 1 0 133800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_269
timestamp 1603391777
transform 0 -1 39593 1 0 129800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_275
timestamp 1603391777
transform 0 -1 39593 1 0 153800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_274
timestamp 1603391777
transform 0 -1 39593 1 0 149800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_273
timestamp 1603391777
transform 0 -1 39593 1 0 145800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_272
timestamp 1603391777
transform 0 -1 39593 1 0 141800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_279
timestamp 1603391777
transform 0 -1 39593 1 0 159200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_278
timestamp 1603391777
transform 0 -1 39593 1 0 159000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_277
timestamp 1603391777
transform 0 -1 39593 1 0 158800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_276
timestamp 1603391777
transform 0 -1 39593 1 0 157800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[19\]
timestamp 1603391777
transform 0 -1 39593 1 0 159400
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_530
timestamp 1603391777
transform 0 1 600407 -1 0 139200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_531
timestamp 1603391777
transform 0 1 600407 -1 0 143200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_532
timestamp 1603391777
transform 0 1 600407 -1 0 147200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_533
timestamp 1603391777
transform 0 1 600407 -1 0 151200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_534
timestamp 1603391777
transform 0 1 600407 -1 0 155200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1603391777
transform 0 1 600407 -1 0 159200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1603391777
transform 0 1 600407 -1 0 163200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_537
timestamp 1603391777
transform 0 1 600407 -1 0 165200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_281
timestamp 1603391777
transform 0 -1 39593 1 0 175400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_282
timestamp 1603391777
transform 0 -1 39593 1 0 179400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_283
timestamp 1603391777
transform 0 -1 39593 1 0 183400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_284
timestamp 1603391777
transform 0 -1 39593 1 0 187400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_285
timestamp 1603391777
transform 0 -1 39593 1 0 191400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_286
timestamp 1603391777
transform 0 -1 39593 1 0 195400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_287
timestamp 1603391777
transform 0 -1 39593 1 0 199400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_288
timestamp 1603391777
transform 0 -1 39593 1 0 203400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_541
timestamp 1603391777
transform 0 1 600407 -1 0 166800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_540
timestamp 1603391777
transform 0 1 600407 -1 0 166600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_539
timestamp 1603391777
transform 0 1 600407 -1 0 166400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_538
timestamp 1603391777
transform 0 1 600407 -1 0 166200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[2\]
timestamp 1603391777
transform 0 1 600407 -1 0 182800
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1603391777
transform 0 1 600407 -1 0 198800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1603391777
transform 0 1 600407 -1 0 194800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_544
timestamp 1603391777
transform 0 1 600407 -1 0 190800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_543
timestamp 1603391777
transform 0 1 600407 -1 0 186800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_548
timestamp 1603391777
transform 0 1 600407 -1 0 206800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_547
timestamp 1603391777
transform 0 1 600407 -1 0 202800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_291
timestamp 1603391777
transform 0 -1 39593 1 0 204800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_290
timestamp 1603391777
transform 0 -1 39593 1 0 204600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_289
timestamp 1603391777
transform 0 -1 39593 1 0 204400
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[18\]
timestamp 1603391777
transform 0 -1 39593 1 0 205000
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_296
timestamp 1603391777
transform 0 -1 39593 1 0 233000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_295
timestamp 1603391777
transform 0 -1 39593 1 0 229000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_294
timestamp 1603391777
transform 0 -1 39593 1 0 225000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_293
timestamp 1603391777
transform 0 -1 39593 1 0 221000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_298
timestamp 1603391777
transform 0 -1 39593 1 0 241000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_297
timestamp 1603391777
transform 0 -1 39593 1 0 237000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_554
timestamp 1603391777
transform 0 1 600407 -1 0 214400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_553
timestamp 1603391777
transform 0 1 600407 -1 0 214200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_552
timestamp 1603391777
transform 0 1 600407 -1 0 214000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_551
timestamp 1603391777
transform 0 1 600407 -1 0 213800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_550
timestamp 1603391777
transform 0 1 600407 -1 0 212800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_549
timestamp 1603391777
transform 0 1 600407 -1 0 210800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[3\]
timestamp 1603391777
transform 0 1 600407 -1 0 230400
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_557
timestamp 1603391777
transform 0 1 600407 -1 0 238400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1603391777
transform 0 1 600407 -1 0 234400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_559
timestamp 1603391777
transform 0 1 600407 -1 0 246400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_558
timestamp 1603391777
transform 0 1 600407 -1 0 242400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_302
timestamp 1603391777
transform 0 -1 39593 1 0 250200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_301
timestamp 1603391777
transform 0 -1 39593 1 0 250000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_300
timestamp 1603391777
transform 0 -1 39593 1 0 249000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_299
timestamp 1603391777
transform 0 -1 39593 1 0 245000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[17\]
timestamp 1603391777
transform 0 -1 39593 1 0 250400
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_306
timestamp 1603391777
transform 0 -1 39593 1 0 274400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_305
timestamp 1603391777
transform 0 -1 39593 1 0 270400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_304
timestamp 1603391777
transform 0 -1 39593 1 0 266400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_308
timestamp 1603391777
transform 0 -1 39593 1 0 282400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_307
timestamp 1603391777
transform 0 -1 39593 1 0 278400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_564
timestamp 1603391777
transform 0 1 600407 -1 0 261400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_563
timestamp 1603391777
transform 0 1 600407 -1 0 260400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_562
timestamp 1603391777
transform 0 1 600407 -1 0 258400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_561
timestamp 1603391777
transform 0 1 600407 -1 0 254400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_560
timestamp 1603391777
transform 0 1 600407 -1 0 250400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_567
timestamp 1603391777
transform 0 1 600407 -1 0 262000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_566
timestamp 1603391777
transform 0 1 600407 -1 0 261800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_565
timestamp 1603391777
transform 0 1 600407 -1 0 261600
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[4\]
timestamp 1603391777
transform 0 1 600407 -1 0 278000
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_570
timestamp 1603391777
transform 0 1 600407 -1 0 286000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_569
timestamp 1603391777
transform 0 1 600407 -1 0 282000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_314
timestamp 1603391777
transform 0 -1 39593 1 0 295800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_313
timestamp 1603391777
transform 0 -1 39593 1 0 295600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_312
timestamp 1603391777
transform 0 -1 39593 1 0 295400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_311
timestamp 1603391777
transform 0 -1 39593 1 0 294400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_310
timestamp 1603391777
transform 0 -1 39593 1 0 290400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_309
timestamp 1603391777
transform 0 -1 39593 1 0 286400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[16\]
timestamp 1603391777
transform 0 -1 39593 1 0 296000
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_317
timestamp 1603391777
transform 0 -1 39593 1 0 316000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_316
timestamp 1603391777
transform 0 -1 39593 1 0 312000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_319
timestamp 1603391777
transform 0 -1 39593 1 0 324000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_318
timestamp 1603391777
transform 0 -1 39593 1 0 320000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_574
timestamp 1603391777
transform 0 1 600407 -1 0 302000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_573
timestamp 1603391777
transform 0 1 600407 -1 0 298000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_572
timestamp 1603391777
transform 0 1 600407 -1 0 294000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_571
timestamp 1603391777
transform 0 1 600407 -1 0 290000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_580
timestamp 1603391777
transform 0 1 600407 -1 0 309600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_579
timestamp 1603391777
transform 0 1 600407 -1 0 309400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_578
timestamp 1603391777
transform 0 1 600407 -1 0 309200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_577
timestamp 1603391777
transform 0 1 600407 -1 0 309000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_576
timestamp 1603391777
transform 0 1 600407 -1 0 308000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1603391777
transform 0 1 600407 -1 0 306000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[5\]
timestamp 1603391777
transform 0 1 600407 -1 0 325600
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_582
timestamp 1603391777
transform 0 1 600407 -1 0 329600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_326
timestamp 1603391777
transform 0 -1 39593 1 0 341400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_325
timestamp 1603391777
transform 0 -1 39593 1 0 341200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_324
timestamp 1603391777
transform 0 -1 39593 1 0 341000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_323
timestamp 1603391777
transform 0 -1 39593 1 0 340000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_322
timestamp 1603391777
transform 0 -1 39593 1 0 336000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_321
timestamp 1603391777
transform 0 -1 39593 1 0 332000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_320
timestamp 1603391777
transform 0 -1 39593 1 0 328000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[15\]
timestamp 1603391777
transform 0 -1 39593 1 0 341600
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_328
timestamp 1603391777
transform 0 -1 39593 1 0 357600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_330
timestamp 1603391777
transform 0 -1 39593 1 0 365600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_329
timestamp 1603391777
transform 0 -1 39593 1 0 361600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1603391777
transform 0 1 600407 -1 0 345600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1603391777
transform 0 1 600407 -1 0 341600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_584
timestamp 1603391777
transform 0 1 600407 -1 0 337600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_583
timestamp 1603391777
transform 0 1 600407 -1 0 333600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_594
timestamp 1603391777
transform 0 1 600407 -1 0 357400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_593
timestamp 1603391777
transform 0 1 600407 -1 0 357200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_592
timestamp 1603391777
transform 0 1 600407 -1 0 357000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_591
timestamp 1603391777
transform 0 1 600407 -1 0 356800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_590
timestamp 1603391777
transform 0 1 600407 -1 0 356600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_589
timestamp 1603391777
transform 0 1 600407 -1 0 355600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_588
timestamp 1603391777
transform 0 1 600407 -1 0 353600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_587
timestamp 1603391777
transform 0 1 600407 -1 0 349600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[6\]
timestamp 1603391777
transform 0 1 600407 -1 0 373400
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_334
timestamp 1603391777
transform 0 -1 39593 1 0 381600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_333
timestamp 1603391777
transform 0 -1 39593 1 0 377600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_332
timestamp 1603391777
transform 0 -1 39593 1 0 373600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_331
timestamp 1603391777
transform 0 -1 39593 1 0 369600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_338
timestamp 1603391777
transform 0 -1 39593 1 0 387000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_337
timestamp 1603391777
transform 0 -1 39593 1 0 386800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_336
timestamp 1603391777
transform 0 -1 39593 1 0 386600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_335
timestamp 1603391777
transform 0 -1 39593 1 0 385600
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[14\]
timestamp 1603391777
transform 0 -1 39593 1 0 387200
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_341
timestamp 1603391777
transform 0 -1 39593 1 0 407200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_340
timestamp 1603391777
transform 0 -1 39593 1 0 403200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_598
timestamp 1603391777
transform 0 1 600407 -1 0 385400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_597
timestamp 1603391777
transform 0 1 600407 -1 0 381400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1603391777
transform 0 1 600407 -1 0 377400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_601
timestamp 1603391777
transform 0 1 600407 -1 0 397400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_600
timestamp 1603391777
transform 0 1 600407 -1 0 393400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_599
timestamp 1603391777
transform 0 1 600407 -1 0 389400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_607
timestamp 1603391777
transform 0 1 600407 -1 0 405000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_606
timestamp 1603391777
transform 0 1 600407 -1 0 404800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_605
timestamp 1603391777
transform 0 1 600407 -1 0 404600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_604
timestamp 1603391777
transform 0 1 600407 -1 0 404400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_603
timestamp 1603391777
transform 0 1 600407 -1 0 403400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_602
timestamp 1603391777
transform 0 1 600407 -1 0 401400
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1603391777
transform 0 1 600407 -1 0 420000
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_344
timestamp 1603391777
transform 0 -1 39593 1 0 419200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_343
timestamp 1603391777
transform 0 -1 39593 1 0 415200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_342
timestamp 1603391777
transform 0 -1 39593 1 0 411200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_349
timestamp 1603391777
transform 0 -1 39593 1 0 432400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_348
timestamp 1603391777
transform 0 -1 39593 1 0 432200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_347
timestamp 1603391777
transform 0 -1 39593 1 0 431200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_346
timestamp 1603391777
transform 0 -1 39593 1 0 427200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_345
timestamp 1603391777
transform 0 -1 39593 1 0 423200
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_pad  user2_vssd_lvclmap_pad
timestamp 1603391777
transform 0 -1 39593 1 0 432600
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_351
timestamp 1603391777
transform 0 -1 39593 1 0 447600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_609
timestamp 1603391777
transform 0 1 600407 -1 0 424000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_610
timestamp 1603391777
transform 0 1 600407 -1 0 428000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_611
timestamp 1603391777
transform 0 1 600407 -1 0 432000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_612
timestamp 1603391777
transform 0 1 600407 -1 0 436000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_613
timestamp 1603391777
transform 0 1 600407 -1 0 440000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_614
timestamp 1603391777
transform 0 1 600407 -1 0 444000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1603391777
transform 0 1 600407 -1 0 448000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_616
timestamp 1603391777
transform 0 1 600407 -1 0 450000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_355
timestamp 1603391777
transform 0 -1 39593 1 0 463600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_354
timestamp 1603391777
transform 0 -1 39593 1 0 459600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_353
timestamp 1603391777
transform 0 -1 39593 1 0 455600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_352
timestamp 1603391777
transform 0 -1 39593 1 0 451600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_361
timestamp 1603391777
transform 0 -1 39593 1 0 477000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_360
timestamp 1603391777
transform 0 -1 39593 1 0 476800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_359
timestamp 1603391777
transform 0 -1 39593 1 0 476600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_358
timestamp 1603391777
transform 0 -1 39593 1 0 475600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_357
timestamp 1603391777
transform 0 -1 39593 1 0 471600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_356
timestamp 1603391777
transform 0 -1 39593 1 0 467600
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user2_vdda_hvclamp_pad
timestamp 1603391777
transform 0 -1 39593 1 0 477200
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_620
timestamp 1603391777
transform 0 1 600407 -1 0 451600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_619
timestamp 1603391777
transform 0 1 600407 -1 0 451400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_618
timestamp 1603391777
transform 0 1 600407 -1 0 451200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_617
timestamp 1603391777
transform 0 1 600407 -1 0 451000
box 0 0 1000 39593
use sky130_ef_io__vssd_lvc_pad  user1_vssd_lvclmap_pad
timestamp 1603391777
transform 0 1 600407 -1 0 466600
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_625
timestamp 1603391777
transform 0 1 600407 -1 0 482600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1603391777
transform 0 1 600407 -1 0 478600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_623
timestamp 1603391777
transform 0 1 600407 -1 0 474600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_622
timestamp 1603391777
transform 0 1 600407 -1 0 470600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_627
timestamp 1603391777
transform 0 1 600407 -1 0 490600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_626
timestamp 1603391777
transform 0 1 600407 -1 0 486600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_366
timestamp 1603391777
transform 0 -1 39593 1 0 504200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_365
timestamp 1603391777
transform 0 -1 39593 1 0 500200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_364
timestamp 1603391777
transform 0 -1 39593 1 0 496200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_363
timestamp 1603391777
transform 0 -1 39593 1 0 492200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_373
timestamp 1603391777
transform 0 -1 39593 1 0 521600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_372
timestamp 1603391777
transform 0 -1 39593 1 0 521400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_371
timestamp 1603391777
transform 0 -1 39593 1 0 521200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_370
timestamp 1603391777
transform 0 -1 39593 1 0 520200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_369
timestamp 1603391777
transform 0 -1 39593 1 0 516200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_368
timestamp 1603391777
transform 0 -1 39593 1 0 512200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_367
timestamp 1603391777
transform 0 -1 39593 1 0 508200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[13\]
timestamp 1603391777
transform 0 -1 39593 1 0 521800
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_633
timestamp 1603391777
transform 0 1 600407 -1 0 498200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_632
timestamp 1603391777
transform 0 1 600407 -1 0 498000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_631
timestamp 1603391777
transform 0 1 600407 -1 0 497800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_630
timestamp 1603391777
transform 0 1 600407 -1 0 497600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_629
timestamp 1603391777
transform 0 1 600407 -1 0 496600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1603391777
transform 0 1 600407 -1 0 494600
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1603391777
transform 0 1 600407 -1 0 513200
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_636
timestamp 1603391777
transform 0 1 600407 -1 0 521200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_635
timestamp 1603391777
transform 0 1 600407 -1 0 517200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_639
timestamp 1603391777
transform 0 1 600407 -1 0 533200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_638
timestamp 1603391777
transform 0 1 600407 -1 0 529200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1603391777
transform 0 1 600407 -1 0 525200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_377
timestamp 1603391777
transform 0 -1 39593 1 0 545800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_376
timestamp 1603391777
transform 0 -1 39593 1 0 541800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1603391777
transform 0 -1 39593 1 0 537800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_381
timestamp 1603391777
transform 0 -1 39593 1 0 561800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_380
timestamp 1603391777
transform 0 -1 39593 1 0 557800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_379
timestamp 1603391777
transform 0 -1 39593 1 0 553800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_378
timestamp 1603391777
transform 0 -1 39593 1 0 549800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_385
timestamp 1603391777
transform 0 -1 39593 1 0 567200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_384
timestamp 1603391777
transform 0 -1 39593 1 0 567000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_383
timestamp 1603391777
transform 0 -1 39593 1 0 566800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_382
timestamp 1603391777
transform 0 -1 39593 1 0 565800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[12\]
timestamp 1603391777
transform 0 -1 39593 1 0 567400
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_646
timestamp 1603391777
transform 0 1 600407 -1 0 544800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_645
timestamp 1603391777
transform 0 1 600407 -1 0 544600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_644
timestamp 1603391777
transform 0 1 600407 -1 0 544400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_643
timestamp 1603391777
transform 0 1 600407 -1 0 544200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_642
timestamp 1603391777
transform 0 1 600407 -1 0 543200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_641
timestamp 1603391777
transform 0 1 600407 -1 0 541200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_640
timestamp 1603391777
transform 0 1 600407 -1 0 537200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[7\]
timestamp 1603391777
transform 0 1 600407 -1 0 560800
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_648
timestamp 1603391777
transform 0 1 600407 -1 0 564800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_650
timestamp 1603391777
transform 0 1 600407 -1 0 572800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_649
timestamp 1603391777
transform 0 1 600407 -1 0 568800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_387
timestamp 1603391777
transform 0 -1 39593 1 0 583400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_388
timestamp 1603391777
transform 0 -1 39593 1 0 587400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_389
timestamp 1603391777
transform 0 -1 39593 1 0 591400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_390
timestamp 1603391777
transform 0 -1 39593 1 0 595400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_391
timestamp 1603391777
transform 0 -1 39593 1 0 599400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_392
timestamp 1603391777
transform 0 -1 39593 1 0 603400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_393
timestamp 1603391777
transform 0 -1 39593 1 0 607400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_394
timestamp 1603391777
transform 0 -1 39593 1 0 611400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_654
timestamp 1603391777
transform 0 1 600407 -1 0 588800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_653
timestamp 1603391777
transform 0 1 600407 -1 0 584800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_652
timestamp 1603391777
transform 0 1 600407 -1 0 580800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_651
timestamp 1603391777
transform 0 1 600407 -1 0 576800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_659
timestamp 1603391777
transform 0 1 600407 -1 0 592400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_658
timestamp 1603391777
transform 0 1 600407 -1 0 592200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_657
timestamp 1603391777
transform 0 1 600407 -1 0 592000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_656
timestamp 1603391777
transform 0 1 600407 -1 0 591800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_655
timestamp 1603391777
transform 0 1 600407 -1 0 590800
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[8\]
timestamp 1603391777
transform 0 1 600407 -1 0 608400
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_661
timestamp 1603391777
transform 0 1 600407 -1 0 612400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_397
timestamp 1603391777
transform 0 -1 39593 1 0 612800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_396
timestamp 1603391777
transform 0 -1 39593 1 0 612600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_395
timestamp 1603391777
transform 0 -1 39593 1 0 612400
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[11\]
timestamp 1603391777
transform 0 -1 39593 1 0 613000
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_402
timestamp 1603391777
transform 0 -1 39593 1 0 641000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_401
timestamp 1603391777
transform 0 -1 39593 1 0 637000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_400
timestamp 1603391777
transform 0 -1 39593 1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_399
timestamp 1603391777
transform 0 -1 39593 1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_404
timestamp 1603391777
transform 0 -1 39593 1 0 649000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_403
timestamp 1603391777
transform 0 -1 39593 1 0 645000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1603391777
transform 0 1 600407 -1 0 628400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_664
timestamp 1603391777
transform 0 1 600407 -1 0 624400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_663
timestamp 1603391777
transform 0 1 600407 -1 0 620400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1603391777
transform 0 1 600407 -1 0 616400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_672
timestamp 1603391777
transform 0 1 600407 -1 0 640000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_671
timestamp 1603391777
transform 0 1 600407 -1 0 639800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_670
timestamp 1603391777
transform 0 1 600407 -1 0 639600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_669
timestamp 1603391777
transform 0 1 600407 -1 0 639400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_668
timestamp 1603391777
transform 0 1 600407 -1 0 638400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_667
timestamp 1603391777
transform 0 1 600407 -1 0 636400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1603391777
transform 0 1 600407 -1 0 632400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[9\]
timestamp 1603391777
transform 0 1 600407 -1 0 656000
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_408
timestamp 1603391777
transform 0 -1 39593 1 0 658200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_407
timestamp 1603391777
transform 0 -1 39593 1 0 658000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_406
timestamp 1603391777
transform 0 -1 39593 1 0 657000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1603391777
transform 0 -1 39593 1 0 653000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[10\]
timestamp 1603391777
transform 0 -1 39593 1 0 658400
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_412
timestamp 1603391777
transform 0 -1 39593 1 0 682400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_411
timestamp 1603391777
transform 0 -1 39593 1 0 678400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_410
timestamp 1603391777
transform 0 -1 39593 1 0 674400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_414
timestamp 1603391777
transform 0 -1 39593 1 0 690400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_413
timestamp 1603391777
transform 0 -1 39593 1 0 686400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_677
timestamp 1603391777
transform 0 1 600407 -1 0 672000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_676
timestamp 1603391777
transform 0 1 600407 -1 0 668000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1603391777
transform 0 1 600407 -1 0 664000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_674
timestamp 1603391777
transform 0 1 600407 -1 0 660000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_681
timestamp 1603391777
transform 0 1 600407 -1 0 686000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_680
timestamp 1603391777
transform 0 1 600407 -1 0 684000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_679
timestamp 1603391777
transform 0 1 600407 -1 0 680000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_678
timestamp 1603391777
transform 0 1 600407 -1 0 676000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_686
timestamp 1603391777
transform 0 1 600407 -1 0 687800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_685
timestamp 1603391777
transform 0 1 600407 -1 0 687600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_684
timestamp 1603391777
transform 0 1 600407 -1 0 687400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_683
timestamp 1603391777
transform 0 1 600407 -1 0 687200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_682
timestamp 1603391777
transform 0 1 600407 -1 0 687000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[10\]
timestamp 1603391777
transform 0 1 600407 -1 0 703800
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_420
timestamp 1603391777
transform 0 -1 39593 1 0 703800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_419
timestamp 1603391777
transform 0 -1 39593 1 0 703600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_418
timestamp 1603391777
transform 0 -1 39593 1 0 703400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_417
timestamp 1603391777
transform 0 -1 39593 1 0 702400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1603391777
transform 0 -1 39593 1 0 698400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1603391777
transform 0 -1 39593 1 0 694400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[9\]
timestamp 1603391777
transform 0 -1 39593 1 0 704000
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_423
timestamp 1603391777
transform 0 -1 39593 1 0 724000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_422
timestamp 1603391777
transform 0 -1 39593 1 0 720000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1603391777
transform 0 -1 39593 1 0 732000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_424
timestamp 1603391777
transform 0 -1 39593 1 0 728000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_688
timestamp 1603391777
transform 0 1 600407 -1 0 707800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_689
timestamp 1603391777
transform 0 1 600407 -1 0 711800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1603391777
transform 0 1 600407 -1 0 715800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_691
timestamp 1603391777
transform 0 1 600407 -1 0 719800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_692
timestamp 1603391777
transform 0 1 600407 -1 0 723800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1603391777
transform 0 1 600407 -1 0 727800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1603391777
transform 0 1 600407 -1 0 731800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_695
timestamp 1603391777
transform 0 1 600407 -1 0 733800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_696
timestamp 1603391777
transform 0 1 600407 -1 0 734800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_432
timestamp 1603391777
transform 0 -1 39593 1 0 749400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_431
timestamp 1603391777
transform 0 -1 39593 1 0 749200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_430
timestamp 1603391777
transform 0 -1 39593 1 0 749000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_429
timestamp 1603391777
transform 0 -1 39593 1 0 748000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_428
timestamp 1603391777
transform 0 -1 39593 1 0 744000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_427
timestamp 1603391777
transform 0 -1 39593 1 0 740000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1603391777
transform 0 -1 39593 1 0 736000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[8\]
timestamp 1603391777
transform 0 -1 39593 1 0 749600
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_434
timestamp 1603391777
transform 0 -1 39593 1 0 765600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1603391777
transform 0 -1 39593 1 0 773600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1603391777
transform 0 -1 39593 1 0 769600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_699
timestamp 1603391777
transform 0 1 600407 -1 0 735400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_698
timestamp 1603391777
transform 0 1 600407 -1 0 735200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_697
timestamp 1603391777
transform 0 1 600407 -1 0 735000
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[11\]
timestamp 1603391777
transform 0 1 600407 -1 0 751400
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_704
timestamp 1603391777
transform 0 1 600407 -1 0 767400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1603391777
transform 0 1 600407 -1 0 763400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_702
timestamp 1603391777
transform 0 1 600407 -1 0 759400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_701
timestamp 1603391777
transform 0 1 600407 -1 0 755400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_706
timestamp 1603391777
transform 0 1 600407 -1 0 775400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_705
timestamp 1603391777
transform 0 1 600407 -1 0 771400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_440
timestamp 1603391777
transform 0 -1 39593 1 0 789600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_439
timestamp 1603391777
transform 0 -1 39593 1 0 785600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_438
timestamp 1603391777
transform 0 -1 39593 1 0 781600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_437
timestamp 1603391777
transform 0 -1 39593 1 0 777600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_444
timestamp 1603391777
transform 0 -1 39593 1 0 795000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_443
timestamp 1603391777
transform 0 -1 39593 1 0 794800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_442
timestamp 1603391777
transform 0 -1 39593 1 0 794600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_441
timestamp 1603391777
transform 0 -1 39593 1 0 793600
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[7\]
timestamp 1603391777
transform 0 -1 39593 1 0 795200
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_447
timestamp 1603391777
transform 0 -1 39593 1 0 815200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1603391777
transform 0 -1 39593 1 0 811200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_712
timestamp 1603391777
transform 0 1 600407 -1 0 783000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_711
timestamp 1603391777
transform 0 1 600407 -1 0 782800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_710
timestamp 1603391777
transform 0 1 600407 -1 0 782600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_709
timestamp 1603391777
transform 0 1 600407 -1 0 782400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_708
timestamp 1603391777
transform 0 1 600407 -1 0 781400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_707
timestamp 1603391777
transform 0 1 600407 -1 0 779400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[12\]
timestamp 1603391777
transform 0 1 600407 -1 0 799000
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_716
timestamp 1603391777
transform 0 1 600407 -1 0 811000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_715
timestamp 1603391777
transform 0 1 600407 -1 0 807000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_714
timestamp 1603391777
transform 0 1 600407 -1 0 803000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1603391777
transform 0 1 600407 -1 0 819000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_717
timestamp 1603391777
transform 0 1 600407 -1 0 815000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_450
timestamp 1603391777
transform 0 -1 39593 1 0 827200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_449
timestamp 1603391777
transform 0 -1 39593 1 0 823200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_448
timestamp 1603391777
transform 0 -1 39593 1 0 819200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_455
timestamp 1603391777
transform 0 -1 39593 1 0 840400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_454
timestamp 1603391777
transform 0 -1 39593 1 0 840200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_453
timestamp 1603391777
transform 0 -1 39593 1 0 839200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_452
timestamp 1603391777
transform 0 -1 39593 1 0 835200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_451
timestamp 1603391777
transform 0 -1 39593 1 0 831200
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user2_vssa_hvclamp_pad
timestamp 1603391777
transform 0 -1 39593 1 0 840600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_457
timestamp 1603391777
transform 0 -1 39593 1 0 855600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_725
timestamp 1603391777
transform 0 1 600407 -1 0 830600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_724
timestamp 1603391777
transform 0 1 600407 -1 0 830400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_723
timestamp 1603391777
transform 0 1 600407 -1 0 830200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_722
timestamp 1603391777
transform 0 1 600407 -1 0 830000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_721
timestamp 1603391777
transform 0 1 600407 -1 0 829000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_720
timestamp 1603391777
transform 0 1 600407 -1 0 827000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_719
timestamp 1603391777
transform 0 1 600407 -1 0 823000
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1603391777
transform 0 1 600407 -1 0 845600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_727
timestamp 1603391777
transform 0 1 600407 -1 0 849600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_729
timestamp 1603391777
transform 0 1 600407 -1 0 857600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1603391777
transform 0 1 600407 -1 0 853600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_461
timestamp 1603391777
transform 0 -1 39593 1 0 871600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_460
timestamp 1603391777
transform 0 -1 39593 1 0 867600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_459
timestamp 1603391777
transform 0 -1 39593 1 0 863600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_458
timestamp 1603391777
transform 0 -1 39593 1 0 859600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_467
timestamp 1603391777
transform 0 -1 39593 1 0 885000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_466
timestamp 1603391777
transform 0 -1 39593 1 0 884800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_465
timestamp 1603391777
transform 0 -1 39593 1 0 884600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_464
timestamp 1603391777
transform 0 -1 39593 1 0 883600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_463
timestamp 1603391777
transform 0 -1 39593 1 0 879600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_462
timestamp 1603391777
transform 0 -1 39593 1 0 875600
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1603391777
transform 0 -1 39593 1 0 885200
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_733
timestamp 1603391777
transform 0 1 600407 -1 0 873600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_732
timestamp 1603391777
transform 0 1 600407 -1 0 869600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1603391777
transform 0 1 600407 -1 0 865600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_730
timestamp 1603391777
transform 0 1 600407 -1 0 861600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_738
timestamp 1603391777
transform 0 1 600407 -1 0 877200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_737
timestamp 1603391777
transform 0 1 600407 -1 0 877000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_736
timestamp 1603391777
transform 0 1 600407 -1 0 876800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_735
timestamp 1603391777
transform 0 1 600407 -1 0 876600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_734
timestamp 1603391777
transform 0 1 600407 -1 0 875600
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[13\]
timestamp 1603391777
transform 0 1 600407 -1 0 893200
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1603391777
transform 0 1 600407 -1 0 901200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1603391777
transform 0 1 600407 -1 0 897200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_472
timestamp 1603391777
transform 0 -1 39593 1 0 912200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_471
timestamp 1603391777
transform 0 -1 39593 1 0 908200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_470
timestamp 1603391777
transform 0 -1 39593 1 0 904200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_469
timestamp 1603391777
transform 0 -1 39593 1 0 900200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1603391777
transform 0 -1 39593 1 0 924200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_474
timestamp 1603391777
transform 0 -1 39593 1 0 920200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_473
timestamp 1603391777
transform 0 -1 39593 1 0 916200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_479
timestamp 1603391777
transform 0 -1 39593 1 0 929600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_478
timestamp 1603391777
transform 0 -1 39593 1 0 929400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_477
timestamp 1603391777
transform 0 -1 39593 1 0 929200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_476
timestamp 1603391777
transform 0 -1 39593 1 0 928200
box 0 0 1000 39593
use sky130_ef_io__vccd_lvc_pad  user2_vccd_lvclamp_pad
timestamp 1603391777
transform 0 -1 39593 1 0 929800
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_744
timestamp 1603391777
transform 0 1 600407 -1 0 913200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_743
timestamp 1603391777
transform 0 1 600407 -1 0 909200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_742
timestamp 1603391777
transform 0 1 600407 -1 0 905200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_751
timestamp 1603391777
transform 0 1 600407 -1 0 924800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_750
timestamp 1603391777
transform 0 1 600407 -1 0 924600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_749
timestamp 1603391777
transform 0 1 600407 -1 0 924400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_748
timestamp 1603391777
transform 0 1 600407 -1 0 924200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_747
timestamp 1603391777
transform 0 1 600407 -1 0 923200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_746
timestamp 1603391777
transform 0 1 600407 -1 0 921200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_745
timestamp 1603391777
transform 0 1 600407 -1 0 917200
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  user1_vccd_lvclamp_pad
timestamp 1603391777
transform 0 1 600407 -1 0 939800
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_483
timestamp 1603391777
transform 0 -1 39593 1 0 952800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_482
timestamp 1603391777
transform 0 -1 39593 1 0 948800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_481
timestamp 1603391777
transform 0 -1 39593 1 0 944800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_487
timestamp 1603391777
transform 0 -1 39593 1 0 968800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1603391777
transform 0 -1 39593 1 0 964800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1603391777
transform 0 -1 39593 1 0 960800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_484
timestamp 1603391777
transform 0 -1 39593 1 0 956800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_491
timestamp 1603391777
transform 0 -1 39593 1 0 974200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_490
timestamp 1603391777
transform 0 -1 39593 1 0 974000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_489
timestamp 1603391777
transform 0 -1 39593 1 0 973800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_488
timestamp 1603391777
transform 0 -1 39593 1 0 972800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[6\]
timestamp 1603391777
transform 0 -1 39593 1 0 974400
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1603391777
transform 0 1 600407 -1 0 955800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_755
timestamp 1603391777
transform 0 1 600407 -1 0 951800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_754
timestamp 1603391777
transform 0 1 600407 -1 0 947800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_753
timestamp 1603391777
transform 0 1 600407 -1 0 943800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_761
timestamp 1603391777
transform 0 1 600407 -1 0 970800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_760
timestamp 1603391777
transform 0 1 600407 -1 0 969800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1603391777
transform 0 1 600407 -1 0 967800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_758
timestamp 1603391777
transform 0 1 600407 -1 0 963800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_757
timestamp 1603391777
transform 0 1 600407 -1 0 959800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_764
timestamp 1603391777
transform 0 1 600407 -1 0 971400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_763
timestamp 1603391777
transform 0 1 600407 -1 0 971200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_762
timestamp 1603391777
transform 0 1 600407 -1 0 971000
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[14\]
timestamp 1603391777
transform 0 1 600407 -1 0 987400
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1603391777
transform 0 -1 39593 1 0 998400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_494
timestamp 1603391777
transform 0 -1 39593 1 0 994400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_493
timestamp 1603391777
transform 0 -1 39593 1 0 990400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_503
timestamp 1603391777
transform 0 -1 39593 1 0 1019800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_502
timestamp 1603391777
transform 0 -1 39593 1 0 1019600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_501
timestamp 1603391777
transform 0 -1 39593 1 0 1019400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_500
timestamp 1603391777
transform 0 -1 39593 1 0 1018400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_499
timestamp 1603391777
transform 0 -1 39593 1 0 1014400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_498
timestamp 1603391777
transform 0 -1 39593 1 0 1010400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_497
timestamp 1603391777
transform 0 -1 39593 1 0 1006400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1603391777
transform 0 -1 39593 1 0 1002400
box 0 0 4000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1603391777
transform 0 -1 40800 1 0 1020000
box 0 0 40000 40800
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[5\]
timestamp 1603391777
transform 1 0 72800 0 1 1020407
box 0 -407 16000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[4\]
timestamp 1603391777
transform 1 0 121000 0 1 1020407
box 0 -407 16000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[3\]
timestamp 1603391777
transform 1 0 169000 0 1 1020407
box 0 -407 16000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[2\]
timestamp 1603391777
transform 1 0 217200 0 1 1020407
box 0 -407 16000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[1\]
timestamp 1603391777
transform 1 0 265200 0 1 1020407
box 0 -407 16000 39593
use sky130_ef_io__vssio_hvc_pad  mgmt_vssio_hvclamp_pad\[0\]
timestamp 1603391777
transform 1 0 313400 0 1 1020407
box 0 -407 15000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area2_io_pad\[0\]
timestamp 1603391777
transform 1 0 360400 0 1 1020407
box 0 -407 16000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[17\]
timestamp 1603391777
transform 1 0 408600 0 1 1020407
box 0 -407 16000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[16\]
timestamp 1603391777
transform 1 0 456600 0 1 1020407
box 0 -407 16000 39593
use sky130_ef_io__vssa_hvc_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1603391777
transform 1 0 504800 0 1 1020407
box 0 -407 15000 39593
use sky130_ef_io__gpiov2_pad  mprj_pads/area1_io_pad\[15\]
timestamp 1603391777
transform 1 0 551800 0 1 1020407
box 0 -407 16000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1603391777
transform 0 1 600407 -1 0 1003400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_768
timestamp 1603391777
transform 0 1 600407 -1 0 999400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_767
timestamp 1603391777
transform 0 1 600407 -1 0 995400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_766
timestamp 1603391777
transform 0 1 600407 -1 0 991400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_778
timestamp 1603391777
transform 0 1 600407 -1 0 1019200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_777
timestamp 1603391777
transform 0 1 600407 -1 0 1019000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_776
timestamp 1603391777
transform 0 1 600407 -1 0 1018800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_775
timestamp 1603391777
transform 0 1 600407 -1 0 1018600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_774
timestamp 1603391777
transform 0 1 600407 -1 0 1018400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_773
timestamp 1603391777
transform 0 1 600407 -1 0 1017400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_772
timestamp 1603391777
transform 0 1 600407 -1 0 1015400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_771
timestamp 1603391777
transform 0 1 600407 -1 0 1011400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_770
timestamp 1603391777
transform 0 1 600407 -1 0 1007400
box 0 0 4000 39593
use sky130_ef_io__corner_pad  user1_corner
timestamp 1603391777
transform 1 0 600000 0 1 1019200
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_5
timestamp 1603391777
transform 1 0 40800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1603391777
transform 1 0 44800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1603391777
transform 1 0 48800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1603391777
transform 1 0 52800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1603391777
transform 1 0 56800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1603391777
transform 1 0 60800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1603391777
transform 1 0 64800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1603391777
transform 1 0 68800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_14
timestamp 1603391777
transform 1 0 88800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_15
timestamp 1603391777
transform 1 0 92800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_16
timestamp 1603391777
transform 1 0 96800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_17
timestamp 1603391777
transform 1 0 100800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1603391777
transform 1 0 104800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1603391777
transform 1 0 108800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1603391777
transform 1 0 112800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1603391777
transform 1 0 116800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_22
timestamp 1603391777
transform 1 0 120800 0 1 1020407
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1603391777
transform 1 0 137000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1603391777
transform 1 0 141000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_26
timestamp 1603391777
transform 1 0 145000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_27
timestamp 1603391777
transform 1 0 149000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_28
timestamp 1603391777
transform 1 0 153000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_29
timestamp 1603391777
transform 1 0 157000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_30
timestamp 1603391777
transform 1 0 161000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1603391777
transform 1 0 165000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1603391777
transform 1 0 185000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1603391777
transform 1 0 189000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1603391777
transform 1 0 193000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1603391777
transform 1 0 197000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1603391777
transform 1 0 201000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_38
timestamp 1603391777
transform 1 0 205000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_39
timestamp 1603391777
transform 1 0 209000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_40
timestamp 1603391777
transform 1 0 213000 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_41
timestamp 1603391777
transform 1 0 217000 0 1 1020407
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_43
timestamp 1603391777
transform 1 0 233200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1603391777
transform 1 0 237200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1603391777
transform 1 0 241200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1603391777
transform 1 0 245200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_47
timestamp 1603391777
transform 1 0 249200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_48
timestamp 1603391777
transform 1 0 253200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1603391777
transform 1 0 257200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1603391777
transform 1 0 261200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_52
timestamp 1603391777
transform 1 0 281200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_53
timestamp 1603391777
transform 1 0 285200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_54
timestamp 1603391777
transform 1 0 289200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_55
timestamp 1603391777
transform 1 0 293200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_56
timestamp 1603391777
transform 1 0 297200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_57
timestamp 1603391777
transform 1 0 301200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_58
timestamp 1603391777
transform 1 0 305200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_59
timestamp 1603391777
transform 1 0 309200 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_60
timestamp 1603391777
transform 1 0 313200 0 1 1020407
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1603391777
transform 1 0 328400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1603391777
transform 1 0 332400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1603391777
transform 1 0 336400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_65
timestamp 1603391777
transform 1 0 340400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_66
timestamp 1603391777
transform 1 0 344400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_67
timestamp 1603391777
transform 1 0 348400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_68
timestamp 1603391777
transform 1 0 352400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_69
timestamp 1603391777
transform 1 0 356400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1603391777
transform 1 0 376400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1603391777
transform 1 0 380400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1603391777
transform 1 0 384400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_74
timestamp 1603391777
transform 1 0 388400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_75
timestamp 1603391777
transform 1 0 392400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_76
timestamp 1603391777
transform 1 0 396400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_77
timestamp 1603391777
transform 1 0 400400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1603391777
transform 1 0 404400 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_79
timestamp 1603391777
transform 1 0 408400 0 1 1020407
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_81
timestamp 1603391777
transform 1 0 424600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_82
timestamp 1603391777
transform 1 0 428600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_83
timestamp 1603391777
transform 1 0 432600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_84
timestamp 1603391777
transform 1 0 436600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_85
timestamp 1603391777
transform 1 0 440600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1603391777
transform 1 0 444600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1603391777
transform 1 0 448600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1603391777
transform 1 0 452600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1603391777
transform 1 0 472600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1603391777
transform 1 0 476600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_92
timestamp 1603391777
transform 1 0 480600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_93
timestamp 1603391777
transform 1 0 484600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_94
timestamp 1603391777
transform 1 0 488600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_95
timestamp 1603391777
transform 1 0 492600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_96
timestamp 1603391777
transform 1 0 496600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_97
timestamp 1603391777
transform 1 0 500600 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_98
timestamp 1603391777
transform 1 0 504600 0 1 1020407
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1603391777
transform 1 0 519800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1603391777
transform 1 0 523800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1603391777
transform 1 0 527800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1603391777
transform 1 0 531800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1603391777
transform 1 0 535800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_105
timestamp 1603391777
transform 1 0 539800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_106
timestamp 1603391777
transform 1 0 543800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_107
timestamp 1603391777
transform 1 0 547800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_109
timestamp 1603391777
transform 1 0 567800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_110
timestamp 1603391777
transform 1 0 571800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1603391777
transform 1 0 575800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1603391777
transform 1 0 579800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1603391777
transform 1 0 583800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1603391777
transform 1 0 587800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1603391777
transform 1 0 591800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_116
timestamp 1603391777
transform 1 0 595800 0 1 1020407
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_117
timestamp 1603391777
transform 1 0 599800 0 1 1020407
box 0 0 200 39593
<< labels >>
rlabel metal5 s 168240 6598 180760 19088 6 clock
port 0 nsew default input
rlabel metal3 s 167086 2088 167152 40000 6 clock_core
port 1 nsew default tristate
rlabel metal5 s 312240 6598 324760 19088 6 flash_clk
port 2 nsew default tristate
rlabel metal2 s 322477 38715 322529 39999 6 flash_clk_core
port 3 nsew default input
rlabel metal2 s 317899 38982 317951 40000 6 flash_clk_ieb_core
port 4 nsew default input
rlabel metal2 s 326279 39105 326325 39999 6 flash_clk_oeb_core
port 5 nsew default input
rlabel metal5 s 263840 6598 276360 19088 6 flash_csb
port 6 nsew default tristate
rlabel metal2 s 274077 38715 274129 39999 6 flash_csb_core
port 7 nsew default input
rlabel metal2 s 269499 38982 269551 40000 6 flash_csb_ieb_core
port 8 nsew default input
rlabel metal2 s 277879 39105 277925 39999 6 flash_csb_oeb_core
port 9 nsew default input
rlabel metal5 s 360640 6598 373160 19088 6 flash_io0
port 10 nsew default bidirectional
rlabel metal3 s 359486 2088 359552 40000 6 flash_io0_di_core
port 11 nsew default tristate
rlabel metal2 s 370877 38715 370929 39999 6 flash_io0_do_core
port 12 nsew default input
rlabel metal2 s 366299 38982 366351 40000 6 flash_io0_ieb_core
port 13 nsew default input
rlabel metal2 s 374679 39105 374725 39999 6 flash_io0_oeb_core
port 14 nsew default input
rlabel metal5 s 409040 6598 421560 19088 6 flash_io1
port 15 nsew default bidirectional
rlabel metal3 s 407886 2088 407952 40000 6 flash_io1_di_core
port 16 nsew default tristate
rlabel metal2 s 419277 38715 419329 39999 6 flash_io1_do_core
port 17 nsew default input
rlabel metal2 s 414699 38982 414751 40000 6 flash_io1_ieb_core
port 18 nsew default input
rlabel metal2 s 423079 39105 423125 39999 6 flash_io1_oeb_core
port 19 nsew default input
rlabel metal5 s 457240 6598 469760 19088 6 gpio
port 20 nsew default bidirectional
rlabel metal3 s 456086 2088 456152 40000 6 gpio_in_core
port 21 nsew default tristate
rlabel metal2 s 462899 38982 462951 40000 6 gpio_inenb_core
port 22 nsew default input
rlabel metal2 s 461977 39891 462029 39999 6 gpio_mode0_core
port 23 nsew default input
rlabel metal2 s 466250 39186 466302 40000 6 gpio_mode1_core
port 24 nsew default input
rlabel metal2 s 467477 38715 467529 39999 6 gpio_out_core
port 25 nsew default input
rlabel metal2 s 471279 39105 471325 39999 6 gpio_outenb_core
port 26 nsew default input
rlabel metal5 s 620912 72840 633402 85360 6 mprj_io[0]
port 27 nsew default bidirectional
rlabel metal5 s 620912 689040 633402 701560 6 mprj_io[10]
port 28 nsew default bidirectional
rlabel metal5 s 620912 736640 633402 749160 6 mprj_io[11]
port 29 nsew default bidirectional
rlabel metal5 s 620912 784240 633402 796760 6 mprj_io[12]
port 30 nsew default bidirectional
rlabel metal5 s 620912 878440 633402 890960 6 mprj_io[13]
port 31 nsew default bidirectional
rlabel metal5 s 620912 972640 633402 985160 6 mprj_io[14]
port 32 nsew default bidirectional
rlabel metal5 s 554040 1040912 566560 1053402 6 mprj_io[15]
port 33 nsew default bidirectional
rlabel metal5 s 458840 1040912 471360 1053402 6 mprj_io[16]
port 34 nsew default bidirectional
rlabel metal5 s 410840 1040912 423360 1053402 6 mprj_io[17]
port 35 nsew default bidirectional
rlabel metal5 s 362640 1040912 375160 1053402 6 mprj_io[18]
port 36 nsew default bidirectional
rlabel metal5 s 267440 1040912 279960 1053402 6 mprj_io[19]
port 37 nsew default bidirectional
rlabel metal5 s 620912 120440 633402 132960 6 mprj_io[1]
port 38 nsew default bidirectional
rlabel metal5 s 219440 1040912 231960 1053402 6 mprj_io[20]
port 39 nsew default bidirectional
rlabel metal5 s 171240 1040912 183760 1053402 6 mprj_io[21]
port 40 nsew default bidirectional
rlabel metal5 s 123240 1040912 135760 1053402 6 mprj_io[22]
port 41 nsew default bidirectional
rlabel metal5 s 75040 1040912 87560 1053402 6 mprj_io[23]
port 42 nsew default bidirectional
rlabel metal5 s 6598 976640 19088 989160 6 mprj_io[24]
port 43 nsew default bidirectional
rlabel metal5 s 6598 797440 19088 809960 6 mprj_io[25]
port 44 nsew default bidirectional
rlabel metal5 s 6598 751840 19088 764360 6 mprj_io[26]
port 45 nsew default bidirectional
rlabel metal5 s 6598 706240 19088 718760 6 mprj_io[27]
port 46 nsew default bidirectional
rlabel metal5 s 6598 660640 19088 673160 6 mprj_io[28]
port 47 nsew default bidirectional
rlabel metal5 s 6598 615240 19088 627760 6 mprj_io[29]
port 48 nsew default bidirectional
rlabel metal5 s 620912 168040 633402 180560 6 mprj_io[2]
port 49 nsew default bidirectional
rlabel metal5 s 6598 569640 19088 582160 6 mprj_io[30]
port 50 nsew default bidirectional
rlabel metal5 s 6598 524040 19088 536560 6 mprj_io[31]
port 51 nsew default bidirectional
rlabel metal5 s 6598 389440 19088 401960 6 mprj_io[32]
port 52 nsew default bidirectional
rlabel metal5 s 6598 343840 19088 356360 6 mprj_io[33]
port 53 nsew default bidirectional
rlabel metal5 s 6598 298240 19088 310760 6 mprj_io[34]
port 54 nsew default bidirectional
rlabel metal5 s 6598 252640 19088 265160 6 mprj_io[35]
port 55 nsew default bidirectional
rlabel metal5 s 6598 207240 19088 219760 6 mprj_io[36]
port 56 nsew default bidirectional
rlabel metal5 s 6598 161640 19088 174160 6 mprj_io[37]
port 57 nsew default bidirectional
rlabel metal5 s 620912 215640 633402 228160 6 mprj_io[3]
port 58 nsew default bidirectional
rlabel metal5 s 620912 263240 633402 275760 6 mprj_io[4]
port 59 nsew default bidirectional
rlabel metal5 s 620912 310840 633402 323360 6 mprj_io[5]
port 60 nsew default bidirectional
rlabel metal5 s 620912 358640 633402 371160 6 mprj_io[6]
port 61 nsew default bidirectional
rlabel metal5 s 620912 546040 633402 558560 6 mprj_io[7]
port 62 nsew default bidirectional
rlabel metal5 s 620912 593640 633402 606160 6 mprj_io[8]
port 63 nsew default bidirectional
rlabel metal5 s 620912 641240 633402 653760 6 mprj_io[9]
port 64 nsew default bidirectional
rlabel metal1 s 600000 75062 600260 75114 6 mprj_io_analog_en[0]
port 65 nsew default input
rlabel metal1 s 600000 691262 600260 691314 6 mprj_io_analog_en[10]
port 66 nsew default input
rlabel metal1 s 600000 738862 600260 738914 6 mprj_io_analog_en[11]
port 67 nsew default input
rlabel metal1 s 600000 786462 600260 786514 6 mprj_io_analog_en[12]
port 68 nsew default input
rlabel metal1 s 600000 880662 600260 880714 6 mprj_io_analog_en[13]
port 69 nsew default input
rlabel metal1 s 600000 974862 600260 974914 6 mprj_io_analog_en[14]
port 70 nsew default input
rlabel metal1 s 564286 1020000 564338 1020260 6 mprj_io_analog_en[15]
port 71 nsew default input
rlabel metal1 s 469086 1020000 469138 1020260 6 mprj_io_analog_en[16]
port 72 nsew default input
rlabel metal1 s 421086 1020000 421138 1020260 6 mprj_io_analog_en[17]
port 73 nsew default input
rlabel metal1 s 372886 1020000 372938 1020260 6 mprj_io_analog_en[18]
port 74 nsew default input
rlabel metal1 s 277686 1020000 277738 1020260 6 mprj_io_analog_en[19]
port 75 nsew default input
rlabel metal1 s 600000 122662 600260 122714 6 mprj_io_analog_en[1]
port 76 nsew default input
rlabel metal1 s 229686 1020000 229738 1020260 6 mprj_io_analog_en[20]
port 77 nsew default input
rlabel metal1 s 181486 1020000 181538 1020260 6 mprj_io_analog_en[21]
port 78 nsew default input
rlabel metal1 s 133486 1020000 133538 1020260 6 mprj_io_analog_en[22]
port 79 nsew default input
rlabel metal1 s 85286 1020000 85338 1020260 6 mprj_io_analog_en[23]
port 80 nsew default input
rlabel metal1 s 39739 986886 39999 986938 6 mprj_io_analog_en[24]
port 81 nsew default input
rlabel metal1 s 39739 807686 39999 807738 6 mprj_io_analog_en[25]
port 82 nsew default input
rlabel metal1 s 39739 762086 39999 762138 6 mprj_io_analog_en[26]
port 83 nsew default input
rlabel metal1 s 39739 716486 39999 716538 6 mprj_io_analog_en[27]
port 84 nsew default input
rlabel metal1 s 39739 670886 39999 670938 6 mprj_io_analog_en[28]
port 85 nsew default input
rlabel metal1 s 39739 625486 39999 625538 6 mprj_io_analog_en[29]
port 86 nsew default input
rlabel metal1 s 600000 170262 600260 170314 6 mprj_io_analog_en[2]
port 87 nsew default input
rlabel metal1 s 39739 579886 39999 579938 6 mprj_io_analog_en[30]
port 88 nsew default input
rlabel metal1 s 39739 534286 39999 534338 6 mprj_io_analog_en[31]
port 89 nsew default input
rlabel metal1 s 39739 399686 39999 399738 6 mprj_io_analog_en[32]
port 90 nsew default input
rlabel metal1 s 39739 354086 39999 354138 6 mprj_io_analog_en[33]
port 91 nsew default input
rlabel metal1 s 39739 308486 39999 308538 6 mprj_io_analog_en[34]
port 92 nsew default input
rlabel metal1 s 39739 262886 39999 262938 6 mprj_io_analog_en[35]
port 93 nsew default input
rlabel metal1 s 39739 217486 39999 217538 6 mprj_io_analog_en[36]
port 94 nsew default input
rlabel metal1 s 39739 171886 39999 171938 6 mprj_io_analog_en[37]
port 95 nsew default input
rlabel metal1 s 600000 217862 600260 217914 6 mprj_io_analog_en[3]
port 96 nsew default input
rlabel metal1 s 600000 265462 600260 265514 6 mprj_io_analog_en[4]
port 97 nsew default input
rlabel metal1 s 600000 313062 600260 313114 6 mprj_io_analog_en[5]
port 98 nsew default input
rlabel metal1 s 600000 360862 600260 360914 6 mprj_io_analog_en[6]
port 99 nsew default input
rlabel metal1 s 600000 548262 600260 548314 6 mprj_io_analog_en[7]
port 100 nsew default input
rlabel metal1 s 600000 595862 600260 595914 6 mprj_io_analog_en[8]
port 101 nsew default input
rlabel metal1 s 600000 643462 600260 643514 6 mprj_io_analog_en[9]
port 102 nsew default input
rlabel metal3 s 600000 78361 607360 78427 6 mprj_io_analog_pol[0]
port 103 nsew default input
rlabel metal3 s 600000 694561 607360 694627 6 mprj_io_analog_pol[10]
port 104 nsew default input
rlabel metal3 s 600000 742161 607360 742227 6 mprj_io_analog_pol[11]
port 105 nsew default input
rlabel metal3 s 600000 789761 607360 789827 6 mprj_io_analog_pol[12]
port 106 nsew default input
rlabel metal3 s 600000 883961 607360 884027 6 mprj_io_analog_pol[13]
port 107 nsew default input
rlabel metal3 s 600000 978161 607360 978227 6 mprj_io_analog_pol[14]
port 108 nsew default input
rlabel metal3 s 560973 1020000 561039 1027360 6 mprj_io_analog_pol[15]
port 109 nsew default input
rlabel metal3 s 465773 1020000 465839 1027360 6 mprj_io_analog_pol[16]
port 110 nsew default input
rlabel metal3 s 417773 1020000 417839 1027360 6 mprj_io_analog_pol[17]
port 111 nsew default input
rlabel metal3 s 369573 1020000 369639 1027360 6 mprj_io_analog_pol[18]
port 112 nsew default input
rlabel metal3 s 274373 1020000 274439 1027360 6 mprj_io_analog_pol[19]
port 113 nsew default input
rlabel metal3 s 600000 125961 607360 126027 6 mprj_io_analog_pol[1]
port 114 nsew default input
rlabel metal3 s 226373 1020000 226439 1027360 6 mprj_io_analog_pol[20]
port 115 nsew default input
rlabel metal3 s 178173 1020000 178239 1027360 6 mprj_io_analog_pol[21]
port 116 nsew default input
rlabel metal3 s 130173 1020000 130239 1027360 6 mprj_io_analog_pol[22]
port 117 nsew default input
rlabel metal3 s 81973 1020000 82039 1027360 6 mprj_io_analog_pol[23]
port 118 nsew default input
rlabel metal3 s 32639 983573 39999 983639 6 mprj_io_analog_pol[24]
port 119 nsew default input
rlabel metal3 s 32639 804373 39999 804439 6 mprj_io_analog_pol[25]
port 120 nsew default input
rlabel metal3 s 32639 758773 39999 758839 6 mprj_io_analog_pol[26]
port 121 nsew default input
rlabel metal3 s 32639 713173 39999 713239 6 mprj_io_analog_pol[27]
port 122 nsew default input
rlabel metal3 s 32639 667573 39999 667639 6 mprj_io_analog_pol[28]
port 123 nsew default input
rlabel metal3 s 32639 622173 39999 622239 6 mprj_io_analog_pol[29]
port 124 nsew default input
rlabel metal3 s 600000 173561 607360 173627 6 mprj_io_analog_pol[2]
port 125 nsew default input
rlabel metal3 s 32639 576573 39999 576639 6 mprj_io_analog_pol[30]
port 126 nsew default input
rlabel metal3 s 32639 530973 39999 531039 6 mprj_io_analog_pol[31]
port 127 nsew default input
rlabel metal3 s 32639 396373 39999 396439 6 mprj_io_analog_pol[32]
port 128 nsew default input
rlabel metal3 s 32639 350773 39999 350839 6 mprj_io_analog_pol[33]
port 129 nsew default input
rlabel metal3 s 32639 305173 39999 305239 6 mprj_io_analog_pol[34]
port 130 nsew default input
rlabel metal3 s 32639 259573 39999 259639 6 mprj_io_analog_pol[35]
port 131 nsew default input
rlabel metal3 s 32639 214173 39999 214239 6 mprj_io_analog_pol[36]
port 132 nsew default input
rlabel metal3 s 32639 168573 39999 168639 6 mprj_io_analog_pol[37]
port 133 nsew default input
rlabel metal3 s 600000 221161 607360 221227 6 mprj_io_analog_pol[3]
port 134 nsew default input
rlabel metal3 s 600000 268761 607360 268827 6 mprj_io_analog_pol[4]
port 135 nsew default input
rlabel metal3 s 600000 316361 607360 316427 6 mprj_io_analog_pol[5]
port 136 nsew default input
rlabel metal3 s 600000 364161 607360 364227 6 mprj_io_analog_pol[6]
port 137 nsew default input
rlabel metal3 s 600000 551561 607360 551627 6 mprj_io_analog_pol[7]
port 138 nsew default input
rlabel metal3 s 600000 599161 607360 599227 6 mprj_io_analog_pol[8]
port 139 nsew default input
rlabel metal3 s 600000 646761 607360 646827 6 mprj_io_analog_pol[9]
port 140 nsew default input
rlabel metal2 s 600000 81398 600452 81450 6 mprj_io_analog_sel[0]
port 141 nsew default input
rlabel metal2 s 600000 697598 600452 697650 6 mprj_io_analog_sel[10]
port 142 nsew default input
rlabel metal2 s 600000 745198 600452 745250 6 mprj_io_analog_sel[11]
port 143 nsew default input
rlabel metal2 s 600000 792798 600452 792850 6 mprj_io_analog_sel[12]
port 144 nsew default input
rlabel metal2 s 600000 886998 600452 887050 6 mprj_io_analog_sel[13]
port 145 nsew default input
rlabel metal2 s 600000 981198 600452 981250 6 mprj_io_analog_sel[14]
port 146 nsew default input
rlabel metal2 s 557950 1020000 558002 1020452 6 mprj_io_analog_sel[15]
port 147 nsew default input
rlabel metal2 s 462750 1020000 462802 1020452 6 mprj_io_analog_sel[16]
port 148 nsew default input
rlabel metal2 s 414750 1020000 414802 1020452 6 mprj_io_analog_sel[17]
port 149 nsew default input
rlabel metal2 s 366550 1020000 366602 1020452 6 mprj_io_analog_sel[18]
port 150 nsew default input
rlabel metal2 s 271350 1020000 271402 1020452 6 mprj_io_analog_sel[19]
port 151 nsew default input
rlabel metal2 s 600000 128998 600452 129050 6 mprj_io_analog_sel[1]
port 152 nsew default input
rlabel metal2 s 223350 1020000 223402 1020452 6 mprj_io_analog_sel[20]
port 153 nsew default input
rlabel metal2 s 175150 1020000 175202 1020452 6 mprj_io_analog_sel[21]
port 154 nsew default input
rlabel metal2 s 127150 1020000 127202 1020452 6 mprj_io_analog_sel[22]
port 155 nsew default input
rlabel metal2 s 78950 1020000 79002 1020452 6 mprj_io_analog_sel[23]
port 156 nsew default input
rlabel metal2 s 39547 980550 39999 980602 6 mprj_io_analog_sel[24]
port 157 nsew default input
rlabel metal2 s 39547 801350 39999 801402 6 mprj_io_analog_sel[25]
port 158 nsew default input
rlabel metal2 s 39547 755750 39999 755802 6 mprj_io_analog_sel[26]
port 159 nsew default input
rlabel metal2 s 39547 710150 39999 710202 6 mprj_io_analog_sel[27]
port 160 nsew default input
rlabel metal2 s 39547 664550 39999 664602 6 mprj_io_analog_sel[28]
port 161 nsew default input
rlabel metal2 s 39547 619150 39999 619202 6 mprj_io_analog_sel[29]
port 162 nsew default input
rlabel metal2 s 600000 176598 600452 176650 6 mprj_io_analog_sel[2]
port 163 nsew default input
rlabel metal2 s 39547 573550 39999 573602 6 mprj_io_analog_sel[30]
port 164 nsew default input
rlabel metal2 s 39547 527950 39999 528002 6 mprj_io_analog_sel[31]
port 165 nsew default input
rlabel metal2 s 39547 393350 39999 393402 6 mprj_io_analog_sel[32]
port 166 nsew default input
rlabel metal2 s 39547 347750 39999 347802 6 mprj_io_analog_sel[33]
port 167 nsew default input
rlabel metal2 s 39547 302150 39999 302202 6 mprj_io_analog_sel[34]
port 168 nsew default input
rlabel metal2 s 39547 256550 39999 256602 6 mprj_io_analog_sel[35]
port 169 nsew default input
rlabel metal2 s 39547 211150 39999 211202 6 mprj_io_analog_sel[36]
port 170 nsew default input
rlabel metal2 s 39547 165550 39999 165602 6 mprj_io_analog_sel[37]
port 171 nsew default input
rlabel metal2 s 600000 224198 600452 224250 6 mprj_io_analog_sel[3]
port 172 nsew default input
rlabel metal2 s 600000 271798 600452 271850 6 mprj_io_analog_sel[4]
port 173 nsew default input
rlabel metal2 s 600000 319398 600452 319450 6 mprj_io_analog_sel[5]
port 174 nsew default input
rlabel metal2 s 600000 367198 600452 367250 6 mprj_io_analog_sel[6]
port 175 nsew default input
rlabel metal2 s 600000 554598 600452 554650 6 mprj_io_analog_sel[7]
port 176 nsew default input
rlabel metal2 s 600000 602198 600452 602250 6 mprj_io_analog_sel[8]
port 177 nsew default input
rlabel metal2 s 600000 649798 600452 649850 6 mprj_io_analog_sel[9]
port 178 nsew default input
rlabel metal2 s 600000 77577 600108 77629 6 mprj_io_dm[0]
port 179 nsew default input
rlabel metal2 s 39761 354967 39999 355019 6 mprj_io_dm[100]
port 180 nsew default input
rlabel metal2 s 39186 347298 40000 347350 6 mprj_io_dm[101]
port 181 nsew default input
rlabel metal2 s 39891 305971 39999 306023 6 mprj_io_dm[102]
port 182 nsew default input
rlabel metal2 s 39761 309367 39999 309419 6 mprj_io_dm[103]
port 183 nsew default input
rlabel metal2 s 39186 301698 40000 301750 6 mprj_io_dm[104]
port 184 nsew default input
rlabel metal2 s 39891 260371 39999 260423 6 mprj_io_dm[105]
port 185 nsew default input
rlabel metal2 s 39761 263767 39999 263819 6 mprj_io_dm[106]
port 186 nsew default input
rlabel metal2 s 39186 256098 40000 256150 6 mprj_io_dm[107]
port 187 nsew default input
rlabel metal2 s 39891 214971 39999 215023 6 mprj_io_dm[108]
port 188 nsew default input
rlabel metal2 s 39761 218367 39999 218419 6 mprj_io_dm[109]
port 189 nsew default input
rlabel metal2 s 600000 216981 600238 217033 6 mprj_io_dm[10]
port 190 nsew default input
rlabel metal2 s 39186 210698 40000 210750 6 mprj_io_dm[110]
port 191 nsew default input
rlabel metal2 s 39891 169371 39999 169423 6 mprj_io_dm[111]
port 192 nsew default input
rlabel metal2 s 39761 172767 39999 172819 6 mprj_io_dm[112]
port 193 nsew default input
rlabel metal2 s 39186 165098 40000 165150 6 mprj_io_dm[113]
port 194 nsew default input
rlabel metal2 s 600000 224650 600814 224702 6 mprj_io_dm[11]
port 195 nsew default input
rlabel metal2 s 600000 267977 600108 268029 6 mprj_io_dm[12]
port 196 nsew default input
rlabel metal2 s 600000 264581 600238 264633 6 mprj_io_dm[13]
port 197 nsew default input
rlabel metal2 s 600000 272250 600814 272302 6 mprj_io_dm[14]
port 198 nsew default input
rlabel metal2 s 600000 315577 600108 315629 6 mprj_io_dm[15]
port 199 nsew default input
rlabel metal2 s 600000 312181 600238 312233 6 mprj_io_dm[16]
port 200 nsew default input
rlabel metal2 s 600000 319850 600814 319902 6 mprj_io_dm[17]
port 201 nsew default input
rlabel metal2 s 600000 363377 600108 363429 6 mprj_io_dm[18]
port 202 nsew default input
rlabel metal2 s 600000 359981 600238 360033 6 mprj_io_dm[19]
port 203 nsew default input
rlabel metal2 s 600000 74181 600238 74233 6 mprj_io_dm[1]
port 204 nsew default input
rlabel metal2 s 600000 367650 600814 367702 6 mprj_io_dm[20]
port 205 nsew default input
rlabel metal2 s 600000 550777 600108 550829 6 mprj_io_dm[21]
port 206 nsew default input
rlabel metal2 s 600000 547381 600238 547433 6 mprj_io_dm[22]
port 207 nsew default input
rlabel metal2 s 600000 555050 600814 555102 6 mprj_io_dm[23]
port 208 nsew default input
rlabel metal2 s 600000 598377 600108 598429 6 mprj_io_dm[24]
port 209 nsew default input
rlabel metal2 s 600000 594981 600238 595033 6 mprj_io_dm[25]
port 210 nsew default input
rlabel metal2 s 600000 602650 600814 602702 6 mprj_io_dm[26]
port 211 nsew default input
rlabel metal2 s 600000 645977 600108 646029 6 mprj_io_dm[27]
port 212 nsew default input
rlabel metal2 s 600000 642581 600238 642633 6 mprj_io_dm[28]
port 213 nsew default input
rlabel metal2 s 600000 650250 600814 650302 6 mprj_io_dm[29]
port 214 nsew default input
rlabel metal2 s 600000 81850 600814 81902 6 mprj_io_dm[2]
port 215 nsew default input
rlabel metal2 s 600000 693777 600108 693829 6 mprj_io_dm[30]
port 216 nsew default input
rlabel metal2 s 600000 690381 600238 690433 6 mprj_io_dm[31]
port 217 nsew default input
rlabel metal2 s 600000 698050 600814 698102 6 mprj_io_dm[32]
port 218 nsew default input
rlabel metal2 s 600000 741377 600108 741429 6 mprj_io_dm[33]
port 219 nsew default input
rlabel metal2 s 600000 737981 600238 738033 6 mprj_io_dm[34]
port 220 nsew default input
rlabel metal2 s 600000 745650 600814 745702 6 mprj_io_dm[35]
port 221 nsew default input
rlabel metal2 s 600000 788977 600108 789029 6 mprj_io_dm[36]
port 222 nsew default input
rlabel metal2 s 600000 785581 600238 785633 6 mprj_io_dm[37]
port 223 nsew default input
rlabel metal2 s 600000 793250 600814 793302 6 mprj_io_dm[38]
port 224 nsew default input
rlabel metal2 s 600000 883177 600108 883229 6 mprj_io_dm[39]
port 225 nsew default input
rlabel metal2 s 600000 125177 600108 125229 6 mprj_io_dm[3]
port 226 nsew default input
rlabel metal2 s 600000 879781 600238 879833 6 mprj_io_dm[40]
port 227 nsew default input
rlabel metal2 s 600000 887450 600814 887502 6 mprj_io_dm[41]
port 228 nsew default input
rlabel metal2 s 600000 977377 600108 977429 6 mprj_io_dm[42]
port 229 nsew default input
rlabel metal2 s 600000 973981 600238 974033 6 mprj_io_dm[43]
port 230 nsew default input
rlabel metal2 s 600000 981650 600814 981702 6 mprj_io_dm[44]
port 231 nsew default input
rlabel metal2 s 561771 1020000 561823 1020108 6 mprj_io_dm[45]
port 232 nsew default input
rlabel metal2 s 565167 1020000 565219 1020238 6 mprj_io_dm[46]
port 233 nsew default input
rlabel metal2 s 557498 1020000 557550 1020814 6 mprj_io_dm[47]
port 234 nsew default input
rlabel metal2 s 466571 1020000 466623 1020108 6 mprj_io_dm[48]
port 235 nsew default input
rlabel metal2 s 469967 1020000 470019 1020238 6 mprj_io_dm[49]
port 236 nsew default input
rlabel metal2 s 600000 121781 600238 121833 6 mprj_io_dm[4]
port 237 nsew default input
rlabel metal2 s 462298 1020000 462350 1020814 6 mprj_io_dm[50]
port 238 nsew default input
rlabel metal2 s 418571 1020000 418623 1020108 6 mprj_io_dm[51]
port 239 nsew default input
rlabel metal2 s 421967 1020000 422019 1020238 6 mprj_io_dm[52]
port 240 nsew default input
rlabel metal2 s 414298 1020000 414350 1020814 6 mprj_io_dm[53]
port 241 nsew default input
rlabel metal2 s 370371 1020000 370423 1020108 6 mprj_io_dm[54]
port 242 nsew default input
rlabel metal2 s 373767 1020000 373819 1020238 6 mprj_io_dm[55]
port 243 nsew default input
rlabel metal2 s 366098 1020000 366150 1020814 6 mprj_io_dm[56]
port 244 nsew default input
rlabel metal2 s 275171 1020000 275223 1020108 6 mprj_io_dm[57]
port 245 nsew default input
rlabel metal2 s 278567 1020000 278619 1020238 6 mprj_io_dm[58]
port 246 nsew default input
rlabel metal2 s 270898 1020000 270950 1020814 6 mprj_io_dm[59]
port 247 nsew default input
rlabel metal2 s 600000 129450 600814 129502 6 mprj_io_dm[5]
port 248 nsew default input
rlabel metal2 s 227171 1020000 227223 1020108 6 mprj_io_dm[60]
port 249 nsew default input
rlabel metal2 s 230567 1020000 230619 1020238 6 mprj_io_dm[61]
port 250 nsew default input
rlabel metal2 s 222898 1020000 222950 1020814 6 mprj_io_dm[62]
port 251 nsew default input
rlabel metal2 s 178971 1020000 179023 1020108 6 mprj_io_dm[63]
port 252 nsew default input
rlabel metal2 s 182367 1020000 182419 1020238 6 mprj_io_dm[64]
port 253 nsew default input
rlabel metal2 s 174698 1020000 174750 1020814 6 mprj_io_dm[65]
port 254 nsew default input
rlabel metal2 s 130971 1020000 131023 1020108 6 mprj_io_dm[66]
port 255 nsew default input
rlabel metal2 s 134367 1020000 134419 1020238 6 mprj_io_dm[67]
port 256 nsew default input
rlabel metal2 s 126698 1020000 126750 1020814 6 mprj_io_dm[68]
port 257 nsew default input
rlabel metal2 s 82771 1020000 82823 1020108 6 mprj_io_dm[69]
port 258 nsew default input
rlabel metal2 s 600000 172777 600108 172829 6 mprj_io_dm[6]
port 259 nsew default input
rlabel metal2 s 86167 1020000 86219 1020238 6 mprj_io_dm[70]
port 260 nsew default input
rlabel metal2 s 78498 1020000 78550 1020814 6 mprj_io_dm[71]
port 261 nsew default input
rlabel metal2 s 39891 984371 39999 984423 6 mprj_io_dm[72]
port 262 nsew default input
rlabel metal2 s 39761 987767 39999 987819 6 mprj_io_dm[73]
port 263 nsew default input
rlabel metal2 s 39186 980098 40000 980150 6 mprj_io_dm[74]
port 264 nsew default input
rlabel metal2 s 39891 805171 39999 805223 6 mprj_io_dm[75]
port 265 nsew default input
rlabel metal2 s 39761 808567 39999 808619 6 mprj_io_dm[76]
port 266 nsew default input
rlabel metal2 s 39186 800898 40000 800950 6 mprj_io_dm[77]
port 267 nsew default input
rlabel metal2 s 39891 759571 39999 759623 6 mprj_io_dm[78]
port 268 nsew default input
rlabel metal2 s 39761 762967 39999 763019 6 mprj_io_dm[79]
port 269 nsew default input
rlabel metal2 s 600000 169381 600238 169433 6 mprj_io_dm[7]
port 270 nsew default input
rlabel metal2 s 39186 755298 40000 755350 6 mprj_io_dm[80]
port 271 nsew default input
rlabel metal2 s 39891 713971 39999 714023 6 mprj_io_dm[81]
port 272 nsew default input
rlabel metal2 s 39761 717367 39999 717419 6 mprj_io_dm[82]
port 273 nsew default input
rlabel metal2 s 39186 709698 40000 709750 6 mprj_io_dm[83]
port 274 nsew default input
rlabel metal2 s 39891 668371 39999 668423 6 mprj_io_dm[84]
port 275 nsew default input
rlabel metal2 s 39761 671767 39999 671819 6 mprj_io_dm[85]
port 276 nsew default input
rlabel metal2 s 39186 664098 40000 664150 6 mprj_io_dm[86]
port 277 nsew default input
rlabel metal2 s 39891 622971 39999 623023 6 mprj_io_dm[87]
port 278 nsew default input
rlabel metal2 s 39761 626367 39999 626419 6 mprj_io_dm[88]
port 279 nsew default input
rlabel metal2 s 39186 618698 40000 618750 6 mprj_io_dm[89]
port 280 nsew default input
rlabel metal2 s 600000 177050 600814 177102 6 mprj_io_dm[8]
port 281 nsew default input
rlabel metal2 s 39891 577371 39999 577423 6 mprj_io_dm[90]
port 282 nsew default input
rlabel metal2 s 39761 580767 39999 580819 6 mprj_io_dm[91]
port 283 nsew default input
rlabel metal2 s 39186 573098 40000 573150 6 mprj_io_dm[92]
port 284 nsew default input
rlabel metal2 s 39891 531771 39999 531823 6 mprj_io_dm[93]
port 285 nsew default input
rlabel metal2 s 39761 535167 39999 535219 6 mprj_io_dm[94]
port 286 nsew default input
rlabel metal2 s 39186 527498 40000 527550 6 mprj_io_dm[95]
port 287 nsew default input
rlabel metal2 s 39891 397171 39999 397223 6 mprj_io_dm[96]
port 288 nsew default input
rlabel metal2 s 39761 400567 39999 400619 6 mprj_io_dm[97]
port 289 nsew default input
rlabel metal2 s 39186 392898 40000 392950 6 mprj_io_dm[98]
port 290 nsew default input
rlabel metal2 s 39891 351571 39999 351623 6 mprj_io_dm[99]
port 291 nsew default input
rlabel metal2 s 600000 220377 600108 220429 6 mprj_io_dm[9]
port 292 nsew default input
rlabel metal2 s 600000 80456 600310 80508 6 mprj_io_enh[0]
port 293 nsew default input
rlabel metal2 s 600000 696656 600310 696708 6 mprj_io_enh[10]
port 294 nsew default input
rlabel metal2 s 600000 744256 600310 744308 6 mprj_io_enh[11]
port 295 nsew default input
rlabel metal2 s 600000 791856 600310 791908 6 mprj_io_enh[12]
port 296 nsew default input
rlabel metal2 s 600000 886056 600310 886108 6 mprj_io_enh[13]
port 297 nsew default input
rlabel metal2 s 600000 980256 600310 980308 6 mprj_io_enh[14]
port 298 nsew default input
rlabel metal2 s 558892 1020000 558944 1020310 6 mprj_io_enh[15]
port 299 nsew default input
rlabel metal2 s 463692 1020000 463744 1020310 6 mprj_io_enh[16]
port 300 nsew default input
rlabel metal2 s 415692 1020000 415744 1020310 6 mprj_io_enh[17]
port 301 nsew default input
rlabel metal2 s 367492 1020000 367544 1020310 6 mprj_io_enh[18]
port 302 nsew default input
rlabel metal2 s 272292 1020000 272344 1020310 6 mprj_io_enh[19]
port 303 nsew default input
rlabel metal2 s 600000 128056 600310 128108 6 mprj_io_enh[1]
port 304 nsew default input
rlabel metal2 s 224292 1020000 224344 1020310 6 mprj_io_enh[20]
port 305 nsew default input
rlabel metal2 s 176092 1020000 176144 1020310 6 mprj_io_enh[21]
port 306 nsew default input
rlabel metal2 s 128092 1020000 128144 1020310 6 mprj_io_enh[22]
port 307 nsew default input
rlabel metal2 s 79892 1020000 79944 1020310 6 mprj_io_enh[23]
port 308 nsew default input
rlabel metal2 s 39690 981492 40000 981544 6 mprj_io_enh[24]
port 309 nsew default input
rlabel metal2 s 39690 802292 40000 802344 6 mprj_io_enh[25]
port 310 nsew default input
rlabel metal2 s 39690 756692 40000 756744 6 mprj_io_enh[26]
port 311 nsew default input
rlabel metal2 s 39690 711092 40000 711144 6 mprj_io_enh[27]
port 312 nsew default input
rlabel metal2 s 39690 665492 40000 665544 6 mprj_io_enh[28]
port 313 nsew default input
rlabel metal2 s 39690 620092 40000 620144 6 mprj_io_enh[29]
port 314 nsew default input
rlabel metal2 s 600000 175656 600310 175708 6 mprj_io_enh[2]
port 315 nsew default input
rlabel metal2 s 39690 574492 40000 574544 6 mprj_io_enh[30]
port 316 nsew default input
rlabel metal2 s 39690 528892 40000 528944 6 mprj_io_enh[31]
port 317 nsew default input
rlabel metal2 s 39690 394292 40000 394344 6 mprj_io_enh[32]
port 318 nsew default input
rlabel metal2 s 39690 348692 40000 348744 6 mprj_io_enh[33]
port 319 nsew default input
rlabel metal2 s 39690 303092 40000 303144 6 mprj_io_enh[34]
port 320 nsew default input
rlabel metal2 s 39690 257492 40000 257544 6 mprj_io_enh[35]
port 321 nsew default input
rlabel metal2 s 39690 212092 40000 212144 6 mprj_io_enh[36]
port 322 nsew default input
rlabel metal2 s 39690 166492 40000 166544 6 mprj_io_enh[37]
port 323 nsew default input
rlabel metal2 s 600000 223256 600310 223308 6 mprj_io_enh[3]
port 324 nsew default input
rlabel metal2 s 600000 270856 600310 270908 6 mprj_io_enh[4]
port 325 nsew default input
rlabel metal2 s 600000 318456 600310 318508 6 mprj_io_enh[5]
port 326 nsew default input
rlabel metal2 s 600000 366256 600310 366308 6 mprj_io_enh[6]
port 327 nsew default input
rlabel metal2 s 600000 553656 600310 553708 6 mprj_io_enh[7]
port 328 nsew default input
rlabel metal2 s 600000 601256 600310 601308 6 mprj_io_enh[8]
port 329 nsew default input
rlabel metal2 s 600000 648856 600310 648908 6 mprj_io_enh[9]
port 330 nsew default input
rlabel metal2 s 600000 81185 600668 81237 6 mprj_io_hldh_n[0]
port 331 nsew default input
rlabel metal2 s 600000 697385 600668 697437 6 mprj_io_hldh_n[10]
port 332 nsew default input
rlabel metal2 s 600000 744985 600668 745037 6 mprj_io_hldh_n[11]
port 333 nsew default input
rlabel metal2 s 600000 792585 600668 792637 6 mprj_io_hldh_n[12]
port 334 nsew default input
rlabel metal2 s 600000 886785 600668 886837 6 mprj_io_hldh_n[13]
port 335 nsew default input
rlabel metal2 s 600000 980985 600668 981037 6 mprj_io_hldh_n[14]
port 336 nsew default input
rlabel metal2 s 558163 1020000 558215 1020668 6 mprj_io_hldh_n[15]
port 337 nsew default input
rlabel metal2 s 462963 1020000 463015 1020668 6 mprj_io_hldh_n[16]
port 338 nsew default input
rlabel metal2 s 414963 1020000 415015 1020668 6 mprj_io_hldh_n[17]
port 339 nsew default input
rlabel metal2 s 366763 1020000 366815 1020668 6 mprj_io_hldh_n[18]
port 340 nsew default input
rlabel metal2 s 271563 1020000 271615 1020668 6 mprj_io_hldh_n[19]
port 341 nsew default input
rlabel metal2 s 600000 128785 600668 128837 6 mprj_io_hldh_n[1]
port 342 nsew default input
rlabel metal2 s 223563 1020000 223615 1020668 6 mprj_io_hldh_n[20]
port 343 nsew default input
rlabel metal2 s 175363 1020000 175415 1020668 6 mprj_io_hldh_n[21]
port 344 nsew default input
rlabel metal2 s 127363 1020000 127415 1020668 6 mprj_io_hldh_n[22]
port 345 nsew default input
rlabel metal2 s 79163 1020000 79215 1020668 6 mprj_io_hldh_n[23]
port 346 nsew default input
rlabel metal2 s 39332 980763 40000 980815 6 mprj_io_hldh_n[24]
port 347 nsew default input
rlabel metal2 s 39332 801563 40000 801615 6 mprj_io_hldh_n[25]
port 348 nsew default input
rlabel metal2 s 39332 755963 40000 756015 6 mprj_io_hldh_n[26]
port 349 nsew default input
rlabel metal2 s 39332 710363 40000 710415 6 mprj_io_hldh_n[27]
port 350 nsew default input
rlabel metal2 s 39332 664763 40000 664815 6 mprj_io_hldh_n[28]
port 351 nsew default input
rlabel metal2 s 39332 619363 40000 619415 6 mprj_io_hldh_n[29]
port 352 nsew default input
rlabel metal2 s 600000 176385 600668 176437 6 mprj_io_hldh_n[2]
port 353 nsew default input
rlabel metal2 s 39332 573763 40000 573815 6 mprj_io_hldh_n[30]
port 354 nsew default input
rlabel metal2 s 39332 528163 40000 528215 6 mprj_io_hldh_n[31]
port 355 nsew default input
rlabel metal2 s 39332 393563 40000 393615 6 mprj_io_hldh_n[32]
port 356 nsew default input
rlabel metal2 s 39332 347963 40000 348015 6 mprj_io_hldh_n[33]
port 357 nsew default input
rlabel metal2 s 39332 302363 40000 302415 6 mprj_io_hldh_n[34]
port 358 nsew default input
rlabel metal2 s 39332 256763 40000 256815 6 mprj_io_hldh_n[35]
port 359 nsew default input
rlabel metal2 s 39332 211363 40000 211415 6 mprj_io_hldh_n[36]
port 360 nsew default input
rlabel metal2 s 39332 165763 40000 165815 6 mprj_io_hldh_n[37]
port 361 nsew default input
rlabel metal2 s 600000 223985 600668 224037 6 mprj_io_hldh_n[3]
port 362 nsew default input
rlabel metal2 s 600000 271585 600668 271637 6 mprj_io_hldh_n[4]
port 363 nsew default input
rlabel metal2 s 600000 319185 600668 319237 6 mprj_io_hldh_n[5]
port 364 nsew default input
rlabel metal2 s 600000 366985 600668 367037 6 mprj_io_hldh_n[6]
port 365 nsew default input
rlabel metal2 s 600000 554385 600668 554437 6 mprj_io_hldh_n[7]
port 366 nsew default input
rlabel metal2 s 600000 601985 600668 602037 6 mprj_io_hldh_n[8]
port 367 nsew default input
rlabel metal2 s 600000 649585 600668 649637 6 mprj_io_hldh_n[9]
port 368 nsew default input
rlabel metal2 s 600000 82228 600540 82280 6 mprj_io_holdover[0]
port 369 nsew default input
rlabel metal2 s 600000 698428 600540 698480 6 mprj_io_holdover[10]
port 370 nsew default input
rlabel metal2 s 600000 746028 600540 746080 6 mprj_io_holdover[11]
port 371 nsew default input
rlabel metal2 s 600000 793628 600540 793680 6 mprj_io_holdover[12]
port 372 nsew default input
rlabel metal2 s 600000 887828 600540 887880 6 mprj_io_holdover[13]
port 373 nsew default input
rlabel metal2 s 600000 982028 600540 982080 6 mprj_io_holdover[14]
port 374 nsew default input
rlabel metal2 s 557120 1020000 557172 1020540 6 mprj_io_holdover[15]
port 375 nsew default input
rlabel metal2 s 461920 1020000 461972 1020540 6 mprj_io_holdover[16]
port 376 nsew default input
rlabel metal2 s 413920 1020000 413972 1020540 6 mprj_io_holdover[17]
port 377 nsew default input
rlabel metal2 s 365720 1020000 365772 1020540 6 mprj_io_holdover[18]
port 378 nsew default input
rlabel metal2 s 270520 1020000 270572 1020540 6 mprj_io_holdover[19]
port 379 nsew default input
rlabel metal2 s 600000 129828 600540 129880 6 mprj_io_holdover[1]
port 380 nsew default input
rlabel metal2 s 222520 1020000 222572 1020540 6 mprj_io_holdover[20]
port 381 nsew default input
rlabel metal2 s 174320 1020000 174372 1020540 6 mprj_io_holdover[21]
port 382 nsew default input
rlabel metal2 s 126320 1020000 126372 1020540 6 mprj_io_holdover[22]
port 383 nsew default input
rlabel metal2 s 78120 1020000 78172 1020540 6 mprj_io_holdover[23]
port 384 nsew default input
rlabel metal2 s 39459 979720 39999 979772 6 mprj_io_holdover[24]
port 385 nsew default input
rlabel metal2 s 39459 800520 39999 800572 6 mprj_io_holdover[25]
port 386 nsew default input
rlabel metal2 s 39459 754920 39999 754972 6 mprj_io_holdover[26]
port 387 nsew default input
rlabel metal2 s 39459 709320 39999 709372 6 mprj_io_holdover[27]
port 388 nsew default input
rlabel metal2 s 39459 663720 39999 663772 6 mprj_io_holdover[28]
port 389 nsew default input
rlabel metal2 s 39459 618320 39999 618372 6 mprj_io_holdover[29]
port 390 nsew default input
rlabel metal2 s 600000 177428 600540 177480 6 mprj_io_holdover[2]
port 391 nsew default input
rlabel metal2 s 39459 572720 39999 572772 6 mprj_io_holdover[30]
port 392 nsew default input
rlabel metal2 s 39459 527120 39999 527172 6 mprj_io_holdover[31]
port 393 nsew default input
rlabel metal2 s 39459 392520 39999 392572 6 mprj_io_holdover[32]
port 394 nsew default input
rlabel metal2 s 39459 346920 39999 346972 6 mprj_io_holdover[33]
port 395 nsew default input
rlabel metal2 s 39459 301320 39999 301372 6 mprj_io_holdover[34]
port 396 nsew default input
rlabel metal2 s 39459 255720 39999 255772 6 mprj_io_holdover[35]
port 397 nsew default input
rlabel metal2 s 39459 210320 39999 210372 6 mprj_io_holdover[36]
port 398 nsew default input
rlabel metal2 s 39459 164720 39999 164772 6 mprj_io_holdover[37]
port 399 nsew default input
rlabel metal2 s 600000 225028 600540 225080 6 mprj_io_holdover[3]
port 400 nsew default input
rlabel metal2 s 600000 272628 600540 272680 6 mprj_io_holdover[4]
port 401 nsew default input
rlabel metal2 s 600000 320228 600540 320280 6 mprj_io_holdover[5]
port 402 nsew default input
rlabel metal2 s 600000 368028 600540 368080 6 mprj_io_holdover[6]
port 403 nsew default input
rlabel metal2 s 600000 555428 600540 555480 6 mprj_io_holdover[7]
port 404 nsew default input
rlabel metal2 s 600000 603028 600540 603080 6 mprj_io_holdover[8]
port 405 nsew default input
rlabel metal2 s 600000 650628 600540 650680 6 mprj_io_holdover[9]
port 406 nsew default input
rlabel metal2 s 600000 86470 600894 86516 6 mprj_io_ib_mode_sel[0]
port 407 nsew default input
rlabel metal2 s 600000 702670 600894 702716 6 mprj_io_ib_mode_sel[10]
port 408 nsew default input
rlabel metal2 s 600000 750270 600894 750316 6 mprj_io_ib_mode_sel[11]
port 409 nsew default input
rlabel metal2 s 600000 797870 600894 797916 6 mprj_io_ib_mode_sel[12]
port 410 nsew default input
rlabel metal2 s 600000 892070 600894 892116 6 mprj_io_ib_mode_sel[13]
port 411 nsew default input
rlabel metal2 s 600000 986270 600894 986316 6 mprj_io_ib_mode_sel[14]
port 412 nsew default input
rlabel metal2 s 552884 1020000 552930 1020894 6 mprj_io_ib_mode_sel[15]
port 413 nsew default input
rlabel metal2 s 457684 1020000 457730 1020894 6 mprj_io_ib_mode_sel[16]
port 414 nsew default input
rlabel metal2 s 409684 1020000 409730 1020894 6 mprj_io_ib_mode_sel[17]
port 415 nsew default input
rlabel metal2 s 361484 1020000 361530 1020894 6 mprj_io_ib_mode_sel[18]
port 416 nsew default input
rlabel metal2 s 266284 1020000 266330 1020894 6 mprj_io_ib_mode_sel[19]
port 417 nsew default input
rlabel metal2 s 600000 134070 600894 134116 6 mprj_io_ib_mode_sel[1]
port 418 nsew default input
rlabel metal2 s 218284 1020000 218330 1020894 6 mprj_io_ib_mode_sel[20]
port 419 nsew default input
rlabel metal2 s 170084 1020000 170130 1020894 6 mprj_io_ib_mode_sel[21]
port 420 nsew default input
rlabel metal2 s 122084 1020000 122130 1020894 6 mprj_io_ib_mode_sel[22]
port 421 nsew default input
rlabel metal2 s 73884 1020000 73930 1020894 6 mprj_io_ib_mode_sel[23]
port 422 nsew default input
rlabel metal2 s 39105 975484 39999 975530 6 mprj_io_ib_mode_sel[24]
port 423 nsew default input
rlabel metal2 s 39105 796284 39999 796330 6 mprj_io_ib_mode_sel[25]
port 424 nsew default input
rlabel metal2 s 39105 750684 39999 750730 6 mprj_io_ib_mode_sel[26]
port 425 nsew default input
rlabel metal2 s 39105 705084 39999 705130 6 mprj_io_ib_mode_sel[27]
port 426 nsew default input
rlabel metal2 s 39105 659484 39999 659530 6 mprj_io_ib_mode_sel[28]
port 427 nsew default input
rlabel metal2 s 39105 614084 39999 614130 6 mprj_io_ib_mode_sel[29]
port 428 nsew default input
rlabel metal2 s 600000 181670 600894 181716 6 mprj_io_ib_mode_sel[2]
port 429 nsew default input
rlabel metal2 s 39105 568484 39999 568530 6 mprj_io_ib_mode_sel[30]
port 430 nsew default input
rlabel metal2 s 39105 522884 39999 522930 6 mprj_io_ib_mode_sel[31]
port 431 nsew default input
rlabel metal2 s 39105 388284 39999 388330 6 mprj_io_ib_mode_sel[32]
port 432 nsew default input
rlabel metal2 s 39105 342684 39999 342730 6 mprj_io_ib_mode_sel[33]
port 433 nsew default input
rlabel metal2 s 39105 297084 39999 297130 6 mprj_io_ib_mode_sel[34]
port 434 nsew default input
rlabel metal2 s 39105 251484 39999 251530 6 mprj_io_ib_mode_sel[35]
port 435 nsew default input
rlabel metal2 s 39105 206084 39999 206130 6 mprj_io_ib_mode_sel[36]
port 436 nsew default input
rlabel metal2 s 39105 160484 39999 160530 6 mprj_io_ib_mode_sel[37]
port 437 nsew default input
rlabel metal2 s 600000 229270 600894 229316 6 mprj_io_ib_mode_sel[3]
port 438 nsew default input
rlabel metal2 s 600000 276870 600894 276916 6 mprj_io_ib_mode_sel[4]
port 439 nsew default input
rlabel metal2 s 600000 324470 600894 324516 6 mprj_io_ib_mode_sel[5]
port 440 nsew default input
rlabel metal2 s 600000 372270 600894 372316 6 mprj_io_ib_mode_sel[6]
port 441 nsew default input
rlabel metal2 s 600000 559670 600894 559716 6 mprj_io_ib_mode_sel[7]
port 442 nsew default input
rlabel metal2 s 600000 607270 600894 607316 6 mprj_io_ib_mode_sel[8]
port 443 nsew default input
rlabel metal2 s 600000 654870 600894 654916 6 mprj_io_ib_mode_sel[9]
port 444 nsew default input
rlabel metal3 s 600000 71686 637912 71752 6 mprj_io_in[0]
port 445 nsew default tristate
rlabel metal3 s 600000 687886 637912 687952 6 mprj_io_in[10]
port 446 nsew default tristate
rlabel metal3 s 600000 735486 637912 735552 6 mprj_io_in[11]
port 447 nsew default tristate
rlabel metal3 s 600000 783086 637912 783152 6 mprj_io_in[12]
port 448 nsew default tristate
rlabel metal3 s 600000 877286 637912 877352 6 mprj_io_in[13]
port 449 nsew default tristate
rlabel metal3 s 600000 971486 637912 971552 6 mprj_io_in[14]
port 450 nsew default tristate
rlabel metal3 s 567648 1020000 567714 1057912 6 mprj_io_in[15]
port 451 nsew default tristate
rlabel metal3 s 472448 1020000 472514 1057912 6 mprj_io_in[16]
port 452 nsew default tristate
rlabel metal3 s 424448 1020000 424514 1057912 6 mprj_io_in[17]
port 453 nsew default tristate
rlabel metal3 s 376248 1020000 376314 1057912 6 mprj_io_in[18]
port 454 nsew default tristate
rlabel metal3 s 281048 1020000 281114 1057912 6 mprj_io_in[19]
port 455 nsew default tristate
rlabel metal3 s 600000 119286 637912 119352 6 mprj_io_in[1]
port 456 nsew default tristate
rlabel metal3 s 233048 1020000 233114 1057912 6 mprj_io_in[20]
port 457 nsew default tristate
rlabel metal3 s 184848 1020000 184914 1057912 6 mprj_io_in[21]
port 458 nsew default tristate
rlabel metal3 s 136848 1020000 136914 1057912 6 mprj_io_in[22]
port 459 nsew default tristate
rlabel metal3 s 88648 1020000 88714 1057912 6 mprj_io_in[23]
port 460 nsew default tristate
rlabel metal3 s 2088 990248 40000 990314 6 mprj_io_in[24]
port 461 nsew default tristate
rlabel metal3 s 2088 811048 40000 811114 6 mprj_io_in[25]
port 462 nsew default tristate
rlabel metal3 s 2088 765448 40000 765514 6 mprj_io_in[26]
port 463 nsew default tristate
rlabel metal3 s 2088 719848 40000 719914 6 mprj_io_in[27]
port 464 nsew default tristate
rlabel metal3 s 2088 674248 40000 674314 6 mprj_io_in[28]
port 465 nsew default tristate
rlabel metal3 s 2088 628848 40000 628914 6 mprj_io_in[29]
port 466 nsew default tristate
rlabel metal3 s 600000 166886 637912 166952 6 mprj_io_in[2]
port 467 nsew default tristate
rlabel metal3 s 2088 583248 40000 583314 6 mprj_io_in[30]
port 468 nsew default tristate
rlabel metal3 s 2088 537648 40000 537714 6 mprj_io_in[31]
port 469 nsew default tristate
rlabel metal3 s 2088 403048 40000 403114 6 mprj_io_in[32]
port 470 nsew default tristate
rlabel metal3 s 2088 357448 40000 357514 6 mprj_io_in[33]
port 471 nsew default tristate
rlabel metal3 s 2088 311848 40000 311914 6 mprj_io_in[34]
port 472 nsew default tristate
rlabel metal3 s 2088 266248 40000 266314 6 mprj_io_in[35]
port 473 nsew default tristate
rlabel metal3 s 2088 220848 40000 220914 6 mprj_io_in[36]
port 474 nsew default tristate
rlabel metal3 s 2088 175248 40000 175314 6 mprj_io_in[37]
port 475 nsew default tristate
rlabel metal3 s 600000 214486 637912 214552 6 mprj_io_in[3]
port 476 nsew default tristate
rlabel metal3 s 600000 262086 637912 262152 6 mprj_io_in[4]
port 477 nsew default tristate
rlabel metal3 s 600000 309686 637912 309752 6 mprj_io_in[5]
port 478 nsew default tristate
rlabel metal3 s 600000 357486 637912 357552 6 mprj_io_in[6]
port 479 nsew default tristate
rlabel metal3 s 600000 544886 637912 544952 6 mprj_io_in[7]
port 480 nsew default tristate
rlabel metal3 s 600000 592486 637912 592552 6 mprj_io_in[8]
port 481 nsew default tristate
rlabel metal3 s 600000 640086 637912 640152 6 mprj_io_in[9]
port 482 nsew default tristate
rlabel metal2 s 600000 78499 601018 78551 6 mprj_io_inp_dis[0]
port 483 nsew default input
rlabel metal2 s 600000 694699 601018 694751 6 mprj_io_inp_dis[10]
port 484 nsew default input
rlabel metal2 s 600000 742299 601018 742351 6 mprj_io_inp_dis[11]
port 485 nsew default input
rlabel metal2 s 600000 789899 601018 789951 6 mprj_io_inp_dis[12]
port 486 nsew default input
rlabel metal2 s 600000 884099 601018 884151 6 mprj_io_inp_dis[13]
port 487 nsew default input
rlabel metal2 s 600000 978299 601018 978351 6 mprj_io_inp_dis[14]
port 488 nsew default input
rlabel metal2 s 560849 1020000 560901 1021018 6 mprj_io_inp_dis[15]
port 489 nsew default input
rlabel metal2 s 465649 1020000 465701 1021018 6 mprj_io_inp_dis[16]
port 490 nsew default input
rlabel metal2 s 417649 1020000 417701 1021018 6 mprj_io_inp_dis[17]
port 491 nsew default input
rlabel metal2 s 369449 1020000 369501 1021018 6 mprj_io_inp_dis[18]
port 492 nsew default input
rlabel metal2 s 274249 1020000 274301 1021018 6 mprj_io_inp_dis[19]
port 493 nsew default input
rlabel metal2 s 600000 126099 601018 126151 6 mprj_io_inp_dis[1]
port 494 nsew default input
rlabel metal2 s 226249 1020000 226301 1021018 6 mprj_io_inp_dis[20]
port 495 nsew default input
rlabel metal2 s 178049 1020000 178101 1021018 6 mprj_io_inp_dis[21]
port 496 nsew default input
rlabel metal2 s 130049 1020000 130101 1021018 6 mprj_io_inp_dis[22]
port 497 nsew default input
rlabel metal2 s 81849 1020000 81901 1021018 6 mprj_io_inp_dis[23]
port 498 nsew default input
rlabel metal2 s 38982 983449 40000 983501 6 mprj_io_inp_dis[24]
port 499 nsew default input
rlabel metal2 s 38982 804249 40000 804301 6 mprj_io_inp_dis[25]
port 500 nsew default input
rlabel metal2 s 38982 758649 40000 758701 6 mprj_io_inp_dis[26]
port 501 nsew default input
rlabel metal2 s 38982 713049 40000 713101 6 mprj_io_inp_dis[27]
port 502 nsew default input
rlabel metal2 s 38982 667449 40000 667501 6 mprj_io_inp_dis[28]
port 503 nsew default input
rlabel metal2 s 38982 622049 40000 622101 6 mprj_io_inp_dis[29]
port 504 nsew default input
rlabel metal2 s 600000 173699 601018 173751 6 mprj_io_inp_dis[2]
port 505 nsew default input
rlabel metal2 s 38982 576449 40000 576501 6 mprj_io_inp_dis[30]
port 506 nsew default input
rlabel metal2 s 38982 530849 40000 530901 6 mprj_io_inp_dis[31]
port 507 nsew default input
rlabel metal2 s 38982 396249 40000 396301 6 mprj_io_inp_dis[32]
port 508 nsew default input
rlabel metal2 s 38982 350649 40000 350701 6 mprj_io_inp_dis[33]
port 509 nsew default input
rlabel metal2 s 38982 305049 40000 305101 6 mprj_io_inp_dis[34]
port 510 nsew default input
rlabel metal2 s 38982 259449 40000 259501 6 mprj_io_inp_dis[35]
port 511 nsew default input
rlabel metal2 s 38982 214049 40000 214101 6 mprj_io_inp_dis[36]
port 512 nsew default input
rlabel metal2 s 38982 168449 40000 168501 6 mprj_io_inp_dis[37]
port 513 nsew default input
rlabel metal2 s 600000 221299 601018 221351 6 mprj_io_inp_dis[3]
port 514 nsew default input
rlabel metal2 s 600000 268899 601018 268951 6 mprj_io_inp_dis[4]
port 515 nsew default input
rlabel metal2 s 600000 316499 601018 316551 6 mprj_io_inp_dis[5]
port 516 nsew default input
rlabel metal2 s 600000 364299 601018 364351 6 mprj_io_inp_dis[6]
port 517 nsew default input
rlabel metal2 s 600000 551699 601018 551751 6 mprj_io_inp_dis[7]
port 518 nsew default input
rlabel metal2 s 600000 599299 601018 599351 6 mprj_io_inp_dis[8]
port 519 nsew default input
rlabel metal2 s 600000 646899 601018 646951 6 mprj_io_inp_dis[9]
port 520 nsew default input
rlabel metal2 s 600000 86879 600894 86925 6 mprj_io_oeb[0]
port 521 nsew default input
rlabel metal2 s 600000 703079 600894 703125 6 mprj_io_oeb[10]
port 522 nsew default input
rlabel metal2 s 600000 750679 600894 750725 6 mprj_io_oeb[11]
port 523 nsew default input
rlabel metal2 s 600000 798279 600894 798325 6 mprj_io_oeb[12]
port 524 nsew default input
rlabel metal2 s 600000 892479 600894 892525 6 mprj_io_oeb[13]
port 525 nsew default input
rlabel metal2 s 600000 986679 600894 986725 6 mprj_io_oeb[14]
port 526 nsew default input
rlabel metal2 s 552475 1020000 552521 1020894 6 mprj_io_oeb[15]
port 527 nsew default input
rlabel metal2 s 457275 1020000 457321 1020894 6 mprj_io_oeb[16]
port 528 nsew default input
rlabel metal2 s 409275 1020000 409321 1020894 6 mprj_io_oeb[17]
port 529 nsew default input
rlabel metal2 s 361075 1020000 361121 1020894 6 mprj_io_oeb[18]
port 530 nsew default input
rlabel metal2 s 265875 1020000 265921 1020894 6 mprj_io_oeb[19]
port 531 nsew default input
rlabel metal2 s 600000 134479 600894 134525 6 mprj_io_oeb[1]
port 532 nsew default input
rlabel metal2 s 217875 1020000 217921 1020894 6 mprj_io_oeb[20]
port 533 nsew default input
rlabel metal2 s 169675 1020000 169721 1020894 6 mprj_io_oeb[21]
port 534 nsew default input
rlabel metal2 s 121675 1020000 121721 1020894 6 mprj_io_oeb[22]
port 535 nsew default input
rlabel metal2 s 73475 1020000 73521 1020894 6 mprj_io_oeb[23]
port 536 nsew default input
rlabel metal2 s 39105 975075 39999 975121 6 mprj_io_oeb[24]
port 537 nsew default input
rlabel metal2 s 39105 795875 39999 795921 6 mprj_io_oeb[25]
port 538 nsew default input
rlabel metal2 s 39105 750275 39999 750321 6 mprj_io_oeb[26]
port 539 nsew default input
rlabel metal2 s 39105 704675 39999 704721 6 mprj_io_oeb[27]
port 540 nsew default input
rlabel metal2 s 39105 659075 39999 659121 6 mprj_io_oeb[28]
port 541 nsew default input
rlabel metal2 s 39105 613675 39999 613721 6 mprj_io_oeb[29]
port 542 nsew default input
rlabel metal2 s 600000 182079 600894 182125 6 mprj_io_oeb[2]
port 543 nsew default input
rlabel metal2 s 39105 568075 39999 568121 6 mprj_io_oeb[30]
port 544 nsew default input
rlabel metal2 s 39105 522475 39999 522521 6 mprj_io_oeb[31]
port 545 nsew default input
rlabel metal2 s 39105 387875 39999 387921 6 mprj_io_oeb[32]
port 546 nsew default input
rlabel metal2 s 39105 342275 39999 342321 6 mprj_io_oeb[33]
port 547 nsew default input
rlabel metal2 s 39105 296675 39999 296721 6 mprj_io_oeb[34]
port 548 nsew default input
rlabel metal2 s 39105 251075 39999 251121 6 mprj_io_oeb[35]
port 549 nsew default input
rlabel metal2 s 39105 205675 39999 205721 6 mprj_io_oeb[36]
port 550 nsew default input
rlabel metal2 s 39105 160075 39999 160121 6 mprj_io_oeb[37]
port 551 nsew default input
rlabel metal2 s 600000 229679 600894 229725 6 mprj_io_oeb[3]
port 552 nsew default input
rlabel metal2 s 600000 277279 600894 277325 6 mprj_io_oeb[4]
port 553 nsew default input
rlabel metal2 s 600000 324879 600894 324925 6 mprj_io_oeb[5]
port 554 nsew default input
rlabel metal2 s 600000 372679 600894 372725 6 mprj_io_oeb[6]
port 555 nsew default input
rlabel metal2 s 600000 560079 600894 560125 6 mprj_io_oeb[7]
port 556 nsew default input
rlabel metal2 s 600000 607679 600894 607725 6 mprj_io_oeb[8]
port 557 nsew default input
rlabel metal2 s 600000 655279 600894 655325 6 mprj_io_oeb[9]
port 558 nsew default input
rlabel metal2 s 600000 83077 601284 83129 6 mprj_io_out[0]
port 559 nsew default input
rlabel metal2 s 600000 699277 601284 699329 6 mprj_io_out[10]
port 560 nsew default input
rlabel metal2 s 600000 746877 601284 746929 6 mprj_io_out[11]
port 561 nsew default input
rlabel metal2 s 600000 794477 601284 794529 6 mprj_io_out[12]
port 562 nsew default input
rlabel metal2 s 600000 888677 601284 888729 6 mprj_io_out[13]
port 563 nsew default input
rlabel metal2 s 600000 982877 601284 982929 6 mprj_io_out[14]
port 564 nsew default input
rlabel metal2 s 556271 1020000 556323 1021284 6 mprj_io_out[15]
port 565 nsew default input
rlabel metal2 s 461071 1020000 461123 1021284 6 mprj_io_out[16]
port 566 nsew default input
rlabel metal2 s 413071 1020000 413123 1021284 6 mprj_io_out[17]
port 567 nsew default input
rlabel metal2 s 364871 1020000 364923 1021284 6 mprj_io_out[18]
port 568 nsew default input
rlabel metal2 s 269671 1020000 269723 1021284 6 mprj_io_out[19]
port 569 nsew default input
rlabel metal2 s 600000 130677 601284 130729 6 mprj_io_out[1]
port 570 nsew default input
rlabel metal2 s 221671 1020000 221723 1021284 6 mprj_io_out[20]
port 571 nsew default input
rlabel metal2 s 173471 1020000 173523 1021284 6 mprj_io_out[21]
port 572 nsew default input
rlabel metal2 s 125471 1020000 125523 1021284 6 mprj_io_out[22]
port 573 nsew default input
rlabel metal2 s 77271 1020000 77323 1021284 6 mprj_io_out[23]
port 574 nsew default input
rlabel metal2 s 38715 978871 39999 978923 6 mprj_io_out[24]
port 575 nsew default input
rlabel metal2 s 38715 799671 39999 799723 6 mprj_io_out[25]
port 576 nsew default input
rlabel metal2 s 38715 754071 39999 754123 6 mprj_io_out[26]
port 577 nsew default input
rlabel metal2 s 38715 708471 39999 708523 6 mprj_io_out[27]
port 578 nsew default input
rlabel metal2 s 38715 662871 39999 662923 6 mprj_io_out[28]
port 579 nsew default input
rlabel metal2 s 38715 617471 39999 617523 6 mprj_io_out[29]
port 580 nsew default input
rlabel metal2 s 600000 178277 601284 178329 6 mprj_io_out[2]
port 581 nsew default input
rlabel metal2 s 38715 571871 39999 571923 6 mprj_io_out[30]
port 582 nsew default input
rlabel metal2 s 38715 526271 39999 526323 6 mprj_io_out[31]
port 583 nsew default input
rlabel metal2 s 38715 391671 39999 391723 6 mprj_io_out[32]
port 584 nsew default input
rlabel metal2 s 38715 346071 39999 346123 6 mprj_io_out[33]
port 585 nsew default input
rlabel metal2 s 38715 300471 39999 300523 6 mprj_io_out[34]
port 586 nsew default input
rlabel metal2 s 38715 254871 39999 254923 6 mprj_io_out[35]
port 587 nsew default input
rlabel metal2 s 38715 209471 39999 209523 6 mprj_io_out[36]
port 588 nsew default input
rlabel metal2 s 38715 163871 39999 163923 6 mprj_io_out[37]
port 589 nsew default input
rlabel metal2 s 600000 225877 601284 225929 6 mprj_io_out[3]
port 590 nsew default input
rlabel metal2 s 600000 273477 601284 273529 6 mprj_io_out[4]
port 591 nsew default input
rlabel metal2 s 600000 321077 601284 321129 6 mprj_io_out[5]
port 592 nsew default input
rlabel metal2 s 600000 368877 601284 368929 6 mprj_io_out[6]
port 593 nsew default input
rlabel metal2 s 600000 556277 601284 556329 6 mprj_io_out[7]
port 594 nsew default input
rlabel metal2 s 600000 603877 601284 603929 6 mprj_io_out[8]
port 595 nsew default input
rlabel metal2 s 600000 651477 601284 651529 6 mprj_io_out[9]
port 596 nsew default input
rlabel metal2 s 600000 72026 600236 72078 6 mprj_io_slow_sel[0]
port 597 nsew default input
rlabel metal2 s 600000 688226 600236 688278 6 mprj_io_slow_sel[10]
port 598 nsew default input
rlabel metal2 s 600000 735826 600236 735878 6 mprj_io_slow_sel[11]
port 599 nsew default input
rlabel metal2 s 600000 783426 600236 783478 6 mprj_io_slow_sel[12]
port 600 nsew default input
rlabel metal2 s 600000 877626 600236 877678 6 mprj_io_slow_sel[13]
port 601 nsew default input
rlabel metal2 s 600000 971826 600236 971878 6 mprj_io_slow_sel[14]
port 602 nsew default input
rlabel metal2 s 567322 1020000 567374 1020236 6 mprj_io_slow_sel[15]
port 603 nsew default input
rlabel metal2 s 472122 1020000 472174 1020236 6 mprj_io_slow_sel[16]
port 604 nsew default input
rlabel metal2 s 424122 1020000 424174 1020236 6 mprj_io_slow_sel[17]
port 605 nsew default input
rlabel metal2 s 375922 1020000 375974 1020236 6 mprj_io_slow_sel[18]
port 606 nsew default input
rlabel metal2 s 280722 1020000 280774 1020236 6 mprj_io_slow_sel[19]
port 607 nsew default input
rlabel metal2 s 600000 119626 600236 119678 6 mprj_io_slow_sel[1]
port 608 nsew default input
rlabel metal2 s 232722 1020000 232774 1020236 6 mprj_io_slow_sel[20]
port 609 nsew default input
rlabel metal2 s 184522 1020000 184574 1020236 6 mprj_io_slow_sel[21]
port 610 nsew default input
rlabel metal2 s 136522 1020000 136574 1020236 6 mprj_io_slow_sel[22]
port 611 nsew default input
rlabel metal2 s 88322 1020000 88374 1020236 6 mprj_io_slow_sel[23]
port 612 nsew default input
rlabel metal2 s 39763 989922 39999 989974 6 mprj_io_slow_sel[24]
port 613 nsew default input
rlabel metal2 s 39763 810722 39999 810774 6 mprj_io_slow_sel[25]
port 614 nsew default input
rlabel metal2 s 39763 765122 39999 765174 6 mprj_io_slow_sel[26]
port 615 nsew default input
rlabel metal2 s 39763 719522 39999 719574 6 mprj_io_slow_sel[27]
port 616 nsew default input
rlabel metal2 s 39763 673922 39999 673974 6 mprj_io_slow_sel[28]
port 617 nsew default input
rlabel metal2 s 39763 628522 39999 628574 6 mprj_io_slow_sel[29]
port 618 nsew default input
rlabel metal2 s 600000 167226 600236 167278 6 mprj_io_slow_sel[2]
port 619 nsew default input
rlabel metal2 s 39763 582922 39999 582974 6 mprj_io_slow_sel[30]
port 620 nsew default input
rlabel metal2 s 39763 537322 39999 537374 6 mprj_io_slow_sel[31]
port 621 nsew default input
rlabel metal2 s 39763 402722 39999 402774 6 mprj_io_slow_sel[32]
port 622 nsew default input
rlabel metal2 s 39763 357122 39999 357174 6 mprj_io_slow_sel[33]
port 623 nsew default input
rlabel metal2 s 39763 311522 39999 311574 6 mprj_io_slow_sel[34]
port 624 nsew default input
rlabel metal2 s 39763 265922 39999 265974 6 mprj_io_slow_sel[35]
port 625 nsew default input
rlabel metal2 s 39763 220522 39999 220574 6 mprj_io_slow_sel[36]
port 626 nsew default input
rlabel metal2 s 39763 174922 39999 174974 6 mprj_io_slow_sel[37]
port 627 nsew default input
rlabel metal2 s 600000 214826 600236 214878 6 mprj_io_slow_sel[3]
port 628 nsew default input
rlabel metal2 s 600000 262426 600236 262478 6 mprj_io_slow_sel[4]
port 629 nsew default input
rlabel metal2 s 600000 310026 600236 310078 6 mprj_io_slow_sel[5]
port 630 nsew default input
rlabel metal2 s 600000 357826 600236 357878 6 mprj_io_slow_sel[6]
port 631 nsew default input
rlabel metal2 s 600000 545226 600236 545278 6 mprj_io_slow_sel[7]
port 632 nsew default input
rlabel metal2 s 600000 592826 600236 592878 6 mprj_io_slow_sel[8]
port 633 nsew default input
rlabel metal2 s 600000 640426 600236 640478 6 mprj_io_slow_sel[9]
port 634 nsew default input
rlabel metal2 s 600000 86322 600310 86374 6 mprj_io_vtrip_sel[0]
port 635 nsew default input
rlabel metal2 s 600000 702522 600310 702574 6 mprj_io_vtrip_sel[10]
port 636 nsew default input
rlabel metal2 s 600000 750122 600310 750174 6 mprj_io_vtrip_sel[11]
port 637 nsew default input
rlabel metal2 s 600000 797722 600310 797774 6 mprj_io_vtrip_sel[12]
port 638 nsew default input
rlabel metal2 s 600000 891922 600310 891974 6 mprj_io_vtrip_sel[13]
port 639 nsew default input
rlabel metal2 s 600000 986122 600310 986174 6 mprj_io_vtrip_sel[14]
port 640 nsew default input
rlabel metal2 s 553026 1020000 553078 1020310 6 mprj_io_vtrip_sel[15]
port 641 nsew default input
rlabel metal2 s 457826 1020000 457878 1020310 6 mprj_io_vtrip_sel[16]
port 642 nsew default input
rlabel metal2 s 409826 1020000 409878 1020310 6 mprj_io_vtrip_sel[17]
port 643 nsew default input
rlabel metal2 s 361626 1020000 361678 1020310 6 mprj_io_vtrip_sel[18]
port 644 nsew default input
rlabel metal2 s 266426 1020000 266478 1020310 6 mprj_io_vtrip_sel[19]
port 645 nsew default input
rlabel metal2 s 600000 133922 600310 133974 6 mprj_io_vtrip_sel[1]
port 646 nsew default input
rlabel metal2 s 218426 1020000 218478 1020310 6 mprj_io_vtrip_sel[20]
port 647 nsew default input
rlabel metal2 s 170226 1020000 170278 1020310 6 mprj_io_vtrip_sel[21]
port 648 nsew default input
rlabel metal2 s 122226 1020000 122278 1020310 6 mprj_io_vtrip_sel[22]
port 649 nsew default input
rlabel metal2 s 74026 1020000 74078 1020310 6 mprj_io_vtrip_sel[23]
port 650 nsew default input
rlabel metal2 s 39690 975626 40000 975678 6 mprj_io_vtrip_sel[24]
port 651 nsew default input
rlabel metal2 s 39690 796426 40000 796478 6 mprj_io_vtrip_sel[25]
port 652 nsew default input
rlabel metal2 s 39690 750826 40000 750878 6 mprj_io_vtrip_sel[26]
port 653 nsew default input
rlabel metal2 s 39690 705226 40000 705278 6 mprj_io_vtrip_sel[27]
port 654 nsew default input
rlabel metal2 s 39690 659626 40000 659678 6 mprj_io_vtrip_sel[28]
port 655 nsew default input
rlabel metal2 s 39690 614226 40000 614278 6 mprj_io_vtrip_sel[29]
port 656 nsew default input
rlabel metal2 s 600000 181522 600310 181574 6 mprj_io_vtrip_sel[2]
port 657 nsew default input
rlabel metal2 s 39690 568626 40000 568678 6 mprj_io_vtrip_sel[30]
port 658 nsew default input
rlabel metal2 s 39690 523026 40000 523078 6 mprj_io_vtrip_sel[31]
port 659 nsew default input
rlabel metal2 s 39690 388426 40000 388478 6 mprj_io_vtrip_sel[32]
port 660 nsew default input
rlabel metal2 s 39690 342826 40000 342878 6 mprj_io_vtrip_sel[33]
port 661 nsew default input
rlabel metal2 s 39690 297226 40000 297278 6 mprj_io_vtrip_sel[34]
port 662 nsew default input
rlabel metal2 s 39690 251626 40000 251678 6 mprj_io_vtrip_sel[35]
port 663 nsew default input
rlabel metal2 s 39690 206226 40000 206278 6 mprj_io_vtrip_sel[36]
port 664 nsew default input
rlabel metal2 s 39690 160626 40000 160678 6 mprj_io_vtrip_sel[37]
port 665 nsew default input
rlabel metal2 s 600000 229122 600310 229174 6 mprj_io_vtrip_sel[3]
port 666 nsew default input
rlabel metal2 s 600000 276722 600310 276774 6 mprj_io_vtrip_sel[4]
port 667 nsew default input
rlabel metal2 s 600000 324322 600310 324374 6 mprj_io_vtrip_sel[5]
port 668 nsew default input
rlabel metal2 s 600000 372122 600310 372174 6 mprj_io_vtrip_sel[6]
port 669 nsew default input
rlabel metal2 s 600000 559522 600310 559574 6 mprj_io_vtrip_sel[7]
port 670 nsew default input
rlabel metal2 s 600000 607122 600310 607174 6 mprj_io_vtrip_sel[8]
port 671 nsew default input
rlabel metal2 s 600000 654722 600310 654774 6 mprj_io_vtrip_sel[9]
port 672 nsew default input
rlabel metal2 s 173899 38982 173951 40000 6 por
port 673 nsew default input
rlabel metal2 s 132091 39706 132143 40000 6 porb_h
port 674 nsew default input
rlabel metal5 s 120840 6675 133380 19197 6 resetb
port 675 nsew default input
rlabel metal3 s 128667 38031 128813 39999 6 resetb_core_h
port 676 nsew default tristate
rlabel metal5 s 6086 72063 19572 83391 6 vccd
port 677 nsew default bidirectional
rlabel metal5 s 620428 926609 633914 937937 6 vccd1
port 678 nsew default bidirectional
rlabel metal5 s 6086 931663 19572 942991 6 vccd2
port 679 nsew default bidirectional
rlabel metal5 s 553040 6675 565580 19197 6 vdda
port 680 nsew default bidirectional
rlabel metal5 s 620802 831840 633324 844380 6 vdda1
port 681 nsew default bidirectional
rlabel metal5 s 6675 478420 19197 490960 6 vdda2
port 682 nsew default bidirectional
rlabel metal5 s 6675 116020 19197 128560 6 vddio
port 683 nsew default bidirectional
rlabel metal5 s 73440 6675 85980 19197 6 vssa
port 684 nsew default bidirectional
rlabel metal5 s 506020 1040802 518560 1053324 6 vssa1
port 685 nsew default bidirectional
rlabel metal5 s 6675 841820 19197 854360 6 vssa2
port 686 nsew default bidirectional
rlabel metal5 s 217209 6086 228537 19572 6 vssd
port 687 nsew default bidirectional
rlabel metal5 s 620428 453409 633914 464737 6 vssd1
port 688 nsew default bidirectional
rlabel metal5 s 6086 434463 19572 445791 6 vssd2
port 689 nsew default bidirectional
rlabel metal5 s 314620 1040802 327160 1053324 6 vssio
port 690 nsew default bidirectional
<< properties >>
string FIXED_BBOX 0 0 640000 1060000
<< end >>
