magic
tech sky130A
magscale 1 2
timestamp 1606431493
<< metal3 >>
rect -5928 3222 -2056 3250
rect -5928 78 -2140 3222
rect -2076 78 -2056 3222
rect -5928 50 -2056 78
rect -1936 3222 1936 3250
rect -1936 78 1852 3222
rect 1916 78 1936 3222
rect -1936 50 1936 78
rect 2056 3222 5928 3250
rect 2056 78 5844 3222
rect 5908 78 5928 3222
rect 2056 50 5928 78
rect -5928 -78 -2056 -50
rect -5928 -3222 -2140 -78
rect -2076 -3222 -2056 -78
rect -5928 -3250 -2056 -3222
rect -1936 -78 1936 -50
rect -1936 -3222 1852 -78
rect 1916 -3222 1936 -78
rect -1936 -3250 1936 -3222
rect 2056 -78 5928 -50
rect 2056 -3222 5844 -78
rect 5908 -3222 5928 -78
rect 2056 -3250 5928 -3222
<< via3 >>
rect -2140 78 -2076 3222
rect 1852 78 1916 3222
rect 5844 78 5908 3222
rect -2140 -3222 -2076 -78
rect 1852 -3222 1916 -78
rect 5844 -3222 5908 -78
<< mimcap >>
rect -5828 3110 -2328 3150
rect -5828 190 -5788 3110
rect -2368 190 -2328 3110
rect -5828 150 -2328 190
rect -1836 3110 1664 3150
rect -1836 190 -1796 3110
rect 1624 190 1664 3110
rect -1836 150 1664 190
rect 2156 3110 5656 3150
rect 2156 190 2196 3110
rect 5616 190 5656 3110
rect 2156 150 5656 190
rect -5828 -190 -2328 -150
rect -5828 -3110 -5788 -190
rect -2368 -3110 -2328 -190
rect -5828 -3150 -2328 -3110
rect -1836 -190 1664 -150
rect -1836 -3110 -1796 -190
rect 1624 -3110 1664 -190
rect -1836 -3150 1664 -3110
rect 2156 -190 5656 -150
rect 2156 -3110 2196 -190
rect 5616 -3110 5656 -190
rect 2156 -3150 5656 -3110
<< mimcapcontact >>
rect -5788 190 -2368 3110
rect -1796 190 1624 3110
rect 2196 190 5616 3110
rect -5788 -3110 -2368 -190
rect -1796 -3110 1624 -190
rect 2196 -3110 5616 -190
<< metal4 >>
rect -4130 3111 -4026 3300
rect -2160 3222 -2056 3300
rect -5789 3110 -2367 3111
rect -5789 190 -5788 3110
rect -2368 190 -2367 3110
rect -5789 189 -2367 190
rect -4130 -189 -4026 189
rect -2160 78 -2140 3222
rect -2076 78 -2056 3222
rect -138 3111 -34 3300
rect 1832 3222 1936 3300
rect -1797 3110 1625 3111
rect -1797 190 -1796 3110
rect 1624 190 1625 3110
rect -1797 189 1625 190
rect -2160 -78 -2056 78
rect -5789 -190 -2367 -189
rect -5789 -3110 -5788 -190
rect -2368 -3110 -2367 -190
rect -5789 -3111 -2367 -3110
rect -4130 -3300 -4026 -3111
rect -2160 -3222 -2140 -78
rect -2076 -3222 -2056 -78
rect -138 -189 -34 189
rect 1832 78 1852 3222
rect 1916 78 1936 3222
rect 3854 3111 3958 3300
rect 5824 3222 5928 3300
rect 2195 3110 5617 3111
rect 2195 190 2196 3110
rect 5616 190 5617 3110
rect 2195 189 5617 190
rect 1832 -78 1936 78
rect -1797 -190 1625 -189
rect -1797 -3110 -1796 -190
rect 1624 -3110 1625 -190
rect -1797 -3111 1625 -3110
rect -2160 -3300 -2056 -3222
rect -138 -3300 -34 -3111
rect 1832 -3222 1852 -78
rect 1916 -3222 1936 -78
rect 3854 -189 3958 189
rect 5824 78 5844 3222
rect 5908 78 5928 3222
rect 5824 -78 5928 78
rect 2195 -190 5617 -189
rect 2195 -3110 2196 -190
rect 5616 -3110 5617 -190
rect 2195 -3111 5617 -3110
rect 1832 -3300 1936 -3222
rect 3854 -3300 3958 -3111
rect 5824 -3222 5844 -78
rect 5908 -3222 5928 -78
rect 5824 -3300 5928 -3222
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 2056 50 5756 3250
string parameters w 17.5 l 15 val 273.55 carea 1.00 cperi 0.17 nx 3 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string library sky130
<< end >>
