magic
tech sky130A
magscale 1 2
timestamp 1622459969
<< obsli1 >>
rect 1104 1071 13892 15793
<< obsm1 >>
rect 474 1040 13892 15824
<< metal2 >>
rect 478 16200 534 17000
rect 1858 16200 1914 17000
rect 3238 16200 3294 17000
rect 4618 16200 4674 17000
rect 5998 16200 6054 17000
rect 6918 16200 6974 17000
rect 8298 16200 8354 17000
rect 9678 16200 9734 17000
rect 11058 16200 11114 17000
rect 12438 16200 12494 17000
rect 13818 16200 13874 17000
rect 478 0 534 800
rect 1398 0 1454 800
rect 2778 0 2834 800
rect 4158 0 4214 800
rect 5538 0 5594 800
rect 6918 0 6974 800
rect 8298 0 8354 800
rect 9678 0 9734 800
rect 11058 0 11114 800
rect 12438 0 12494 800
rect 13818 0 13874 800
<< obsm2 >>
rect 590 16144 1802 16200
rect 1970 16144 3182 16200
rect 3350 16144 4562 16200
rect 4730 16144 5942 16200
rect 6110 16144 6862 16200
rect 7030 16144 8242 16200
rect 8410 16144 9622 16200
rect 9790 16144 11002 16200
rect 11170 16144 12382 16200
rect 12550 16144 13762 16200
rect 480 856 13874 16144
rect 590 800 1342 856
rect 1510 800 2722 856
rect 2890 800 4102 856
rect 4270 800 5482 856
rect 5650 800 6862 856
rect 7030 800 8242 856
rect 8410 800 9622 856
rect 9790 800 11002 856
rect 11170 800 12382 856
rect 12550 800 13762 856
<< metal3 >>
rect 14200 14968 15000 15088
rect 0 14288 800 14408
rect 14200 12928 15000 13048
rect 0 12248 800 12368
rect 14200 10888 15000 11008
rect 0 10208 800 10328
rect 14200 8848 15000 8968
rect 0 8168 800 8288
rect 14200 6808 15000 6928
rect 0 6128 800 6248
rect 14200 4768 15000 4888
rect 0 4088 800 4208
rect 14200 3408 15000 3528
rect 0 2048 800 2168
rect 14200 1368 15000 1488
<< obsm3 >>
rect 800 15168 14200 15809
rect 800 14888 14120 15168
rect 800 14488 14200 14888
rect 880 14208 14200 14488
rect 800 13128 14200 14208
rect 800 12848 14120 13128
rect 800 12448 14200 12848
rect 880 12168 14200 12448
rect 800 11088 14200 12168
rect 800 10808 14120 11088
rect 800 10408 14200 10808
rect 880 10128 14200 10408
rect 800 9048 14200 10128
rect 800 8768 14120 9048
rect 800 8368 14200 8768
rect 880 8088 14200 8368
rect 800 7008 14200 8088
rect 800 6728 14120 7008
rect 800 6328 14200 6728
rect 880 6048 14200 6328
rect 800 4968 14200 6048
rect 800 4688 14120 4968
rect 800 4288 14200 4688
rect 880 4008 14200 4288
rect 800 3608 14200 4008
rect 800 3328 14120 3608
rect 800 2248 14200 3328
rect 880 1968 14200 2248
rect 800 1568 14200 1968
rect 800 1288 14120 1568
rect 800 1055 14200 1288
<< metal4 >>
rect 4208 1040 4528 15824
rect 8208 1040 8528 15824
rect 12208 1040 12528 15824
<< labels >>
rlabel metal2 s 5538 0 5594 800 6 clockp[0]
port 1 nsew signal output
rlabel metal2 s 5998 16200 6054 17000 6 clockp[1]
port 2 nsew signal output
rlabel metal2 s 8298 16200 8354 17000 6 dco
port 3 nsew signal input
rlabel metal2 s 11058 16200 11114 17000 6 div[0]
port 4 nsew signal input
rlabel metal3 s 14200 3408 15000 3528 6 div[1]
port 5 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 div[2]
port 6 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 div[3]
port 7 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 div[4]
port 8 nsew signal input
rlabel metal2 s 13818 16200 13874 17000 6 enable
port 9 nsew signal input
rlabel metal2 s 6918 16200 6974 17000 6 ext_trim[0]
port 10 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 ext_trim[10]
port 11 nsew signal input
rlabel metal2 s 478 0 534 800 6 ext_trim[11]
port 12 nsew signal input
rlabel metal2 s 3238 16200 3294 17000 6 ext_trim[12]
port 13 nsew signal input
rlabel metal2 s 4618 16200 4674 17000 6 ext_trim[13]
port 14 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 ext_trim[14]
port 15 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 ext_trim[15]
port 16 nsew signal input
rlabel metal3 s 14200 8848 15000 8968 6 ext_trim[16]
port 17 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 ext_trim[17]
port 18 nsew signal input
rlabel metal3 s 14200 1368 15000 1488 6 ext_trim[18]
port 19 nsew signal input
rlabel metal2 s 12438 16200 12494 17000 6 ext_trim[19]
port 20 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 ext_trim[1]
port 21 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 ext_trim[20]
port 22 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 ext_trim[21]
port 23 nsew signal input
rlabel metal3 s 14200 12928 15000 13048 6 ext_trim[22]
port 24 nsew signal input
rlabel metal2 s 1858 16200 1914 17000 6 ext_trim[23]
port 25 nsew signal input
rlabel metal2 s 478 16200 534 17000 6 ext_trim[24]
port 26 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 ext_trim[25]
port 27 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 ext_trim[2]
port 28 nsew signal input
rlabel metal2 s 9678 16200 9734 17000 6 ext_trim[3]
port 29 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 ext_trim[4]
port 30 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 ext_trim[5]
port 31 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 ext_trim[6]
port 32 nsew signal input
rlabel metal3 s 14200 10888 15000 11008 6 ext_trim[7]
port 33 nsew signal input
rlabel metal3 s 14200 4768 15000 4888 6 ext_trim[8]
port 34 nsew signal input
rlabel metal3 s 14200 14968 15000 15088 6 ext_trim[9]
port 35 nsew signal input
rlabel metal3 s 14200 6808 15000 6928 6 osc
port 36 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 resetb
port 37 nsew signal input
rlabel metal4 s 12208 1040 12528 15824 6 VPWR
port 38 nsew power bidirectional
rlabel metal4 s 4208 1040 4528 15824 6 VPWR
port 39 nsew power bidirectional
rlabel metal4 s 8208 1040 8528 15824 6 VGND
port 40 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 15000 17000
string LEFview TRUE
string GDS_FILE ../gds/digital_pll.gds
string GDS_END 1103108
string GDS_START 339452
<< end >>

