magic
tech sky130A
magscale 12 1
timestamp 1598765816
<< metal5 >>
rect 0 90 45 105
rect 15 15 30 90
rect 0 0 45 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
