* SPICE NETLIST
***************************************

.SUBCKT MN g s d b
.ENDS
***************************************
.SUBCKT MP g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT condiodeHvPsub pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20nativevhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT n20nativevhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT p20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808678
** N=22 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808675
** N=61 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808679
** N=22 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808662
** N=60 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808663
** N=120 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_5595914180851
** N=17 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 2 3
** N=9 EP=2 IP=6 FDC=1
*.SEEDPROM
M0 2 3 2 2 nhv L=4 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 r=1.25 sa=2e+06 sb=2e+06 a=20 p=18 mult=1 $X=0 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT sky130_fd_io__sio_clamp_pcap_4x5 2 3
** N=83 EP=2 IP=6 FDC=1
*.SEEDPROM
X0 2 3 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 $T=1145 720 0 0 $X=700 $Y=540
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s2__example_55959141808676
** N=90 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__esd_rcclamp_nfetcap 2 3
** N=122 EP=2 IP=6 FDC=1
*.SEEDPROM
M0 2 3 2 2 nhv L=8 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 r=0.625 sa=4e+06 sb=4e+06 a=40 p=26 mult=1 $X=895 $Y=630 $D=49
.ENDS
***************************************
.SUBCKT ICV_2 2 3
** N=167 EP=2 IP=188 FDC=2
*.SEEDPROM
X0 2 3 sky130_fd_io__esd_rcclamp_nfetcap $T=-9760 0 0 0 $X=-10010 $Y=-90
X1 2 3 sky130_fd_io__esd_rcclamp_nfetcap $T=0 0 0 0 $X=-250 $Y=-90
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808671
** N=119 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s2__example_55959141808672
** N=177 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808670
** N=23 EP=0 IP=30 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808673
** N=27 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808336
** N=22 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808666
** N=23 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_3
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_4
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_5
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_6
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808665 2 3 4
** N=254 EP=3 IP=16 FDC=50
*.SEEDPROM
M0 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 r=14 sa=250000 sb=250020 a=3.5 p=15 mult=1 $X=0 $Y=0 $D=109
M1 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250001 sb=250020 a=3.5 p=15 mult=1 $X=780 $Y=0 $D=109
M2 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250020 a=3.5 p=15 mult=1 $X=1560 $Y=0 $D=109
M3 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250020 a=3.5 p=15 mult=1 $X=2340 $Y=0 $D=109
M4 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250003 sb=250020 a=3.5 p=15 mult=1 $X=3120 $Y=0 $D=109
M5 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250004 sb=250020 a=3.5 p=15 mult=1 $X=3900 $Y=0 $D=109
M6 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250020 a=3.5 p=15 mult=1 $X=4680 $Y=0 $D=109
M7 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250020 a=3.5 p=15 mult=1 $X=5460 $Y=0 $D=109
M8 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250006 sb=250020 a=3.5 p=15 mult=1 $X=6240 $Y=0 $D=109
M9 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250007 sb=250020 a=3.5 p=15 mult=1 $X=7020 $Y=0 $D=109
M10 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250008 sb=250020 a=3.5 p=15 mult=1 $X=7800 $Y=0 $D=109
M11 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250020 a=3.5 p=15 mult=1 $X=8580 $Y=0 $D=109
M12 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250020 a=3.5 p=15 mult=1 $X=9360 $Y=0 $D=109
M13 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250010 sb=250020 a=3.5 p=15 mult=1 $X=10140 $Y=0 $D=109
M14 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250011 sb=250020 a=3.5 p=15 mult=1 $X=10920 $Y=0 $D=109
M15 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250012 sb=250020 a=3.5 p=15 mult=1 $X=11700 $Y=0 $D=109
M16 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250012 sb=250020 a=3.5 p=15 mult=1 $X=12480 $Y=0 $D=109
M17 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250013 sb=250020 a=3.5 p=15 mult=1 $X=13260 $Y=0 $D=109
M18 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250014 sb=250020 a=3.5 p=15 mult=1 $X=14040 $Y=0 $D=109
M19 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250015 sb=250020 a=3.5 p=15 mult=1 $X=14820 $Y=0 $D=109
M20 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250016 sb=250020 a=3.5 p=15 mult=1 $X=15600 $Y=0 $D=109
M21 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250016 sb=250020 a=3.5 p=15 mult=1 $X=16380 $Y=0 $D=109
M22 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250017 sb=250020 a=3.5 p=15 mult=1 $X=17160 $Y=0 $D=109
M23 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250018 sb=250020 a=3.5 p=15 mult=1 $X=17940 $Y=0 $D=109
M24 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250019 sb=250020 a=3.5 p=15 mult=1 $X=18720 $Y=0 $D=109
M25 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250019 a=3.5 p=15 mult=1 $X=19500 $Y=0 $D=109
M26 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250018 a=3.5 p=15 mult=1 $X=20280 $Y=0 $D=109
M27 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250017 a=3.5 p=15 mult=1 $X=21060 $Y=0 $D=109
M28 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250016 a=3.5 p=15 mult=1 $X=21840 $Y=0 $D=109
M29 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250016 a=3.5 p=15 mult=1 $X=22620 $Y=0 $D=109
M30 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250015 a=3.5 p=15 mult=1 $X=23400 $Y=0 $D=109
M31 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250014 a=3.5 p=15 mult=1 $X=24180 $Y=0 $D=109
M32 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250013 a=3.5 p=15 mult=1 $X=24960 $Y=0 $D=109
M33 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250012 a=3.5 p=15 mult=1 $X=25740 $Y=0 $D=109
M34 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250012 a=3.5 p=15 mult=1 $X=26520 $Y=0 $D=109
M35 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250011 a=3.5 p=15 mult=1 $X=27300 $Y=0 $D=109
M36 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250010 a=3.5 p=15 mult=1 $X=28080 $Y=0 $D=109
M37 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250009 a=3.5 p=15 mult=1 $X=28860 $Y=0 $D=109
M38 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250009 a=3.5 p=15 mult=1 $X=29640 $Y=0 $D=109
M39 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250008 a=3.5 p=15 mult=1 $X=30420 $Y=0 $D=109
M40 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250007 a=3.5 p=15 mult=1 $X=31200 $Y=0 $D=109
M41 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250006 a=3.5 p=15 mult=1 $X=31980 $Y=0 $D=109
M42 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250005 a=3.5 p=15 mult=1 $X=32760 $Y=0 $D=109
M43 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250005 a=3.5 p=15 mult=1 $X=33540 $Y=0 $D=109
M44 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250004 a=3.5 p=15 mult=1 $X=34320 $Y=0 $D=109
M45 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250003 a=3.5 p=15 mult=1 $X=35100 $Y=0 $D=109
M46 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250002 a=3.5 p=15 mult=1 $X=35880 $Y=0 $D=109
M47 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250002 a=3.5 p=15 mult=1 $X=36660 $Y=0 $D=109
M48 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250001 a=3.5 p=15 mult=1 $X=37440 $Y=0 $D=109
M49 2 3 4 2 phv L=0.5 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250000 a=3.5 p=15 mult=1 $X=38220 $Y=0 $D=109
.ENDS
***************************************
.SUBCKT sky130_ef_io__vssa_hvc_clamped_pad VSSD VSSA VDDA VDDIO VCCHIB VCCD VSSIO VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
** N=14084 EP=12 IP=1840 FDC=241
M0 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=15885 $Y=45145 $D=49
M1 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=15885 $Y=137145 $D=49
M2 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=15885 $Y=160145 $D=49
M3 VDDA 8 VSSA VSSA nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250001 sb=250020 a=5 p=21 mult=1 $X=15885 $Y=183145 $D=49
M4 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=17895 $Y=45145 $D=49
M5 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=17895 $Y=137145 $D=49
M6 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=17895 $Y=160145 $D=49
M7 VSSA 8 VDDA VSSA nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250003 sb=250020 a=5 p=21 mult=1 $X=17895 $Y=183145 $D=49
M8 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=20485 $Y=45145 $D=49
M9 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=20485 $Y=137145 $D=49
M10 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=20485 $Y=160145 $D=49
M11 VDDA 8 VSSA VSSA nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250006 sb=250020 a=5 p=21 mult=1 $X=20485 $Y=183145 $D=49
M12 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=22495 $Y=45145 $D=49
M13 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=22495 $Y=137145 $D=49
M14 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=22495 $Y=160145 $D=49
M15 VSSA 8 VDDA VSSA nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250008 sb=250020 a=5 p=21 mult=1 $X=22495 $Y=183145 $D=49
M16 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=45145 $D=49
M17 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=68145 $D=49
M18 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=91145 $D=49
M19 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=114145 $D=49
M20 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=137145 $D=49
M21 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=25085 $Y=160145 $D=49
M22 VDDA 8 VSSA VSSA nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250010 sb=250020 a=5 p=21 mult=1 $X=25085 $Y=183145 $D=49
M23 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=45145 $D=49
M24 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=68145 $D=49
M25 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=91145 $D=49
M26 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=114145 $D=49
M27 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=137145 $D=49
M28 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=27095 $Y=160145 $D=49
M29 VSSA 8 VDDA VSSA nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250012 sb=250020 a=5 p=21 mult=1 $X=27095 $Y=183145 $D=49
M30 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=45145 $D=49
M31 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=68145 $D=49
M32 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=91145 $D=49
M33 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=114145 $D=49
M34 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=137145 $D=49
M35 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=29685 $Y=160145 $D=49
M36 VDDA 8 VSSA VSSA nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250015 sb=250020 a=5 p=21 mult=1 $X=29685 $Y=183145 $D=49
M37 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=45145 $D=49
M38 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=68145 $D=49
M39 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=91145 $D=49
M40 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=114145 $D=49
M41 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=137145 $D=49
M42 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=31695 $Y=160145 $D=49
M43 VSSA 8 VDDA VSSA nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250017 sb=250020 a=5 p=21 mult=1 $X=31695 $Y=183145 $D=49
M44 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=45145 $D=49
M45 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=68145 $D=49
M46 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=91145 $D=49
M47 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=114145 $D=49
M48 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=137145 $D=49
M49 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=34285 $Y=160145 $D=49
M50 VDDA 8 VSSA VSSA nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=34285 $Y=183145 $D=49
M51 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=45145 $D=49
M52 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=68145 $D=49
M53 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=91145 $D=49
M54 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=114145 $D=49
M55 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=137145 $D=49
M56 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=36295 $Y=160145 $D=49
M57 VSSA 8 VDDA VSSA nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=36295 $Y=183145 $D=49
M58 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=45145 $D=49
M59 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=68145 $D=49
M60 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=91145 $D=49
M61 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=114145 $D=49
M62 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=137145 $D=49
M63 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=38885 $Y=160145 $D=49
M64 VDDA 8 VSSA VSSA nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=38885 $Y=183145 $D=49
M65 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=45145 $D=49
M66 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=68145 $D=49
M67 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=91145 $D=49
M68 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=114145 $D=49
M69 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=137145 $D=49
M70 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=40895 $Y=160145 $D=49
M71 VSSA 8 VDDA VSSA nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=40895 $Y=183145 $D=49
M72 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=45145 $D=49
M73 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=68145 $D=49
M74 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=91145 $D=49
M75 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=114145 $D=49
M76 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=137145 $D=49
M77 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=43485 $Y=160145 $D=49
M78 VDDA 8 VSSA VSSA nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=43485 $Y=183145 $D=49
M79 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=45145 $D=49
M80 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=68145 $D=49
M81 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=91145 $D=49
M82 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=114145 $D=49
M83 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=137145 $D=49
M84 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=45495 $Y=160145 $D=49
M85 VSSA 8 VDDA VSSA nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=45495 $Y=183145 $D=49
M86 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=45145 $D=49
M87 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=68145 $D=49
M88 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=91145 $D=49
M89 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=114145 $D=49
M90 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=137145 $D=49
M91 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=48085 $Y=160145 $D=49
M92 VDDA 8 VSSA VSSA nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250017 a=5 p=21 mult=1 $X=48085 $Y=183145 $D=49
M93 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=45145 $D=49
M94 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=68145 $D=49
M95 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=91145 $D=49
M96 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=114145 $D=49
M97 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=137145 $D=49
M98 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=50095 $Y=160145 $D=49
M99 VSSA 8 VDDA VSSA nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250015 a=5 p=21 mult=1 $X=50095 $Y=183145 $D=49
M100 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=45145 $D=49
M101 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=68145 $D=49
M102 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=91145 $D=49
M103 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=114145 $D=49
M104 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=137145 $D=49
M105 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=52685 $Y=160145 $D=49
M106 VDDA 8 VSSA VSSA nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250012 a=5 p=21 mult=1 $X=52685 $Y=183145 $D=49
M107 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=45145 $D=49
M108 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=68145 $D=49
M109 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=91145 $D=49
M110 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=114145 $D=49
M111 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=137145 $D=49
M112 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=54695 $Y=160145 $D=49
M113 VSSA 8 VDDA VSSA nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250010 a=5 p=21 mult=1 $X=54695 $Y=183145 $D=49
M114 8 6 VSSA VSSA nhv L=0.5 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 r=14 sa=250000 sb=250011 a=3.5 p=15 mult=1 $X=54915 $Y=30545 $D=49
M115 VSSA 6 8 VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250001 sb=250010 a=3.5 p=15 mult=1 $X=55695 $Y=30545 $D=49
M116 8 6 VSSA VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250009 a=3.5 p=15 mult=1 $X=56475 $Y=30545 $D=49
M117 VSSA 6 8 VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250009 a=3.5 p=15 mult=1 $X=57255 $Y=30545 $D=49
M118 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=45145 $D=49
M119 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=68145 $D=49
M120 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=91145 $D=49
M121 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=114145 $D=49
M122 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=137145 $D=49
M123 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=57285 $Y=160145 $D=49
M124 VDDA 8 VSSA VSSA nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250008 a=5 p=21 mult=1 $X=57285 $Y=183145 $D=49
M125 8 6 VSSA VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250003 sb=250008 a=3.5 p=15 mult=1 $X=58035 $Y=30545 $D=49
M126 VSSA 6 8 VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250004 sb=250007 a=3.5 p=15 mult=1 $X=58815 $Y=30545 $D=49
M127 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=45145 $D=49
M128 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=68145 $D=49
M129 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=91145 $D=49
M130 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=114145 $D=49
M131 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=137145 $D=49
M132 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=59295 $Y=160145 $D=49
M133 VSSA 8 VDDA VSSA nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250006 a=5 p=21 mult=1 $X=59295 $Y=183145 $D=49
M134 8 6 VSSA VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250006 a=3.5 p=15 mult=1 $X=59595 $Y=30545 $D=49
M135 VSSA 6 8 VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250005 a=3.5 p=15 mult=1 $X=60375 $Y=30545 $D=49
M136 8 6 VSSA VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250006 sb=250005 a=3.5 p=15 mult=1 $X=61155 $Y=30545 $D=49
M137 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=45145 $D=49
M138 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=68145 $D=49
M139 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=91145 $D=49
M140 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=114145 $D=49
M141 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=137145 $D=49
M142 VDDA 8 VSSA VSSA nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=61885 $Y=160145 $D=49
M143 VDDA 8 VSSA VSSA nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250003 a=5 p=21 mult=1 $X=61885 $Y=183145 $D=49
M144 VSSA 6 8 VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250007 sb=250004 a=3.5 p=15 mult=1 $X=61935 $Y=30545 $D=49
M145 8 6 VSSA VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250008 sb=250003 a=3.5 p=15 mult=1 $X=62715 $Y=30545 $D=49
M146 VSSA 6 8 VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250002 a=3.5 p=15 mult=1 $X=63495 $Y=30545 $D=49
M147 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=45145 $D=49
M148 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=68145 $D=49
M149 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=91145 $D=49
M150 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=114145 $D=49
M151 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=137145 $D=49
M152 VSSA 8 VDDA VSSA nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=63895 $Y=160145 $D=49
M153 VSSA 8 VDDA VSSA nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250001 a=5 p=21 mult=1 $X=63895 $Y=183145 $D=49
M154 8 6 VSSA VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250002 a=3.5 p=15 mult=1 $X=64275 $Y=30545 $D=49
M155 VSSA 6 8 VSSA nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250010 sb=250001 a=3.5 p=15 mult=1 $X=65055 $Y=30545 $D=49
M156 8 6 VSSA VSSA nhv L=0.5 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250011 sb=250000 a=3.5 p=15 mult=1 $X=65835 $Y=30545 $D=49
X157 VSSA VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=51225 $Y=19700 $D=150
X158 VSSA VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=51225 $Y=43275 $D=150
X159 VSSA VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=64770 $Y=38800 $D=150
X160 VSSA VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=68375 $Y=195640 $D=150
X161 VSSD VDDIO Dpar a=126.883 p=0 m=1 $[nwdiode] $X=8835 $Y=41140 $D=189
X162 VSSD VDDA Dpar a=376.949 p=101.73 m=1 $[nwdiode] $X=4400 $Y=26890 $D=191
X163 VSSD VDDIO Dpar a=10358.7 p=619.08 m=1 $[dnwdiode_psub] $X=9500 $Y=131800 $D=193
X164 VSSA VDDIO Dpar a=137.463 p=47.72 m=1 $[dnwdiode_pw] $X=53530 $Y=29360 $D=194
X165 VSSA VDDIO Dpar a=8184.99 p=443.22 m=1 $[dnwdiode_pw] $X=10695 $Y=43000 $D=194
X166 VSSA VDDIO Dpar a=1172.63 p=163 m=1 $[dnwdiode_pw] $X=13380 $Y=170 $D=194
R167 5 7 L=1550 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=1070 $Y=41405 $D=257
R168 5 VDDA L=700 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=9500 $Y=72320 $D=257
R169 7 6 L=470 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=70725 $Y=40980 $D=257
R170 VSSA VSSA 0.01 m=1 $[short] $X=6670 $Y=103310 $D=286
X253 VSSA 6 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 $T=61815 25110 0 180 $X=57370 $Y=19930
X254 VSSA 6 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 7170 0 180 $X=13630 $Y=420
X255 VSSA 6 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 13390 0 180 $X=13630 $Y=6640
X256 VSSA 6 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 19610 0 180 $X=13630 $Y=12860
X257 VSSA 6 sky130_fd_io__sio_clamp_pcap_4x5 $T=68720 25830 0 180 $X=62430 $Y=19080
X268 VSSA 6 sky130_fd_io__esd_rcclamp_nfetcap $T=68470 7080 0 180 $X=58430 $Y=420
X269 VSSA 6 sky130_fd_io__esd_rcclamp_nfetcap $T=68470 13300 0 180 $X=58430 $Y=6640
X270 VSSA 6 sky130_fd_io__esd_rcclamp_nfetcap $T=68470 19520 0 180 $X=58430 $Y=12860
X271 VSSA 6 ICV_2 $T=29430 7080 0 180 $X=19390 $Y=420
X272 VSSA 6 ICV_2 $T=29430 13300 0 180 $X=19390 $Y=6640
X273 VSSA 6 ICV_2 $T=29430 19520 0 180 $X=19390 $Y=12860
X274 VSSA 6 ICV_2 $T=48950 7080 0 180 $X=38910 $Y=420
X275 VSSA 6 ICV_2 $T=48950 13300 0 180 $X=38910 $Y=6640
X276 VSSA 6 ICV_2 $T=48950 19520 0 180 $X=38910 $Y=12860
X283 VDDA 6 8 sky130_fd_pr__pfet_01v8__example_55959141808665 $T=6340 27765 0 0 $X=5745 $Y=27435
.ENDS
***************************************
