magic
tech sky130A
magscale 1 2
timestamp 1613304635
<< obsactive >>
rect 1000 1000 76296 90247
<< obsli1 >>
rect 1000 1000 76356 90307
<< obsm1 >>
rect 1000 1000 76356 90307
<< obsm2 >>
rect 1000 1000 76356 90307
<< metal3 >>
rect 71856 90307 72204 90428
rect 76208 90410 77260 90428
rect 76208 90307 76944 90410
rect 0 86557 920 86617
rect 0 85429 920 85489
rect 0 83729 920 83789
rect 0 82601 920 82661
rect 0 80901 920 80961
rect 0 79773 920 79833
rect 0 78073 920 78133
rect 0 20225 920 20285
rect 0 18525 920 18585
rect 76356 90088 76944 90307
rect 77248 90088 77260 90410
rect 76356 90080 77260 90088
rect 76436 89653 77296 89713
rect 76356 88926 76810 88932
rect 76356 88724 76500 88926
rect 76804 88724 76810 88926
rect 76356 88720 76810 88724
rect 76436 29382 77296 29442
rect 76436 27682 77296 27742
rect 76436 26554 77296 26614
rect 76436 24854 77296 24914
rect 76436 23726 77296 23786
rect 76436 22026 77296 22086
rect 76436 20898 77296 20958
<< obsm3 >>
rect 1000 1000 76356 90307
<< via3 >>
rect 76944 90088 77248 90410
rect 76500 88724 76804 88926
<< metal4 >>
rect 18805 90407 18865 91247
rect 20053 90407 20113 91247
rect 21301 90407 21361 91247
rect 22549 90407 22609 91247
rect 23797 90407 23857 91247
rect 25045 90407 25105 91247
rect 26293 90407 26353 91247
rect 27541 90407 27601 91247
rect 28789 90407 28849 91247
rect 30037 90407 30097 91247
rect 31285 90407 31345 91247
rect 32533 90407 32593 91247
rect 33781 90407 33841 91247
rect 35029 90407 35089 91247
rect 36277 90407 36337 91247
rect 37525 90407 37585 91247
rect 38773 90407 38833 91247
rect 40021 90407 40081 91247
rect 41269 90407 41329 91247
rect 42517 90407 42577 91247
rect 43765 90407 43825 91247
rect 45013 90407 45073 91247
rect 46261 90407 46321 91247
rect 47509 90407 47569 91247
rect 48757 90407 48817 91247
rect 50005 90407 50065 91247
rect 51253 90407 51313 91247
rect 52501 90407 52561 91247
rect 53749 90407 53809 91247
rect 54997 90407 55057 91247
rect 56245 90407 56305 91247
rect 57493 90407 57553 91247
rect 68578 90407 68638 91247
rect 73573 90407 73633 91247
rect 76938 90410 77262 90428
rect 76938 90088 76944 90410
rect 77248 90088 77262 90410
rect 76494 88926 76814 88936
rect 76494 88724 76500 88926
rect 76804 88724 76814 88926
rect 3803 0 3863 920
rect 6802 0 6862 920
rect 7970 0 8030 920
rect 9138 0 9198 920
rect 10306 0 10366 920
rect 11474 0 11534 920
rect 12642 0 12702 920
rect 12766 0 12826 920
rect 13810 0 13870 920
rect 13934 0 13994 920
rect 14978 0 15038 920
rect 15102 0 15162 920
rect 16146 0 16206 920
rect 16270 0 16330 920
rect 17314 0 17374 920
rect 17438 0 17498 920
rect 18482 0 18542 920
rect 18606 0 18666 920
rect 19650 0 19710 920
rect 19774 0 19834 920
rect 20818 0 20878 920
rect 20942 0 21002 920
rect 21986 0 22046 920
rect 22110 0 22170 920
rect 23154 0 23214 920
rect 23278 0 23338 920
rect 24322 0 24382 920
rect 24446 0 24506 920
rect 25490 0 25550 920
rect 25614 0 25674 920
rect 26658 0 26718 920
rect 26782 0 26842 920
rect 27826 0 27886 920
rect 27950 0 28010 920
rect 28994 0 29054 920
rect 29118 0 29178 920
rect 30162 0 30222 920
rect 30286 0 30346 920
rect 31330 0 31390 920
rect 31454 0 31514 920
rect 32498 0 32558 920
rect 32622 0 32682 920
rect 33666 0 33726 920
rect 33790 0 33850 920
rect 34834 0 34894 920
rect 34958 0 35018 920
rect 36002 0 36062 920
rect 36126 0 36186 920
rect 37170 0 37230 920
rect 37294 0 37354 920
rect 38338 0 38398 920
rect 38462 0 38522 920
rect 39506 0 39566 920
rect 39630 0 39690 920
rect 40674 0 40734 920
rect 40798 0 40858 920
rect 41842 0 41902 920
rect 41966 0 42026 920
rect 43010 0 43070 920
rect 43134 0 43194 920
rect 44178 0 44238 920
rect 44302 0 44362 920
rect 45346 0 45406 920
rect 45470 0 45530 920
rect 46514 0 46574 920
rect 46638 0 46698 920
rect 47682 0 47742 920
rect 47806 0 47866 920
rect 48850 0 48910 920
rect 48974 0 49034 920
rect 76494 734 76814 88724
rect 76938 812 77262 90088
<< obsm4 >>
rect 1000 1000 76356 90307
<< labels >>
rlabel metal4 s 12642 0 12702 920 6 din0[0]
port 1 nsew default input
rlabel metal4 s 13810 0 13870 920 6 din0[1]
port 2 nsew default input
rlabel metal4 s 14978 0 15038 920 6 din0[2]
port 3 nsew default input
rlabel metal4 s 16146 0 16206 920 6 din0[3]
port 4 nsew default input
rlabel metal4 s 17314 0 17374 920 6 din0[4]
port 5 nsew default input
rlabel metal4 s 18482 0 18542 920 6 din0[5]
port 6 nsew default input
rlabel metal4 s 19650 0 19710 920 6 din0[6]
port 7 nsew default input
rlabel metal4 s 20818 0 20878 920 6 din0[7]
port 8 nsew default input
rlabel metal4 s 21986 0 22046 920 6 din0[8]
port 9 nsew default input
rlabel metal4 s 23154 0 23214 920 6 din0[9]
port 10 nsew default input
rlabel metal4 s 24322 0 24382 920 6 din0[10]
port 11 nsew default input
rlabel metal4 s 25490 0 25550 920 6 din0[11]
port 12 nsew default input
rlabel metal4 s 26658 0 26718 920 6 din0[12]
port 13 nsew default input
rlabel metal4 s 27826 0 27886 920 6 din0[13]
port 14 nsew default input
rlabel metal4 s 28994 0 29054 920 6 din0[14]
port 15 nsew default input
rlabel metal4 s 30162 0 30222 920 6 din0[15]
port 16 nsew default input
rlabel metal4 s 31330 0 31390 920 6 din0[16]
port 17 nsew default input
rlabel metal4 s 32498 0 32558 920 6 din0[17]
port 18 nsew default input
rlabel metal4 s 33666 0 33726 920 6 din0[18]
port 19 nsew default input
rlabel metal4 s 34834 0 34894 920 6 din0[19]
port 20 nsew default input
rlabel metal4 s 36002 0 36062 920 6 din0[20]
port 21 nsew default input
rlabel metal4 s 37170 0 37230 920 6 din0[21]
port 22 nsew default input
rlabel metal4 s 38338 0 38398 920 6 din0[22]
port 23 nsew default input
rlabel metal4 s 39506 0 39566 920 6 din0[23]
port 24 nsew default input
rlabel metal4 s 40674 0 40734 920 6 din0[24]
port 25 nsew default input
rlabel metal4 s 41842 0 41902 920 6 din0[25]
port 26 nsew default input
rlabel metal4 s 43010 0 43070 920 6 din0[26]
port 27 nsew default input
rlabel metal4 s 44178 0 44238 920 6 din0[27]
port 28 nsew default input
rlabel metal4 s 45346 0 45406 920 6 din0[28]
port 29 nsew default input
rlabel metal4 s 46514 0 46574 920 6 din0[29]
port 30 nsew default input
rlabel metal4 s 47682 0 47742 920 6 din0[30]
port 31 nsew default input
rlabel metal4 s 48850 0 48910 920 6 din0[31]
port 32 nsew default input
rlabel metal4 s 6802 0 6862 920 6 addr0[0]
port 33 nsew default input
rlabel metal3 s 0 78073 920 78133 6 addr0[1]
port 34 nsew default input
rlabel metal3 s 0 79773 920 79833 6 addr0[2]
port 35 nsew default input
rlabel metal3 s 0 80901 920 80961 6 addr0[3]
port 36 nsew default input
rlabel metal3 s 0 82601 920 82661 6 addr0[4]
port 37 nsew default input
rlabel metal3 s 0 83729 920 83789 6 addr0[5]
port 38 nsew default input
rlabel metal3 s 0 85429 920 85489 6 addr0[6]
port 39 nsew default input
rlabel metal3 s 0 86557 920 86617 6 addr0[7]
port 40 nsew default input
rlabel metal4 s 68578 90407 68638 91247 6 addr1[0]
port 41 nsew default input
rlabel metal3 s 76436 29382 77296 29442 6 addr1[1]
port 42 nsew default input
rlabel metal3 s 76436 27682 77296 27742 6 addr1[2]
port 43 nsew default input
rlabel metal3 s 76436 26554 77296 26614 6 addr1[3]
port 44 nsew default input
rlabel metal3 s 76436 24854 77296 24914 6 addr1[4]
port 45 nsew default input
rlabel metal3 s 76436 23726 77296 23786 6 addr1[5]
port 46 nsew default input
rlabel metal3 s 76436 22026 77296 22086 6 addr1[6]
port 47 nsew default input
rlabel metal3 s 76436 20898 77296 20958 6 addr1[7]
port 48 nsew default input
rlabel metal3 s 0 18525 920 18585 6 csb0
port 49 nsew default input
rlabel metal3 s 76436 89653 77296 89713 6 csb1
port 50 nsew default input
rlabel metal3 s 0 20225 920 20285 6 web0
port 51 nsew default input
rlabel metal4 s 3803 0 3863 920 6 clk0
port 52 nsew default input
rlabel metal4 s 73573 90407 73633 91247 6 clk1
port 53 nsew default input
rlabel metal4 s 7970 0 8030 920 6 wmask0[0]
port 54 nsew default input
rlabel metal4 s 9138 0 9198 920 6 wmask0[1]
port 55 nsew default input
rlabel metal4 s 10306 0 10366 920 6 wmask0[2]
port 56 nsew default input
rlabel metal4 s 11474 0 11534 920 6 wmask0[3]
port 57 nsew default input
rlabel metal4 s 12766 0 12826 920 6 dout0[0]
port 58 nsew default output
rlabel metal4 s 13934 0 13994 920 6 dout0[1]
port 59 nsew default output
rlabel metal4 s 15102 0 15162 920 6 dout0[2]
port 60 nsew default output
rlabel metal4 s 16270 0 16330 920 6 dout0[3]
port 61 nsew default output
rlabel metal4 s 17438 0 17498 920 6 dout0[4]
port 62 nsew default output
rlabel metal4 s 18606 0 18666 920 6 dout0[5]
port 63 nsew default output
rlabel metal4 s 19774 0 19834 920 6 dout0[6]
port 64 nsew default output
rlabel metal4 s 20942 0 21002 920 6 dout0[7]
port 65 nsew default output
rlabel metal4 s 22110 0 22170 920 6 dout0[8]
port 66 nsew default output
rlabel metal4 s 23278 0 23338 920 6 dout0[9]
port 67 nsew default output
rlabel metal4 s 24446 0 24506 920 6 dout0[10]
port 68 nsew default output
rlabel metal4 s 25614 0 25674 920 6 dout0[11]
port 69 nsew default output
rlabel metal4 s 26782 0 26842 920 6 dout0[12]
port 70 nsew default output
rlabel metal4 s 27950 0 28010 920 6 dout0[13]
port 71 nsew default output
rlabel metal4 s 29118 0 29178 920 6 dout0[14]
port 72 nsew default output
rlabel metal4 s 30286 0 30346 920 6 dout0[15]
port 73 nsew default output
rlabel metal4 s 31454 0 31514 920 6 dout0[16]
port 74 nsew default output
rlabel metal4 s 32622 0 32682 920 6 dout0[17]
port 75 nsew default output
rlabel metal4 s 33790 0 33850 920 6 dout0[18]
port 76 nsew default output
rlabel metal4 s 34958 0 35018 920 6 dout0[19]
port 77 nsew default output
rlabel metal4 s 36126 0 36186 920 6 dout0[20]
port 78 nsew default output
rlabel metal4 s 37294 0 37354 920 6 dout0[21]
port 79 nsew default output
rlabel metal4 s 38462 0 38522 920 6 dout0[22]
port 80 nsew default output
rlabel metal4 s 39630 0 39690 920 6 dout0[23]
port 81 nsew default output
rlabel metal4 s 40798 0 40858 920 6 dout0[24]
port 82 nsew default output
rlabel metal4 s 41966 0 42026 920 6 dout0[25]
port 83 nsew default output
rlabel metal4 s 43134 0 43194 920 6 dout0[26]
port 84 nsew default output
rlabel metal4 s 44302 0 44362 920 6 dout0[27]
port 85 nsew default output
rlabel metal4 s 45470 0 45530 920 6 dout0[28]
port 86 nsew default output
rlabel metal4 s 46638 0 46698 920 6 dout0[29]
port 87 nsew default output
rlabel metal4 s 47806 0 47866 920 6 dout0[30]
port 88 nsew default output
rlabel metal4 s 48974 0 49034 920 6 dout0[31]
port 89 nsew default output
rlabel metal4 s 18805 90407 18865 91247 6 dout1[0]
port 90 nsew default output
rlabel metal4 s 20053 90407 20113 91247 6 dout1[1]
port 91 nsew default output
rlabel metal4 s 21301 90407 21361 91247 6 dout1[2]
port 92 nsew default output
rlabel metal4 s 22549 90407 22609 91247 6 dout1[3]
port 93 nsew default output
rlabel metal4 s 23797 90407 23857 91247 6 dout1[4]
port 94 nsew default output
rlabel metal4 s 25045 90407 25105 91247 6 dout1[5]
port 95 nsew default output
rlabel metal4 s 26293 90407 26353 91247 6 dout1[6]
port 96 nsew default output
rlabel metal4 s 27541 90407 27601 91247 6 dout1[7]
port 97 nsew default output
rlabel metal4 s 28789 90407 28849 91247 6 dout1[8]
port 98 nsew default output
rlabel metal4 s 30037 90407 30097 91247 6 dout1[9]
port 99 nsew default output
rlabel metal4 s 31285 90407 31345 91247 6 dout1[10]
port 100 nsew default output
rlabel metal4 s 32533 90407 32593 91247 6 dout1[11]
port 101 nsew default output
rlabel metal4 s 33781 90407 33841 91247 6 dout1[12]
port 102 nsew default output
rlabel metal4 s 35029 90407 35089 91247 6 dout1[13]
port 103 nsew default output
rlabel metal4 s 36277 90407 36337 91247 6 dout1[14]
port 104 nsew default output
rlabel metal4 s 37525 90407 37585 91247 6 dout1[15]
port 105 nsew default output
rlabel metal4 s 38773 90407 38833 91247 6 dout1[16]
port 106 nsew default output
rlabel metal4 s 40021 90407 40081 91247 6 dout1[17]
port 107 nsew default output
rlabel metal4 s 41269 90407 41329 91247 6 dout1[18]
port 108 nsew default output
rlabel metal4 s 42517 90407 42577 91247 6 dout1[19]
port 109 nsew default output
rlabel metal4 s 43765 90407 43825 91247 6 dout1[20]
port 110 nsew default output
rlabel metal4 s 45013 90407 45073 91247 6 dout1[21]
port 111 nsew default output
rlabel metal4 s 46261 90407 46321 91247 6 dout1[22]
port 112 nsew default output
rlabel metal4 s 47509 90407 47569 91247 6 dout1[23]
port 113 nsew default output
rlabel metal4 s 48757 90407 48817 91247 6 dout1[24]
port 114 nsew default output
rlabel metal4 s 50005 90407 50065 91247 6 dout1[25]
port 115 nsew default output
rlabel metal4 s 51253 90407 51313 91247 6 dout1[26]
port 116 nsew default output
rlabel metal4 s 52501 90407 52561 91247 6 dout1[27]
port 117 nsew default output
rlabel metal4 s 53749 90407 53809 91247 6 dout1[28]
port 118 nsew default output
rlabel metal4 s 54997 90407 55057 91247 6 dout1[29]
port 119 nsew default output
rlabel metal4 s 56245 90407 56305 91247 6 dout1[30]
port 120 nsew default output
rlabel metal4 s 57493 90407 57553 91247 6 dout1[31]
port 121 nsew default output
rlabel metal4 s 76494 734 76814 88936 6 vdd
port 122 nsew power bidirectional
rlabel via3 s 76500 88724 76804 88926 6 vdd
port 122 nsew power bidirectional
rlabel metal3 s 76208 88720 76810 88932 6 vdd
port 122 nsew power bidirectional
rlabel metal3 s 71856 90216 72204 90428 6 gnd
port 123 nsew ground bidirectional
rlabel metal4 s 76938 812 77262 90428 6 gnd
port 123 nsew ground bidirectional
rlabel via3 s 76944 90088 77248 90410 6 gnd
port 123 nsew ground bidirectional
rlabel metal3 s 76208 90080 77260 90428 6 gnd
port 123 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 77296 91247
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE ../gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_END 13299042
string GDS_START 13275442
<< end >>
