magic
tech sky130A
magscale 1 2
timestamp 1608143558
<< obsli1 >>
rect 55873 17940 55907 18003
rect 64429 17969 65659 18003
rect 70133 17969 70351 18003
rect 64429 17940 64463 17969
rect 70317 17940 70351 17969
rect 79885 17969 80195 18003
rect 79885 17940 79919 17969
rect 80161 17940 80195 17969
rect 92581 17969 93075 18003
rect 113097 17969 113959 18003
rect 92581 17940 92615 17969
rect 93041 17940 93075 17969
rect 113925 17940 113959 17969
rect 118617 17940 118651 18003
rect 1104 629 198812 17940
<< obsm1 >>
rect 55861 18000 55919 18009
rect 65613 18000 65671 18009
rect 68830 18000 68894 18012
rect 55861 17972 65472 18000
rect 55861 17963 55919 17972
rect 40770 17940 40834 17944
rect 65337 17940 65395 17941
rect 65444 17940 65472 17972
rect 65613 17972 68894 18000
rect 65613 17963 65671 17972
rect 68830 17960 68894 17972
rect 69106 18000 69170 18012
rect 70121 18000 70179 18009
rect 69106 17972 70179 18000
rect 69106 17960 69170 17972
rect 70121 17963 70179 17972
rect 70210 18000 70274 18012
rect 113085 18000 113143 18009
rect 70210 17972 113143 18000
rect 70210 17960 70274 17972
rect 113085 17963 113143 17972
rect 113174 18000 113238 18012
rect 118605 18000 118663 18009
rect 113174 17972 118663 18000
rect 113174 17960 113238 17972
rect 118605 17963 118663 17972
rect 65521 17940 65579 17941
rect 74718 17940 74782 17944
rect 74810 17940 74874 17944
rect 79873 17940 79931 17941
rect 80149 17940 80207 17941
rect 89717 17940 89775 17941
rect 89806 17940 89870 17944
rect 91922 17940 91986 17944
rect 92017 17940 92075 17941
rect 92753 17940 92811 17941
rect 101398 17940 101462 17944
rect 101858 17940 101922 17944
rect 103698 17940 103762 17944
rect 126330 17940 126394 17944
rect 198 620 199810 17940
<< metal2 >>
rect 202 17940 258 18400
rect 570 17940 626 18400
rect 1030 17940 1086 18400
rect 1490 17940 1546 18400
rect 1858 17940 1914 18400
rect 2318 17940 2374 18400
rect 2778 17940 2834 18400
rect 3238 17940 3294 18400
rect 3606 17940 3662 18400
rect 4066 17940 4122 18400
rect 4526 17940 4582 18400
rect 4986 17940 5042 18400
rect 5354 17940 5410 18400
rect 5814 17940 5870 18400
rect 6274 17940 6330 18400
rect 6734 17940 6790 18400
rect 7102 17940 7158 18400
rect 7562 17940 7618 18400
rect 8022 17940 8078 18400
rect 8390 17940 8446 18400
rect 8850 17940 8906 18400
rect 9310 17940 9366 18400
rect 9770 17940 9826 18400
rect 10138 17940 10194 18400
rect 10598 17940 10654 18400
rect 11058 17940 11114 18400
rect 11518 17940 11574 18400
rect 11886 17940 11942 18400
rect 12346 17940 12402 18400
rect 12806 17940 12862 18400
rect 13266 17940 13322 18400
rect 13634 17940 13690 18400
rect 14094 17940 14150 18400
rect 14554 17940 14610 18400
rect 15014 17940 15070 18400
rect 15382 17940 15438 18400
rect 15842 17940 15898 18400
rect 16302 17940 16358 18400
rect 16670 17940 16726 18400
rect 17130 17940 17186 18400
rect 17590 17940 17646 18400
rect 18050 17940 18106 18400
rect 18418 17940 18474 18400
rect 18878 17940 18934 18400
rect 19338 17940 19394 18400
rect 19798 17940 19854 18400
rect 20166 17940 20222 18400
rect 20626 17940 20682 18400
rect 21086 17940 21142 18400
rect 21546 17940 21602 18400
rect 21914 17940 21970 18400
rect 22374 17940 22430 18400
rect 22834 17940 22890 18400
rect 23294 17940 23350 18400
rect 23662 17940 23718 18400
rect 24122 17940 24178 18400
rect 24582 17940 24638 18400
rect 24950 17940 25006 18400
rect 25410 17940 25466 18400
rect 25870 17940 25926 18400
rect 26330 17940 26386 18400
rect 26698 17940 26754 18400
rect 27158 17940 27214 18400
rect 27618 17940 27674 18400
rect 28078 17940 28134 18400
rect 28446 17940 28502 18400
rect 28906 17940 28962 18400
rect 29366 17940 29422 18400
rect 29826 17940 29882 18400
rect 30194 17940 30250 18400
rect 30654 17940 30710 18400
rect 31114 17940 31170 18400
rect 31574 17940 31630 18400
rect 31942 17940 31998 18400
rect 32402 17940 32458 18400
rect 32862 17940 32918 18400
rect 33230 17940 33286 18400
rect 33690 17940 33746 18400
rect 34150 17940 34206 18400
rect 34610 17940 34666 18400
rect 34978 17940 35034 18400
rect 35438 17940 35494 18400
rect 35898 17940 35954 18400
rect 36358 17940 36414 18400
rect 36726 17940 36782 18400
rect 37186 17940 37242 18400
rect 37646 17940 37702 18400
rect 38106 17940 38162 18400
rect 38474 17940 38530 18400
rect 38934 17940 38990 18400
rect 39394 17940 39450 18400
rect 39854 17940 39910 18400
rect 40222 17940 40278 18400
rect 40682 17940 40738 18400
rect 41142 17940 41198 18400
rect 41510 17940 41566 18400
rect 41970 17940 42026 18400
rect 42430 17940 42486 18400
rect 42890 17940 42946 18400
rect 43258 17940 43314 18400
rect 43718 17940 43774 18400
rect 44178 17940 44234 18400
rect 44638 17940 44694 18400
rect 45006 17940 45062 18400
rect 45466 17940 45522 18400
rect 45926 17940 45982 18400
rect 46386 17940 46442 18400
rect 46754 17940 46810 18400
rect 47214 17940 47270 18400
rect 47674 17940 47730 18400
rect 48134 17940 48190 18400
rect 48502 17940 48558 18400
rect 48962 17940 49018 18400
rect 49422 17940 49478 18400
rect 49790 17940 49846 18400
rect 50250 17940 50306 18400
rect 50710 17940 50766 18400
rect 51170 17940 51226 18400
rect 51538 17940 51594 18400
rect 51998 17940 52054 18400
rect 52458 17940 52514 18400
rect 52918 17940 52974 18400
rect 53286 17940 53342 18400
rect 53746 17940 53802 18400
rect 54206 17940 54262 18400
rect 54666 17940 54722 18400
rect 55034 17940 55090 18400
rect 55494 17940 55550 18400
rect 55954 17940 56010 18400
rect 56322 17940 56378 18400
rect 56782 17940 56838 18400
rect 57242 17940 57298 18400
rect 57702 17940 57758 18400
rect 58070 17940 58126 18400
rect 58530 17940 58586 18400
rect 58990 17940 59046 18400
rect 59450 17940 59506 18400
rect 59818 17940 59874 18400
rect 60278 17940 60334 18400
rect 60738 17940 60794 18400
rect 61198 17940 61254 18400
rect 61566 17940 61622 18400
rect 62026 17940 62082 18400
rect 62486 17940 62542 18400
rect 62946 17940 63002 18400
rect 63314 17940 63370 18400
rect 63774 17940 63830 18400
rect 64234 17940 64290 18400
rect 64602 17940 64658 18400
rect 65062 17940 65118 18400
rect 65522 17940 65578 18400
rect 65982 17940 66038 18400
rect 66350 17940 66406 18400
rect 66810 17940 66866 18400
rect 67270 17940 67326 18400
rect 67730 17940 67786 18400
rect 68098 17940 68154 18400
rect 68558 17940 68614 18400
rect 69018 17940 69074 18400
rect 69478 17940 69534 18400
rect 69846 17940 69902 18400
rect 70306 17940 70362 18400
rect 70766 17940 70822 18400
rect 71226 17940 71282 18400
rect 71594 17940 71650 18400
rect 72054 17940 72110 18400
rect 72514 17940 72570 18400
rect 72882 17940 72938 18400
rect 73342 17940 73398 18400
rect 73802 17940 73858 18400
rect 74262 17940 74318 18400
rect 74630 17940 74686 18400
rect 75090 17940 75146 18400
rect 75550 17940 75606 18400
rect 76010 17940 76066 18400
rect 76378 17940 76434 18400
rect 76838 17940 76894 18400
rect 77298 17940 77354 18400
rect 77758 17940 77814 18400
rect 78126 17940 78182 18400
rect 78586 17940 78642 18400
rect 79046 17940 79102 18400
rect 79506 17940 79562 18400
rect 79874 17940 79930 18400
rect 80334 17940 80390 18400
rect 80794 17940 80850 18400
rect 81162 17940 81218 18400
rect 81622 17940 81678 18400
rect 82082 17940 82138 18400
rect 82542 17940 82598 18400
rect 82910 17940 82966 18400
rect 83370 17940 83426 18400
rect 83830 17940 83886 18400
rect 84290 17940 84346 18400
rect 84658 17940 84714 18400
rect 85118 17940 85174 18400
rect 85578 17940 85634 18400
rect 86038 17940 86094 18400
rect 86406 17940 86462 18400
rect 86866 17940 86922 18400
rect 87326 17940 87382 18400
rect 87786 17940 87842 18400
rect 88154 17940 88210 18400
rect 88614 17940 88670 18400
rect 89074 17940 89130 18400
rect 89442 17940 89498 18400
rect 89902 17940 89958 18400
rect 90362 17940 90418 18400
rect 90822 17940 90878 18400
rect 91190 17940 91246 18400
rect 91650 17940 91706 18400
rect 92110 17940 92166 18400
rect 92570 17940 92626 18400
rect 92938 17940 92994 18400
rect 93398 17940 93454 18400
rect 93858 17940 93914 18400
rect 94318 17940 94374 18400
rect 94686 17940 94742 18400
rect 95146 17940 95202 18400
rect 95606 17940 95662 18400
rect 96066 17940 96122 18400
rect 96434 17940 96490 18400
rect 96894 17940 96950 18400
rect 97354 17940 97410 18400
rect 97722 17940 97778 18400
rect 98182 17940 98238 18400
rect 98642 17940 98698 18400
rect 99102 17940 99158 18400
rect 99470 17940 99526 18400
rect 99930 17940 99986 18400
rect 100390 17940 100446 18400
rect 100850 17940 100906 18400
rect 101218 17940 101274 18400
rect 101678 17940 101734 18400
rect 102138 17940 102194 18400
rect 102598 17940 102654 18400
rect 102966 17940 103022 18400
rect 103426 17940 103482 18400
rect 103886 17940 103942 18400
rect 104254 17940 104310 18400
rect 104714 17940 104770 18400
rect 105174 17940 105230 18400
rect 105634 17940 105690 18400
rect 106002 17940 106058 18400
rect 106462 17940 106518 18400
rect 106922 17940 106978 18400
rect 107382 17940 107438 18400
rect 107750 17940 107806 18400
rect 108210 17940 108266 18400
rect 108670 17940 108726 18400
rect 109130 17940 109186 18400
rect 109498 17940 109554 18400
rect 109958 17940 110014 18400
rect 110418 17940 110474 18400
rect 110878 17940 110934 18400
rect 111246 17940 111302 18400
rect 111706 17940 111762 18400
rect 112166 17940 112222 18400
rect 112534 17940 112590 18400
rect 112994 17940 113050 18400
rect 113454 17940 113510 18400
rect 113914 17940 113970 18400
rect 114282 17940 114338 18400
rect 114742 17940 114798 18400
rect 115202 17940 115258 18400
rect 115662 17940 115718 18400
rect 116030 17940 116086 18400
rect 116490 17940 116546 18400
rect 116950 17940 117006 18400
rect 117410 17940 117466 18400
rect 117778 17940 117834 18400
rect 118238 17940 118294 18400
rect 118698 17940 118754 18400
rect 119158 17940 119214 18400
rect 119526 17940 119582 18400
rect 119986 17940 120042 18400
rect 120446 17940 120502 18400
rect 120814 17940 120870 18400
rect 121274 17940 121330 18400
rect 121734 17940 121790 18400
rect 122194 17940 122250 18400
rect 122562 17940 122618 18400
rect 123022 17940 123078 18400
rect 123482 17940 123538 18400
rect 123942 17940 123998 18400
rect 124310 17940 124366 18400
rect 124770 17940 124826 18400
rect 125230 17940 125286 18400
rect 125690 17940 125746 18400
rect 126058 17940 126114 18400
rect 126518 17940 126574 18400
rect 126978 17940 127034 18400
rect 127438 17940 127494 18400
rect 127806 17940 127862 18400
rect 128266 17940 128322 18400
rect 128726 17940 128782 18400
rect 129094 17940 129150 18400
rect 129554 17940 129610 18400
rect 130014 17940 130070 18400
rect 130474 17940 130530 18400
rect 130842 17940 130898 18400
rect 131302 17940 131358 18400
rect 131762 17940 131818 18400
rect 132222 17940 132278 18400
rect 132590 17940 132646 18400
rect 133050 17940 133106 18400
rect 133510 17940 133566 18400
rect 133970 17940 134026 18400
rect 134338 17940 134394 18400
rect 134798 17940 134854 18400
rect 135258 17940 135314 18400
rect 135718 17940 135774 18400
rect 136086 17940 136142 18400
rect 136546 17940 136602 18400
rect 137006 17940 137062 18400
rect 137374 17940 137430 18400
rect 137834 17940 137890 18400
rect 138294 17940 138350 18400
rect 138754 17940 138810 18400
rect 139122 17940 139178 18400
rect 139582 17940 139638 18400
rect 140042 17940 140098 18400
rect 140502 17940 140558 18400
rect 140870 17940 140926 18400
rect 141330 17940 141386 18400
rect 141790 17940 141846 18400
rect 142250 17940 142306 18400
rect 142618 17940 142674 18400
rect 143078 17940 143134 18400
rect 143538 17940 143594 18400
rect 143998 17940 144054 18400
rect 144366 17940 144422 18400
rect 144826 17940 144882 18400
rect 145286 17940 145342 18400
rect 145654 17940 145710 18400
rect 146114 17940 146170 18400
rect 146574 17940 146630 18400
rect 147034 17940 147090 18400
rect 147402 17940 147458 18400
rect 147862 17940 147918 18400
rect 148322 17940 148378 18400
rect 148782 17940 148838 18400
rect 149150 17940 149206 18400
rect 149610 17940 149666 18400
rect 150070 17940 150126 18400
rect 150530 17940 150586 18400
rect 150898 17940 150954 18400
rect 151358 17940 151414 18400
rect 151818 17940 151874 18400
rect 152186 17940 152242 18400
rect 152646 17940 152702 18400
rect 153106 17940 153162 18400
rect 153566 17940 153622 18400
rect 153934 17940 153990 18400
rect 154394 17940 154450 18400
rect 154854 17940 154910 18400
rect 155314 17940 155370 18400
rect 155682 17940 155738 18400
rect 156142 17940 156198 18400
rect 156602 17940 156658 18400
rect 157062 17940 157118 18400
rect 157430 17940 157486 18400
rect 157890 17940 157946 18400
rect 158350 17940 158406 18400
rect 158810 17940 158866 18400
rect 159178 17940 159234 18400
rect 159638 17940 159694 18400
rect 160098 17940 160154 18400
rect 160466 17940 160522 18400
rect 160926 17940 160982 18400
rect 161386 17940 161442 18400
rect 161846 17940 161902 18400
rect 162214 17940 162270 18400
rect 162674 17940 162730 18400
rect 163134 17940 163190 18400
rect 163594 17940 163650 18400
rect 163962 17940 164018 18400
rect 164422 17940 164478 18400
rect 164882 17940 164938 18400
rect 165342 17940 165398 18400
rect 165710 17940 165766 18400
rect 166170 17940 166226 18400
rect 166630 17940 166686 18400
rect 167090 17940 167146 18400
rect 167458 17940 167514 18400
rect 167918 17940 167974 18400
rect 168378 17940 168434 18400
rect 168746 17940 168802 18400
rect 169206 17940 169262 18400
rect 169666 17940 169722 18400
rect 170126 17940 170182 18400
rect 170494 17940 170550 18400
rect 170954 17940 171010 18400
rect 171414 17940 171470 18400
rect 171874 17940 171930 18400
rect 172242 17940 172298 18400
rect 172702 17940 172758 18400
rect 173162 17940 173218 18400
rect 173622 17940 173678 18400
rect 173990 17940 174046 18400
rect 174450 17940 174506 18400
rect 174910 17940 174966 18400
rect 175370 17940 175426 18400
rect 175738 17940 175794 18400
rect 176198 17940 176254 18400
rect 176658 17940 176714 18400
rect 177026 17940 177082 18400
rect 177486 17940 177542 18400
rect 177946 17940 178002 18400
rect 178406 17940 178462 18400
rect 178774 17940 178830 18400
rect 179234 17940 179290 18400
rect 179694 17940 179750 18400
rect 180154 17940 180210 18400
rect 180522 17940 180578 18400
rect 180982 17940 181038 18400
rect 181442 17940 181498 18400
rect 181902 17940 181958 18400
rect 182270 17940 182326 18400
rect 182730 17940 182786 18400
rect 183190 17940 183246 18400
rect 183650 17940 183706 18400
rect 184018 17940 184074 18400
rect 184478 17940 184534 18400
rect 184938 17940 184994 18400
rect 185306 17940 185362 18400
rect 185766 17940 185822 18400
rect 186226 17940 186282 18400
rect 186686 17940 186742 18400
rect 187054 17940 187110 18400
rect 187514 17940 187570 18400
rect 187974 17940 188030 18400
rect 188434 17940 188490 18400
rect 188802 17940 188858 18400
rect 189262 17940 189318 18400
rect 189722 17940 189778 18400
rect 190182 17940 190238 18400
rect 190550 17940 190606 18400
rect 191010 17940 191066 18400
rect 191470 17940 191526 18400
rect 191930 17940 191986 18400
rect 192298 17940 192354 18400
rect 192758 17940 192814 18400
rect 193218 17940 193274 18400
rect 193586 17940 193642 18400
rect 194046 17940 194102 18400
rect 194506 17940 194562 18400
rect 194966 17940 195022 18400
rect 195334 17940 195390 18400
rect 195794 17940 195850 18400
rect 196254 17940 196310 18400
rect 196714 17940 196770 18400
rect 197082 17940 197138 18400
rect 197542 17940 197598 18400
rect 198002 17940 198058 18400
rect 198462 17940 198518 18400
rect 198830 17940 198886 18400
rect 199290 17940 199346 18400
rect 199750 17940 199806 18400
rect 202 -400 258 60
rect 570 -400 626 60
rect 1030 -400 1086 60
rect 1490 -400 1546 60
rect 1858 -400 1914 60
rect 2318 -400 2374 60
rect 2778 -400 2834 60
rect 3238 -400 3294 60
rect 3606 -400 3662 60
rect 4066 -400 4122 60
rect 4526 -400 4582 60
rect 4986 -400 5042 60
rect 5354 -400 5410 60
rect 5814 -400 5870 60
rect 6274 -400 6330 60
rect 6734 -400 6790 60
rect 7102 -400 7158 60
rect 7562 -400 7618 60
rect 8022 -400 8078 60
rect 8390 -400 8446 60
rect 8850 -400 8906 60
rect 9310 -400 9366 60
rect 9770 -400 9826 60
rect 10138 -400 10194 60
rect 10598 -400 10654 60
rect 11058 -400 11114 60
rect 11518 -400 11574 60
rect 11886 -400 11942 60
rect 12346 -400 12402 60
rect 12806 -400 12862 60
rect 13266 -400 13322 60
rect 13634 -400 13690 60
rect 14094 -400 14150 60
rect 14554 -400 14610 60
rect 15014 -400 15070 60
rect 15382 -400 15438 60
rect 15842 -400 15898 60
rect 16302 -400 16358 60
rect 16670 -400 16726 60
rect 17130 -400 17186 60
rect 17590 -400 17646 60
rect 18050 -400 18106 60
rect 18418 -400 18474 60
rect 18878 -400 18934 60
rect 19338 -400 19394 60
rect 19798 -400 19854 60
rect 20166 -400 20222 60
rect 20626 -400 20682 60
rect 21086 -400 21142 60
rect 21546 -400 21602 60
rect 21914 -400 21970 60
rect 22374 -400 22430 60
rect 22834 -400 22890 60
rect 23294 -400 23350 60
rect 23662 -400 23718 60
rect 24122 -400 24178 60
rect 24582 -400 24638 60
rect 24950 -400 25006 60
rect 25410 -400 25466 60
rect 25870 -400 25926 60
rect 26330 -400 26386 60
rect 26698 -400 26754 60
rect 27158 -400 27214 60
rect 27618 -400 27674 60
rect 28078 -400 28134 60
rect 28446 -400 28502 60
rect 28906 -400 28962 60
rect 29366 -400 29422 60
rect 29826 -400 29882 60
rect 30194 -400 30250 60
rect 30654 -400 30710 60
rect 31114 -400 31170 60
rect 31574 -400 31630 60
rect 31942 -400 31998 60
rect 32402 -400 32458 60
rect 32862 -400 32918 60
rect 33230 -400 33286 60
rect 33690 -400 33746 60
rect 34150 -400 34206 60
rect 34610 -400 34666 60
rect 34978 -400 35034 60
rect 35438 -400 35494 60
rect 35898 -400 35954 60
rect 36358 -400 36414 60
rect 36726 -400 36782 60
rect 37186 -400 37242 60
rect 37646 -400 37702 60
rect 38106 -400 38162 60
rect 38474 -400 38530 60
rect 38934 -400 38990 60
rect 39394 -400 39450 60
rect 39854 -400 39910 60
rect 40222 -400 40278 60
rect 40682 -400 40738 60
rect 41142 -400 41198 60
rect 41510 -400 41566 60
rect 41970 -400 42026 60
rect 42430 -400 42486 60
rect 42890 -400 42946 60
rect 43258 -400 43314 60
rect 43718 -400 43774 60
rect 44178 -400 44234 60
rect 44638 -400 44694 60
rect 45006 -400 45062 60
rect 45466 -400 45522 60
rect 45926 -400 45982 60
rect 46386 -400 46442 60
rect 46754 -400 46810 60
rect 47214 -400 47270 60
rect 47674 -400 47730 60
rect 48134 -400 48190 60
rect 48502 -400 48558 60
rect 48962 -400 49018 60
rect 49422 -400 49478 60
rect 49790 -400 49846 60
rect 50250 -400 50306 60
rect 50710 -400 50766 60
rect 51170 -400 51226 60
rect 51538 -400 51594 60
rect 51998 -400 52054 60
rect 52458 -400 52514 60
rect 52918 -400 52974 60
rect 53286 -400 53342 60
rect 53746 -400 53802 60
rect 54206 -400 54262 60
rect 54666 -400 54722 60
rect 55034 -400 55090 60
rect 55494 -400 55550 60
rect 55954 -400 56010 60
rect 56322 -400 56378 60
rect 56782 -400 56838 60
rect 57242 -400 57298 60
rect 57702 -400 57758 60
rect 58070 -400 58126 60
rect 58530 -400 58586 60
rect 58990 -400 59046 60
rect 59450 -400 59506 60
rect 59818 -400 59874 60
rect 60278 -400 60334 60
rect 60738 -400 60794 60
rect 61198 -400 61254 60
rect 61566 -400 61622 60
rect 62026 -400 62082 60
rect 62486 -400 62542 60
rect 62946 -400 63002 60
rect 63314 -400 63370 60
rect 63774 -400 63830 60
rect 64234 -400 64290 60
rect 64602 -400 64658 60
rect 65062 -400 65118 60
rect 65522 -400 65578 60
rect 65982 -400 66038 60
rect 66350 -400 66406 60
rect 66810 -400 66866 60
rect 67270 -400 67326 60
rect 67730 -400 67786 60
rect 68098 -400 68154 60
rect 68558 -400 68614 60
rect 69018 -400 69074 60
rect 69478 -400 69534 60
rect 69846 -400 69902 60
rect 70306 -400 70362 60
rect 70766 -400 70822 60
rect 71226 -400 71282 60
rect 71594 -400 71650 60
rect 72054 -400 72110 60
rect 72514 -400 72570 60
rect 72882 -400 72938 60
rect 73342 -400 73398 60
rect 73802 -400 73858 60
rect 74262 -400 74318 60
rect 74630 -400 74686 60
rect 75090 -400 75146 60
rect 75550 -400 75606 60
rect 76010 -400 76066 60
rect 76378 -400 76434 60
rect 76838 -400 76894 60
rect 77298 -400 77354 60
rect 77758 -400 77814 60
rect 78126 -400 78182 60
rect 78586 -400 78642 60
rect 79046 -400 79102 60
rect 79506 -400 79562 60
rect 79874 -400 79930 60
rect 80334 -400 80390 60
rect 80794 -400 80850 60
rect 81162 -400 81218 60
rect 81622 -400 81678 60
rect 82082 -400 82138 60
rect 82542 -400 82598 60
rect 82910 -400 82966 60
rect 83370 -400 83426 60
rect 83830 -400 83886 60
rect 84290 -400 84346 60
rect 84658 -400 84714 60
rect 85118 -400 85174 60
rect 85578 -400 85634 60
rect 86038 -400 86094 60
rect 86406 -400 86462 60
rect 86866 -400 86922 60
rect 87326 -400 87382 60
rect 87786 -400 87842 60
rect 88154 -400 88210 60
rect 88614 -400 88670 60
rect 89074 -400 89130 60
rect 89442 -400 89498 60
rect 89902 -400 89958 60
rect 90362 -400 90418 60
rect 90822 -400 90878 60
rect 91190 -400 91246 60
rect 91650 -400 91706 60
rect 92110 -400 92166 60
rect 92570 -400 92626 60
rect 92938 -400 92994 60
rect 93398 -400 93454 60
rect 93858 -400 93914 60
rect 94318 -400 94374 60
rect 94686 -400 94742 60
rect 95146 -400 95202 60
rect 95606 -400 95662 60
rect 96066 -400 96122 60
rect 96434 -400 96490 60
rect 96894 -400 96950 60
rect 97354 -400 97410 60
rect 97722 -400 97778 60
rect 98182 -400 98238 60
rect 98642 -400 98698 60
rect 99102 -400 99158 60
rect 99470 -400 99526 60
rect 99930 -400 99986 60
rect 100390 -400 100446 60
rect 100850 -400 100906 60
rect 101218 -400 101274 60
rect 101678 -400 101734 60
rect 102138 -400 102194 60
rect 102598 -400 102654 60
rect 102966 -400 103022 60
rect 103426 -400 103482 60
rect 103886 -400 103942 60
rect 104254 -400 104310 60
rect 104714 -400 104770 60
rect 105174 -400 105230 60
rect 105634 -400 105690 60
rect 106002 -400 106058 60
rect 106462 -400 106518 60
rect 106922 -400 106978 60
rect 107382 -400 107438 60
rect 107750 -400 107806 60
rect 108210 -400 108266 60
rect 108670 -400 108726 60
rect 109130 -400 109186 60
rect 109498 -400 109554 60
rect 109958 -400 110014 60
rect 110418 -400 110474 60
rect 110878 -400 110934 60
rect 111246 -400 111302 60
rect 111706 -400 111762 60
rect 112166 -400 112222 60
rect 112534 -400 112590 60
rect 112994 -400 113050 60
rect 113454 -400 113510 60
rect 113914 -400 113970 60
rect 114282 -400 114338 60
rect 114742 -400 114798 60
rect 115202 -400 115258 60
rect 115662 -400 115718 60
rect 116030 -400 116086 60
rect 116490 -400 116546 60
rect 116950 -400 117006 60
rect 117410 -400 117466 60
rect 117778 -400 117834 60
rect 118238 -400 118294 60
rect 118698 -400 118754 60
rect 119158 -400 119214 60
rect 119526 -400 119582 60
rect 119986 -400 120042 60
rect 120446 -400 120502 60
rect 120814 -400 120870 60
rect 121274 -400 121330 60
rect 121734 -400 121790 60
rect 122194 -400 122250 60
rect 122562 -400 122618 60
rect 123022 -400 123078 60
rect 123482 -400 123538 60
rect 123942 -400 123998 60
rect 124310 -400 124366 60
rect 124770 -400 124826 60
rect 125230 -400 125286 60
rect 125690 -400 125746 60
rect 126058 -400 126114 60
rect 126518 -400 126574 60
rect 126978 -400 127034 60
rect 127438 -400 127494 60
rect 127806 -400 127862 60
rect 128266 -400 128322 60
rect 128726 -400 128782 60
rect 129094 -400 129150 60
rect 129554 -400 129610 60
rect 130014 -400 130070 60
rect 130474 -400 130530 60
rect 130842 -400 130898 60
rect 131302 -400 131358 60
rect 131762 -400 131818 60
rect 132222 -400 132278 60
rect 132590 -400 132646 60
rect 133050 -400 133106 60
rect 133510 -400 133566 60
rect 133970 -400 134026 60
rect 134338 -400 134394 60
rect 134798 -400 134854 60
rect 135258 -400 135314 60
rect 135718 -400 135774 60
rect 136086 -400 136142 60
rect 136546 -400 136602 60
rect 137006 -400 137062 60
rect 137374 -400 137430 60
rect 137834 -400 137890 60
rect 138294 -400 138350 60
rect 138754 -400 138810 60
rect 139122 -400 139178 60
rect 139582 -400 139638 60
rect 140042 -400 140098 60
rect 140502 -400 140558 60
rect 140870 -400 140926 60
rect 141330 -400 141386 60
rect 141790 -400 141846 60
rect 142250 -400 142306 60
rect 142618 -400 142674 60
rect 143078 -400 143134 60
rect 143538 -400 143594 60
rect 143998 -400 144054 60
rect 144366 -400 144422 60
rect 144826 -400 144882 60
rect 145286 -400 145342 60
rect 145654 -400 145710 60
rect 146114 -400 146170 60
rect 146574 -400 146630 60
rect 147034 -400 147090 60
rect 147402 -400 147458 60
rect 147862 -400 147918 60
rect 148322 -400 148378 60
rect 148782 -400 148838 60
rect 149150 -400 149206 60
rect 149610 -400 149666 60
rect 150070 -400 150126 60
rect 150530 -400 150586 60
rect 150898 -400 150954 60
rect 151358 -400 151414 60
rect 151818 -400 151874 60
rect 152186 -400 152242 60
rect 152646 -400 152702 60
rect 153106 -400 153162 60
rect 153566 -400 153622 60
rect 153934 -400 153990 60
rect 154394 -400 154450 60
rect 154854 -400 154910 60
rect 155314 -400 155370 60
rect 155682 -400 155738 60
rect 156142 -400 156198 60
rect 156602 -400 156658 60
rect 157062 -400 157118 60
rect 157430 -400 157486 60
rect 157890 -400 157946 60
rect 158350 -400 158406 60
rect 158810 -400 158866 60
rect 159178 -400 159234 60
rect 159638 -400 159694 60
rect 160098 -400 160154 60
rect 160466 -400 160522 60
rect 160926 -400 160982 60
rect 161386 -400 161442 60
rect 161846 -400 161902 60
rect 162214 -400 162270 60
rect 162674 -400 162730 60
rect 163134 -400 163190 60
rect 163594 -400 163650 60
rect 163962 -400 164018 60
rect 164422 -400 164478 60
rect 164882 -400 164938 60
rect 165342 -400 165398 60
rect 165710 -400 165766 60
rect 166170 -400 166226 60
rect 166630 -400 166686 60
rect 167090 -400 167146 60
rect 167458 -400 167514 60
rect 167918 -400 167974 60
rect 168378 -400 168434 60
rect 168746 -400 168802 60
rect 169206 -400 169262 60
rect 169666 -400 169722 60
rect 170126 -400 170182 60
rect 170494 -400 170550 60
rect 170954 -400 171010 60
rect 171414 -400 171470 60
rect 171874 -400 171930 60
rect 172242 -400 172298 60
rect 172702 -400 172758 60
rect 173162 -400 173218 60
rect 173622 -400 173678 60
rect 173990 -400 174046 60
rect 174450 -400 174506 60
rect 174910 -400 174966 60
rect 175370 -400 175426 60
rect 175738 -400 175794 60
rect 176198 -400 176254 60
rect 176658 -400 176714 60
rect 177026 -400 177082 60
rect 177486 -400 177542 60
rect 177946 -400 178002 60
rect 178406 -400 178462 60
rect 178774 -400 178830 60
rect 179234 -400 179290 60
rect 179694 -400 179750 60
rect 180154 -400 180210 60
rect 180522 -400 180578 60
rect 180982 -400 181038 60
rect 181442 -400 181498 60
rect 181902 -400 181958 60
rect 182270 -400 182326 60
rect 182730 -400 182786 60
rect 183190 -400 183246 60
rect 183650 -400 183706 60
rect 184018 -400 184074 60
rect 184478 -400 184534 60
rect 184938 -400 184994 60
rect 185306 -400 185362 60
rect 185766 -400 185822 60
rect 186226 -400 186282 60
rect 186686 -400 186742 60
rect 187054 -400 187110 60
rect 187514 -400 187570 60
rect 187974 -400 188030 60
rect 188434 -400 188490 60
rect 188802 -400 188858 60
rect 189262 -400 189318 60
rect 189722 -400 189778 60
rect 190182 -400 190238 60
rect 190550 -400 190606 60
rect 191010 -400 191066 60
rect 191470 -400 191526 60
rect 191930 -400 191986 60
rect 192298 -400 192354 60
rect 192758 -400 192814 60
rect 193218 -400 193274 60
rect 193586 -400 193642 60
rect 194046 -400 194102 60
rect 194506 -400 194562 60
rect 194966 -400 195022 60
rect 195334 -400 195390 60
rect 195794 -400 195850 60
rect 196254 -400 196310 60
rect 196714 -400 196770 60
rect 197082 -400 197138 60
rect 197542 -400 197598 60
rect 198002 -400 198058 60
rect 198462 -400 198518 60
rect 198830 -400 198886 60
rect 199290 -400 199346 60
rect 199750 -400 199806 60
<< obsm2 >>
rect 40776 17940 40828 17950
rect 68836 17954 68888 18018
rect 68848 17940 68876 17954
rect 69112 17954 69164 18018
rect 69124 17940 69152 17954
rect 70216 17954 70268 18018
rect 70228 17940 70256 17954
rect 74724 17940 74776 17950
rect 74816 17940 74868 17950
rect 89812 17940 89864 17950
rect 91928 17940 91980 17950
rect 101404 17940 101456 17950
rect 101864 17940 101916 17950
rect 103704 17940 103756 17950
rect 113180 17954 113232 18018
rect 113192 17940 113220 17954
rect 126336 17940 126388 17950
rect 202 60 199806 17940
<< metal3 >>
rect -2762 20712 202678 20730
rect -2762 20648 -2744 20712
rect -2680 20648 -2664 20712
rect -2600 20648 22312 20712
rect 22376 20648 22392 20712
rect 22456 20648 52312 20712
rect 52376 20648 52392 20712
rect 52456 20648 82312 20712
rect 82376 20648 82392 20712
rect 82456 20648 112312 20712
rect 112376 20648 112392 20712
rect 112456 20648 142312 20712
rect 142376 20648 142392 20712
rect 142456 20648 172312 20712
rect 172376 20648 172392 20712
rect 172456 20648 202516 20712
rect 202580 20648 202596 20712
rect 202660 20648 202678 20712
rect -2762 20632 202678 20648
rect -2762 20568 -2744 20632
rect -2680 20568 -2664 20632
rect -2600 20568 22312 20632
rect 22376 20568 22392 20632
rect 22456 20568 52312 20632
rect 52376 20568 52392 20632
rect 52456 20568 82312 20632
rect 82376 20568 82392 20632
rect 82456 20568 112312 20632
rect 112376 20568 112392 20632
rect 112456 20568 142312 20632
rect 142376 20568 142392 20632
rect 142456 20568 172312 20632
rect 172376 20568 172392 20632
rect 172456 20568 202516 20632
rect 202580 20568 202596 20632
rect 202660 20568 202678 20632
rect -2762 20550 202678 20568
rect -2498 20448 202414 20466
rect -2498 20384 -2480 20448
rect -2416 20384 -2400 20448
rect -2336 20384 7312 20448
rect 7376 20384 7392 20448
rect 7456 20384 37312 20448
rect 37376 20384 37392 20448
rect 37456 20384 67312 20448
rect 67376 20384 67392 20448
rect 67456 20384 97312 20448
rect 97376 20384 97392 20448
rect 97456 20384 127312 20448
rect 127376 20384 127392 20448
rect 127456 20384 157312 20448
rect 157376 20384 157392 20448
rect 157456 20384 187312 20448
rect 187376 20384 187392 20448
rect 187456 20384 202252 20448
rect 202316 20384 202332 20448
rect 202396 20384 202414 20448
rect -2498 20368 202414 20384
rect -2498 20304 -2480 20368
rect -2416 20304 -2400 20368
rect -2336 20304 7312 20368
rect 7376 20304 7392 20368
rect 7456 20304 37312 20368
rect 37376 20304 37392 20368
rect 37456 20304 67312 20368
rect 67376 20304 67392 20368
rect 67456 20304 97312 20368
rect 97376 20304 97392 20368
rect 97456 20304 127312 20368
rect 127376 20304 127392 20368
rect 127456 20304 157312 20368
rect 157376 20304 157392 20368
rect 157456 20304 187312 20368
rect 187376 20304 187392 20368
rect 187456 20304 202252 20368
rect 202316 20304 202332 20368
rect 202396 20304 202414 20368
rect -2498 20286 202414 20304
rect -2234 20184 202150 20202
rect -2234 20120 -2216 20184
rect -2152 20120 -2136 20184
rect -2072 20120 21492 20184
rect 21556 20120 21572 20184
rect 21636 20120 51492 20184
rect 51556 20120 51572 20184
rect 51636 20120 81492 20184
rect 81556 20120 81572 20184
rect 81636 20120 111492 20184
rect 111556 20120 111572 20184
rect 111636 20120 141492 20184
rect 141556 20120 141572 20184
rect 141636 20120 171492 20184
rect 171556 20120 171572 20184
rect 171636 20120 201988 20184
rect 202052 20120 202068 20184
rect 202132 20120 202150 20184
rect -2234 20104 202150 20120
rect -2234 20040 -2216 20104
rect -2152 20040 -2136 20104
rect -2072 20040 21492 20104
rect 21556 20040 21572 20104
rect 21636 20040 51492 20104
rect 51556 20040 51572 20104
rect 51636 20040 81492 20104
rect 81556 20040 81572 20104
rect 81636 20040 111492 20104
rect 111556 20040 111572 20104
rect 111636 20040 141492 20104
rect 141556 20040 141572 20104
rect 141636 20040 171492 20104
rect 171556 20040 171572 20104
rect 171636 20040 201988 20104
rect 202052 20040 202068 20104
rect 202132 20040 202150 20104
rect -2234 20022 202150 20040
rect -1970 19920 201886 19938
rect -1970 19856 -1952 19920
rect -1888 19856 -1872 19920
rect -1808 19856 6492 19920
rect 6556 19856 6572 19920
rect 6636 19856 36492 19920
rect 36556 19856 36572 19920
rect 36636 19856 66492 19920
rect 66556 19856 66572 19920
rect 66636 19856 96492 19920
rect 96556 19856 96572 19920
rect 96636 19856 126492 19920
rect 126556 19856 126572 19920
rect 126636 19856 156492 19920
rect 156556 19856 156572 19920
rect 156636 19856 186492 19920
rect 186556 19856 186572 19920
rect 186636 19856 201724 19920
rect 201788 19856 201804 19920
rect 201868 19856 201886 19920
rect -1970 19840 201886 19856
rect -1970 19776 -1952 19840
rect -1888 19776 -1872 19840
rect -1808 19776 6492 19840
rect 6556 19776 6572 19840
rect 6636 19776 36492 19840
rect 36556 19776 36572 19840
rect 36636 19776 66492 19840
rect 66556 19776 66572 19840
rect 66636 19776 96492 19840
rect 96556 19776 96572 19840
rect 96636 19776 126492 19840
rect 126556 19776 126572 19840
rect 126636 19776 156492 19840
rect 156556 19776 156572 19840
rect 156636 19776 186492 19840
rect 186556 19776 186572 19840
rect 186636 19776 201724 19840
rect 201788 19776 201804 19840
rect 201868 19776 201886 19840
rect -1970 19758 201886 19776
rect -1706 19656 201622 19674
rect -1706 19592 -1688 19656
rect -1624 19592 -1608 19656
rect -1544 19592 20672 19656
rect 20736 19592 20752 19656
rect 20816 19592 50672 19656
rect 50736 19592 50752 19656
rect 50816 19592 80672 19656
rect 80736 19592 80752 19656
rect 80816 19592 110672 19656
rect 110736 19592 110752 19656
rect 110816 19592 140672 19656
rect 140736 19592 140752 19656
rect 140816 19592 170672 19656
rect 170736 19592 170752 19656
rect 170816 19592 201460 19656
rect 201524 19592 201540 19656
rect 201604 19592 201622 19656
rect -1706 19576 201622 19592
rect -1706 19512 -1688 19576
rect -1624 19512 -1608 19576
rect -1544 19512 20672 19576
rect 20736 19512 20752 19576
rect 20816 19512 50672 19576
rect 50736 19512 50752 19576
rect 50816 19512 80672 19576
rect 80736 19512 80752 19576
rect 80816 19512 110672 19576
rect 110736 19512 110752 19576
rect 110816 19512 140672 19576
rect 140736 19512 140752 19576
rect 140816 19512 170672 19576
rect 170736 19512 170752 19576
rect 170816 19512 201460 19576
rect 201524 19512 201540 19576
rect 201604 19512 201622 19576
rect -1706 19494 201622 19512
rect -1442 19392 201358 19410
rect -1442 19328 -1424 19392
rect -1360 19328 -1344 19392
rect -1280 19328 5672 19392
rect 5736 19328 5752 19392
rect 5816 19328 35672 19392
rect 35736 19328 35752 19392
rect 35816 19328 65672 19392
rect 65736 19328 65752 19392
rect 65816 19328 95672 19392
rect 95736 19328 95752 19392
rect 95816 19328 125672 19392
rect 125736 19328 125752 19392
rect 125816 19328 155672 19392
rect 155736 19328 155752 19392
rect 155816 19328 185672 19392
rect 185736 19328 185752 19392
rect 185816 19328 201196 19392
rect 201260 19328 201276 19392
rect 201340 19328 201358 19392
rect -1442 19312 201358 19328
rect -1442 19248 -1424 19312
rect -1360 19248 -1344 19312
rect -1280 19248 5672 19312
rect 5736 19248 5752 19312
rect 5816 19248 35672 19312
rect 35736 19248 35752 19312
rect 35816 19248 65672 19312
rect 65736 19248 65752 19312
rect 65816 19248 95672 19312
rect 95736 19248 95752 19312
rect 95816 19248 125672 19312
rect 125736 19248 125752 19312
rect 125816 19248 155672 19312
rect 155736 19248 155752 19312
rect 155816 19248 185672 19312
rect 185736 19248 185752 19312
rect 185816 19248 201196 19312
rect 201260 19248 201276 19312
rect 201340 19248 201358 19312
rect -1442 19230 201358 19248
rect -1178 19128 201094 19146
rect -1178 19064 -1160 19128
rect -1096 19064 -1080 19128
rect -1016 19064 19852 19128
rect 19916 19064 19932 19128
rect 19996 19064 49852 19128
rect 49916 19064 49932 19128
rect 49996 19064 79852 19128
rect 79916 19064 79932 19128
rect 79996 19064 109852 19128
rect 109916 19064 109932 19128
rect 109996 19064 139852 19128
rect 139916 19064 139932 19128
rect 139996 19064 169852 19128
rect 169916 19064 169932 19128
rect 169996 19064 200932 19128
rect 200996 19064 201012 19128
rect 201076 19064 201094 19128
rect -1178 19048 201094 19064
rect -1178 18984 -1160 19048
rect -1096 18984 -1080 19048
rect -1016 18984 19852 19048
rect 19916 18984 19932 19048
rect 19996 18984 49852 19048
rect 49916 18984 49932 19048
rect 49996 18984 79852 19048
rect 79916 18984 79932 19048
rect 79996 18984 109852 19048
rect 109916 18984 109932 19048
rect 109996 18984 139852 19048
rect 139916 18984 139932 19048
rect 139996 18984 169852 19048
rect 169916 18984 169932 19048
rect 169996 18984 200932 19048
rect 200996 18984 201012 19048
rect 201076 18984 201094 19048
rect -1178 18966 201094 18984
rect -914 18864 200830 18882
rect -914 18800 -896 18864
rect -832 18800 -816 18864
rect -752 18800 4852 18864
rect 4916 18800 4932 18864
rect 4996 18800 34852 18864
rect 34916 18800 34932 18864
rect 34996 18800 64852 18864
rect 64916 18800 64932 18864
rect 64996 18800 94852 18864
rect 94916 18800 94932 18864
rect 94996 18800 124852 18864
rect 124916 18800 124932 18864
rect 124996 18800 154852 18864
rect 154916 18800 154932 18864
rect 154996 18800 184852 18864
rect 184916 18800 184932 18864
rect 184996 18800 200668 18864
rect 200732 18800 200748 18864
rect 200812 18800 200830 18864
rect -914 18784 200830 18800
rect -914 18720 -896 18784
rect -832 18720 -816 18784
rect -752 18720 4852 18784
rect 4916 18720 4932 18784
rect 4996 18720 34852 18784
rect 34916 18720 34932 18784
rect 34996 18720 64852 18784
rect 64916 18720 64932 18784
rect 64996 18720 94852 18784
rect 94916 18720 94932 18784
rect 94996 18720 124852 18784
rect 124916 18720 124932 18784
rect 124996 18720 154852 18784
rect 154916 18720 154932 18784
rect 154996 18720 184852 18784
rect 184916 18720 184932 18784
rect 184996 18720 200668 18784
rect 200732 18720 200748 18784
rect 200812 18720 200830 18784
rect -914 18702 200830 18720
rect -650 18600 200566 18618
rect -650 18536 -632 18600
rect -568 18536 -552 18600
rect -488 18536 19032 18600
rect 19096 18536 19112 18600
rect 19176 18536 49032 18600
rect 49096 18536 49112 18600
rect 49176 18536 79032 18600
rect 79096 18536 79112 18600
rect 79176 18536 109032 18600
rect 109096 18536 109112 18600
rect 109176 18536 139032 18600
rect 139096 18536 139112 18600
rect 139176 18536 169032 18600
rect 169096 18536 169112 18600
rect 169176 18536 200404 18600
rect 200468 18536 200484 18600
rect 200548 18536 200566 18600
rect -650 18520 200566 18536
rect -650 18456 -632 18520
rect -568 18456 -552 18520
rect -488 18456 19032 18520
rect 19096 18456 19112 18520
rect 19176 18456 49032 18520
rect 49096 18456 49112 18520
rect 49176 18456 79032 18520
rect 79096 18456 79112 18520
rect 79176 18456 109032 18520
rect 109096 18456 109112 18520
rect 109176 18456 139032 18520
rect 139096 18456 139112 18520
rect 139176 18456 169032 18520
rect 169096 18456 169112 18520
rect 169176 18456 200404 18520
rect 200468 18456 200484 18520
rect 200548 18456 200566 18520
rect -650 18438 200566 18456
rect -386 18336 200302 18354
rect -386 18272 -368 18336
rect -304 18272 -288 18336
rect -224 18272 4032 18336
rect 4096 18272 4112 18336
rect 4176 18272 34032 18336
rect 34096 18272 34112 18336
rect 34176 18272 64032 18336
rect 64096 18272 64112 18336
rect 64176 18272 94032 18336
rect 94096 18272 94112 18336
rect 94176 18272 124032 18336
rect 124096 18272 124112 18336
rect 124176 18272 154032 18336
rect 154096 18272 154112 18336
rect 154176 18272 184032 18336
rect 184096 18272 184112 18336
rect 184176 18272 200140 18336
rect 200204 18272 200220 18336
rect 200284 18272 200302 18336
rect -386 18256 200302 18272
rect -386 18192 -368 18256
rect -304 18192 -288 18256
rect -224 18192 4032 18256
rect 4096 18192 4112 18256
rect 4176 18192 34032 18256
rect 34096 18192 34112 18256
rect 34176 18192 64032 18256
rect 64096 18192 64112 18256
rect 64176 18192 94032 18256
rect 94096 18192 94112 18256
rect 94176 18192 124032 18256
rect 124096 18192 124112 18256
rect 124176 18192 154032 18256
rect 154096 18192 154112 18256
rect 154176 18192 184032 18256
rect 184096 18192 184112 18256
rect 184176 18192 200140 18256
rect 200204 18192 200220 18256
rect 200284 18192 200302 18256
rect -386 18174 200302 18192
rect -400 14968 60 15088
rect -400 8984 60 9104
rect -400 3000 60 3120
rect -386 -240 200302 -222
rect -386 -304 -368 -240
rect -304 -304 -288 -240
rect -224 -304 4032 -240
rect 4096 -304 4112 -240
rect 4176 -304 34032 -240
rect 34096 -304 34112 -240
rect 34176 -304 64032 -240
rect 64096 -304 64112 -240
rect 64176 -304 94032 -240
rect 94096 -304 94112 -240
rect 94176 -304 124032 -240
rect 124096 -304 124112 -240
rect 124176 -304 154032 -240
rect 154096 -304 154112 -240
rect 154176 -304 184032 -240
rect 184096 -304 184112 -240
rect 184176 -304 200140 -240
rect 200204 -304 200220 -240
rect 200284 -304 200302 -240
rect -386 -320 200302 -304
rect -386 -384 -368 -320
rect -304 -384 -288 -320
rect -224 -384 4032 -320
rect 4096 -384 4112 -320
rect 4176 -384 34032 -320
rect 34096 -384 34112 -320
rect 34176 -384 64032 -320
rect 64096 -384 64112 -320
rect 64176 -384 94032 -320
rect 94096 -384 94112 -320
rect 94176 -384 124032 -320
rect 124096 -384 124112 -320
rect 124176 -384 154032 -320
rect 154096 -384 154112 -320
rect 154176 -384 184032 -320
rect 184096 -384 184112 -320
rect 184176 -384 200140 -320
rect 200204 -384 200220 -320
rect 200284 -384 200302 -320
rect -386 -402 200302 -384
rect -650 -504 200566 -486
rect -650 -568 -632 -504
rect -568 -568 -552 -504
rect -488 -568 19032 -504
rect 19096 -568 19112 -504
rect 19176 -568 49032 -504
rect 49096 -568 49112 -504
rect 49176 -568 79032 -504
rect 79096 -568 79112 -504
rect 79176 -568 109032 -504
rect 109096 -568 109112 -504
rect 109176 -568 139032 -504
rect 139096 -568 139112 -504
rect 139176 -568 169032 -504
rect 169096 -568 169112 -504
rect 169176 -568 200404 -504
rect 200468 -568 200484 -504
rect 200548 -568 200566 -504
rect -650 -584 200566 -568
rect -650 -648 -632 -584
rect -568 -648 -552 -584
rect -488 -648 19032 -584
rect 19096 -648 19112 -584
rect 19176 -648 49032 -584
rect 49096 -648 49112 -584
rect 49176 -648 79032 -584
rect 79096 -648 79112 -584
rect 79176 -648 109032 -584
rect 109096 -648 109112 -584
rect 109176 -648 139032 -584
rect 139096 -648 139112 -584
rect 139176 -648 169032 -584
rect 169096 -648 169112 -584
rect 169176 -648 200404 -584
rect 200468 -648 200484 -584
rect 200548 -648 200566 -584
rect -650 -666 200566 -648
rect -914 -768 200830 -750
rect -914 -832 -896 -768
rect -832 -832 -816 -768
rect -752 -832 4852 -768
rect 4916 -832 4932 -768
rect 4996 -832 34852 -768
rect 34916 -832 34932 -768
rect 34996 -832 64852 -768
rect 64916 -832 64932 -768
rect 64996 -832 94852 -768
rect 94916 -832 94932 -768
rect 94996 -832 124852 -768
rect 124916 -832 124932 -768
rect 124996 -832 154852 -768
rect 154916 -832 154932 -768
rect 154996 -832 184852 -768
rect 184916 -832 184932 -768
rect 184996 -832 200668 -768
rect 200732 -832 200748 -768
rect 200812 -832 200830 -768
rect -914 -848 200830 -832
rect -914 -912 -896 -848
rect -832 -912 -816 -848
rect -752 -912 4852 -848
rect 4916 -912 4932 -848
rect 4996 -912 34852 -848
rect 34916 -912 34932 -848
rect 34996 -912 64852 -848
rect 64916 -912 64932 -848
rect 64996 -912 94852 -848
rect 94916 -912 94932 -848
rect 94996 -912 124852 -848
rect 124916 -912 124932 -848
rect 124996 -912 154852 -848
rect 154916 -912 154932 -848
rect 154996 -912 184852 -848
rect 184916 -912 184932 -848
rect 184996 -912 200668 -848
rect 200732 -912 200748 -848
rect 200812 -912 200830 -848
rect -914 -930 200830 -912
rect -1178 -1032 201094 -1014
rect -1178 -1096 -1160 -1032
rect -1096 -1096 -1080 -1032
rect -1016 -1096 19852 -1032
rect 19916 -1096 19932 -1032
rect 19996 -1096 49852 -1032
rect 49916 -1096 49932 -1032
rect 49996 -1096 79852 -1032
rect 79916 -1096 79932 -1032
rect 79996 -1096 109852 -1032
rect 109916 -1096 109932 -1032
rect 109996 -1096 139852 -1032
rect 139916 -1096 139932 -1032
rect 139996 -1096 169852 -1032
rect 169916 -1096 169932 -1032
rect 169996 -1096 200932 -1032
rect 200996 -1096 201012 -1032
rect 201076 -1096 201094 -1032
rect -1178 -1112 201094 -1096
rect -1178 -1176 -1160 -1112
rect -1096 -1176 -1080 -1112
rect -1016 -1176 19852 -1112
rect 19916 -1176 19932 -1112
rect 19996 -1176 49852 -1112
rect 49916 -1176 49932 -1112
rect 49996 -1176 79852 -1112
rect 79916 -1176 79932 -1112
rect 79996 -1176 109852 -1112
rect 109916 -1176 109932 -1112
rect 109996 -1176 139852 -1112
rect 139916 -1176 139932 -1112
rect 139996 -1176 169852 -1112
rect 169916 -1176 169932 -1112
rect 169996 -1176 200932 -1112
rect 200996 -1176 201012 -1112
rect 201076 -1176 201094 -1112
rect -1178 -1194 201094 -1176
rect -1442 -1296 201358 -1278
rect -1442 -1360 -1424 -1296
rect -1360 -1360 -1344 -1296
rect -1280 -1360 5672 -1296
rect 5736 -1360 5752 -1296
rect 5816 -1360 35672 -1296
rect 35736 -1360 35752 -1296
rect 35816 -1360 65672 -1296
rect 65736 -1360 65752 -1296
rect 65816 -1360 95672 -1296
rect 95736 -1360 95752 -1296
rect 95816 -1360 125672 -1296
rect 125736 -1360 125752 -1296
rect 125816 -1360 155672 -1296
rect 155736 -1360 155752 -1296
rect 155816 -1360 185672 -1296
rect 185736 -1360 185752 -1296
rect 185816 -1360 201196 -1296
rect 201260 -1360 201276 -1296
rect 201340 -1360 201358 -1296
rect -1442 -1376 201358 -1360
rect -1442 -1440 -1424 -1376
rect -1360 -1440 -1344 -1376
rect -1280 -1440 5672 -1376
rect 5736 -1440 5752 -1376
rect 5816 -1440 35672 -1376
rect 35736 -1440 35752 -1376
rect 35816 -1440 65672 -1376
rect 65736 -1440 65752 -1376
rect 65816 -1440 95672 -1376
rect 95736 -1440 95752 -1376
rect 95816 -1440 125672 -1376
rect 125736 -1440 125752 -1376
rect 125816 -1440 155672 -1376
rect 155736 -1440 155752 -1376
rect 155816 -1440 185672 -1376
rect 185736 -1440 185752 -1376
rect 185816 -1440 201196 -1376
rect 201260 -1440 201276 -1376
rect 201340 -1440 201358 -1376
rect -1442 -1458 201358 -1440
rect -1706 -1560 201622 -1542
rect -1706 -1624 -1688 -1560
rect -1624 -1624 -1608 -1560
rect -1544 -1624 20672 -1560
rect 20736 -1624 20752 -1560
rect 20816 -1624 50672 -1560
rect 50736 -1624 50752 -1560
rect 50816 -1624 80672 -1560
rect 80736 -1624 80752 -1560
rect 80816 -1624 110672 -1560
rect 110736 -1624 110752 -1560
rect 110816 -1624 140672 -1560
rect 140736 -1624 140752 -1560
rect 140816 -1624 170672 -1560
rect 170736 -1624 170752 -1560
rect 170816 -1624 201460 -1560
rect 201524 -1624 201540 -1560
rect 201604 -1624 201622 -1560
rect -1706 -1640 201622 -1624
rect -1706 -1704 -1688 -1640
rect -1624 -1704 -1608 -1640
rect -1544 -1704 20672 -1640
rect 20736 -1704 20752 -1640
rect 20816 -1704 50672 -1640
rect 50736 -1704 50752 -1640
rect 50816 -1704 80672 -1640
rect 80736 -1704 80752 -1640
rect 80816 -1704 110672 -1640
rect 110736 -1704 110752 -1640
rect 110816 -1704 140672 -1640
rect 140736 -1704 140752 -1640
rect 140816 -1704 170672 -1640
rect 170736 -1704 170752 -1640
rect 170816 -1704 201460 -1640
rect 201524 -1704 201540 -1640
rect 201604 -1704 201622 -1640
rect -1706 -1722 201622 -1704
rect -1970 -1824 201886 -1806
rect -1970 -1888 -1952 -1824
rect -1888 -1888 -1872 -1824
rect -1808 -1888 6492 -1824
rect 6556 -1888 6572 -1824
rect 6636 -1888 36492 -1824
rect 36556 -1888 36572 -1824
rect 36636 -1888 66492 -1824
rect 66556 -1888 66572 -1824
rect 66636 -1888 96492 -1824
rect 96556 -1888 96572 -1824
rect 96636 -1888 126492 -1824
rect 126556 -1888 126572 -1824
rect 126636 -1888 156492 -1824
rect 156556 -1888 156572 -1824
rect 156636 -1888 186492 -1824
rect 186556 -1888 186572 -1824
rect 186636 -1888 201724 -1824
rect 201788 -1888 201804 -1824
rect 201868 -1888 201886 -1824
rect -1970 -1904 201886 -1888
rect -1970 -1968 -1952 -1904
rect -1888 -1968 -1872 -1904
rect -1808 -1968 6492 -1904
rect 6556 -1968 6572 -1904
rect 6636 -1968 36492 -1904
rect 36556 -1968 36572 -1904
rect 36636 -1968 66492 -1904
rect 66556 -1968 66572 -1904
rect 66636 -1968 96492 -1904
rect 96556 -1968 96572 -1904
rect 96636 -1968 126492 -1904
rect 126556 -1968 126572 -1904
rect 126636 -1968 156492 -1904
rect 156556 -1968 156572 -1904
rect 156636 -1968 186492 -1904
rect 186556 -1968 186572 -1904
rect 186636 -1968 201724 -1904
rect 201788 -1968 201804 -1904
rect 201868 -1968 201886 -1904
rect -1970 -1986 201886 -1968
rect -2234 -2088 202150 -2070
rect -2234 -2152 -2216 -2088
rect -2152 -2152 -2136 -2088
rect -2072 -2152 21492 -2088
rect 21556 -2152 21572 -2088
rect 21636 -2152 51492 -2088
rect 51556 -2152 51572 -2088
rect 51636 -2152 81492 -2088
rect 81556 -2152 81572 -2088
rect 81636 -2152 111492 -2088
rect 111556 -2152 111572 -2088
rect 111636 -2152 141492 -2088
rect 141556 -2152 141572 -2088
rect 141636 -2152 171492 -2088
rect 171556 -2152 171572 -2088
rect 171636 -2152 201988 -2088
rect 202052 -2152 202068 -2088
rect 202132 -2152 202150 -2088
rect -2234 -2168 202150 -2152
rect -2234 -2232 -2216 -2168
rect -2152 -2232 -2136 -2168
rect -2072 -2232 21492 -2168
rect 21556 -2232 21572 -2168
rect 21636 -2232 51492 -2168
rect 51556 -2232 51572 -2168
rect 51636 -2232 81492 -2168
rect 81556 -2232 81572 -2168
rect 81636 -2232 111492 -2168
rect 111556 -2232 111572 -2168
rect 111636 -2232 141492 -2168
rect 141556 -2232 141572 -2168
rect 141636 -2232 171492 -2168
rect 171556 -2232 171572 -2168
rect 171636 -2232 201988 -2168
rect 202052 -2232 202068 -2168
rect 202132 -2232 202150 -2168
rect -2234 -2250 202150 -2232
rect -2498 -2352 202414 -2334
rect -2498 -2416 -2480 -2352
rect -2416 -2416 -2400 -2352
rect -2336 -2416 7312 -2352
rect 7376 -2416 7392 -2352
rect 7456 -2416 37312 -2352
rect 37376 -2416 37392 -2352
rect 37456 -2416 67312 -2352
rect 67376 -2416 67392 -2352
rect 67456 -2416 97312 -2352
rect 97376 -2416 97392 -2352
rect 97456 -2416 127312 -2352
rect 127376 -2416 127392 -2352
rect 127456 -2416 157312 -2352
rect 157376 -2416 157392 -2352
rect 157456 -2416 187312 -2352
rect 187376 -2416 187392 -2352
rect 187456 -2416 202252 -2352
rect 202316 -2416 202332 -2352
rect 202396 -2416 202414 -2352
rect -2498 -2432 202414 -2416
rect -2498 -2496 -2480 -2432
rect -2416 -2496 -2400 -2432
rect -2336 -2496 7312 -2432
rect 7376 -2496 7392 -2432
rect 7456 -2496 37312 -2432
rect 37376 -2496 37392 -2432
rect 37456 -2496 67312 -2432
rect 67376 -2496 67392 -2432
rect 67456 -2496 97312 -2432
rect 97376 -2496 97392 -2432
rect 97456 -2496 127312 -2432
rect 127376 -2496 127392 -2432
rect 127456 -2496 157312 -2432
rect 157376 -2496 157392 -2432
rect 157456 -2496 187312 -2432
rect 187376 -2496 187392 -2432
rect 187456 -2496 202252 -2432
rect 202316 -2496 202332 -2432
rect 202396 -2496 202414 -2432
rect -2498 -2514 202414 -2496
rect -2762 -2616 202678 -2598
rect -2762 -2680 -2744 -2616
rect -2680 -2680 -2664 -2616
rect -2600 -2680 22312 -2616
rect 22376 -2680 22392 -2616
rect 22456 -2680 52312 -2616
rect 52376 -2680 52392 -2616
rect 52456 -2680 82312 -2616
rect 82376 -2680 82392 -2616
rect 82456 -2680 112312 -2616
rect 112376 -2680 112392 -2616
rect 112456 -2680 142312 -2616
rect 142376 -2680 142392 -2616
rect 142456 -2680 172312 -2616
rect 172376 -2680 172392 -2616
rect 172456 -2680 202516 -2616
rect 202580 -2680 202596 -2616
rect 202660 -2680 202678 -2616
rect -2762 -2696 202678 -2680
rect -2762 -2760 -2744 -2696
rect -2680 -2760 -2664 -2696
rect -2600 -2760 22312 -2696
rect 22376 -2760 22392 -2696
rect 22456 -2760 52312 -2696
rect 52376 -2760 52392 -2696
rect 52456 -2760 82312 -2696
rect 82376 -2760 82392 -2696
rect 82456 -2760 112312 -2696
rect 112376 -2760 112392 -2696
rect 112456 -2760 142312 -2696
rect 142376 -2760 142392 -2696
rect 142456 -2760 172312 -2696
rect 172376 -2760 172392 -2696
rect 172456 -2760 202516 -2696
rect 202580 -2760 202596 -2696
rect 202660 -2760 202678 -2696
rect -2762 -2778 202678 -2760
<< obsm3 >>
rect 60 851 194659 17917
<< via3 >>
rect -2744 20648 -2680 20712
rect -2664 20648 -2600 20712
rect 22312 20648 22376 20712
rect 22392 20648 22456 20712
rect 52312 20648 52376 20712
rect 52392 20648 52456 20712
rect 82312 20648 82376 20712
rect 82392 20648 82456 20712
rect 112312 20648 112376 20712
rect 112392 20648 112456 20712
rect 142312 20648 142376 20712
rect 142392 20648 142456 20712
rect 172312 20648 172376 20712
rect 172392 20648 172456 20712
rect 202516 20648 202580 20712
rect 202596 20648 202660 20712
rect -2744 20568 -2680 20632
rect -2664 20568 -2600 20632
rect 22312 20568 22376 20632
rect 22392 20568 22456 20632
rect 52312 20568 52376 20632
rect 52392 20568 52456 20632
rect 82312 20568 82376 20632
rect 82392 20568 82456 20632
rect 112312 20568 112376 20632
rect 112392 20568 112456 20632
rect 142312 20568 142376 20632
rect 142392 20568 142456 20632
rect 172312 20568 172376 20632
rect 172392 20568 172456 20632
rect 202516 20568 202580 20632
rect 202596 20568 202660 20632
rect -2480 20384 -2416 20448
rect -2400 20384 -2336 20448
rect 7312 20384 7376 20448
rect 7392 20384 7456 20448
rect 37312 20384 37376 20448
rect 37392 20384 37456 20448
rect 67312 20384 67376 20448
rect 67392 20384 67456 20448
rect 97312 20384 97376 20448
rect 97392 20384 97456 20448
rect 127312 20384 127376 20448
rect 127392 20384 127456 20448
rect 157312 20384 157376 20448
rect 157392 20384 157456 20448
rect 187312 20384 187376 20448
rect 187392 20384 187456 20448
rect 202252 20384 202316 20448
rect 202332 20384 202396 20448
rect -2480 20304 -2416 20368
rect -2400 20304 -2336 20368
rect 7312 20304 7376 20368
rect 7392 20304 7456 20368
rect 37312 20304 37376 20368
rect 37392 20304 37456 20368
rect 67312 20304 67376 20368
rect 67392 20304 67456 20368
rect 97312 20304 97376 20368
rect 97392 20304 97456 20368
rect 127312 20304 127376 20368
rect 127392 20304 127456 20368
rect 157312 20304 157376 20368
rect 157392 20304 157456 20368
rect 187312 20304 187376 20368
rect 187392 20304 187456 20368
rect 202252 20304 202316 20368
rect 202332 20304 202396 20368
rect -2216 20120 -2152 20184
rect -2136 20120 -2072 20184
rect 21492 20120 21556 20184
rect 21572 20120 21636 20184
rect 51492 20120 51556 20184
rect 51572 20120 51636 20184
rect 81492 20120 81556 20184
rect 81572 20120 81636 20184
rect 111492 20120 111556 20184
rect 111572 20120 111636 20184
rect 141492 20120 141556 20184
rect 141572 20120 141636 20184
rect 171492 20120 171556 20184
rect 171572 20120 171636 20184
rect 201988 20120 202052 20184
rect 202068 20120 202132 20184
rect -2216 20040 -2152 20104
rect -2136 20040 -2072 20104
rect 21492 20040 21556 20104
rect 21572 20040 21636 20104
rect 51492 20040 51556 20104
rect 51572 20040 51636 20104
rect 81492 20040 81556 20104
rect 81572 20040 81636 20104
rect 111492 20040 111556 20104
rect 111572 20040 111636 20104
rect 141492 20040 141556 20104
rect 141572 20040 141636 20104
rect 171492 20040 171556 20104
rect 171572 20040 171636 20104
rect 201988 20040 202052 20104
rect 202068 20040 202132 20104
rect -1952 19856 -1888 19920
rect -1872 19856 -1808 19920
rect 6492 19856 6556 19920
rect 6572 19856 6636 19920
rect 36492 19856 36556 19920
rect 36572 19856 36636 19920
rect 66492 19856 66556 19920
rect 66572 19856 66636 19920
rect 96492 19856 96556 19920
rect 96572 19856 96636 19920
rect 126492 19856 126556 19920
rect 126572 19856 126636 19920
rect 156492 19856 156556 19920
rect 156572 19856 156636 19920
rect 186492 19856 186556 19920
rect 186572 19856 186636 19920
rect 201724 19856 201788 19920
rect 201804 19856 201868 19920
rect -1952 19776 -1888 19840
rect -1872 19776 -1808 19840
rect 6492 19776 6556 19840
rect 6572 19776 6636 19840
rect 36492 19776 36556 19840
rect 36572 19776 36636 19840
rect 66492 19776 66556 19840
rect 66572 19776 66636 19840
rect 96492 19776 96556 19840
rect 96572 19776 96636 19840
rect 126492 19776 126556 19840
rect 126572 19776 126636 19840
rect 156492 19776 156556 19840
rect 156572 19776 156636 19840
rect 186492 19776 186556 19840
rect 186572 19776 186636 19840
rect 201724 19776 201788 19840
rect 201804 19776 201868 19840
rect -1688 19592 -1624 19656
rect -1608 19592 -1544 19656
rect 20672 19592 20736 19656
rect 20752 19592 20816 19656
rect 50672 19592 50736 19656
rect 50752 19592 50816 19656
rect 80672 19592 80736 19656
rect 80752 19592 80816 19656
rect 110672 19592 110736 19656
rect 110752 19592 110816 19656
rect 140672 19592 140736 19656
rect 140752 19592 140816 19656
rect 170672 19592 170736 19656
rect 170752 19592 170816 19656
rect 201460 19592 201524 19656
rect 201540 19592 201604 19656
rect -1688 19512 -1624 19576
rect -1608 19512 -1544 19576
rect 20672 19512 20736 19576
rect 20752 19512 20816 19576
rect 50672 19512 50736 19576
rect 50752 19512 50816 19576
rect 80672 19512 80736 19576
rect 80752 19512 80816 19576
rect 110672 19512 110736 19576
rect 110752 19512 110816 19576
rect 140672 19512 140736 19576
rect 140752 19512 140816 19576
rect 170672 19512 170736 19576
rect 170752 19512 170816 19576
rect 201460 19512 201524 19576
rect 201540 19512 201604 19576
rect -1424 19328 -1360 19392
rect -1344 19328 -1280 19392
rect 5672 19328 5736 19392
rect 5752 19328 5816 19392
rect 35672 19328 35736 19392
rect 35752 19328 35816 19392
rect 65672 19328 65736 19392
rect 65752 19328 65816 19392
rect 95672 19328 95736 19392
rect 95752 19328 95816 19392
rect 125672 19328 125736 19392
rect 125752 19328 125816 19392
rect 155672 19328 155736 19392
rect 155752 19328 155816 19392
rect 185672 19328 185736 19392
rect 185752 19328 185816 19392
rect 201196 19328 201260 19392
rect 201276 19328 201340 19392
rect -1424 19248 -1360 19312
rect -1344 19248 -1280 19312
rect 5672 19248 5736 19312
rect 5752 19248 5816 19312
rect 35672 19248 35736 19312
rect 35752 19248 35816 19312
rect 65672 19248 65736 19312
rect 65752 19248 65816 19312
rect 95672 19248 95736 19312
rect 95752 19248 95816 19312
rect 125672 19248 125736 19312
rect 125752 19248 125816 19312
rect 155672 19248 155736 19312
rect 155752 19248 155816 19312
rect 185672 19248 185736 19312
rect 185752 19248 185816 19312
rect 201196 19248 201260 19312
rect 201276 19248 201340 19312
rect -1160 19064 -1096 19128
rect -1080 19064 -1016 19128
rect 19852 19064 19916 19128
rect 19932 19064 19996 19128
rect 49852 19064 49916 19128
rect 49932 19064 49996 19128
rect 79852 19064 79916 19128
rect 79932 19064 79996 19128
rect 109852 19064 109916 19128
rect 109932 19064 109996 19128
rect 139852 19064 139916 19128
rect 139932 19064 139996 19128
rect 169852 19064 169916 19128
rect 169932 19064 169996 19128
rect 200932 19064 200996 19128
rect 201012 19064 201076 19128
rect -1160 18984 -1096 19048
rect -1080 18984 -1016 19048
rect 19852 18984 19916 19048
rect 19932 18984 19996 19048
rect 49852 18984 49916 19048
rect 49932 18984 49996 19048
rect 79852 18984 79916 19048
rect 79932 18984 79996 19048
rect 109852 18984 109916 19048
rect 109932 18984 109996 19048
rect 139852 18984 139916 19048
rect 139932 18984 139996 19048
rect 169852 18984 169916 19048
rect 169932 18984 169996 19048
rect 200932 18984 200996 19048
rect 201012 18984 201076 19048
rect -896 18800 -832 18864
rect -816 18800 -752 18864
rect 4852 18800 4916 18864
rect 4932 18800 4996 18864
rect 34852 18800 34916 18864
rect 34932 18800 34996 18864
rect 64852 18800 64916 18864
rect 64932 18800 64996 18864
rect 94852 18800 94916 18864
rect 94932 18800 94996 18864
rect 124852 18800 124916 18864
rect 124932 18800 124996 18864
rect 154852 18800 154916 18864
rect 154932 18800 154996 18864
rect 184852 18800 184916 18864
rect 184932 18800 184996 18864
rect 200668 18800 200732 18864
rect 200748 18800 200812 18864
rect -896 18720 -832 18784
rect -816 18720 -752 18784
rect 4852 18720 4916 18784
rect 4932 18720 4996 18784
rect 34852 18720 34916 18784
rect 34932 18720 34996 18784
rect 64852 18720 64916 18784
rect 64932 18720 64996 18784
rect 94852 18720 94916 18784
rect 94932 18720 94996 18784
rect 124852 18720 124916 18784
rect 124932 18720 124996 18784
rect 154852 18720 154916 18784
rect 154932 18720 154996 18784
rect 184852 18720 184916 18784
rect 184932 18720 184996 18784
rect 200668 18720 200732 18784
rect 200748 18720 200812 18784
rect -632 18536 -568 18600
rect -552 18536 -488 18600
rect 19032 18536 19096 18600
rect 19112 18536 19176 18600
rect 49032 18536 49096 18600
rect 49112 18536 49176 18600
rect 79032 18536 79096 18600
rect 79112 18536 79176 18600
rect 109032 18536 109096 18600
rect 109112 18536 109176 18600
rect 139032 18536 139096 18600
rect 139112 18536 139176 18600
rect 169032 18536 169096 18600
rect 169112 18536 169176 18600
rect 200404 18536 200468 18600
rect 200484 18536 200548 18600
rect -632 18456 -568 18520
rect -552 18456 -488 18520
rect 19032 18456 19096 18520
rect 19112 18456 19176 18520
rect 49032 18456 49096 18520
rect 49112 18456 49176 18520
rect 79032 18456 79096 18520
rect 79112 18456 79176 18520
rect 109032 18456 109096 18520
rect 109112 18456 109176 18520
rect 139032 18456 139096 18520
rect 139112 18456 139176 18520
rect 169032 18456 169096 18520
rect 169112 18456 169176 18520
rect 200404 18456 200468 18520
rect 200484 18456 200548 18520
rect -368 18272 -304 18336
rect -288 18272 -224 18336
rect 4032 18272 4096 18336
rect 4112 18272 4176 18336
rect 34032 18272 34096 18336
rect 34112 18272 34176 18336
rect 64032 18272 64096 18336
rect 64112 18272 64176 18336
rect 94032 18272 94096 18336
rect 94112 18272 94176 18336
rect 124032 18272 124096 18336
rect 124112 18272 124176 18336
rect 154032 18272 154096 18336
rect 154112 18272 154176 18336
rect 184032 18272 184096 18336
rect 184112 18272 184176 18336
rect 200140 18272 200204 18336
rect 200220 18272 200284 18336
rect -368 18192 -304 18256
rect -288 18192 -224 18256
rect 4032 18192 4096 18256
rect 4112 18192 4176 18256
rect 34032 18192 34096 18256
rect 34112 18192 34176 18256
rect 64032 18192 64096 18256
rect 64112 18192 64176 18256
rect 94032 18192 94096 18256
rect 94112 18192 94176 18256
rect 124032 18192 124096 18256
rect 124112 18192 124176 18256
rect 154032 18192 154096 18256
rect 154112 18192 154176 18256
rect 184032 18192 184096 18256
rect 184112 18192 184176 18256
rect 200140 18192 200204 18256
rect 200220 18192 200284 18256
rect -368 -304 -304 -240
rect -288 -304 -224 -240
rect 4032 -304 4096 -240
rect 4112 -304 4176 -240
rect 34032 -304 34096 -240
rect 34112 -304 34176 -240
rect 64032 -304 64096 -240
rect 64112 -304 64176 -240
rect 94032 -304 94096 -240
rect 94112 -304 94176 -240
rect 124032 -304 124096 -240
rect 124112 -304 124176 -240
rect 154032 -304 154096 -240
rect 154112 -304 154176 -240
rect 184032 -304 184096 -240
rect 184112 -304 184176 -240
rect 200140 -304 200204 -240
rect 200220 -304 200284 -240
rect -368 -384 -304 -320
rect -288 -384 -224 -320
rect 4032 -384 4096 -320
rect 4112 -384 4176 -320
rect 34032 -384 34096 -320
rect 34112 -384 34176 -320
rect 64032 -384 64096 -320
rect 64112 -384 64176 -320
rect 94032 -384 94096 -320
rect 94112 -384 94176 -320
rect 124032 -384 124096 -320
rect 124112 -384 124176 -320
rect 154032 -384 154096 -320
rect 154112 -384 154176 -320
rect 184032 -384 184096 -320
rect 184112 -384 184176 -320
rect 200140 -384 200204 -320
rect 200220 -384 200284 -320
rect -632 -568 -568 -504
rect -552 -568 -488 -504
rect 19032 -568 19096 -504
rect 19112 -568 19176 -504
rect 49032 -568 49096 -504
rect 49112 -568 49176 -504
rect 79032 -568 79096 -504
rect 79112 -568 79176 -504
rect 109032 -568 109096 -504
rect 109112 -568 109176 -504
rect 139032 -568 139096 -504
rect 139112 -568 139176 -504
rect 169032 -568 169096 -504
rect 169112 -568 169176 -504
rect 200404 -568 200468 -504
rect 200484 -568 200548 -504
rect -632 -648 -568 -584
rect -552 -648 -488 -584
rect 19032 -648 19096 -584
rect 19112 -648 19176 -584
rect 49032 -648 49096 -584
rect 49112 -648 49176 -584
rect 79032 -648 79096 -584
rect 79112 -648 79176 -584
rect 109032 -648 109096 -584
rect 109112 -648 109176 -584
rect 139032 -648 139096 -584
rect 139112 -648 139176 -584
rect 169032 -648 169096 -584
rect 169112 -648 169176 -584
rect 200404 -648 200468 -584
rect 200484 -648 200548 -584
rect -896 -832 -832 -768
rect -816 -832 -752 -768
rect 4852 -832 4916 -768
rect 4932 -832 4996 -768
rect 34852 -832 34916 -768
rect 34932 -832 34996 -768
rect 64852 -832 64916 -768
rect 64932 -832 64996 -768
rect 94852 -832 94916 -768
rect 94932 -832 94996 -768
rect 124852 -832 124916 -768
rect 124932 -832 124996 -768
rect 154852 -832 154916 -768
rect 154932 -832 154996 -768
rect 184852 -832 184916 -768
rect 184932 -832 184996 -768
rect 200668 -832 200732 -768
rect 200748 -832 200812 -768
rect -896 -912 -832 -848
rect -816 -912 -752 -848
rect 4852 -912 4916 -848
rect 4932 -912 4996 -848
rect 34852 -912 34916 -848
rect 34932 -912 34996 -848
rect 64852 -912 64916 -848
rect 64932 -912 64996 -848
rect 94852 -912 94916 -848
rect 94932 -912 94996 -848
rect 124852 -912 124916 -848
rect 124932 -912 124996 -848
rect 154852 -912 154916 -848
rect 154932 -912 154996 -848
rect 184852 -912 184916 -848
rect 184932 -912 184996 -848
rect 200668 -912 200732 -848
rect 200748 -912 200812 -848
rect -1160 -1096 -1096 -1032
rect -1080 -1096 -1016 -1032
rect 19852 -1096 19916 -1032
rect 19932 -1096 19996 -1032
rect 49852 -1096 49916 -1032
rect 49932 -1096 49996 -1032
rect 79852 -1096 79916 -1032
rect 79932 -1096 79996 -1032
rect 109852 -1096 109916 -1032
rect 109932 -1096 109996 -1032
rect 139852 -1096 139916 -1032
rect 139932 -1096 139996 -1032
rect 169852 -1096 169916 -1032
rect 169932 -1096 169996 -1032
rect 200932 -1096 200996 -1032
rect 201012 -1096 201076 -1032
rect -1160 -1176 -1096 -1112
rect -1080 -1176 -1016 -1112
rect 19852 -1176 19916 -1112
rect 19932 -1176 19996 -1112
rect 49852 -1176 49916 -1112
rect 49932 -1176 49996 -1112
rect 79852 -1176 79916 -1112
rect 79932 -1176 79996 -1112
rect 109852 -1176 109916 -1112
rect 109932 -1176 109996 -1112
rect 139852 -1176 139916 -1112
rect 139932 -1176 139996 -1112
rect 169852 -1176 169916 -1112
rect 169932 -1176 169996 -1112
rect 200932 -1176 200996 -1112
rect 201012 -1176 201076 -1112
rect -1424 -1360 -1360 -1296
rect -1344 -1360 -1280 -1296
rect 5672 -1360 5736 -1296
rect 5752 -1360 5816 -1296
rect 35672 -1360 35736 -1296
rect 35752 -1360 35816 -1296
rect 65672 -1360 65736 -1296
rect 65752 -1360 65816 -1296
rect 95672 -1360 95736 -1296
rect 95752 -1360 95816 -1296
rect 125672 -1360 125736 -1296
rect 125752 -1360 125816 -1296
rect 155672 -1360 155736 -1296
rect 155752 -1360 155816 -1296
rect 185672 -1360 185736 -1296
rect 185752 -1360 185816 -1296
rect 201196 -1360 201260 -1296
rect 201276 -1360 201340 -1296
rect -1424 -1440 -1360 -1376
rect -1344 -1440 -1280 -1376
rect 5672 -1440 5736 -1376
rect 5752 -1440 5816 -1376
rect 35672 -1440 35736 -1376
rect 35752 -1440 35816 -1376
rect 65672 -1440 65736 -1376
rect 65752 -1440 65816 -1376
rect 95672 -1440 95736 -1376
rect 95752 -1440 95816 -1376
rect 125672 -1440 125736 -1376
rect 125752 -1440 125816 -1376
rect 155672 -1440 155736 -1376
rect 155752 -1440 155816 -1376
rect 185672 -1440 185736 -1376
rect 185752 -1440 185816 -1376
rect 201196 -1440 201260 -1376
rect 201276 -1440 201340 -1376
rect -1688 -1624 -1624 -1560
rect -1608 -1624 -1544 -1560
rect 20672 -1624 20736 -1560
rect 20752 -1624 20816 -1560
rect 50672 -1624 50736 -1560
rect 50752 -1624 50816 -1560
rect 80672 -1624 80736 -1560
rect 80752 -1624 80816 -1560
rect 110672 -1624 110736 -1560
rect 110752 -1624 110816 -1560
rect 140672 -1624 140736 -1560
rect 140752 -1624 140816 -1560
rect 170672 -1624 170736 -1560
rect 170752 -1624 170816 -1560
rect 201460 -1624 201524 -1560
rect 201540 -1624 201604 -1560
rect -1688 -1704 -1624 -1640
rect -1608 -1704 -1544 -1640
rect 20672 -1704 20736 -1640
rect 20752 -1704 20816 -1640
rect 50672 -1704 50736 -1640
rect 50752 -1704 50816 -1640
rect 80672 -1704 80736 -1640
rect 80752 -1704 80816 -1640
rect 110672 -1704 110736 -1640
rect 110752 -1704 110816 -1640
rect 140672 -1704 140736 -1640
rect 140752 -1704 140816 -1640
rect 170672 -1704 170736 -1640
rect 170752 -1704 170816 -1640
rect 201460 -1704 201524 -1640
rect 201540 -1704 201604 -1640
rect -1952 -1888 -1888 -1824
rect -1872 -1888 -1808 -1824
rect 6492 -1888 6556 -1824
rect 6572 -1888 6636 -1824
rect 36492 -1888 36556 -1824
rect 36572 -1888 36636 -1824
rect 66492 -1888 66556 -1824
rect 66572 -1888 66636 -1824
rect 96492 -1888 96556 -1824
rect 96572 -1888 96636 -1824
rect 126492 -1888 126556 -1824
rect 126572 -1888 126636 -1824
rect 156492 -1888 156556 -1824
rect 156572 -1888 156636 -1824
rect 186492 -1888 186556 -1824
rect 186572 -1888 186636 -1824
rect 201724 -1888 201788 -1824
rect 201804 -1888 201868 -1824
rect -1952 -1968 -1888 -1904
rect -1872 -1968 -1808 -1904
rect 6492 -1968 6556 -1904
rect 6572 -1968 6636 -1904
rect 36492 -1968 36556 -1904
rect 36572 -1968 36636 -1904
rect 66492 -1968 66556 -1904
rect 66572 -1968 66636 -1904
rect 96492 -1968 96556 -1904
rect 96572 -1968 96636 -1904
rect 126492 -1968 126556 -1904
rect 126572 -1968 126636 -1904
rect 156492 -1968 156556 -1904
rect 156572 -1968 156636 -1904
rect 186492 -1968 186556 -1904
rect 186572 -1968 186636 -1904
rect 201724 -1968 201788 -1904
rect 201804 -1968 201868 -1904
rect -2216 -2152 -2152 -2088
rect -2136 -2152 -2072 -2088
rect 21492 -2152 21556 -2088
rect 21572 -2152 21636 -2088
rect 51492 -2152 51556 -2088
rect 51572 -2152 51636 -2088
rect 81492 -2152 81556 -2088
rect 81572 -2152 81636 -2088
rect 111492 -2152 111556 -2088
rect 111572 -2152 111636 -2088
rect 141492 -2152 141556 -2088
rect 141572 -2152 141636 -2088
rect 171492 -2152 171556 -2088
rect 171572 -2152 171636 -2088
rect 201988 -2152 202052 -2088
rect 202068 -2152 202132 -2088
rect -2216 -2232 -2152 -2168
rect -2136 -2232 -2072 -2168
rect 21492 -2232 21556 -2168
rect 21572 -2232 21636 -2168
rect 51492 -2232 51556 -2168
rect 51572 -2232 51636 -2168
rect 81492 -2232 81556 -2168
rect 81572 -2232 81636 -2168
rect 111492 -2232 111556 -2168
rect 111572 -2232 111636 -2168
rect 141492 -2232 141556 -2168
rect 141572 -2232 141636 -2168
rect 171492 -2232 171556 -2168
rect 171572 -2232 171636 -2168
rect 201988 -2232 202052 -2168
rect 202068 -2232 202132 -2168
rect -2480 -2416 -2416 -2352
rect -2400 -2416 -2336 -2352
rect 7312 -2416 7376 -2352
rect 7392 -2416 7456 -2352
rect 37312 -2416 37376 -2352
rect 37392 -2416 37456 -2352
rect 67312 -2416 67376 -2352
rect 67392 -2416 67456 -2352
rect 97312 -2416 97376 -2352
rect 97392 -2416 97456 -2352
rect 127312 -2416 127376 -2352
rect 127392 -2416 127456 -2352
rect 157312 -2416 157376 -2352
rect 157392 -2416 157456 -2352
rect 187312 -2416 187376 -2352
rect 187392 -2416 187456 -2352
rect 202252 -2416 202316 -2352
rect 202332 -2416 202396 -2352
rect -2480 -2496 -2416 -2432
rect -2400 -2496 -2336 -2432
rect 7312 -2496 7376 -2432
rect 7392 -2496 7456 -2432
rect 37312 -2496 37376 -2432
rect 37392 -2496 37456 -2432
rect 67312 -2496 67376 -2432
rect 67392 -2496 67456 -2432
rect 97312 -2496 97376 -2432
rect 97392 -2496 97456 -2432
rect 127312 -2496 127376 -2432
rect 127392 -2496 127456 -2432
rect 157312 -2496 157376 -2432
rect 157392 -2496 157456 -2432
rect 187312 -2496 187376 -2432
rect 187392 -2496 187456 -2432
rect 202252 -2496 202316 -2432
rect 202332 -2496 202396 -2432
rect -2744 -2680 -2680 -2616
rect -2664 -2680 -2600 -2616
rect 22312 -2680 22376 -2616
rect 22392 -2680 22456 -2616
rect 52312 -2680 52376 -2616
rect 52392 -2680 52456 -2616
rect 82312 -2680 82376 -2616
rect 82392 -2680 82456 -2616
rect 112312 -2680 112376 -2616
rect 112392 -2680 112456 -2616
rect 142312 -2680 142376 -2616
rect 142392 -2680 142456 -2616
rect 172312 -2680 172376 -2616
rect 172392 -2680 172456 -2616
rect 202516 -2680 202580 -2616
rect 202596 -2680 202660 -2616
rect -2744 -2760 -2680 -2696
rect -2664 -2760 -2600 -2696
rect 22312 -2760 22376 -2696
rect 22392 -2760 22456 -2696
rect 52312 -2760 52376 -2696
rect 52392 -2760 52456 -2696
rect 82312 -2760 82376 -2696
rect 82392 -2760 82456 -2696
rect 112312 -2760 112376 -2696
rect 112392 -2760 112456 -2696
rect 142312 -2760 142376 -2696
rect 142392 -2760 142456 -2696
rect 172312 -2760 172376 -2696
rect 172392 -2760 172456 -2696
rect 202516 -2760 202580 -2696
rect 202596 -2760 202660 -2696
<< metal4 >>
rect -2762 20712 -2582 20730
rect -2762 20648 -2744 20712
rect -2680 20648 -2664 20712
rect -2600 20648 -2582 20712
rect -2762 20632 -2582 20648
rect -2762 20568 -2744 20632
rect -2680 20568 -2664 20632
rect -2600 20568 -2582 20632
rect -2762 -2616 -2582 20568
rect -2498 20448 -2318 20466
rect -2498 20384 -2480 20448
rect -2416 20384 -2400 20448
rect -2336 20384 -2318 20448
rect -2498 20368 -2318 20384
rect -2498 20304 -2480 20368
rect -2416 20304 -2400 20368
rect -2336 20304 -2318 20368
rect -2498 -2352 -2318 20304
rect 7294 20448 7474 20730
rect 7294 20384 7312 20448
rect 7376 20384 7392 20448
rect 7456 20384 7474 20448
rect 7294 20368 7474 20384
rect 7294 20304 7312 20368
rect 7376 20304 7392 20368
rect 7456 20304 7474 20368
rect -2234 20184 -2054 20202
rect -2234 20120 -2216 20184
rect -2152 20120 -2136 20184
rect -2072 20120 -2054 20184
rect -2234 20104 -2054 20120
rect -2234 20040 -2216 20104
rect -2152 20040 -2136 20104
rect -2072 20040 -2054 20104
rect -2234 -2088 -2054 20040
rect -1970 19920 -1790 19938
rect -1970 19856 -1952 19920
rect -1888 19856 -1872 19920
rect -1808 19856 -1790 19920
rect -1970 19840 -1790 19856
rect -1970 19776 -1952 19840
rect -1888 19776 -1872 19840
rect -1808 19776 -1790 19840
rect -1970 -1824 -1790 19776
rect 6474 19920 6654 20202
rect 6474 19856 6492 19920
rect 6556 19856 6572 19920
rect 6636 19856 6654 19920
rect 6474 19840 6654 19856
rect 6474 19776 6492 19840
rect 6556 19776 6572 19840
rect 6636 19776 6654 19840
rect -1706 19656 -1526 19674
rect -1706 19592 -1688 19656
rect -1624 19592 -1608 19656
rect -1544 19592 -1526 19656
rect -1706 19576 -1526 19592
rect -1706 19512 -1688 19576
rect -1624 19512 -1608 19576
rect -1544 19512 -1526 19576
rect -1706 -1560 -1526 19512
rect -1442 19392 -1262 19410
rect -1442 19328 -1424 19392
rect -1360 19328 -1344 19392
rect -1280 19328 -1262 19392
rect -1442 19312 -1262 19328
rect -1442 19248 -1424 19312
rect -1360 19248 -1344 19312
rect -1280 19248 -1262 19312
rect -1442 -1296 -1262 19248
rect 5654 19392 5834 19674
rect 5654 19328 5672 19392
rect 5736 19328 5752 19392
rect 5816 19328 5834 19392
rect 5654 19312 5834 19328
rect 5654 19248 5672 19312
rect 5736 19248 5752 19312
rect 5816 19248 5834 19312
rect -1178 19128 -998 19146
rect -1178 19064 -1160 19128
rect -1096 19064 -1080 19128
rect -1016 19064 -998 19128
rect -1178 19048 -998 19064
rect -1178 18984 -1160 19048
rect -1096 18984 -1080 19048
rect -1016 18984 -998 19048
rect -1178 -1032 -998 18984
rect -914 18864 -734 18882
rect -914 18800 -896 18864
rect -832 18800 -816 18864
rect -752 18800 -734 18864
rect -914 18784 -734 18800
rect -914 18720 -896 18784
rect -832 18720 -816 18784
rect -752 18720 -734 18784
rect -914 -768 -734 18720
rect 4834 18864 5014 19146
rect 4834 18800 4852 18864
rect 4916 18800 4932 18864
rect 4996 18800 5014 18864
rect 4834 18784 5014 18800
rect 4834 18720 4852 18784
rect 4916 18720 4932 18784
rect 4996 18720 5014 18784
rect -650 18600 -470 18618
rect -650 18536 -632 18600
rect -568 18536 -552 18600
rect -488 18536 -470 18600
rect -650 18520 -470 18536
rect -650 18456 -632 18520
rect -568 18456 -552 18520
rect -488 18456 -470 18520
rect -650 -504 -470 18456
rect -386 18336 -206 18354
rect -386 18272 -368 18336
rect -304 18272 -288 18336
rect -224 18272 -206 18336
rect -386 18256 -206 18272
rect -386 18192 -368 18256
rect -304 18192 -288 18256
rect -224 18192 -206 18256
rect -386 -240 -206 18192
rect -386 -304 -368 -240
rect -304 -304 -288 -240
rect -224 -304 -206 -240
rect -386 -320 -206 -304
rect -386 -384 -368 -320
rect -304 -384 -288 -320
rect -224 -384 -206 -320
rect -386 -402 -206 -384
rect 4014 18336 4194 18618
rect 4014 18272 4032 18336
rect 4096 18272 4112 18336
rect 4176 18272 4194 18336
rect 4014 18256 4194 18272
rect 4014 18192 4032 18256
rect 4096 18192 4112 18256
rect 4176 18192 4194 18256
rect 4014 17940 4194 18192
rect 4834 17940 5014 18720
rect 5654 17940 5834 19248
rect 6474 17940 6654 19776
rect 7294 17940 7474 20304
rect 22294 20712 22474 20730
rect 22294 20648 22312 20712
rect 22376 20648 22392 20712
rect 22456 20648 22474 20712
rect 22294 20632 22474 20648
rect 22294 20568 22312 20632
rect 22376 20568 22392 20632
rect 22456 20568 22474 20632
rect 21474 20184 21654 20202
rect 21474 20120 21492 20184
rect 21556 20120 21572 20184
rect 21636 20120 21654 20184
rect 21474 20104 21654 20120
rect 21474 20040 21492 20104
rect 21556 20040 21572 20104
rect 21636 20040 21654 20104
rect 20654 19656 20834 19674
rect 20654 19592 20672 19656
rect 20736 19592 20752 19656
rect 20816 19592 20834 19656
rect 20654 19576 20834 19592
rect 20654 19512 20672 19576
rect 20736 19512 20752 19576
rect 20816 19512 20834 19576
rect 19834 19128 20014 19146
rect 19834 19064 19852 19128
rect 19916 19064 19932 19128
rect 19996 19064 20014 19128
rect 19834 19048 20014 19064
rect 19834 18984 19852 19048
rect 19916 18984 19932 19048
rect 19996 18984 20014 19048
rect 19014 18600 19194 18618
rect 19014 18536 19032 18600
rect 19096 18536 19112 18600
rect 19176 18536 19194 18600
rect 19014 18520 19194 18536
rect 19014 18456 19032 18520
rect 19096 18456 19112 18520
rect 19176 18456 19194 18520
rect 19014 17940 19194 18456
rect 19834 17940 20014 18984
rect 20654 17940 20834 19512
rect 21474 17940 21654 20040
rect 22294 17940 22474 20568
rect 37294 20448 37474 20730
rect 37294 20384 37312 20448
rect 37376 20384 37392 20448
rect 37456 20384 37474 20448
rect 37294 20368 37474 20384
rect 37294 20304 37312 20368
rect 37376 20304 37392 20368
rect 37456 20304 37474 20368
rect 36474 19920 36654 20202
rect 36474 19856 36492 19920
rect 36556 19856 36572 19920
rect 36636 19856 36654 19920
rect 36474 19840 36654 19856
rect 36474 19776 36492 19840
rect 36556 19776 36572 19840
rect 36636 19776 36654 19840
rect 35654 19392 35834 19674
rect 35654 19328 35672 19392
rect 35736 19328 35752 19392
rect 35816 19328 35834 19392
rect 35654 19312 35834 19328
rect 35654 19248 35672 19312
rect 35736 19248 35752 19312
rect 35816 19248 35834 19312
rect 34834 18864 35014 19146
rect 34834 18800 34852 18864
rect 34916 18800 34932 18864
rect 34996 18800 35014 18864
rect 34834 18784 35014 18800
rect 34834 18720 34852 18784
rect 34916 18720 34932 18784
rect 34996 18720 35014 18784
rect 34014 18336 34194 18618
rect 34014 18272 34032 18336
rect 34096 18272 34112 18336
rect 34176 18272 34194 18336
rect 34014 18256 34194 18272
rect 34014 18192 34032 18256
rect 34096 18192 34112 18256
rect 34176 18192 34194 18256
rect 34014 17940 34194 18192
rect 34834 17940 35014 18720
rect 35654 17940 35834 19248
rect 36474 17940 36654 19776
rect 37294 17940 37474 20304
rect 52294 20712 52474 20730
rect 52294 20648 52312 20712
rect 52376 20648 52392 20712
rect 52456 20648 52474 20712
rect 52294 20632 52474 20648
rect 52294 20568 52312 20632
rect 52376 20568 52392 20632
rect 52456 20568 52474 20632
rect 51474 20184 51654 20202
rect 51474 20120 51492 20184
rect 51556 20120 51572 20184
rect 51636 20120 51654 20184
rect 51474 20104 51654 20120
rect 51474 20040 51492 20104
rect 51556 20040 51572 20104
rect 51636 20040 51654 20104
rect 50654 19656 50834 19674
rect 50654 19592 50672 19656
rect 50736 19592 50752 19656
rect 50816 19592 50834 19656
rect 50654 19576 50834 19592
rect 50654 19512 50672 19576
rect 50736 19512 50752 19576
rect 50816 19512 50834 19576
rect 49834 19128 50014 19146
rect 49834 19064 49852 19128
rect 49916 19064 49932 19128
rect 49996 19064 50014 19128
rect 49834 19048 50014 19064
rect 49834 18984 49852 19048
rect 49916 18984 49932 19048
rect 49996 18984 50014 19048
rect 49014 18600 49194 18618
rect 49014 18536 49032 18600
rect 49096 18536 49112 18600
rect 49176 18536 49194 18600
rect 49014 18520 49194 18536
rect 49014 18456 49032 18520
rect 49096 18456 49112 18520
rect 49176 18456 49194 18520
rect 49014 17940 49194 18456
rect 49834 17940 50014 18984
rect 50654 17940 50834 19512
rect 51474 17940 51654 20040
rect 52294 17940 52474 20568
rect 67294 20448 67474 20730
rect 67294 20384 67312 20448
rect 67376 20384 67392 20448
rect 67456 20384 67474 20448
rect 67294 20368 67474 20384
rect 67294 20304 67312 20368
rect 67376 20304 67392 20368
rect 67456 20304 67474 20368
rect 66474 19920 66654 20202
rect 66474 19856 66492 19920
rect 66556 19856 66572 19920
rect 66636 19856 66654 19920
rect 66474 19840 66654 19856
rect 66474 19776 66492 19840
rect 66556 19776 66572 19840
rect 66636 19776 66654 19840
rect 65654 19392 65834 19674
rect 65654 19328 65672 19392
rect 65736 19328 65752 19392
rect 65816 19328 65834 19392
rect 65654 19312 65834 19328
rect 65654 19248 65672 19312
rect 65736 19248 65752 19312
rect 65816 19248 65834 19312
rect 64834 18864 65014 19146
rect 64834 18800 64852 18864
rect 64916 18800 64932 18864
rect 64996 18800 65014 18864
rect 64834 18784 65014 18800
rect 64834 18720 64852 18784
rect 64916 18720 64932 18784
rect 64996 18720 65014 18784
rect 64014 18336 64194 18618
rect 64014 18272 64032 18336
rect 64096 18272 64112 18336
rect 64176 18272 64194 18336
rect 64014 18256 64194 18272
rect 64014 18192 64032 18256
rect 64096 18192 64112 18256
rect 64176 18192 64194 18256
rect 64014 17940 64194 18192
rect 64834 17940 65014 18720
rect 65654 17940 65834 19248
rect 66474 17940 66654 19776
rect 67294 17940 67474 20304
rect 82294 20712 82474 20730
rect 82294 20648 82312 20712
rect 82376 20648 82392 20712
rect 82456 20648 82474 20712
rect 82294 20632 82474 20648
rect 82294 20568 82312 20632
rect 82376 20568 82392 20632
rect 82456 20568 82474 20632
rect 81474 20184 81654 20202
rect 81474 20120 81492 20184
rect 81556 20120 81572 20184
rect 81636 20120 81654 20184
rect 81474 20104 81654 20120
rect 81474 20040 81492 20104
rect 81556 20040 81572 20104
rect 81636 20040 81654 20104
rect 80654 19656 80834 19674
rect 80654 19592 80672 19656
rect 80736 19592 80752 19656
rect 80816 19592 80834 19656
rect 80654 19576 80834 19592
rect 80654 19512 80672 19576
rect 80736 19512 80752 19576
rect 80816 19512 80834 19576
rect 79834 19128 80014 19146
rect 79834 19064 79852 19128
rect 79916 19064 79932 19128
rect 79996 19064 80014 19128
rect 79834 19048 80014 19064
rect 79834 18984 79852 19048
rect 79916 18984 79932 19048
rect 79996 18984 80014 19048
rect 79014 18600 79194 18618
rect 79014 18536 79032 18600
rect 79096 18536 79112 18600
rect 79176 18536 79194 18600
rect 79014 18520 79194 18536
rect 79014 18456 79032 18520
rect 79096 18456 79112 18520
rect 79176 18456 79194 18520
rect 79014 17940 79194 18456
rect 79834 17940 80014 18984
rect 80654 17940 80834 19512
rect 81474 17940 81654 20040
rect 82294 17940 82474 20568
rect 97294 20448 97474 20730
rect 97294 20384 97312 20448
rect 97376 20384 97392 20448
rect 97456 20384 97474 20448
rect 97294 20368 97474 20384
rect 97294 20304 97312 20368
rect 97376 20304 97392 20368
rect 97456 20304 97474 20368
rect 96474 19920 96654 20202
rect 96474 19856 96492 19920
rect 96556 19856 96572 19920
rect 96636 19856 96654 19920
rect 96474 19840 96654 19856
rect 96474 19776 96492 19840
rect 96556 19776 96572 19840
rect 96636 19776 96654 19840
rect 95654 19392 95834 19674
rect 95654 19328 95672 19392
rect 95736 19328 95752 19392
rect 95816 19328 95834 19392
rect 95654 19312 95834 19328
rect 95654 19248 95672 19312
rect 95736 19248 95752 19312
rect 95816 19248 95834 19312
rect 94834 18864 95014 19146
rect 94834 18800 94852 18864
rect 94916 18800 94932 18864
rect 94996 18800 95014 18864
rect 94834 18784 95014 18800
rect 94834 18720 94852 18784
rect 94916 18720 94932 18784
rect 94996 18720 95014 18784
rect 94014 18336 94194 18618
rect 94014 18272 94032 18336
rect 94096 18272 94112 18336
rect 94176 18272 94194 18336
rect 94014 18256 94194 18272
rect 94014 18192 94032 18256
rect 94096 18192 94112 18256
rect 94176 18192 94194 18256
rect 94014 17940 94194 18192
rect 94834 17940 95014 18720
rect 95654 17940 95834 19248
rect 96474 17940 96654 19776
rect 97294 17940 97474 20304
rect 112294 20712 112474 20730
rect 112294 20648 112312 20712
rect 112376 20648 112392 20712
rect 112456 20648 112474 20712
rect 112294 20632 112474 20648
rect 112294 20568 112312 20632
rect 112376 20568 112392 20632
rect 112456 20568 112474 20632
rect 111474 20184 111654 20202
rect 111474 20120 111492 20184
rect 111556 20120 111572 20184
rect 111636 20120 111654 20184
rect 111474 20104 111654 20120
rect 111474 20040 111492 20104
rect 111556 20040 111572 20104
rect 111636 20040 111654 20104
rect 110654 19656 110834 19674
rect 110654 19592 110672 19656
rect 110736 19592 110752 19656
rect 110816 19592 110834 19656
rect 110654 19576 110834 19592
rect 110654 19512 110672 19576
rect 110736 19512 110752 19576
rect 110816 19512 110834 19576
rect 109834 19128 110014 19146
rect 109834 19064 109852 19128
rect 109916 19064 109932 19128
rect 109996 19064 110014 19128
rect 109834 19048 110014 19064
rect 109834 18984 109852 19048
rect 109916 18984 109932 19048
rect 109996 18984 110014 19048
rect 109014 18600 109194 18618
rect 109014 18536 109032 18600
rect 109096 18536 109112 18600
rect 109176 18536 109194 18600
rect 109014 18520 109194 18536
rect 109014 18456 109032 18520
rect 109096 18456 109112 18520
rect 109176 18456 109194 18520
rect 109014 17940 109194 18456
rect 109834 17940 110014 18984
rect 110654 17940 110834 19512
rect 111474 17940 111654 20040
rect 112294 17940 112474 20568
rect 127294 20448 127474 20730
rect 127294 20384 127312 20448
rect 127376 20384 127392 20448
rect 127456 20384 127474 20448
rect 127294 20368 127474 20384
rect 127294 20304 127312 20368
rect 127376 20304 127392 20368
rect 127456 20304 127474 20368
rect 126474 19920 126654 20202
rect 126474 19856 126492 19920
rect 126556 19856 126572 19920
rect 126636 19856 126654 19920
rect 126474 19840 126654 19856
rect 126474 19776 126492 19840
rect 126556 19776 126572 19840
rect 126636 19776 126654 19840
rect 125654 19392 125834 19674
rect 125654 19328 125672 19392
rect 125736 19328 125752 19392
rect 125816 19328 125834 19392
rect 125654 19312 125834 19328
rect 125654 19248 125672 19312
rect 125736 19248 125752 19312
rect 125816 19248 125834 19312
rect 124834 18864 125014 19146
rect 124834 18800 124852 18864
rect 124916 18800 124932 18864
rect 124996 18800 125014 18864
rect 124834 18784 125014 18800
rect 124834 18720 124852 18784
rect 124916 18720 124932 18784
rect 124996 18720 125014 18784
rect 124014 18336 124194 18618
rect 124014 18272 124032 18336
rect 124096 18272 124112 18336
rect 124176 18272 124194 18336
rect 124014 18256 124194 18272
rect 124014 18192 124032 18256
rect 124096 18192 124112 18256
rect 124176 18192 124194 18256
rect 124014 17940 124194 18192
rect 124834 17940 125014 18720
rect 125654 17940 125834 19248
rect 126474 17940 126654 19776
rect 127294 17940 127474 20304
rect 142294 20712 142474 20730
rect 142294 20648 142312 20712
rect 142376 20648 142392 20712
rect 142456 20648 142474 20712
rect 142294 20632 142474 20648
rect 142294 20568 142312 20632
rect 142376 20568 142392 20632
rect 142456 20568 142474 20632
rect 141474 20184 141654 20202
rect 141474 20120 141492 20184
rect 141556 20120 141572 20184
rect 141636 20120 141654 20184
rect 141474 20104 141654 20120
rect 141474 20040 141492 20104
rect 141556 20040 141572 20104
rect 141636 20040 141654 20104
rect 140654 19656 140834 19674
rect 140654 19592 140672 19656
rect 140736 19592 140752 19656
rect 140816 19592 140834 19656
rect 140654 19576 140834 19592
rect 140654 19512 140672 19576
rect 140736 19512 140752 19576
rect 140816 19512 140834 19576
rect 139834 19128 140014 19146
rect 139834 19064 139852 19128
rect 139916 19064 139932 19128
rect 139996 19064 140014 19128
rect 139834 19048 140014 19064
rect 139834 18984 139852 19048
rect 139916 18984 139932 19048
rect 139996 18984 140014 19048
rect 139014 18600 139194 18618
rect 139014 18536 139032 18600
rect 139096 18536 139112 18600
rect 139176 18536 139194 18600
rect 139014 18520 139194 18536
rect 139014 18456 139032 18520
rect 139096 18456 139112 18520
rect 139176 18456 139194 18520
rect 139014 17940 139194 18456
rect 139834 17940 140014 18984
rect 140654 17940 140834 19512
rect 141474 17940 141654 20040
rect 142294 17940 142474 20568
rect 157294 20448 157474 20730
rect 157294 20384 157312 20448
rect 157376 20384 157392 20448
rect 157456 20384 157474 20448
rect 157294 20368 157474 20384
rect 157294 20304 157312 20368
rect 157376 20304 157392 20368
rect 157456 20304 157474 20368
rect 156474 19920 156654 20202
rect 156474 19856 156492 19920
rect 156556 19856 156572 19920
rect 156636 19856 156654 19920
rect 156474 19840 156654 19856
rect 156474 19776 156492 19840
rect 156556 19776 156572 19840
rect 156636 19776 156654 19840
rect 155654 19392 155834 19674
rect 155654 19328 155672 19392
rect 155736 19328 155752 19392
rect 155816 19328 155834 19392
rect 155654 19312 155834 19328
rect 155654 19248 155672 19312
rect 155736 19248 155752 19312
rect 155816 19248 155834 19312
rect 154834 18864 155014 19146
rect 154834 18800 154852 18864
rect 154916 18800 154932 18864
rect 154996 18800 155014 18864
rect 154834 18784 155014 18800
rect 154834 18720 154852 18784
rect 154916 18720 154932 18784
rect 154996 18720 155014 18784
rect 154014 18336 154194 18618
rect 154014 18272 154032 18336
rect 154096 18272 154112 18336
rect 154176 18272 154194 18336
rect 154014 18256 154194 18272
rect 154014 18192 154032 18256
rect 154096 18192 154112 18256
rect 154176 18192 154194 18256
rect 154014 17940 154194 18192
rect 154834 17940 155014 18720
rect 155654 17940 155834 19248
rect 156474 17940 156654 19776
rect 157294 17940 157474 20304
rect 172294 20712 172474 20730
rect 172294 20648 172312 20712
rect 172376 20648 172392 20712
rect 172456 20648 172474 20712
rect 172294 20632 172474 20648
rect 172294 20568 172312 20632
rect 172376 20568 172392 20632
rect 172456 20568 172474 20632
rect 171474 20184 171654 20202
rect 171474 20120 171492 20184
rect 171556 20120 171572 20184
rect 171636 20120 171654 20184
rect 171474 20104 171654 20120
rect 171474 20040 171492 20104
rect 171556 20040 171572 20104
rect 171636 20040 171654 20104
rect 170654 19656 170834 19674
rect 170654 19592 170672 19656
rect 170736 19592 170752 19656
rect 170816 19592 170834 19656
rect 170654 19576 170834 19592
rect 170654 19512 170672 19576
rect 170736 19512 170752 19576
rect 170816 19512 170834 19576
rect 169834 19128 170014 19146
rect 169834 19064 169852 19128
rect 169916 19064 169932 19128
rect 169996 19064 170014 19128
rect 169834 19048 170014 19064
rect 169834 18984 169852 19048
rect 169916 18984 169932 19048
rect 169996 18984 170014 19048
rect 169014 18600 169194 18618
rect 169014 18536 169032 18600
rect 169096 18536 169112 18600
rect 169176 18536 169194 18600
rect 169014 18520 169194 18536
rect 169014 18456 169032 18520
rect 169096 18456 169112 18520
rect 169176 18456 169194 18520
rect 169014 17940 169194 18456
rect 169834 17940 170014 18984
rect 170654 17940 170834 19512
rect 171474 17940 171654 20040
rect 172294 17940 172474 20568
rect 187294 20448 187474 20730
rect 202498 20712 202678 20730
rect 202498 20648 202516 20712
rect 202580 20648 202596 20712
rect 202660 20648 202678 20712
rect 202498 20632 202678 20648
rect 202498 20568 202516 20632
rect 202580 20568 202596 20632
rect 202660 20568 202678 20632
rect 187294 20384 187312 20448
rect 187376 20384 187392 20448
rect 187456 20384 187474 20448
rect 187294 20368 187474 20384
rect 187294 20304 187312 20368
rect 187376 20304 187392 20368
rect 187456 20304 187474 20368
rect 186474 19920 186654 20202
rect 186474 19856 186492 19920
rect 186556 19856 186572 19920
rect 186636 19856 186654 19920
rect 186474 19840 186654 19856
rect 186474 19776 186492 19840
rect 186556 19776 186572 19840
rect 186636 19776 186654 19840
rect 185654 19392 185834 19674
rect 185654 19328 185672 19392
rect 185736 19328 185752 19392
rect 185816 19328 185834 19392
rect 185654 19312 185834 19328
rect 185654 19248 185672 19312
rect 185736 19248 185752 19312
rect 185816 19248 185834 19312
rect 184834 18864 185014 19146
rect 184834 18800 184852 18864
rect 184916 18800 184932 18864
rect 184996 18800 185014 18864
rect 184834 18784 185014 18800
rect 184834 18720 184852 18784
rect 184916 18720 184932 18784
rect 184996 18720 185014 18784
rect 184014 18336 184194 18618
rect 184014 18272 184032 18336
rect 184096 18272 184112 18336
rect 184176 18272 184194 18336
rect 184014 18256 184194 18272
rect 184014 18192 184032 18256
rect 184096 18192 184112 18256
rect 184176 18192 184194 18256
rect 184014 17940 184194 18192
rect 184834 17940 185014 18720
rect 185654 17940 185834 19248
rect 186474 17940 186654 19776
rect 187294 17940 187474 20304
rect 202234 20448 202414 20466
rect 202234 20384 202252 20448
rect 202316 20384 202332 20448
rect 202396 20384 202414 20448
rect 202234 20368 202414 20384
rect 202234 20304 202252 20368
rect 202316 20304 202332 20368
rect 202396 20304 202414 20368
rect 201970 20184 202150 20202
rect 201970 20120 201988 20184
rect 202052 20120 202068 20184
rect 202132 20120 202150 20184
rect 201970 20104 202150 20120
rect 201970 20040 201988 20104
rect 202052 20040 202068 20104
rect 202132 20040 202150 20104
rect 201706 19920 201886 19938
rect 201706 19856 201724 19920
rect 201788 19856 201804 19920
rect 201868 19856 201886 19920
rect 201706 19840 201886 19856
rect 201706 19776 201724 19840
rect 201788 19776 201804 19840
rect 201868 19776 201886 19840
rect 201442 19656 201622 19674
rect 201442 19592 201460 19656
rect 201524 19592 201540 19656
rect 201604 19592 201622 19656
rect 201442 19576 201622 19592
rect 201442 19512 201460 19576
rect 201524 19512 201540 19576
rect 201604 19512 201622 19576
rect 201178 19392 201358 19410
rect 201178 19328 201196 19392
rect 201260 19328 201276 19392
rect 201340 19328 201358 19392
rect 201178 19312 201358 19328
rect 201178 19248 201196 19312
rect 201260 19248 201276 19312
rect 201340 19248 201358 19312
rect 200914 19128 201094 19146
rect 200914 19064 200932 19128
rect 200996 19064 201012 19128
rect 201076 19064 201094 19128
rect 200914 19048 201094 19064
rect 200914 18984 200932 19048
rect 200996 18984 201012 19048
rect 201076 18984 201094 19048
rect 200650 18864 200830 18882
rect 200650 18800 200668 18864
rect 200732 18800 200748 18864
rect 200812 18800 200830 18864
rect 200650 18784 200830 18800
rect 200650 18720 200668 18784
rect 200732 18720 200748 18784
rect 200812 18720 200830 18784
rect 200386 18600 200566 18618
rect 200386 18536 200404 18600
rect 200468 18536 200484 18600
rect 200548 18536 200566 18600
rect 200386 18520 200566 18536
rect 200386 18456 200404 18520
rect 200468 18456 200484 18520
rect 200548 18456 200566 18520
rect 200122 18336 200302 18354
rect 200122 18272 200140 18336
rect 200204 18272 200220 18336
rect 200284 18272 200302 18336
rect 200122 18256 200302 18272
rect 200122 18192 200140 18256
rect 200204 18192 200220 18256
rect 200284 18192 200302 18256
rect 4014 -240 4194 60
rect 4014 -304 4032 -240
rect 4096 -304 4112 -240
rect 4176 -304 4194 -240
rect 4014 -320 4194 -304
rect 4014 -384 4032 -320
rect 4096 -384 4112 -320
rect 4176 -384 4194 -320
rect -650 -568 -632 -504
rect -568 -568 -552 -504
rect -488 -568 -470 -504
rect -650 -584 -470 -568
rect -650 -648 -632 -584
rect -568 -648 -552 -584
rect -488 -648 -470 -584
rect -650 -666 -470 -648
rect 4014 -666 4194 -384
rect -914 -832 -896 -768
rect -832 -832 -816 -768
rect -752 -832 -734 -768
rect -914 -848 -734 -832
rect -914 -912 -896 -848
rect -832 -912 -816 -848
rect -752 -912 -734 -848
rect -914 -930 -734 -912
rect 4834 -768 5014 60
rect 4834 -832 4852 -768
rect 4916 -832 4932 -768
rect 4996 -832 5014 -768
rect 4834 -848 5014 -832
rect 4834 -912 4852 -848
rect 4916 -912 4932 -848
rect 4996 -912 5014 -848
rect -1178 -1096 -1160 -1032
rect -1096 -1096 -1080 -1032
rect -1016 -1096 -998 -1032
rect -1178 -1112 -998 -1096
rect -1178 -1176 -1160 -1112
rect -1096 -1176 -1080 -1112
rect -1016 -1176 -998 -1112
rect -1178 -1194 -998 -1176
rect 4834 -1194 5014 -912
rect -1442 -1360 -1424 -1296
rect -1360 -1360 -1344 -1296
rect -1280 -1360 -1262 -1296
rect -1442 -1376 -1262 -1360
rect -1442 -1440 -1424 -1376
rect -1360 -1440 -1344 -1376
rect -1280 -1440 -1262 -1376
rect -1442 -1458 -1262 -1440
rect 5654 -1296 5834 60
rect 5654 -1360 5672 -1296
rect 5736 -1360 5752 -1296
rect 5816 -1360 5834 -1296
rect 5654 -1376 5834 -1360
rect 5654 -1440 5672 -1376
rect 5736 -1440 5752 -1376
rect 5816 -1440 5834 -1376
rect -1706 -1624 -1688 -1560
rect -1624 -1624 -1608 -1560
rect -1544 -1624 -1526 -1560
rect -1706 -1640 -1526 -1624
rect -1706 -1704 -1688 -1640
rect -1624 -1704 -1608 -1640
rect -1544 -1704 -1526 -1640
rect -1706 -1722 -1526 -1704
rect 5654 -1722 5834 -1440
rect -1970 -1888 -1952 -1824
rect -1888 -1888 -1872 -1824
rect -1808 -1888 -1790 -1824
rect -1970 -1904 -1790 -1888
rect -1970 -1968 -1952 -1904
rect -1888 -1968 -1872 -1904
rect -1808 -1968 -1790 -1904
rect -1970 -1986 -1790 -1968
rect 6474 -1824 6654 60
rect 6474 -1888 6492 -1824
rect 6556 -1888 6572 -1824
rect 6636 -1888 6654 -1824
rect 6474 -1904 6654 -1888
rect 6474 -1968 6492 -1904
rect 6556 -1968 6572 -1904
rect 6636 -1968 6654 -1904
rect -2234 -2152 -2216 -2088
rect -2152 -2152 -2136 -2088
rect -2072 -2152 -2054 -2088
rect -2234 -2168 -2054 -2152
rect -2234 -2232 -2216 -2168
rect -2152 -2232 -2136 -2168
rect -2072 -2232 -2054 -2168
rect -2234 -2250 -2054 -2232
rect 6474 -2250 6654 -1968
rect -2498 -2416 -2480 -2352
rect -2416 -2416 -2400 -2352
rect -2336 -2416 -2318 -2352
rect -2498 -2432 -2318 -2416
rect -2498 -2496 -2480 -2432
rect -2416 -2496 -2400 -2432
rect -2336 -2496 -2318 -2432
rect -2498 -2514 -2318 -2496
rect 7294 -2352 7474 60
rect 19014 -504 19194 60
rect 19014 -568 19032 -504
rect 19096 -568 19112 -504
rect 19176 -568 19194 -504
rect 19014 -584 19194 -568
rect 19014 -648 19032 -584
rect 19096 -648 19112 -584
rect 19176 -648 19194 -584
rect 19014 -666 19194 -648
rect 19834 -1032 20014 60
rect 19834 -1096 19852 -1032
rect 19916 -1096 19932 -1032
rect 19996 -1096 20014 -1032
rect 19834 -1112 20014 -1096
rect 19834 -1176 19852 -1112
rect 19916 -1176 19932 -1112
rect 19996 -1176 20014 -1112
rect 19834 -1194 20014 -1176
rect 20654 -1560 20834 60
rect 20654 -1624 20672 -1560
rect 20736 -1624 20752 -1560
rect 20816 -1624 20834 -1560
rect 20654 -1640 20834 -1624
rect 20654 -1704 20672 -1640
rect 20736 -1704 20752 -1640
rect 20816 -1704 20834 -1640
rect 20654 -1722 20834 -1704
rect 21474 -2088 21654 60
rect 21474 -2152 21492 -2088
rect 21556 -2152 21572 -2088
rect 21636 -2152 21654 -2088
rect 21474 -2168 21654 -2152
rect 21474 -2232 21492 -2168
rect 21556 -2232 21572 -2168
rect 21636 -2232 21654 -2168
rect 21474 -2250 21654 -2232
rect 7294 -2416 7312 -2352
rect 7376 -2416 7392 -2352
rect 7456 -2416 7474 -2352
rect 7294 -2432 7474 -2416
rect 7294 -2496 7312 -2432
rect 7376 -2496 7392 -2432
rect 7456 -2496 7474 -2432
rect -2762 -2680 -2744 -2616
rect -2680 -2680 -2664 -2616
rect -2600 -2680 -2582 -2616
rect -2762 -2696 -2582 -2680
rect -2762 -2760 -2744 -2696
rect -2680 -2760 -2664 -2696
rect -2600 -2760 -2582 -2696
rect -2762 -2778 -2582 -2760
rect 7294 -2778 7474 -2496
rect 22294 -2616 22474 60
rect 34014 -240 34194 60
rect 34014 -304 34032 -240
rect 34096 -304 34112 -240
rect 34176 -304 34194 -240
rect 34014 -320 34194 -304
rect 34014 -384 34032 -320
rect 34096 -384 34112 -320
rect 34176 -384 34194 -320
rect 34014 -666 34194 -384
rect 34834 -768 35014 60
rect 34834 -832 34852 -768
rect 34916 -832 34932 -768
rect 34996 -832 35014 -768
rect 34834 -848 35014 -832
rect 34834 -912 34852 -848
rect 34916 -912 34932 -848
rect 34996 -912 35014 -848
rect 34834 -1194 35014 -912
rect 35654 -1296 35834 60
rect 35654 -1360 35672 -1296
rect 35736 -1360 35752 -1296
rect 35816 -1360 35834 -1296
rect 35654 -1376 35834 -1360
rect 35654 -1440 35672 -1376
rect 35736 -1440 35752 -1376
rect 35816 -1440 35834 -1376
rect 35654 -1722 35834 -1440
rect 36474 -1824 36654 60
rect 36474 -1888 36492 -1824
rect 36556 -1888 36572 -1824
rect 36636 -1888 36654 -1824
rect 36474 -1904 36654 -1888
rect 36474 -1968 36492 -1904
rect 36556 -1968 36572 -1904
rect 36636 -1968 36654 -1904
rect 36474 -2250 36654 -1968
rect 22294 -2680 22312 -2616
rect 22376 -2680 22392 -2616
rect 22456 -2680 22474 -2616
rect 22294 -2696 22474 -2680
rect 22294 -2760 22312 -2696
rect 22376 -2760 22392 -2696
rect 22456 -2760 22474 -2696
rect 22294 -2778 22474 -2760
rect 37294 -2352 37474 60
rect 49014 -504 49194 60
rect 49014 -568 49032 -504
rect 49096 -568 49112 -504
rect 49176 -568 49194 -504
rect 49014 -584 49194 -568
rect 49014 -648 49032 -584
rect 49096 -648 49112 -584
rect 49176 -648 49194 -584
rect 49014 -666 49194 -648
rect 49834 -1032 50014 60
rect 49834 -1096 49852 -1032
rect 49916 -1096 49932 -1032
rect 49996 -1096 50014 -1032
rect 49834 -1112 50014 -1096
rect 49834 -1176 49852 -1112
rect 49916 -1176 49932 -1112
rect 49996 -1176 50014 -1112
rect 49834 -1194 50014 -1176
rect 50654 -1560 50834 60
rect 50654 -1624 50672 -1560
rect 50736 -1624 50752 -1560
rect 50816 -1624 50834 -1560
rect 50654 -1640 50834 -1624
rect 50654 -1704 50672 -1640
rect 50736 -1704 50752 -1640
rect 50816 -1704 50834 -1640
rect 50654 -1722 50834 -1704
rect 51474 -2088 51654 60
rect 51474 -2152 51492 -2088
rect 51556 -2152 51572 -2088
rect 51636 -2152 51654 -2088
rect 51474 -2168 51654 -2152
rect 51474 -2232 51492 -2168
rect 51556 -2232 51572 -2168
rect 51636 -2232 51654 -2168
rect 51474 -2250 51654 -2232
rect 37294 -2416 37312 -2352
rect 37376 -2416 37392 -2352
rect 37456 -2416 37474 -2352
rect 37294 -2432 37474 -2416
rect 37294 -2496 37312 -2432
rect 37376 -2496 37392 -2432
rect 37456 -2496 37474 -2432
rect 37294 -2778 37474 -2496
rect 52294 -2616 52474 60
rect 64014 -240 64194 60
rect 64014 -304 64032 -240
rect 64096 -304 64112 -240
rect 64176 -304 64194 -240
rect 64014 -320 64194 -304
rect 64014 -384 64032 -320
rect 64096 -384 64112 -320
rect 64176 -384 64194 -320
rect 64014 -666 64194 -384
rect 64834 -768 65014 60
rect 64834 -832 64852 -768
rect 64916 -832 64932 -768
rect 64996 -832 65014 -768
rect 64834 -848 65014 -832
rect 64834 -912 64852 -848
rect 64916 -912 64932 -848
rect 64996 -912 65014 -848
rect 64834 -1194 65014 -912
rect 65654 -1296 65834 60
rect 65654 -1360 65672 -1296
rect 65736 -1360 65752 -1296
rect 65816 -1360 65834 -1296
rect 65654 -1376 65834 -1360
rect 65654 -1440 65672 -1376
rect 65736 -1440 65752 -1376
rect 65816 -1440 65834 -1376
rect 65654 -1722 65834 -1440
rect 66474 -1824 66654 60
rect 66474 -1888 66492 -1824
rect 66556 -1888 66572 -1824
rect 66636 -1888 66654 -1824
rect 66474 -1904 66654 -1888
rect 66474 -1968 66492 -1904
rect 66556 -1968 66572 -1904
rect 66636 -1968 66654 -1904
rect 66474 -2250 66654 -1968
rect 52294 -2680 52312 -2616
rect 52376 -2680 52392 -2616
rect 52456 -2680 52474 -2616
rect 52294 -2696 52474 -2680
rect 52294 -2760 52312 -2696
rect 52376 -2760 52392 -2696
rect 52456 -2760 52474 -2696
rect 52294 -2778 52474 -2760
rect 67294 -2352 67474 60
rect 79014 -504 79194 60
rect 79014 -568 79032 -504
rect 79096 -568 79112 -504
rect 79176 -568 79194 -504
rect 79014 -584 79194 -568
rect 79014 -648 79032 -584
rect 79096 -648 79112 -584
rect 79176 -648 79194 -584
rect 79014 -666 79194 -648
rect 79834 -1032 80014 60
rect 79834 -1096 79852 -1032
rect 79916 -1096 79932 -1032
rect 79996 -1096 80014 -1032
rect 79834 -1112 80014 -1096
rect 79834 -1176 79852 -1112
rect 79916 -1176 79932 -1112
rect 79996 -1176 80014 -1112
rect 79834 -1194 80014 -1176
rect 80654 -1560 80834 60
rect 80654 -1624 80672 -1560
rect 80736 -1624 80752 -1560
rect 80816 -1624 80834 -1560
rect 80654 -1640 80834 -1624
rect 80654 -1704 80672 -1640
rect 80736 -1704 80752 -1640
rect 80816 -1704 80834 -1640
rect 80654 -1722 80834 -1704
rect 81474 -2088 81654 60
rect 81474 -2152 81492 -2088
rect 81556 -2152 81572 -2088
rect 81636 -2152 81654 -2088
rect 81474 -2168 81654 -2152
rect 81474 -2232 81492 -2168
rect 81556 -2232 81572 -2168
rect 81636 -2232 81654 -2168
rect 81474 -2250 81654 -2232
rect 67294 -2416 67312 -2352
rect 67376 -2416 67392 -2352
rect 67456 -2416 67474 -2352
rect 67294 -2432 67474 -2416
rect 67294 -2496 67312 -2432
rect 67376 -2496 67392 -2432
rect 67456 -2496 67474 -2432
rect 67294 -2778 67474 -2496
rect 82294 -2616 82474 60
rect 94014 -240 94194 60
rect 94014 -304 94032 -240
rect 94096 -304 94112 -240
rect 94176 -304 94194 -240
rect 94014 -320 94194 -304
rect 94014 -384 94032 -320
rect 94096 -384 94112 -320
rect 94176 -384 94194 -320
rect 94014 -666 94194 -384
rect 94834 -768 95014 60
rect 94834 -832 94852 -768
rect 94916 -832 94932 -768
rect 94996 -832 95014 -768
rect 94834 -848 95014 -832
rect 94834 -912 94852 -848
rect 94916 -912 94932 -848
rect 94996 -912 95014 -848
rect 94834 -1194 95014 -912
rect 95654 -1296 95834 60
rect 95654 -1360 95672 -1296
rect 95736 -1360 95752 -1296
rect 95816 -1360 95834 -1296
rect 95654 -1376 95834 -1360
rect 95654 -1440 95672 -1376
rect 95736 -1440 95752 -1376
rect 95816 -1440 95834 -1376
rect 95654 -1722 95834 -1440
rect 96474 -1824 96654 60
rect 96474 -1888 96492 -1824
rect 96556 -1888 96572 -1824
rect 96636 -1888 96654 -1824
rect 96474 -1904 96654 -1888
rect 96474 -1968 96492 -1904
rect 96556 -1968 96572 -1904
rect 96636 -1968 96654 -1904
rect 96474 -2250 96654 -1968
rect 82294 -2680 82312 -2616
rect 82376 -2680 82392 -2616
rect 82456 -2680 82474 -2616
rect 82294 -2696 82474 -2680
rect 82294 -2760 82312 -2696
rect 82376 -2760 82392 -2696
rect 82456 -2760 82474 -2696
rect 82294 -2778 82474 -2760
rect 97294 -2352 97474 60
rect 109014 -504 109194 60
rect 109014 -568 109032 -504
rect 109096 -568 109112 -504
rect 109176 -568 109194 -504
rect 109014 -584 109194 -568
rect 109014 -648 109032 -584
rect 109096 -648 109112 -584
rect 109176 -648 109194 -584
rect 109014 -666 109194 -648
rect 109834 -1032 110014 60
rect 109834 -1096 109852 -1032
rect 109916 -1096 109932 -1032
rect 109996 -1096 110014 -1032
rect 109834 -1112 110014 -1096
rect 109834 -1176 109852 -1112
rect 109916 -1176 109932 -1112
rect 109996 -1176 110014 -1112
rect 109834 -1194 110014 -1176
rect 110654 -1560 110834 60
rect 110654 -1624 110672 -1560
rect 110736 -1624 110752 -1560
rect 110816 -1624 110834 -1560
rect 110654 -1640 110834 -1624
rect 110654 -1704 110672 -1640
rect 110736 -1704 110752 -1640
rect 110816 -1704 110834 -1640
rect 110654 -1722 110834 -1704
rect 111474 -2088 111654 60
rect 111474 -2152 111492 -2088
rect 111556 -2152 111572 -2088
rect 111636 -2152 111654 -2088
rect 111474 -2168 111654 -2152
rect 111474 -2232 111492 -2168
rect 111556 -2232 111572 -2168
rect 111636 -2232 111654 -2168
rect 111474 -2250 111654 -2232
rect 97294 -2416 97312 -2352
rect 97376 -2416 97392 -2352
rect 97456 -2416 97474 -2352
rect 97294 -2432 97474 -2416
rect 97294 -2496 97312 -2432
rect 97376 -2496 97392 -2432
rect 97456 -2496 97474 -2432
rect 97294 -2778 97474 -2496
rect 112294 -2616 112474 60
rect 124014 -240 124194 60
rect 124014 -304 124032 -240
rect 124096 -304 124112 -240
rect 124176 -304 124194 -240
rect 124014 -320 124194 -304
rect 124014 -384 124032 -320
rect 124096 -384 124112 -320
rect 124176 -384 124194 -320
rect 124014 -666 124194 -384
rect 124834 -768 125014 60
rect 124834 -832 124852 -768
rect 124916 -832 124932 -768
rect 124996 -832 125014 -768
rect 124834 -848 125014 -832
rect 124834 -912 124852 -848
rect 124916 -912 124932 -848
rect 124996 -912 125014 -848
rect 124834 -1194 125014 -912
rect 125654 -1296 125834 60
rect 125654 -1360 125672 -1296
rect 125736 -1360 125752 -1296
rect 125816 -1360 125834 -1296
rect 125654 -1376 125834 -1360
rect 125654 -1440 125672 -1376
rect 125736 -1440 125752 -1376
rect 125816 -1440 125834 -1376
rect 125654 -1722 125834 -1440
rect 126474 -1824 126654 60
rect 126474 -1888 126492 -1824
rect 126556 -1888 126572 -1824
rect 126636 -1888 126654 -1824
rect 126474 -1904 126654 -1888
rect 126474 -1968 126492 -1904
rect 126556 -1968 126572 -1904
rect 126636 -1968 126654 -1904
rect 126474 -2250 126654 -1968
rect 112294 -2680 112312 -2616
rect 112376 -2680 112392 -2616
rect 112456 -2680 112474 -2616
rect 112294 -2696 112474 -2680
rect 112294 -2760 112312 -2696
rect 112376 -2760 112392 -2696
rect 112456 -2760 112474 -2696
rect 112294 -2778 112474 -2760
rect 127294 -2352 127474 60
rect 139014 -504 139194 60
rect 139014 -568 139032 -504
rect 139096 -568 139112 -504
rect 139176 -568 139194 -504
rect 139014 -584 139194 -568
rect 139014 -648 139032 -584
rect 139096 -648 139112 -584
rect 139176 -648 139194 -584
rect 139014 -666 139194 -648
rect 139834 -1032 140014 60
rect 139834 -1096 139852 -1032
rect 139916 -1096 139932 -1032
rect 139996 -1096 140014 -1032
rect 139834 -1112 140014 -1096
rect 139834 -1176 139852 -1112
rect 139916 -1176 139932 -1112
rect 139996 -1176 140014 -1112
rect 139834 -1194 140014 -1176
rect 140654 -1560 140834 60
rect 140654 -1624 140672 -1560
rect 140736 -1624 140752 -1560
rect 140816 -1624 140834 -1560
rect 140654 -1640 140834 -1624
rect 140654 -1704 140672 -1640
rect 140736 -1704 140752 -1640
rect 140816 -1704 140834 -1640
rect 140654 -1722 140834 -1704
rect 141474 -2088 141654 60
rect 141474 -2152 141492 -2088
rect 141556 -2152 141572 -2088
rect 141636 -2152 141654 -2088
rect 141474 -2168 141654 -2152
rect 141474 -2232 141492 -2168
rect 141556 -2232 141572 -2168
rect 141636 -2232 141654 -2168
rect 141474 -2250 141654 -2232
rect 127294 -2416 127312 -2352
rect 127376 -2416 127392 -2352
rect 127456 -2416 127474 -2352
rect 127294 -2432 127474 -2416
rect 127294 -2496 127312 -2432
rect 127376 -2496 127392 -2432
rect 127456 -2496 127474 -2432
rect 127294 -2778 127474 -2496
rect 142294 -2616 142474 60
rect 154014 -240 154194 60
rect 154014 -304 154032 -240
rect 154096 -304 154112 -240
rect 154176 -304 154194 -240
rect 154014 -320 154194 -304
rect 154014 -384 154032 -320
rect 154096 -384 154112 -320
rect 154176 -384 154194 -320
rect 154014 -666 154194 -384
rect 154834 -768 155014 60
rect 154834 -832 154852 -768
rect 154916 -832 154932 -768
rect 154996 -832 155014 -768
rect 154834 -848 155014 -832
rect 154834 -912 154852 -848
rect 154916 -912 154932 -848
rect 154996 -912 155014 -848
rect 154834 -1194 155014 -912
rect 155654 -1296 155834 60
rect 155654 -1360 155672 -1296
rect 155736 -1360 155752 -1296
rect 155816 -1360 155834 -1296
rect 155654 -1376 155834 -1360
rect 155654 -1440 155672 -1376
rect 155736 -1440 155752 -1376
rect 155816 -1440 155834 -1376
rect 155654 -1722 155834 -1440
rect 156474 -1824 156654 60
rect 156474 -1888 156492 -1824
rect 156556 -1888 156572 -1824
rect 156636 -1888 156654 -1824
rect 156474 -1904 156654 -1888
rect 156474 -1968 156492 -1904
rect 156556 -1968 156572 -1904
rect 156636 -1968 156654 -1904
rect 156474 -2250 156654 -1968
rect 142294 -2680 142312 -2616
rect 142376 -2680 142392 -2616
rect 142456 -2680 142474 -2616
rect 142294 -2696 142474 -2680
rect 142294 -2760 142312 -2696
rect 142376 -2760 142392 -2696
rect 142456 -2760 142474 -2696
rect 142294 -2778 142474 -2760
rect 157294 -2352 157474 60
rect 169014 -504 169194 60
rect 169014 -568 169032 -504
rect 169096 -568 169112 -504
rect 169176 -568 169194 -504
rect 169014 -584 169194 -568
rect 169014 -648 169032 -584
rect 169096 -648 169112 -584
rect 169176 -648 169194 -584
rect 169014 -666 169194 -648
rect 169834 -1032 170014 60
rect 169834 -1096 169852 -1032
rect 169916 -1096 169932 -1032
rect 169996 -1096 170014 -1032
rect 169834 -1112 170014 -1096
rect 169834 -1176 169852 -1112
rect 169916 -1176 169932 -1112
rect 169996 -1176 170014 -1112
rect 169834 -1194 170014 -1176
rect 170654 -1560 170834 60
rect 170654 -1624 170672 -1560
rect 170736 -1624 170752 -1560
rect 170816 -1624 170834 -1560
rect 170654 -1640 170834 -1624
rect 170654 -1704 170672 -1640
rect 170736 -1704 170752 -1640
rect 170816 -1704 170834 -1640
rect 170654 -1722 170834 -1704
rect 171474 -2088 171654 60
rect 171474 -2152 171492 -2088
rect 171556 -2152 171572 -2088
rect 171636 -2152 171654 -2088
rect 171474 -2168 171654 -2152
rect 171474 -2232 171492 -2168
rect 171556 -2232 171572 -2168
rect 171636 -2232 171654 -2168
rect 171474 -2250 171654 -2232
rect 157294 -2416 157312 -2352
rect 157376 -2416 157392 -2352
rect 157456 -2416 157474 -2352
rect 157294 -2432 157474 -2416
rect 157294 -2496 157312 -2432
rect 157376 -2496 157392 -2432
rect 157456 -2496 157474 -2432
rect 157294 -2778 157474 -2496
rect 172294 -2616 172474 60
rect 184014 -240 184194 60
rect 184014 -304 184032 -240
rect 184096 -304 184112 -240
rect 184176 -304 184194 -240
rect 184014 -320 184194 -304
rect 184014 -384 184032 -320
rect 184096 -384 184112 -320
rect 184176 -384 184194 -320
rect 184014 -666 184194 -384
rect 184834 -768 185014 60
rect 184834 -832 184852 -768
rect 184916 -832 184932 -768
rect 184996 -832 185014 -768
rect 184834 -848 185014 -832
rect 184834 -912 184852 -848
rect 184916 -912 184932 -848
rect 184996 -912 185014 -848
rect 184834 -1194 185014 -912
rect 185654 -1296 185834 60
rect 185654 -1360 185672 -1296
rect 185736 -1360 185752 -1296
rect 185816 -1360 185834 -1296
rect 185654 -1376 185834 -1360
rect 185654 -1440 185672 -1376
rect 185736 -1440 185752 -1376
rect 185816 -1440 185834 -1376
rect 185654 -1722 185834 -1440
rect 186474 -1824 186654 60
rect 186474 -1888 186492 -1824
rect 186556 -1888 186572 -1824
rect 186636 -1888 186654 -1824
rect 186474 -1904 186654 -1888
rect 186474 -1968 186492 -1904
rect 186556 -1968 186572 -1904
rect 186636 -1968 186654 -1904
rect 186474 -2250 186654 -1968
rect 172294 -2680 172312 -2616
rect 172376 -2680 172392 -2616
rect 172456 -2680 172474 -2616
rect 172294 -2696 172474 -2680
rect 172294 -2760 172312 -2696
rect 172376 -2760 172392 -2696
rect 172456 -2760 172474 -2696
rect 172294 -2778 172474 -2760
rect 187294 -2352 187474 60
rect 200122 -240 200302 18192
rect 200122 -304 200140 -240
rect 200204 -304 200220 -240
rect 200284 -304 200302 -240
rect 200122 -320 200302 -304
rect 200122 -384 200140 -320
rect 200204 -384 200220 -320
rect 200284 -384 200302 -320
rect 200122 -402 200302 -384
rect 200386 -504 200566 18456
rect 200386 -568 200404 -504
rect 200468 -568 200484 -504
rect 200548 -568 200566 -504
rect 200386 -584 200566 -568
rect 200386 -648 200404 -584
rect 200468 -648 200484 -584
rect 200548 -648 200566 -584
rect 200386 -666 200566 -648
rect 200650 -768 200830 18720
rect 200650 -832 200668 -768
rect 200732 -832 200748 -768
rect 200812 -832 200830 -768
rect 200650 -848 200830 -832
rect 200650 -912 200668 -848
rect 200732 -912 200748 -848
rect 200812 -912 200830 -848
rect 200650 -930 200830 -912
rect 200914 -1032 201094 18984
rect 200914 -1096 200932 -1032
rect 200996 -1096 201012 -1032
rect 201076 -1096 201094 -1032
rect 200914 -1112 201094 -1096
rect 200914 -1176 200932 -1112
rect 200996 -1176 201012 -1112
rect 201076 -1176 201094 -1112
rect 200914 -1194 201094 -1176
rect 201178 -1296 201358 19248
rect 201178 -1360 201196 -1296
rect 201260 -1360 201276 -1296
rect 201340 -1360 201358 -1296
rect 201178 -1376 201358 -1360
rect 201178 -1440 201196 -1376
rect 201260 -1440 201276 -1376
rect 201340 -1440 201358 -1376
rect 201178 -1458 201358 -1440
rect 201442 -1560 201622 19512
rect 201442 -1624 201460 -1560
rect 201524 -1624 201540 -1560
rect 201604 -1624 201622 -1560
rect 201442 -1640 201622 -1624
rect 201442 -1704 201460 -1640
rect 201524 -1704 201540 -1640
rect 201604 -1704 201622 -1640
rect 201442 -1722 201622 -1704
rect 201706 -1824 201886 19776
rect 201706 -1888 201724 -1824
rect 201788 -1888 201804 -1824
rect 201868 -1888 201886 -1824
rect 201706 -1904 201886 -1888
rect 201706 -1968 201724 -1904
rect 201788 -1968 201804 -1904
rect 201868 -1968 201886 -1904
rect 201706 -1986 201886 -1968
rect 201970 -2088 202150 20040
rect 201970 -2152 201988 -2088
rect 202052 -2152 202068 -2088
rect 202132 -2152 202150 -2088
rect 201970 -2168 202150 -2152
rect 201970 -2232 201988 -2168
rect 202052 -2232 202068 -2168
rect 202132 -2232 202150 -2168
rect 201970 -2250 202150 -2232
rect 187294 -2416 187312 -2352
rect 187376 -2416 187392 -2352
rect 187456 -2416 187474 -2352
rect 187294 -2432 187474 -2416
rect 187294 -2496 187312 -2432
rect 187376 -2496 187392 -2432
rect 187456 -2496 187474 -2432
rect 187294 -2778 187474 -2496
rect 202234 -2352 202414 20304
rect 202234 -2416 202252 -2352
rect 202316 -2416 202332 -2352
rect 202396 -2416 202414 -2352
rect 202234 -2432 202414 -2416
rect 202234 -2496 202252 -2432
rect 202316 -2496 202332 -2432
rect 202396 -2496 202414 -2432
rect 202234 -2514 202414 -2496
rect 202498 -2616 202678 20568
rect 202498 -2680 202516 -2616
rect 202580 -2680 202596 -2616
rect 202660 -2680 202678 -2616
rect 202498 -2696 202678 -2680
rect 202498 -2760 202516 -2696
rect 202580 -2760 202596 -2696
rect 202660 -2760 202678 -2696
rect 202498 -2778 202678 -2760
<< obsm4 >>
rect 4014 60 193141 17940
<< labels >>
rlabel metal3 s -400 3000 60 3120 4 caravel_clk
port 1 nsew signal input
rlabel metal3 s -400 8984 60 9104 4 caravel_clk2
port 2 nsew signal input
rlabel metal3 s -400 14968 60 15088 4 caravel_rstn
port 3 nsew signal input
rlabel metal2 s 1858 17940 1914 18400 6 la_data_in_core[0]
port 4 nsew signal output
rlabel metal2 s 45466 17940 45522 18400 6 la_data_in_core[100]
port 5 nsew signal output
rlabel metal2 s 45926 17940 45982 18400 6 la_data_in_core[101]
port 6 nsew signal output
rlabel metal2 s 46386 17940 46442 18400 6 la_data_in_core[102]
port 7 nsew signal output
rlabel metal2 s 46754 17940 46810 18400 6 la_data_in_core[103]
port 8 nsew signal output
rlabel metal2 s 47214 17940 47270 18400 6 la_data_in_core[104]
port 9 nsew signal output
rlabel metal2 s 47674 17940 47730 18400 6 la_data_in_core[105]
port 10 nsew signal output
rlabel metal2 s 48134 17940 48190 18400 6 la_data_in_core[106]
port 11 nsew signal output
rlabel metal2 s 48502 17940 48558 18400 6 la_data_in_core[107]
port 12 nsew signal output
rlabel metal2 s 48962 17940 49018 18400 6 la_data_in_core[108]
port 13 nsew signal output
rlabel metal2 s 49422 17940 49478 18400 6 la_data_in_core[109]
port 14 nsew signal output
rlabel metal2 s 6274 17940 6330 18400 6 la_data_in_core[10]
port 15 nsew signal output
rlabel metal2 s 49790 17940 49846 18400 6 la_data_in_core[110]
port 16 nsew signal output
rlabel metal2 s 50250 17940 50306 18400 6 la_data_in_core[111]
port 17 nsew signal output
rlabel metal2 s 50710 17940 50766 18400 6 la_data_in_core[112]
port 18 nsew signal output
rlabel metal2 s 51170 17940 51226 18400 6 la_data_in_core[113]
port 19 nsew signal output
rlabel metal2 s 51538 17940 51594 18400 6 la_data_in_core[114]
port 20 nsew signal output
rlabel metal2 s 51998 17940 52054 18400 6 la_data_in_core[115]
port 21 nsew signal output
rlabel metal2 s 52458 17940 52514 18400 6 la_data_in_core[116]
port 22 nsew signal output
rlabel metal2 s 52918 17940 52974 18400 6 la_data_in_core[117]
port 23 nsew signal output
rlabel metal2 s 53286 17940 53342 18400 6 la_data_in_core[118]
port 24 nsew signal output
rlabel metal2 s 53746 17940 53802 18400 6 la_data_in_core[119]
port 25 nsew signal output
rlabel metal2 s 6734 17940 6790 18400 6 la_data_in_core[11]
port 26 nsew signal output
rlabel metal2 s 54206 17940 54262 18400 6 la_data_in_core[120]
port 27 nsew signal output
rlabel metal2 s 54666 17940 54722 18400 6 la_data_in_core[121]
port 28 nsew signal output
rlabel metal2 s 55034 17940 55090 18400 6 la_data_in_core[122]
port 29 nsew signal output
rlabel metal2 s 55494 17940 55550 18400 6 la_data_in_core[123]
port 30 nsew signal output
rlabel metal2 s 55954 17940 56010 18400 6 la_data_in_core[124]
port 31 nsew signal output
rlabel metal2 s 56322 17940 56378 18400 6 la_data_in_core[125]
port 32 nsew signal output
rlabel metal2 s 56782 17940 56838 18400 6 la_data_in_core[126]
port 33 nsew signal output
rlabel metal2 s 57242 17940 57298 18400 6 la_data_in_core[127]
port 34 nsew signal output
rlabel metal2 s 7102 17940 7158 18400 6 la_data_in_core[12]
port 35 nsew signal output
rlabel metal2 s 7562 17940 7618 18400 6 la_data_in_core[13]
port 36 nsew signal output
rlabel metal2 s 8022 17940 8078 18400 6 la_data_in_core[14]
port 37 nsew signal output
rlabel metal2 s 8390 17940 8446 18400 6 la_data_in_core[15]
port 38 nsew signal output
rlabel metal2 s 8850 17940 8906 18400 6 la_data_in_core[16]
port 39 nsew signal output
rlabel metal2 s 9310 17940 9366 18400 6 la_data_in_core[17]
port 40 nsew signal output
rlabel metal2 s 9770 17940 9826 18400 6 la_data_in_core[18]
port 41 nsew signal output
rlabel metal2 s 10138 17940 10194 18400 6 la_data_in_core[19]
port 42 nsew signal output
rlabel metal2 s 2318 17940 2374 18400 6 la_data_in_core[1]
port 43 nsew signal output
rlabel metal2 s 10598 17940 10654 18400 6 la_data_in_core[20]
port 44 nsew signal output
rlabel metal2 s 11058 17940 11114 18400 6 la_data_in_core[21]
port 45 nsew signal output
rlabel metal2 s 11518 17940 11574 18400 6 la_data_in_core[22]
port 46 nsew signal output
rlabel metal2 s 11886 17940 11942 18400 6 la_data_in_core[23]
port 47 nsew signal output
rlabel metal2 s 12346 17940 12402 18400 6 la_data_in_core[24]
port 48 nsew signal output
rlabel metal2 s 12806 17940 12862 18400 6 la_data_in_core[25]
port 49 nsew signal output
rlabel metal2 s 13266 17940 13322 18400 6 la_data_in_core[26]
port 50 nsew signal output
rlabel metal2 s 13634 17940 13690 18400 6 la_data_in_core[27]
port 51 nsew signal output
rlabel metal2 s 14094 17940 14150 18400 6 la_data_in_core[28]
port 52 nsew signal output
rlabel metal2 s 14554 17940 14610 18400 6 la_data_in_core[29]
port 53 nsew signal output
rlabel metal2 s 2778 17940 2834 18400 6 la_data_in_core[2]
port 54 nsew signal output
rlabel metal2 s 15014 17940 15070 18400 6 la_data_in_core[30]
port 55 nsew signal output
rlabel metal2 s 15382 17940 15438 18400 6 la_data_in_core[31]
port 56 nsew signal output
rlabel metal2 s 15842 17940 15898 18400 6 la_data_in_core[32]
port 57 nsew signal output
rlabel metal2 s 16302 17940 16358 18400 6 la_data_in_core[33]
port 58 nsew signal output
rlabel metal2 s 16670 17940 16726 18400 6 la_data_in_core[34]
port 59 nsew signal output
rlabel metal2 s 17130 17940 17186 18400 6 la_data_in_core[35]
port 60 nsew signal output
rlabel metal2 s 17590 17940 17646 18400 6 la_data_in_core[36]
port 61 nsew signal output
rlabel metal2 s 18050 17940 18106 18400 6 la_data_in_core[37]
port 62 nsew signal output
rlabel metal2 s 18418 17940 18474 18400 6 la_data_in_core[38]
port 63 nsew signal output
rlabel metal2 s 18878 17940 18934 18400 6 la_data_in_core[39]
port 64 nsew signal output
rlabel metal2 s 3238 17940 3294 18400 6 la_data_in_core[3]
port 65 nsew signal output
rlabel metal2 s 19338 17940 19394 18400 6 la_data_in_core[40]
port 66 nsew signal output
rlabel metal2 s 19798 17940 19854 18400 6 la_data_in_core[41]
port 67 nsew signal output
rlabel metal2 s 20166 17940 20222 18400 6 la_data_in_core[42]
port 68 nsew signal output
rlabel metal2 s 20626 17940 20682 18400 6 la_data_in_core[43]
port 69 nsew signal output
rlabel metal2 s 21086 17940 21142 18400 6 la_data_in_core[44]
port 70 nsew signal output
rlabel metal2 s 21546 17940 21602 18400 6 la_data_in_core[45]
port 71 nsew signal output
rlabel metal2 s 21914 17940 21970 18400 6 la_data_in_core[46]
port 72 nsew signal output
rlabel metal2 s 22374 17940 22430 18400 6 la_data_in_core[47]
port 73 nsew signal output
rlabel metal2 s 22834 17940 22890 18400 6 la_data_in_core[48]
port 74 nsew signal output
rlabel metal2 s 23294 17940 23350 18400 6 la_data_in_core[49]
port 75 nsew signal output
rlabel metal2 s 3606 17940 3662 18400 6 la_data_in_core[4]
port 76 nsew signal output
rlabel metal2 s 23662 17940 23718 18400 6 la_data_in_core[50]
port 77 nsew signal output
rlabel metal2 s 24122 17940 24178 18400 6 la_data_in_core[51]
port 78 nsew signal output
rlabel metal2 s 24582 17940 24638 18400 6 la_data_in_core[52]
port 79 nsew signal output
rlabel metal2 s 24950 17940 25006 18400 6 la_data_in_core[53]
port 80 nsew signal output
rlabel metal2 s 25410 17940 25466 18400 6 la_data_in_core[54]
port 81 nsew signal output
rlabel metal2 s 25870 17940 25926 18400 6 la_data_in_core[55]
port 82 nsew signal output
rlabel metal2 s 26330 17940 26386 18400 6 la_data_in_core[56]
port 83 nsew signal output
rlabel metal2 s 26698 17940 26754 18400 6 la_data_in_core[57]
port 84 nsew signal output
rlabel metal2 s 27158 17940 27214 18400 6 la_data_in_core[58]
port 85 nsew signal output
rlabel metal2 s 27618 17940 27674 18400 6 la_data_in_core[59]
port 86 nsew signal output
rlabel metal2 s 4066 17940 4122 18400 6 la_data_in_core[5]
port 87 nsew signal output
rlabel metal2 s 28078 17940 28134 18400 6 la_data_in_core[60]
port 88 nsew signal output
rlabel metal2 s 28446 17940 28502 18400 6 la_data_in_core[61]
port 89 nsew signal output
rlabel metal2 s 28906 17940 28962 18400 6 la_data_in_core[62]
port 90 nsew signal output
rlabel metal2 s 29366 17940 29422 18400 6 la_data_in_core[63]
port 91 nsew signal output
rlabel metal2 s 29826 17940 29882 18400 6 la_data_in_core[64]
port 92 nsew signal output
rlabel metal2 s 30194 17940 30250 18400 6 la_data_in_core[65]
port 93 nsew signal output
rlabel metal2 s 30654 17940 30710 18400 6 la_data_in_core[66]
port 94 nsew signal output
rlabel metal2 s 31114 17940 31170 18400 6 la_data_in_core[67]
port 95 nsew signal output
rlabel metal2 s 31574 17940 31630 18400 6 la_data_in_core[68]
port 96 nsew signal output
rlabel metal2 s 31942 17940 31998 18400 6 la_data_in_core[69]
port 97 nsew signal output
rlabel metal2 s 4526 17940 4582 18400 6 la_data_in_core[6]
port 98 nsew signal output
rlabel metal2 s 32402 17940 32458 18400 6 la_data_in_core[70]
port 99 nsew signal output
rlabel metal2 s 32862 17940 32918 18400 6 la_data_in_core[71]
port 100 nsew signal output
rlabel metal2 s 33230 17940 33286 18400 6 la_data_in_core[72]
port 101 nsew signal output
rlabel metal2 s 33690 17940 33746 18400 6 la_data_in_core[73]
port 102 nsew signal output
rlabel metal2 s 34150 17940 34206 18400 6 la_data_in_core[74]
port 103 nsew signal output
rlabel metal2 s 34610 17940 34666 18400 6 la_data_in_core[75]
port 104 nsew signal output
rlabel metal2 s 34978 17940 35034 18400 6 la_data_in_core[76]
port 105 nsew signal output
rlabel metal2 s 35438 17940 35494 18400 6 la_data_in_core[77]
port 106 nsew signal output
rlabel metal2 s 35898 17940 35954 18400 6 la_data_in_core[78]
port 107 nsew signal output
rlabel metal2 s 36358 17940 36414 18400 6 la_data_in_core[79]
port 108 nsew signal output
rlabel metal2 s 4986 17940 5042 18400 6 la_data_in_core[7]
port 109 nsew signal output
rlabel metal2 s 36726 17940 36782 18400 6 la_data_in_core[80]
port 110 nsew signal output
rlabel metal2 s 37186 17940 37242 18400 6 la_data_in_core[81]
port 111 nsew signal output
rlabel metal2 s 37646 17940 37702 18400 6 la_data_in_core[82]
port 112 nsew signal output
rlabel metal2 s 38106 17940 38162 18400 6 la_data_in_core[83]
port 113 nsew signal output
rlabel metal2 s 38474 17940 38530 18400 6 la_data_in_core[84]
port 114 nsew signal output
rlabel metal2 s 38934 17940 38990 18400 6 la_data_in_core[85]
port 115 nsew signal output
rlabel metal2 s 39394 17940 39450 18400 6 la_data_in_core[86]
port 116 nsew signal output
rlabel metal2 s 39854 17940 39910 18400 6 la_data_in_core[87]
port 117 nsew signal output
rlabel metal2 s 40222 17940 40278 18400 6 la_data_in_core[88]
port 118 nsew signal output
rlabel metal2 s 40682 17940 40738 18400 6 la_data_in_core[89]
port 119 nsew signal output
rlabel metal2 s 5354 17940 5410 18400 6 la_data_in_core[8]
port 120 nsew signal output
rlabel metal2 s 41142 17940 41198 18400 6 la_data_in_core[90]
port 121 nsew signal output
rlabel metal2 s 41510 17940 41566 18400 6 la_data_in_core[91]
port 122 nsew signal output
rlabel metal2 s 41970 17940 42026 18400 6 la_data_in_core[92]
port 123 nsew signal output
rlabel metal2 s 42430 17940 42486 18400 6 la_data_in_core[93]
port 124 nsew signal output
rlabel metal2 s 42890 17940 42946 18400 6 la_data_in_core[94]
port 125 nsew signal output
rlabel metal2 s 43258 17940 43314 18400 6 la_data_in_core[95]
port 126 nsew signal output
rlabel metal2 s 43718 17940 43774 18400 6 la_data_in_core[96]
port 127 nsew signal output
rlabel metal2 s 44178 17940 44234 18400 6 la_data_in_core[97]
port 128 nsew signal output
rlabel metal2 s 44638 17940 44694 18400 6 la_data_in_core[98]
port 129 nsew signal output
rlabel metal2 s 45006 17940 45062 18400 6 la_data_in_core[99]
port 130 nsew signal output
rlabel metal2 s 5814 17940 5870 18400 6 la_data_in_core[9]
port 131 nsew signal output
rlabel metal2 s 55954 -400 56010 60 8 la_data_in_mprj[0]
port 132 nsew signal output
rlabel metal2 s 99470 -400 99526 60 8 la_data_in_mprj[100]
port 133 nsew signal output
rlabel metal2 s 99930 -400 99986 60 8 la_data_in_mprj[101]
port 134 nsew signal output
rlabel metal2 s 100390 -400 100446 60 8 la_data_in_mprj[102]
port 135 nsew signal output
rlabel metal2 s 100850 -400 100906 60 8 la_data_in_mprj[103]
port 136 nsew signal output
rlabel metal2 s 101218 -400 101274 60 8 la_data_in_mprj[104]
port 137 nsew signal output
rlabel metal2 s 101678 -400 101734 60 8 la_data_in_mprj[105]
port 138 nsew signal output
rlabel metal2 s 102138 -400 102194 60 8 la_data_in_mprj[106]
port 139 nsew signal output
rlabel metal2 s 102598 -400 102654 60 8 la_data_in_mprj[107]
port 140 nsew signal output
rlabel metal2 s 102966 -400 103022 60 8 la_data_in_mprj[108]
port 141 nsew signal output
rlabel metal2 s 103426 -400 103482 60 8 la_data_in_mprj[109]
port 142 nsew signal output
rlabel metal2 s 60278 -400 60334 60 8 la_data_in_mprj[10]
port 143 nsew signal output
rlabel metal2 s 103886 -400 103942 60 8 la_data_in_mprj[110]
port 144 nsew signal output
rlabel metal2 s 104254 -400 104310 60 8 la_data_in_mprj[111]
port 145 nsew signal output
rlabel metal2 s 104714 -400 104770 60 8 la_data_in_mprj[112]
port 146 nsew signal output
rlabel metal2 s 105174 -400 105230 60 8 la_data_in_mprj[113]
port 147 nsew signal output
rlabel metal2 s 105634 -400 105690 60 8 la_data_in_mprj[114]
port 148 nsew signal output
rlabel metal2 s 106002 -400 106058 60 8 la_data_in_mprj[115]
port 149 nsew signal output
rlabel metal2 s 106462 -400 106518 60 8 la_data_in_mprj[116]
port 150 nsew signal output
rlabel metal2 s 106922 -400 106978 60 8 la_data_in_mprj[117]
port 151 nsew signal output
rlabel metal2 s 107382 -400 107438 60 8 la_data_in_mprj[118]
port 152 nsew signal output
rlabel metal2 s 107750 -400 107806 60 8 la_data_in_mprj[119]
port 153 nsew signal output
rlabel metal2 s 60738 -400 60794 60 8 la_data_in_mprj[11]
port 154 nsew signal output
rlabel metal2 s 108210 -400 108266 60 8 la_data_in_mprj[120]
port 155 nsew signal output
rlabel metal2 s 108670 -400 108726 60 8 la_data_in_mprj[121]
port 156 nsew signal output
rlabel metal2 s 109130 -400 109186 60 8 la_data_in_mprj[122]
port 157 nsew signal output
rlabel metal2 s 109498 -400 109554 60 8 la_data_in_mprj[123]
port 158 nsew signal output
rlabel metal2 s 109958 -400 110014 60 8 la_data_in_mprj[124]
port 159 nsew signal output
rlabel metal2 s 110418 -400 110474 60 8 la_data_in_mprj[125]
port 160 nsew signal output
rlabel metal2 s 110878 -400 110934 60 8 la_data_in_mprj[126]
port 161 nsew signal output
rlabel metal2 s 111246 -400 111302 60 8 la_data_in_mprj[127]
port 162 nsew signal output
rlabel metal2 s 61198 -400 61254 60 8 la_data_in_mprj[12]
port 163 nsew signal output
rlabel metal2 s 61566 -400 61622 60 8 la_data_in_mprj[13]
port 164 nsew signal output
rlabel metal2 s 62026 -400 62082 60 8 la_data_in_mprj[14]
port 165 nsew signal output
rlabel metal2 s 62486 -400 62542 60 8 la_data_in_mprj[15]
port 166 nsew signal output
rlabel metal2 s 62946 -400 63002 60 8 la_data_in_mprj[16]
port 167 nsew signal output
rlabel metal2 s 63314 -400 63370 60 8 la_data_in_mprj[17]
port 168 nsew signal output
rlabel metal2 s 63774 -400 63830 60 8 la_data_in_mprj[18]
port 169 nsew signal output
rlabel metal2 s 64234 -400 64290 60 8 la_data_in_mprj[19]
port 170 nsew signal output
rlabel metal2 s 56322 -400 56378 60 8 la_data_in_mprj[1]
port 171 nsew signal output
rlabel metal2 s 64602 -400 64658 60 8 la_data_in_mprj[20]
port 172 nsew signal output
rlabel metal2 s 65062 -400 65118 60 8 la_data_in_mprj[21]
port 173 nsew signal output
rlabel metal2 s 65522 -400 65578 60 8 la_data_in_mprj[22]
port 174 nsew signal output
rlabel metal2 s 65982 -400 66038 60 8 la_data_in_mprj[23]
port 175 nsew signal output
rlabel metal2 s 66350 -400 66406 60 8 la_data_in_mprj[24]
port 176 nsew signal output
rlabel metal2 s 66810 -400 66866 60 8 la_data_in_mprj[25]
port 177 nsew signal output
rlabel metal2 s 67270 -400 67326 60 8 la_data_in_mprj[26]
port 178 nsew signal output
rlabel metal2 s 67730 -400 67786 60 8 la_data_in_mprj[27]
port 179 nsew signal output
rlabel metal2 s 68098 -400 68154 60 8 la_data_in_mprj[28]
port 180 nsew signal output
rlabel metal2 s 68558 -400 68614 60 8 la_data_in_mprj[29]
port 181 nsew signal output
rlabel metal2 s 56782 -400 56838 60 8 la_data_in_mprj[2]
port 182 nsew signal output
rlabel metal2 s 69018 -400 69074 60 8 la_data_in_mprj[30]
port 183 nsew signal output
rlabel metal2 s 69478 -400 69534 60 8 la_data_in_mprj[31]
port 184 nsew signal output
rlabel metal2 s 69846 -400 69902 60 8 la_data_in_mprj[32]
port 185 nsew signal output
rlabel metal2 s 70306 -400 70362 60 8 la_data_in_mprj[33]
port 186 nsew signal output
rlabel metal2 s 70766 -400 70822 60 8 la_data_in_mprj[34]
port 187 nsew signal output
rlabel metal2 s 71226 -400 71282 60 8 la_data_in_mprj[35]
port 188 nsew signal output
rlabel metal2 s 71594 -400 71650 60 8 la_data_in_mprj[36]
port 189 nsew signal output
rlabel metal2 s 72054 -400 72110 60 8 la_data_in_mprj[37]
port 190 nsew signal output
rlabel metal2 s 72514 -400 72570 60 8 la_data_in_mprj[38]
port 191 nsew signal output
rlabel metal2 s 72882 -400 72938 60 8 la_data_in_mprj[39]
port 192 nsew signal output
rlabel metal2 s 57242 -400 57298 60 8 la_data_in_mprj[3]
port 193 nsew signal output
rlabel metal2 s 73342 -400 73398 60 8 la_data_in_mprj[40]
port 194 nsew signal output
rlabel metal2 s 73802 -400 73858 60 8 la_data_in_mprj[41]
port 195 nsew signal output
rlabel metal2 s 74262 -400 74318 60 8 la_data_in_mprj[42]
port 196 nsew signal output
rlabel metal2 s 74630 -400 74686 60 8 la_data_in_mprj[43]
port 197 nsew signal output
rlabel metal2 s 75090 -400 75146 60 8 la_data_in_mprj[44]
port 198 nsew signal output
rlabel metal2 s 75550 -400 75606 60 8 la_data_in_mprj[45]
port 199 nsew signal output
rlabel metal2 s 76010 -400 76066 60 8 la_data_in_mprj[46]
port 200 nsew signal output
rlabel metal2 s 76378 -400 76434 60 8 la_data_in_mprj[47]
port 201 nsew signal output
rlabel metal2 s 76838 -400 76894 60 8 la_data_in_mprj[48]
port 202 nsew signal output
rlabel metal2 s 77298 -400 77354 60 8 la_data_in_mprj[49]
port 203 nsew signal output
rlabel metal2 s 57702 -400 57758 60 8 la_data_in_mprj[4]
port 204 nsew signal output
rlabel metal2 s 77758 -400 77814 60 8 la_data_in_mprj[50]
port 205 nsew signal output
rlabel metal2 s 78126 -400 78182 60 8 la_data_in_mprj[51]
port 206 nsew signal output
rlabel metal2 s 78586 -400 78642 60 8 la_data_in_mprj[52]
port 207 nsew signal output
rlabel metal2 s 79046 -400 79102 60 8 la_data_in_mprj[53]
port 208 nsew signal output
rlabel metal2 s 79506 -400 79562 60 8 la_data_in_mprj[54]
port 209 nsew signal output
rlabel metal2 s 79874 -400 79930 60 8 la_data_in_mprj[55]
port 210 nsew signal output
rlabel metal2 s 80334 -400 80390 60 8 la_data_in_mprj[56]
port 211 nsew signal output
rlabel metal2 s 80794 -400 80850 60 8 la_data_in_mprj[57]
port 212 nsew signal output
rlabel metal2 s 81162 -400 81218 60 8 la_data_in_mprj[58]
port 213 nsew signal output
rlabel metal2 s 81622 -400 81678 60 8 la_data_in_mprj[59]
port 214 nsew signal output
rlabel metal2 s 58070 -400 58126 60 8 la_data_in_mprj[5]
port 215 nsew signal output
rlabel metal2 s 82082 -400 82138 60 8 la_data_in_mprj[60]
port 216 nsew signal output
rlabel metal2 s 82542 -400 82598 60 8 la_data_in_mprj[61]
port 217 nsew signal output
rlabel metal2 s 82910 -400 82966 60 8 la_data_in_mprj[62]
port 218 nsew signal output
rlabel metal2 s 83370 -400 83426 60 8 la_data_in_mprj[63]
port 219 nsew signal output
rlabel metal2 s 83830 -400 83886 60 8 la_data_in_mprj[64]
port 220 nsew signal output
rlabel metal2 s 84290 -400 84346 60 8 la_data_in_mprj[65]
port 221 nsew signal output
rlabel metal2 s 84658 -400 84714 60 8 la_data_in_mprj[66]
port 222 nsew signal output
rlabel metal2 s 85118 -400 85174 60 8 la_data_in_mprj[67]
port 223 nsew signal output
rlabel metal2 s 85578 -400 85634 60 8 la_data_in_mprj[68]
port 224 nsew signal output
rlabel metal2 s 86038 -400 86094 60 8 la_data_in_mprj[69]
port 225 nsew signal output
rlabel metal2 s 58530 -400 58586 60 8 la_data_in_mprj[6]
port 226 nsew signal output
rlabel metal2 s 86406 -400 86462 60 8 la_data_in_mprj[70]
port 227 nsew signal output
rlabel metal2 s 86866 -400 86922 60 8 la_data_in_mprj[71]
port 228 nsew signal output
rlabel metal2 s 87326 -400 87382 60 8 la_data_in_mprj[72]
port 229 nsew signal output
rlabel metal2 s 87786 -400 87842 60 8 la_data_in_mprj[73]
port 230 nsew signal output
rlabel metal2 s 88154 -400 88210 60 8 la_data_in_mprj[74]
port 231 nsew signal output
rlabel metal2 s 88614 -400 88670 60 8 la_data_in_mprj[75]
port 232 nsew signal output
rlabel metal2 s 89074 -400 89130 60 8 la_data_in_mprj[76]
port 233 nsew signal output
rlabel metal2 s 89442 -400 89498 60 8 la_data_in_mprj[77]
port 234 nsew signal output
rlabel metal2 s 89902 -400 89958 60 8 la_data_in_mprj[78]
port 235 nsew signal output
rlabel metal2 s 90362 -400 90418 60 8 la_data_in_mprj[79]
port 236 nsew signal output
rlabel metal2 s 58990 -400 59046 60 8 la_data_in_mprj[7]
port 237 nsew signal output
rlabel metal2 s 90822 -400 90878 60 8 la_data_in_mprj[80]
port 238 nsew signal output
rlabel metal2 s 91190 -400 91246 60 8 la_data_in_mprj[81]
port 239 nsew signal output
rlabel metal2 s 91650 -400 91706 60 8 la_data_in_mprj[82]
port 240 nsew signal output
rlabel metal2 s 92110 -400 92166 60 8 la_data_in_mprj[83]
port 241 nsew signal output
rlabel metal2 s 92570 -400 92626 60 8 la_data_in_mprj[84]
port 242 nsew signal output
rlabel metal2 s 92938 -400 92994 60 8 la_data_in_mprj[85]
port 243 nsew signal output
rlabel metal2 s 93398 -400 93454 60 8 la_data_in_mprj[86]
port 244 nsew signal output
rlabel metal2 s 93858 -400 93914 60 8 la_data_in_mprj[87]
port 245 nsew signal output
rlabel metal2 s 94318 -400 94374 60 8 la_data_in_mprj[88]
port 246 nsew signal output
rlabel metal2 s 94686 -400 94742 60 8 la_data_in_mprj[89]
port 247 nsew signal output
rlabel metal2 s 59450 -400 59506 60 8 la_data_in_mprj[8]
port 248 nsew signal output
rlabel metal2 s 95146 -400 95202 60 8 la_data_in_mprj[90]
port 249 nsew signal output
rlabel metal2 s 95606 -400 95662 60 8 la_data_in_mprj[91]
port 250 nsew signal output
rlabel metal2 s 96066 -400 96122 60 8 la_data_in_mprj[92]
port 251 nsew signal output
rlabel metal2 s 96434 -400 96490 60 8 la_data_in_mprj[93]
port 252 nsew signal output
rlabel metal2 s 96894 -400 96950 60 8 la_data_in_mprj[94]
port 253 nsew signal output
rlabel metal2 s 97354 -400 97410 60 8 la_data_in_mprj[95]
port 254 nsew signal output
rlabel metal2 s 97722 -400 97778 60 8 la_data_in_mprj[96]
port 255 nsew signal output
rlabel metal2 s 98182 -400 98238 60 8 la_data_in_mprj[97]
port 256 nsew signal output
rlabel metal2 s 98642 -400 98698 60 8 la_data_in_mprj[98]
port 257 nsew signal output
rlabel metal2 s 99102 -400 99158 60 8 la_data_in_mprj[99]
port 258 nsew signal output
rlabel metal2 s 59818 -400 59874 60 8 la_data_in_mprj[9]
port 259 nsew signal output
rlabel metal2 s 57702 17940 57758 18400 6 la_data_out_core[0]
port 260 nsew signal input
rlabel metal2 s 101218 17940 101274 18400 6 la_data_out_core[100]
port 261 nsew signal input
rlabel metal2 s 101678 17940 101734 18400 6 la_data_out_core[101]
port 262 nsew signal input
rlabel metal2 s 102138 17940 102194 18400 6 la_data_out_core[102]
port 263 nsew signal input
rlabel metal2 s 102598 17940 102654 18400 6 la_data_out_core[103]
port 264 nsew signal input
rlabel metal2 s 102966 17940 103022 18400 6 la_data_out_core[104]
port 265 nsew signal input
rlabel metal2 s 103426 17940 103482 18400 6 la_data_out_core[105]
port 266 nsew signal input
rlabel metal2 s 103886 17940 103942 18400 6 la_data_out_core[106]
port 267 nsew signal input
rlabel metal2 s 104254 17940 104310 18400 6 la_data_out_core[107]
port 268 nsew signal input
rlabel metal2 s 104714 17940 104770 18400 6 la_data_out_core[108]
port 269 nsew signal input
rlabel metal2 s 105174 17940 105230 18400 6 la_data_out_core[109]
port 270 nsew signal input
rlabel metal2 s 62026 17940 62082 18400 6 la_data_out_core[10]
port 271 nsew signal input
rlabel metal2 s 105634 17940 105690 18400 6 la_data_out_core[110]
port 272 nsew signal input
rlabel metal2 s 106002 17940 106058 18400 6 la_data_out_core[111]
port 273 nsew signal input
rlabel metal2 s 106462 17940 106518 18400 6 la_data_out_core[112]
port 274 nsew signal input
rlabel metal2 s 106922 17940 106978 18400 6 la_data_out_core[113]
port 275 nsew signal input
rlabel metal2 s 107382 17940 107438 18400 6 la_data_out_core[114]
port 276 nsew signal input
rlabel metal2 s 107750 17940 107806 18400 6 la_data_out_core[115]
port 277 nsew signal input
rlabel metal2 s 108210 17940 108266 18400 6 la_data_out_core[116]
port 278 nsew signal input
rlabel metal2 s 108670 17940 108726 18400 6 la_data_out_core[117]
port 279 nsew signal input
rlabel metal2 s 109130 17940 109186 18400 6 la_data_out_core[118]
port 280 nsew signal input
rlabel metal2 s 109498 17940 109554 18400 6 la_data_out_core[119]
port 281 nsew signal input
rlabel metal2 s 62486 17940 62542 18400 6 la_data_out_core[11]
port 282 nsew signal input
rlabel metal2 s 109958 17940 110014 18400 6 la_data_out_core[120]
port 283 nsew signal input
rlabel metal2 s 110418 17940 110474 18400 6 la_data_out_core[121]
port 284 nsew signal input
rlabel metal2 s 110878 17940 110934 18400 6 la_data_out_core[122]
port 285 nsew signal input
rlabel metal2 s 111246 17940 111302 18400 6 la_data_out_core[123]
port 286 nsew signal input
rlabel metal2 s 111706 17940 111762 18400 6 la_data_out_core[124]
port 287 nsew signal input
rlabel metal2 s 112166 17940 112222 18400 6 la_data_out_core[125]
port 288 nsew signal input
rlabel metal2 s 112534 17940 112590 18400 6 la_data_out_core[126]
port 289 nsew signal input
rlabel metal2 s 112994 17940 113050 18400 6 la_data_out_core[127]
port 290 nsew signal input
rlabel metal2 s 62946 17940 63002 18400 6 la_data_out_core[12]
port 291 nsew signal input
rlabel metal2 s 63314 17940 63370 18400 6 la_data_out_core[13]
port 292 nsew signal input
rlabel metal2 s 63774 17940 63830 18400 6 la_data_out_core[14]
port 293 nsew signal input
rlabel metal2 s 64234 17940 64290 18400 6 la_data_out_core[15]
port 294 nsew signal input
rlabel metal2 s 64602 17940 64658 18400 6 la_data_out_core[16]
port 295 nsew signal input
rlabel metal2 s 65062 17940 65118 18400 6 la_data_out_core[17]
port 296 nsew signal input
rlabel metal2 s 65522 17940 65578 18400 6 la_data_out_core[18]
port 297 nsew signal input
rlabel metal2 s 65982 17940 66038 18400 6 la_data_out_core[19]
port 298 nsew signal input
rlabel metal2 s 58070 17940 58126 18400 6 la_data_out_core[1]
port 299 nsew signal input
rlabel metal2 s 66350 17940 66406 18400 6 la_data_out_core[20]
port 300 nsew signal input
rlabel metal2 s 66810 17940 66866 18400 6 la_data_out_core[21]
port 301 nsew signal input
rlabel metal2 s 67270 17940 67326 18400 6 la_data_out_core[22]
port 302 nsew signal input
rlabel metal2 s 67730 17940 67786 18400 6 la_data_out_core[23]
port 303 nsew signal input
rlabel metal2 s 68098 17940 68154 18400 6 la_data_out_core[24]
port 304 nsew signal input
rlabel metal2 s 68558 17940 68614 18400 6 la_data_out_core[25]
port 305 nsew signal input
rlabel metal2 s 69018 17940 69074 18400 6 la_data_out_core[26]
port 306 nsew signal input
rlabel metal2 s 69478 17940 69534 18400 6 la_data_out_core[27]
port 307 nsew signal input
rlabel metal2 s 69846 17940 69902 18400 6 la_data_out_core[28]
port 308 nsew signal input
rlabel metal2 s 70306 17940 70362 18400 6 la_data_out_core[29]
port 309 nsew signal input
rlabel metal2 s 58530 17940 58586 18400 6 la_data_out_core[2]
port 310 nsew signal input
rlabel metal2 s 70766 17940 70822 18400 6 la_data_out_core[30]
port 311 nsew signal input
rlabel metal2 s 71226 17940 71282 18400 6 la_data_out_core[31]
port 312 nsew signal input
rlabel metal2 s 71594 17940 71650 18400 6 la_data_out_core[32]
port 313 nsew signal input
rlabel metal2 s 72054 17940 72110 18400 6 la_data_out_core[33]
port 314 nsew signal input
rlabel metal2 s 72514 17940 72570 18400 6 la_data_out_core[34]
port 315 nsew signal input
rlabel metal2 s 72882 17940 72938 18400 6 la_data_out_core[35]
port 316 nsew signal input
rlabel metal2 s 73342 17940 73398 18400 6 la_data_out_core[36]
port 317 nsew signal input
rlabel metal2 s 73802 17940 73858 18400 6 la_data_out_core[37]
port 318 nsew signal input
rlabel metal2 s 74262 17940 74318 18400 6 la_data_out_core[38]
port 319 nsew signal input
rlabel metal2 s 74630 17940 74686 18400 6 la_data_out_core[39]
port 320 nsew signal input
rlabel metal2 s 58990 17940 59046 18400 6 la_data_out_core[3]
port 321 nsew signal input
rlabel metal2 s 75090 17940 75146 18400 6 la_data_out_core[40]
port 322 nsew signal input
rlabel metal2 s 75550 17940 75606 18400 6 la_data_out_core[41]
port 323 nsew signal input
rlabel metal2 s 76010 17940 76066 18400 6 la_data_out_core[42]
port 324 nsew signal input
rlabel metal2 s 76378 17940 76434 18400 6 la_data_out_core[43]
port 325 nsew signal input
rlabel metal2 s 76838 17940 76894 18400 6 la_data_out_core[44]
port 326 nsew signal input
rlabel metal2 s 77298 17940 77354 18400 6 la_data_out_core[45]
port 327 nsew signal input
rlabel metal2 s 77758 17940 77814 18400 6 la_data_out_core[46]
port 328 nsew signal input
rlabel metal2 s 78126 17940 78182 18400 6 la_data_out_core[47]
port 329 nsew signal input
rlabel metal2 s 78586 17940 78642 18400 6 la_data_out_core[48]
port 330 nsew signal input
rlabel metal2 s 79046 17940 79102 18400 6 la_data_out_core[49]
port 331 nsew signal input
rlabel metal2 s 59450 17940 59506 18400 6 la_data_out_core[4]
port 332 nsew signal input
rlabel metal2 s 79506 17940 79562 18400 6 la_data_out_core[50]
port 333 nsew signal input
rlabel metal2 s 79874 17940 79930 18400 6 la_data_out_core[51]
port 334 nsew signal input
rlabel metal2 s 80334 17940 80390 18400 6 la_data_out_core[52]
port 335 nsew signal input
rlabel metal2 s 80794 17940 80850 18400 6 la_data_out_core[53]
port 336 nsew signal input
rlabel metal2 s 81162 17940 81218 18400 6 la_data_out_core[54]
port 337 nsew signal input
rlabel metal2 s 81622 17940 81678 18400 6 la_data_out_core[55]
port 338 nsew signal input
rlabel metal2 s 82082 17940 82138 18400 6 la_data_out_core[56]
port 339 nsew signal input
rlabel metal2 s 82542 17940 82598 18400 6 la_data_out_core[57]
port 340 nsew signal input
rlabel metal2 s 82910 17940 82966 18400 6 la_data_out_core[58]
port 341 nsew signal input
rlabel metal2 s 83370 17940 83426 18400 6 la_data_out_core[59]
port 342 nsew signal input
rlabel metal2 s 59818 17940 59874 18400 6 la_data_out_core[5]
port 343 nsew signal input
rlabel metal2 s 83830 17940 83886 18400 6 la_data_out_core[60]
port 344 nsew signal input
rlabel metal2 s 84290 17940 84346 18400 6 la_data_out_core[61]
port 345 nsew signal input
rlabel metal2 s 84658 17940 84714 18400 6 la_data_out_core[62]
port 346 nsew signal input
rlabel metal2 s 85118 17940 85174 18400 6 la_data_out_core[63]
port 347 nsew signal input
rlabel metal2 s 85578 17940 85634 18400 6 la_data_out_core[64]
port 348 nsew signal input
rlabel metal2 s 86038 17940 86094 18400 6 la_data_out_core[65]
port 349 nsew signal input
rlabel metal2 s 86406 17940 86462 18400 6 la_data_out_core[66]
port 350 nsew signal input
rlabel metal2 s 86866 17940 86922 18400 6 la_data_out_core[67]
port 351 nsew signal input
rlabel metal2 s 87326 17940 87382 18400 6 la_data_out_core[68]
port 352 nsew signal input
rlabel metal2 s 87786 17940 87842 18400 6 la_data_out_core[69]
port 353 nsew signal input
rlabel metal2 s 60278 17940 60334 18400 6 la_data_out_core[6]
port 354 nsew signal input
rlabel metal2 s 88154 17940 88210 18400 6 la_data_out_core[70]
port 355 nsew signal input
rlabel metal2 s 88614 17940 88670 18400 6 la_data_out_core[71]
port 356 nsew signal input
rlabel metal2 s 89074 17940 89130 18400 6 la_data_out_core[72]
port 357 nsew signal input
rlabel metal2 s 89442 17940 89498 18400 6 la_data_out_core[73]
port 358 nsew signal input
rlabel metal2 s 89902 17940 89958 18400 6 la_data_out_core[74]
port 359 nsew signal input
rlabel metal2 s 90362 17940 90418 18400 6 la_data_out_core[75]
port 360 nsew signal input
rlabel metal2 s 90822 17940 90878 18400 6 la_data_out_core[76]
port 361 nsew signal input
rlabel metal2 s 91190 17940 91246 18400 6 la_data_out_core[77]
port 362 nsew signal input
rlabel metal2 s 91650 17940 91706 18400 6 la_data_out_core[78]
port 363 nsew signal input
rlabel metal2 s 92110 17940 92166 18400 6 la_data_out_core[79]
port 364 nsew signal input
rlabel metal2 s 60738 17940 60794 18400 6 la_data_out_core[7]
port 365 nsew signal input
rlabel metal2 s 92570 17940 92626 18400 6 la_data_out_core[80]
port 366 nsew signal input
rlabel metal2 s 92938 17940 92994 18400 6 la_data_out_core[81]
port 367 nsew signal input
rlabel metal2 s 93398 17940 93454 18400 6 la_data_out_core[82]
port 368 nsew signal input
rlabel metal2 s 93858 17940 93914 18400 6 la_data_out_core[83]
port 369 nsew signal input
rlabel metal2 s 94318 17940 94374 18400 6 la_data_out_core[84]
port 370 nsew signal input
rlabel metal2 s 94686 17940 94742 18400 6 la_data_out_core[85]
port 371 nsew signal input
rlabel metal2 s 95146 17940 95202 18400 6 la_data_out_core[86]
port 372 nsew signal input
rlabel metal2 s 95606 17940 95662 18400 6 la_data_out_core[87]
port 373 nsew signal input
rlabel metal2 s 96066 17940 96122 18400 6 la_data_out_core[88]
port 374 nsew signal input
rlabel metal2 s 96434 17940 96490 18400 6 la_data_out_core[89]
port 375 nsew signal input
rlabel metal2 s 61198 17940 61254 18400 6 la_data_out_core[8]
port 376 nsew signal input
rlabel metal2 s 96894 17940 96950 18400 6 la_data_out_core[90]
port 377 nsew signal input
rlabel metal2 s 97354 17940 97410 18400 6 la_data_out_core[91]
port 378 nsew signal input
rlabel metal2 s 97722 17940 97778 18400 6 la_data_out_core[92]
port 379 nsew signal input
rlabel metal2 s 98182 17940 98238 18400 6 la_data_out_core[93]
port 380 nsew signal input
rlabel metal2 s 98642 17940 98698 18400 6 la_data_out_core[94]
port 381 nsew signal input
rlabel metal2 s 99102 17940 99158 18400 6 la_data_out_core[95]
port 382 nsew signal input
rlabel metal2 s 99470 17940 99526 18400 6 la_data_out_core[96]
port 383 nsew signal input
rlabel metal2 s 99930 17940 99986 18400 6 la_data_out_core[97]
port 384 nsew signal input
rlabel metal2 s 100390 17940 100446 18400 6 la_data_out_core[98]
port 385 nsew signal input
rlabel metal2 s 100850 17940 100906 18400 6 la_data_out_core[99]
port 386 nsew signal input
rlabel metal2 s 61566 17940 61622 18400 6 la_data_out_core[9]
port 387 nsew signal input
rlabel metal2 s 202 -400 258 60 8 la_data_out_mprj[0]
port 388 nsew signal input
rlabel metal2 s 43718 -400 43774 60 8 la_data_out_mprj[100]
port 389 nsew signal input
rlabel metal2 s 44178 -400 44234 60 8 la_data_out_mprj[101]
port 390 nsew signal input
rlabel metal2 s 44638 -400 44694 60 8 la_data_out_mprj[102]
port 391 nsew signal input
rlabel metal2 s 45006 -400 45062 60 8 la_data_out_mprj[103]
port 392 nsew signal input
rlabel metal2 s 45466 -400 45522 60 8 la_data_out_mprj[104]
port 393 nsew signal input
rlabel metal2 s 45926 -400 45982 60 8 la_data_out_mprj[105]
port 394 nsew signal input
rlabel metal2 s 46386 -400 46442 60 8 la_data_out_mprj[106]
port 395 nsew signal input
rlabel metal2 s 46754 -400 46810 60 8 la_data_out_mprj[107]
port 396 nsew signal input
rlabel metal2 s 47214 -400 47270 60 8 la_data_out_mprj[108]
port 397 nsew signal input
rlabel metal2 s 47674 -400 47730 60 8 la_data_out_mprj[109]
port 398 nsew signal input
rlabel metal2 s 4526 -400 4582 60 8 la_data_out_mprj[10]
port 399 nsew signal input
rlabel metal2 s 48134 -400 48190 60 8 la_data_out_mprj[110]
port 400 nsew signal input
rlabel metal2 s 48502 -400 48558 60 8 la_data_out_mprj[111]
port 401 nsew signal input
rlabel metal2 s 48962 -400 49018 60 8 la_data_out_mprj[112]
port 402 nsew signal input
rlabel metal2 s 49422 -400 49478 60 8 la_data_out_mprj[113]
port 403 nsew signal input
rlabel metal2 s 49790 -400 49846 60 8 la_data_out_mprj[114]
port 404 nsew signal input
rlabel metal2 s 50250 -400 50306 60 8 la_data_out_mprj[115]
port 405 nsew signal input
rlabel metal2 s 50710 -400 50766 60 8 la_data_out_mprj[116]
port 406 nsew signal input
rlabel metal2 s 51170 -400 51226 60 8 la_data_out_mprj[117]
port 407 nsew signal input
rlabel metal2 s 51538 -400 51594 60 8 la_data_out_mprj[118]
port 408 nsew signal input
rlabel metal2 s 51998 -400 52054 60 8 la_data_out_mprj[119]
port 409 nsew signal input
rlabel metal2 s 4986 -400 5042 60 8 la_data_out_mprj[11]
port 410 nsew signal input
rlabel metal2 s 52458 -400 52514 60 8 la_data_out_mprj[120]
port 411 nsew signal input
rlabel metal2 s 52918 -400 52974 60 8 la_data_out_mprj[121]
port 412 nsew signal input
rlabel metal2 s 53286 -400 53342 60 8 la_data_out_mprj[122]
port 413 nsew signal input
rlabel metal2 s 53746 -400 53802 60 8 la_data_out_mprj[123]
port 414 nsew signal input
rlabel metal2 s 54206 -400 54262 60 8 la_data_out_mprj[124]
port 415 nsew signal input
rlabel metal2 s 54666 -400 54722 60 8 la_data_out_mprj[125]
port 416 nsew signal input
rlabel metal2 s 55034 -400 55090 60 8 la_data_out_mprj[126]
port 417 nsew signal input
rlabel metal2 s 55494 -400 55550 60 8 la_data_out_mprj[127]
port 418 nsew signal input
rlabel metal2 s 5354 -400 5410 60 8 la_data_out_mprj[12]
port 419 nsew signal input
rlabel metal2 s 5814 -400 5870 60 8 la_data_out_mprj[13]
port 420 nsew signal input
rlabel metal2 s 6274 -400 6330 60 8 la_data_out_mprj[14]
port 421 nsew signal input
rlabel metal2 s 6734 -400 6790 60 8 la_data_out_mprj[15]
port 422 nsew signal input
rlabel metal2 s 7102 -400 7158 60 8 la_data_out_mprj[16]
port 423 nsew signal input
rlabel metal2 s 7562 -400 7618 60 8 la_data_out_mprj[17]
port 424 nsew signal input
rlabel metal2 s 8022 -400 8078 60 8 la_data_out_mprj[18]
port 425 nsew signal input
rlabel metal2 s 8390 -400 8446 60 8 la_data_out_mprj[19]
port 426 nsew signal input
rlabel metal2 s 570 -400 626 60 8 la_data_out_mprj[1]
port 427 nsew signal input
rlabel metal2 s 8850 -400 8906 60 8 la_data_out_mprj[20]
port 428 nsew signal input
rlabel metal2 s 9310 -400 9366 60 8 la_data_out_mprj[21]
port 429 nsew signal input
rlabel metal2 s 9770 -400 9826 60 8 la_data_out_mprj[22]
port 430 nsew signal input
rlabel metal2 s 10138 -400 10194 60 8 la_data_out_mprj[23]
port 431 nsew signal input
rlabel metal2 s 10598 -400 10654 60 8 la_data_out_mprj[24]
port 432 nsew signal input
rlabel metal2 s 11058 -400 11114 60 8 la_data_out_mprj[25]
port 433 nsew signal input
rlabel metal2 s 11518 -400 11574 60 8 la_data_out_mprj[26]
port 434 nsew signal input
rlabel metal2 s 11886 -400 11942 60 8 la_data_out_mprj[27]
port 435 nsew signal input
rlabel metal2 s 12346 -400 12402 60 8 la_data_out_mprj[28]
port 436 nsew signal input
rlabel metal2 s 12806 -400 12862 60 8 la_data_out_mprj[29]
port 437 nsew signal input
rlabel metal2 s 1030 -400 1086 60 8 la_data_out_mprj[2]
port 438 nsew signal input
rlabel metal2 s 13266 -400 13322 60 8 la_data_out_mprj[30]
port 439 nsew signal input
rlabel metal2 s 13634 -400 13690 60 8 la_data_out_mprj[31]
port 440 nsew signal input
rlabel metal2 s 14094 -400 14150 60 8 la_data_out_mprj[32]
port 441 nsew signal input
rlabel metal2 s 14554 -400 14610 60 8 la_data_out_mprj[33]
port 442 nsew signal input
rlabel metal2 s 15014 -400 15070 60 8 la_data_out_mprj[34]
port 443 nsew signal input
rlabel metal2 s 15382 -400 15438 60 8 la_data_out_mprj[35]
port 444 nsew signal input
rlabel metal2 s 15842 -400 15898 60 8 la_data_out_mprj[36]
port 445 nsew signal input
rlabel metal2 s 16302 -400 16358 60 8 la_data_out_mprj[37]
port 446 nsew signal input
rlabel metal2 s 16670 -400 16726 60 8 la_data_out_mprj[38]
port 447 nsew signal input
rlabel metal2 s 17130 -400 17186 60 8 la_data_out_mprj[39]
port 448 nsew signal input
rlabel metal2 s 1490 -400 1546 60 8 la_data_out_mprj[3]
port 449 nsew signal input
rlabel metal2 s 17590 -400 17646 60 8 la_data_out_mprj[40]
port 450 nsew signal input
rlabel metal2 s 18050 -400 18106 60 8 la_data_out_mprj[41]
port 451 nsew signal input
rlabel metal2 s 18418 -400 18474 60 8 la_data_out_mprj[42]
port 452 nsew signal input
rlabel metal2 s 18878 -400 18934 60 8 la_data_out_mprj[43]
port 453 nsew signal input
rlabel metal2 s 19338 -400 19394 60 8 la_data_out_mprj[44]
port 454 nsew signal input
rlabel metal2 s 19798 -400 19854 60 8 la_data_out_mprj[45]
port 455 nsew signal input
rlabel metal2 s 20166 -400 20222 60 8 la_data_out_mprj[46]
port 456 nsew signal input
rlabel metal2 s 20626 -400 20682 60 8 la_data_out_mprj[47]
port 457 nsew signal input
rlabel metal2 s 21086 -400 21142 60 8 la_data_out_mprj[48]
port 458 nsew signal input
rlabel metal2 s 21546 -400 21602 60 8 la_data_out_mprj[49]
port 459 nsew signal input
rlabel metal2 s 1858 -400 1914 60 8 la_data_out_mprj[4]
port 460 nsew signal input
rlabel metal2 s 21914 -400 21970 60 8 la_data_out_mprj[50]
port 461 nsew signal input
rlabel metal2 s 22374 -400 22430 60 8 la_data_out_mprj[51]
port 462 nsew signal input
rlabel metal2 s 22834 -400 22890 60 8 la_data_out_mprj[52]
port 463 nsew signal input
rlabel metal2 s 23294 -400 23350 60 8 la_data_out_mprj[53]
port 464 nsew signal input
rlabel metal2 s 23662 -400 23718 60 8 la_data_out_mprj[54]
port 465 nsew signal input
rlabel metal2 s 24122 -400 24178 60 8 la_data_out_mprj[55]
port 466 nsew signal input
rlabel metal2 s 24582 -400 24638 60 8 la_data_out_mprj[56]
port 467 nsew signal input
rlabel metal2 s 24950 -400 25006 60 8 la_data_out_mprj[57]
port 468 nsew signal input
rlabel metal2 s 25410 -400 25466 60 8 la_data_out_mprj[58]
port 469 nsew signal input
rlabel metal2 s 25870 -400 25926 60 8 la_data_out_mprj[59]
port 470 nsew signal input
rlabel metal2 s 2318 -400 2374 60 8 la_data_out_mprj[5]
port 471 nsew signal input
rlabel metal2 s 26330 -400 26386 60 8 la_data_out_mprj[60]
port 472 nsew signal input
rlabel metal2 s 26698 -400 26754 60 8 la_data_out_mprj[61]
port 473 nsew signal input
rlabel metal2 s 27158 -400 27214 60 8 la_data_out_mprj[62]
port 474 nsew signal input
rlabel metal2 s 27618 -400 27674 60 8 la_data_out_mprj[63]
port 475 nsew signal input
rlabel metal2 s 28078 -400 28134 60 8 la_data_out_mprj[64]
port 476 nsew signal input
rlabel metal2 s 28446 -400 28502 60 8 la_data_out_mprj[65]
port 477 nsew signal input
rlabel metal2 s 28906 -400 28962 60 8 la_data_out_mprj[66]
port 478 nsew signal input
rlabel metal2 s 29366 -400 29422 60 8 la_data_out_mprj[67]
port 479 nsew signal input
rlabel metal2 s 29826 -400 29882 60 8 la_data_out_mprj[68]
port 480 nsew signal input
rlabel metal2 s 30194 -400 30250 60 8 la_data_out_mprj[69]
port 481 nsew signal input
rlabel metal2 s 2778 -400 2834 60 8 la_data_out_mprj[6]
port 482 nsew signal input
rlabel metal2 s 30654 -400 30710 60 8 la_data_out_mprj[70]
port 483 nsew signal input
rlabel metal2 s 31114 -400 31170 60 8 la_data_out_mprj[71]
port 484 nsew signal input
rlabel metal2 s 31574 -400 31630 60 8 la_data_out_mprj[72]
port 485 nsew signal input
rlabel metal2 s 31942 -400 31998 60 8 la_data_out_mprj[73]
port 486 nsew signal input
rlabel metal2 s 32402 -400 32458 60 8 la_data_out_mprj[74]
port 487 nsew signal input
rlabel metal2 s 32862 -400 32918 60 8 la_data_out_mprj[75]
port 488 nsew signal input
rlabel metal2 s 33230 -400 33286 60 8 la_data_out_mprj[76]
port 489 nsew signal input
rlabel metal2 s 33690 -400 33746 60 8 la_data_out_mprj[77]
port 490 nsew signal input
rlabel metal2 s 34150 -400 34206 60 8 la_data_out_mprj[78]
port 491 nsew signal input
rlabel metal2 s 34610 -400 34666 60 8 la_data_out_mprj[79]
port 492 nsew signal input
rlabel metal2 s 3238 -400 3294 60 8 la_data_out_mprj[7]
port 493 nsew signal input
rlabel metal2 s 34978 -400 35034 60 8 la_data_out_mprj[80]
port 494 nsew signal input
rlabel metal2 s 35438 -400 35494 60 8 la_data_out_mprj[81]
port 495 nsew signal input
rlabel metal2 s 35898 -400 35954 60 8 la_data_out_mprj[82]
port 496 nsew signal input
rlabel metal2 s 36358 -400 36414 60 8 la_data_out_mprj[83]
port 497 nsew signal input
rlabel metal2 s 36726 -400 36782 60 8 la_data_out_mprj[84]
port 498 nsew signal input
rlabel metal2 s 37186 -400 37242 60 8 la_data_out_mprj[85]
port 499 nsew signal input
rlabel metal2 s 37646 -400 37702 60 8 la_data_out_mprj[86]
port 500 nsew signal input
rlabel metal2 s 38106 -400 38162 60 8 la_data_out_mprj[87]
port 501 nsew signal input
rlabel metal2 s 38474 -400 38530 60 8 la_data_out_mprj[88]
port 502 nsew signal input
rlabel metal2 s 38934 -400 38990 60 8 la_data_out_mprj[89]
port 503 nsew signal input
rlabel metal2 s 3606 -400 3662 60 8 la_data_out_mprj[8]
port 504 nsew signal input
rlabel metal2 s 39394 -400 39450 60 8 la_data_out_mprj[90]
port 505 nsew signal input
rlabel metal2 s 39854 -400 39910 60 8 la_data_out_mprj[91]
port 506 nsew signal input
rlabel metal2 s 40222 -400 40278 60 8 la_data_out_mprj[92]
port 507 nsew signal input
rlabel metal2 s 40682 -400 40738 60 8 la_data_out_mprj[93]
port 508 nsew signal input
rlabel metal2 s 41142 -400 41198 60 8 la_data_out_mprj[94]
port 509 nsew signal input
rlabel metal2 s 41510 -400 41566 60 8 la_data_out_mprj[95]
port 510 nsew signal input
rlabel metal2 s 41970 -400 42026 60 8 la_data_out_mprj[96]
port 511 nsew signal input
rlabel metal2 s 42430 -400 42486 60 8 la_data_out_mprj[97]
port 512 nsew signal input
rlabel metal2 s 42890 -400 42946 60 8 la_data_out_mprj[98]
port 513 nsew signal input
rlabel metal2 s 43258 -400 43314 60 8 la_data_out_mprj[99]
port 514 nsew signal input
rlabel metal2 s 4066 -400 4122 60 8 la_data_out_mprj[9]
port 515 nsew signal input
rlabel metal2 s 113454 17940 113510 18400 6 la_oen_core[0]
port 516 nsew signal output
rlabel metal2 s 157062 17940 157118 18400 6 la_oen_core[100]
port 517 nsew signal output
rlabel metal2 s 157430 17940 157486 18400 6 la_oen_core[101]
port 518 nsew signal output
rlabel metal2 s 157890 17940 157946 18400 6 la_oen_core[102]
port 519 nsew signal output
rlabel metal2 s 158350 17940 158406 18400 6 la_oen_core[103]
port 520 nsew signal output
rlabel metal2 s 158810 17940 158866 18400 6 la_oen_core[104]
port 521 nsew signal output
rlabel metal2 s 159178 17940 159234 18400 6 la_oen_core[105]
port 522 nsew signal output
rlabel metal2 s 159638 17940 159694 18400 6 la_oen_core[106]
port 523 nsew signal output
rlabel metal2 s 160098 17940 160154 18400 6 la_oen_core[107]
port 524 nsew signal output
rlabel metal2 s 160466 17940 160522 18400 6 la_oen_core[108]
port 525 nsew signal output
rlabel metal2 s 160926 17940 160982 18400 6 la_oen_core[109]
port 526 nsew signal output
rlabel metal2 s 117778 17940 117834 18400 6 la_oen_core[10]
port 527 nsew signal output
rlabel metal2 s 161386 17940 161442 18400 6 la_oen_core[110]
port 528 nsew signal output
rlabel metal2 s 161846 17940 161902 18400 6 la_oen_core[111]
port 529 nsew signal output
rlabel metal2 s 162214 17940 162270 18400 6 la_oen_core[112]
port 530 nsew signal output
rlabel metal2 s 162674 17940 162730 18400 6 la_oen_core[113]
port 531 nsew signal output
rlabel metal2 s 163134 17940 163190 18400 6 la_oen_core[114]
port 532 nsew signal output
rlabel metal2 s 163594 17940 163650 18400 6 la_oen_core[115]
port 533 nsew signal output
rlabel metal2 s 163962 17940 164018 18400 6 la_oen_core[116]
port 534 nsew signal output
rlabel metal2 s 164422 17940 164478 18400 6 la_oen_core[117]
port 535 nsew signal output
rlabel metal2 s 164882 17940 164938 18400 6 la_oen_core[118]
port 536 nsew signal output
rlabel metal2 s 165342 17940 165398 18400 6 la_oen_core[119]
port 537 nsew signal output
rlabel metal2 s 118238 17940 118294 18400 6 la_oen_core[11]
port 538 nsew signal output
rlabel metal2 s 165710 17940 165766 18400 6 la_oen_core[120]
port 539 nsew signal output
rlabel metal2 s 166170 17940 166226 18400 6 la_oen_core[121]
port 540 nsew signal output
rlabel metal2 s 166630 17940 166686 18400 6 la_oen_core[122]
port 541 nsew signal output
rlabel metal2 s 167090 17940 167146 18400 6 la_oen_core[123]
port 542 nsew signal output
rlabel metal2 s 167458 17940 167514 18400 6 la_oen_core[124]
port 543 nsew signal output
rlabel metal2 s 167918 17940 167974 18400 6 la_oen_core[125]
port 544 nsew signal output
rlabel metal2 s 168378 17940 168434 18400 6 la_oen_core[126]
port 545 nsew signal output
rlabel metal2 s 168746 17940 168802 18400 6 la_oen_core[127]
port 546 nsew signal output
rlabel metal2 s 118698 17940 118754 18400 6 la_oen_core[12]
port 547 nsew signal output
rlabel metal2 s 119158 17940 119214 18400 6 la_oen_core[13]
port 548 nsew signal output
rlabel metal2 s 119526 17940 119582 18400 6 la_oen_core[14]
port 549 nsew signal output
rlabel metal2 s 119986 17940 120042 18400 6 la_oen_core[15]
port 550 nsew signal output
rlabel metal2 s 120446 17940 120502 18400 6 la_oen_core[16]
port 551 nsew signal output
rlabel metal2 s 120814 17940 120870 18400 6 la_oen_core[17]
port 552 nsew signal output
rlabel metal2 s 121274 17940 121330 18400 6 la_oen_core[18]
port 553 nsew signal output
rlabel metal2 s 121734 17940 121790 18400 6 la_oen_core[19]
port 554 nsew signal output
rlabel metal2 s 113914 17940 113970 18400 6 la_oen_core[1]
port 555 nsew signal output
rlabel metal2 s 122194 17940 122250 18400 6 la_oen_core[20]
port 556 nsew signal output
rlabel metal2 s 122562 17940 122618 18400 6 la_oen_core[21]
port 557 nsew signal output
rlabel metal2 s 123022 17940 123078 18400 6 la_oen_core[22]
port 558 nsew signal output
rlabel metal2 s 123482 17940 123538 18400 6 la_oen_core[23]
port 559 nsew signal output
rlabel metal2 s 123942 17940 123998 18400 6 la_oen_core[24]
port 560 nsew signal output
rlabel metal2 s 124310 17940 124366 18400 6 la_oen_core[25]
port 561 nsew signal output
rlabel metal2 s 124770 17940 124826 18400 6 la_oen_core[26]
port 562 nsew signal output
rlabel metal2 s 125230 17940 125286 18400 6 la_oen_core[27]
port 563 nsew signal output
rlabel metal2 s 125690 17940 125746 18400 6 la_oen_core[28]
port 564 nsew signal output
rlabel metal2 s 126058 17940 126114 18400 6 la_oen_core[29]
port 565 nsew signal output
rlabel metal2 s 114282 17940 114338 18400 6 la_oen_core[2]
port 566 nsew signal output
rlabel metal2 s 126518 17940 126574 18400 6 la_oen_core[30]
port 567 nsew signal output
rlabel metal2 s 126978 17940 127034 18400 6 la_oen_core[31]
port 568 nsew signal output
rlabel metal2 s 127438 17940 127494 18400 6 la_oen_core[32]
port 569 nsew signal output
rlabel metal2 s 127806 17940 127862 18400 6 la_oen_core[33]
port 570 nsew signal output
rlabel metal2 s 128266 17940 128322 18400 6 la_oen_core[34]
port 571 nsew signal output
rlabel metal2 s 128726 17940 128782 18400 6 la_oen_core[35]
port 572 nsew signal output
rlabel metal2 s 129094 17940 129150 18400 6 la_oen_core[36]
port 573 nsew signal output
rlabel metal2 s 129554 17940 129610 18400 6 la_oen_core[37]
port 574 nsew signal output
rlabel metal2 s 130014 17940 130070 18400 6 la_oen_core[38]
port 575 nsew signal output
rlabel metal2 s 130474 17940 130530 18400 6 la_oen_core[39]
port 576 nsew signal output
rlabel metal2 s 114742 17940 114798 18400 6 la_oen_core[3]
port 577 nsew signal output
rlabel metal2 s 130842 17940 130898 18400 6 la_oen_core[40]
port 578 nsew signal output
rlabel metal2 s 131302 17940 131358 18400 6 la_oen_core[41]
port 579 nsew signal output
rlabel metal2 s 131762 17940 131818 18400 6 la_oen_core[42]
port 580 nsew signal output
rlabel metal2 s 132222 17940 132278 18400 6 la_oen_core[43]
port 581 nsew signal output
rlabel metal2 s 132590 17940 132646 18400 6 la_oen_core[44]
port 582 nsew signal output
rlabel metal2 s 133050 17940 133106 18400 6 la_oen_core[45]
port 583 nsew signal output
rlabel metal2 s 133510 17940 133566 18400 6 la_oen_core[46]
port 584 nsew signal output
rlabel metal2 s 133970 17940 134026 18400 6 la_oen_core[47]
port 585 nsew signal output
rlabel metal2 s 134338 17940 134394 18400 6 la_oen_core[48]
port 586 nsew signal output
rlabel metal2 s 134798 17940 134854 18400 6 la_oen_core[49]
port 587 nsew signal output
rlabel metal2 s 115202 17940 115258 18400 6 la_oen_core[4]
port 588 nsew signal output
rlabel metal2 s 135258 17940 135314 18400 6 la_oen_core[50]
port 589 nsew signal output
rlabel metal2 s 135718 17940 135774 18400 6 la_oen_core[51]
port 590 nsew signal output
rlabel metal2 s 136086 17940 136142 18400 6 la_oen_core[52]
port 591 nsew signal output
rlabel metal2 s 136546 17940 136602 18400 6 la_oen_core[53]
port 592 nsew signal output
rlabel metal2 s 137006 17940 137062 18400 6 la_oen_core[54]
port 593 nsew signal output
rlabel metal2 s 137374 17940 137430 18400 6 la_oen_core[55]
port 594 nsew signal output
rlabel metal2 s 137834 17940 137890 18400 6 la_oen_core[56]
port 595 nsew signal output
rlabel metal2 s 138294 17940 138350 18400 6 la_oen_core[57]
port 596 nsew signal output
rlabel metal2 s 138754 17940 138810 18400 6 la_oen_core[58]
port 597 nsew signal output
rlabel metal2 s 139122 17940 139178 18400 6 la_oen_core[59]
port 598 nsew signal output
rlabel metal2 s 115662 17940 115718 18400 6 la_oen_core[5]
port 599 nsew signal output
rlabel metal2 s 139582 17940 139638 18400 6 la_oen_core[60]
port 600 nsew signal output
rlabel metal2 s 140042 17940 140098 18400 6 la_oen_core[61]
port 601 nsew signal output
rlabel metal2 s 140502 17940 140558 18400 6 la_oen_core[62]
port 602 nsew signal output
rlabel metal2 s 140870 17940 140926 18400 6 la_oen_core[63]
port 603 nsew signal output
rlabel metal2 s 141330 17940 141386 18400 6 la_oen_core[64]
port 604 nsew signal output
rlabel metal2 s 141790 17940 141846 18400 6 la_oen_core[65]
port 605 nsew signal output
rlabel metal2 s 142250 17940 142306 18400 6 la_oen_core[66]
port 606 nsew signal output
rlabel metal2 s 142618 17940 142674 18400 6 la_oen_core[67]
port 607 nsew signal output
rlabel metal2 s 143078 17940 143134 18400 6 la_oen_core[68]
port 608 nsew signal output
rlabel metal2 s 143538 17940 143594 18400 6 la_oen_core[69]
port 609 nsew signal output
rlabel metal2 s 116030 17940 116086 18400 6 la_oen_core[6]
port 610 nsew signal output
rlabel metal2 s 143998 17940 144054 18400 6 la_oen_core[70]
port 611 nsew signal output
rlabel metal2 s 144366 17940 144422 18400 6 la_oen_core[71]
port 612 nsew signal output
rlabel metal2 s 144826 17940 144882 18400 6 la_oen_core[72]
port 613 nsew signal output
rlabel metal2 s 145286 17940 145342 18400 6 la_oen_core[73]
port 614 nsew signal output
rlabel metal2 s 145654 17940 145710 18400 6 la_oen_core[74]
port 615 nsew signal output
rlabel metal2 s 146114 17940 146170 18400 6 la_oen_core[75]
port 616 nsew signal output
rlabel metal2 s 146574 17940 146630 18400 6 la_oen_core[76]
port 617 nsew signal output
rlabel metal2 s 147034 17940 147090 18400 6 la_oen_core[77]
port 618 nsew signal output
rlabel metal2 s 147402 17940 147458 18400 6 la_oen_core[78]
port 619 nsew signal output
rlabel metal2 s 147862 17940 147918 18400 6 la_oen_core[79]
port 620 nsew signal output
rlabel metal2 s 116490 17940 116546 18400 6 la_oen_core[7]
port 621 nsew signal output
rlabel metal2 s 148322 17940 148378 18400 6 la_oen_core[80]
port 622 nsew signal output
rlabel metal2 s 148782 17940 148838 18400 6 la_oen_core[81]
port 623 nsew signal output
rlabel metal2 s 149150 17940 149206 18400 6 la_oen_core[82]
port 624 nsew signal output
rlabel metal2 s 149610 17940 149666 18400 6 la_oen_core[83]
port 625 nsew signal output
rlabel metal2 s 150070 17940 150126 18400 6 la_oen_core[84]
port 626 nsew signal output
rlabel metal2 s 150530 17940 150586 18400 6 la_oen_core[85]
port 627 nsew signal output
rlabel metal2 s 150898 17940 150954 18400 6 la_oen_core[86]
port 628 nsew signal output
rlabel metal2 s 151358 17940 151414 18400 6 la_oen_core[87]
port 629 nsew signal output
rlabel metal2 s 151818 17940 151874 18400 6 la_oen_core[88]
port 630 nsew signal output
rlabel metal2 s 152186 17940 152242 18400 6 la_oen_core[89]
port 631 nsew signal output
rlabel metal2 s 116950 17940 117006 18400 6 la_oen_core[8]
port 632 nsew signal output
rlabel metal2 s 152646 17940 152702 18400 6 la_oen_core[90]
port 633 nsew signal output
rlabel metal2 s 153106 17940 153162 18400 6 la_oen_core[91]
port 634 nsew signal output
rlabel metal2 s 153566 17940 153622 18400 6 la_oen_core[92]
port 635 nsew signal output
rlabel metal2 s 153934 17940 153990 18400 6 la_oen_core[93]
port 636 nsew signal output
rlabel metal2 s 154394 17940 154450 18400 6 la_oen_core[94]
port 637 nsew signal output
rlabel metal2 s 154854 17940 154910 18400 6 la_oen_core[95]
port 638 nsew signal output
rlabel metal2 s 155314 17940 155370 18400 6 la_oen_core[96]
port 639 nsew signal output
rlabel metal2 s 155682 17940 155738 18400 6 la_oen_core[97]
port 640 nsew signal output
rlabel metal2 s 156142 17940 156198 18400 6 la_oen_core[98]
port 641 nsew signal output
rlabel metal2 s 156602 17940 156658 18400 6 la_oen_core[99]
port 642 nsew signal output
rlabel metal2 s 117410 17940 117466 18400 6 la_oen_core[9]
port 643 nsew signal output
rlabel metal2 s 111706 -400 111762 60 8 la_oen_mprj[0]
port 644 nsew signal input
rlabel metal2 s 155314 -400 155370 60 8 la_oen_mprj[100]
port 645 nsew signal input
rlabel metal2 s 155682 -400 155738 60 8 la_oen_mprj[101]
port 646 nsew signal input
rlabel metal2 s 156142 -400 156198 60 8 la_oen_mprj[102]
port 647 nsew signal input
rlabel metal2 s 156602 -400 156658 60 8 la_oen_mprj[103]
port 648 nsew signal input
rlabel metal2 s 157062 -400 157118 60 8 la_oen_mprj[104]
port 649 nsew signal input
rlabel metal2 s 157430 -400 157486 60 8 la_oen_mprj[105]
port 650 nsew signal input
rlabel metal2 s 157890 -400 157946 60 8 la_oen_mprj[106]
port 651 nsew signal input
rlabel metal2 s 158350 -400 158406 60 8 la_oen_mprj[107]
port 652 nsew signal input
rlabel metal2 s 158810 -400 158866 60 8 la_oen_mprj[108]
port 653 nsew signal input
rlabel metal2 s 159178 -400 159234 60 8 la_oen_mprj[109]
port 654 nsew signal input
rlabel metal2 s 116030 -400 116086 60 8 la_oen_mprj[10]
port 655 nsew signal input
rlabel metal2 s 159638 -400 159694 60 8 la_oen_mprj[110]
port 656 nsew signal input
rlabel metal2 s 160098 -400 160154 60 8 la_oen_mprj[111]
port 657 nsew signal input
rlabel metal2 s 160466 -400 160522 60 8 la_oen_mprj[112]
port 658 nsew signal input
rlabel metal2 s 160926 -400 160982 60 8 la_oen_mprj[113]
port 659 nsew signal input
rlabel metal2 s 161386 -400 161442 60 8 la_oen_mprj[114]
port 660 nsew signal input
rlabel metal2 s 161846 -400 161902 60 8 la_oen_mprj[115]
port 661 nsew signal input
rlabel metal2 s 162214 -400 162270 60 8 la_oen_mprj[116]
port 662 nsew signal input
rlabel metal2 s 162674 -400 162730 60 8 la_oen_mprj[117]
port 663 nsew signal input
rlabel metal2 s 163134 -400 163190 60 8 la_oen_mprj[118]
port 664 nsew signal input
rlabel metal2 s 163594 -400 163650 60 8 la_oen_mprj[119]
port 665 nsew signal input
rlabel metal2 s 116490 -400 116546 60 8 la_oen_mprj[11]
port 666 nsew signal input
rlabel metal2 s 163962 -400 164018 60 8 la_oen_mprj[120]
port 667 nsew signal input
rlabel metal2 s 164422 -400 164478 60 8 la_oen_mprj[121]
port 668 nsew signal input
rlabel metal2 s 164882 -400 164938 60 8 la_oen_mprj[122]
port 669 nsew signal input
rlabel metal2 s 165342 -400 165398 60 8 la_oen_mprj[123]
port 670 nsew signal input
rlabel metal2 s 165710 -400 165766 60 8 la_oen_mprj[124]
port 671 nsew signal input
rlabel metal2 s 166170 -400 166226 60 8 la_oen_mprj[125]
port 672 nsew signal input
rlabel metal2 s 166630 -400 166686 60 8 la_oen_mprj[126]
port 673 nsew signal input
rlabel metal2 s 167090 -400 167146 60 8 la_oen_mprj[127]
port 674 nsew signal input
rlabel metal2 s 116950 -400 117006 60 8 la_oen_mprj[12]
port 675 nsew signal input
rlabel metal2 s 117410 -400 117466 60 8 la_oen_mprj[13]
port 676 nsew signal input
rlabel metal2 s 117778 -400 117834 60 8 la_oen_mprj[14]
port 677 nsew signal input
rlabel metal2 s 118238 -400 118294 60 8 la_oen_mprj[15]
port 678 nsew signal input
rlabel metal2 s 118698 -400 118754 60 8 la_oen_mprj[16]
port 679 nsew signal input
rlabel metal2 s 119158 -400 119214 60 8 la_oen_mprj[17]
port 680 nsew signal input
rlabel metal2 s 119526 -400 119582 60 8 la_oen_mprj[18]
port 681 nsew signal input
rlabel metal2 s 119986 -400 120042 60 8 la_oen_mprj[19]
port 682 nsew signal input
rlabel metal2 s 112166 -400 112222 60 8 la_oen_mprj[1]
port 683 nsew signal input
rlabel metal2 s 120446 -400 120502 60 8 la_oen_mprj[20]
port 684 nsew signal input
rlabel metal2 s 120814 -400 120870 60 8 la_oen_mprj[21]
port 685 nsew signal input
rlabel metal2 s 121274 -400 121330 60 8 la_oen_mprj[22]
port 686 nsew signal input
rlabel metal2 s 121734 -400 121790 60 8 la_oen_mprj[23]
port 687 nsew signal input
rlabel metal2 s 122194 -400 122250 60 8 la_oen_mprj[24]
port 688 nsew signal input
rlabel metal2 s 122562 -400 122618 60 8 la_oen_mprj[25]
port 689 nsew signal input
rlabel metal2 s 123022 -400 123078 60 8 la_oen_mprj[26]
port 690 nsew signal input
rlabel metal2 s 123482 -400 123538 60 8 la_oen_mprj[27]
port 691 nsew signal input
rlabel metal2 s 123942 -400 123998 60 8 la_oen_mprj[28]
port 692 nsew signal input
rlabel metal2 s 124310 -400 124366 60 8 la_oen_mprj[29]
port 693 nsew signal input
rlabel metal2 s 112534 -400 112590 60 8 la_oen_mprj[2]
port 694 nsew signal input
rlabel metal2 s 124770 -400 124826 60 8 la_oen_mprj[30]
port 695 nsew signal input
rlabel metal2 s 125230 -400 125286 60 8 la_oen_mprj[31]
port 696 nsew signal input
rlabel metal2 s 125690 -400 125746 60 8 la_oen_mprj[32]
port 697 nsew signal input
rlabel metal2 s 126058 -400 126114 60 8 la_oen_mprj[33]
port 698 nsew signal input
rlabel metal2 s 126518 -400 126574 60 8 la_oen_mprj[34]
port 699 nsew signal input
rlabel metal2 s 126978 -400 127034 60 8 la_oen_mprj[35]
port 700 nsew signal input
rlabel metal2 s 127438 -400 127494 60 8 la_oen_mprj[36]
port 701 nsew signal input
rlabel metal2 s 127806 -400 127862 60 8 la_oen_mprj[37]
port 702 nsew signal input
rlabel metal2 s 128266 -400 128322 60 8 la_oen_mprj[38]
port 703 nsew signal input
rlabel metal2 s 128726 -400 128782 60 8 la_oen_mprj[39]
port 704 nsew signal input
rlabel metal2 s 112994 -400 113050 60 8 la_oen_mprj[3]
port 705 nsew signal input
rlabel metal2 s 129094 -400 129150 60 8 la_oen_mprj[40]
port 706 nsew signal input
rlabel metal2 s 129554 -400 129610 60 8 la_oen_mprj[41]
port 707 nsew signal input
rlabel metal2 s 130014 -400 130070 60 8 la_oen_mprj[42]
port 708 nsew signal input
rlabel metal2 s 130474 -400 130530 60 8 la_oen_mprj[43]
port 709 nsew signal input
rlabel metal2 s 130842 -400 130898 60 8 la_oen_mprj[44]
port 710 nsew signal input
rlabel metal2 s 131302 -400 131358 60 8 la_oen_mprj[45]
port 711 nsew signal input
rlabel metal2 s 131762 -400 131818 60 8 la_oen_mprj[46]
port 712 nsew signal input
rlabel metal2 s 132222 -400 132278 60 8 la_oen_mprj[47]
port 713 nsew signal input
rlabel metal2 s 132590 -400 132646 60 8 la_oen_mprj[48]
port 714 nsew signal input
rlabel metal2 s 133050 -400 133106 60 8 la_oen_mprj[49]
port 715 nsew signal input
rlabel metal2 s 113454 -400 113510 60 8 la_oen_mprj[4]
port 716 nsew signal input
rlabel metal2 s 133510 -400 133566 60 8 la_oen_mprj[50]
port 717 nsew signal input
rlabel metal2 s 133970 -400 134026 60 8 la_oen_mprj[51]
port 718 nsew signal input
rlabel metal2 s 134338 -400 134394 60 8 la_oen_mprj[52]
port 719 nsew signal input
rlabel metal2 s 134798 -400 134854 60 8 la_oen_mprj[53]
port 720 nsew signal input
rlabel metal2 s 135258 -400 135314 60 8 la_oen_mprj[54]
port 721 nsew signal input
rlabel metal2 s 135718 -400 135774 60 8 la_oen_mprj[55]
port 722 nsew signal input
rlabel metal2 s 136086 -400 136142 60 8 la_oen_mprj[56]
port 723 nsew signal input
rlabel metal2 s 136546 -400 136602 60 8 la_oen_mprj[57]
port 724 nsew signal input
rlabel metal2 s 137006 -400 137062 60 8 la_oen_mprj[58]
port 725 nsew signal input
rlabel metal2 s 137374 -400 137430 60 8 la_oen_mprj[59]
port 726 nsew signal input
rlabel metal2 s 113914 -400 113970 60 8 la_oen_mprj[5]
port 727 nsew signal input
rlabel metal2 s 137834 -400 137890 60 8 la_oen_mprj[60]
port 728 nsew signal input
rlabel metal2 s 138294 -400 138350 60 8 la_oen_mprj[61]
port 729 nsew signal input
rlabel metal2 s 138754 -400 138810 60 8 la_oen_mprj[62]
port 730 nsew signal input
rlabel metal2 s 139122 -400 139178 60 8 la_oen_mprj[63]
port 731 nsew signal input
rlabel metal2 s 139582 -400 139638 60 8 la_oen_mprj[64]
port 732 nsew signal input
rlabel metal2 s 140042 -400 140098 60 8 la_oen_mprj[65]
port 733 nsew signal input
rlabel metal2 s 140502 -400 140558 60 8 la_oen_mprj[66]
port 734 nsew signal input
rlabel metal2 s 140870 -400 140926 60 8 la_oen_mprj[67]
port 735 nsew signal input
rlabel metal2 s 141330 -400 141386 60 8 la_oen_mprj[68]
port 736 nsew signal input
rlabel metal2 s 141790 -400 141846 60 8 la_oen_mprj[69]
port 737 nsew signal input
rlabel metal2 s 114282 -400 114338 60 8 la_oen_mprj[6]
port 738 nsew signal input
rlabel metal2 s 142250 -400 142306 60 8 la_oen_mprj[70]
port 739 nsew signal input
rlabel metal2 s 142618 -400 142674 60 8 la_oen_mprj[71]
port 740 nsew signal input
rlabel metal2 s 143078 -400 143134 60 8 la_oen_mprj[72]
port 741 nsew signal input
rlabel metal2 s 143538 -400 143594 60 8 la_oen_mprj[73]
port 742 nsew signal input
rlabel metal2 s 143998 -400 144054 60 8 la_oen_mprj[74]
port 743 nsew signal input
rlabel metal2 s 144366 -400 144422 60 8 la_oen_mprj[75]
port 744 nsew signal input
rlabel metal2 s 144826 -400 144882 60 8 la_oen_mprj[76]
port 745 nsew signal input
rlabel metal2 s 145286 -400 145342 60 8 la_oen_mprj[77]
port 746 nsew signal input
rlabel metal2 s 145654 -400 145710 60 8 la_oen_mprj[78]
port 747 nsew signal input
rlabel metal2 s 146114 -400 146170 60 8 la_oen_mprj[79]
port 748 nsew signal input
rlabel metal2 s 114742 -400 114798 60 8 la_oen_mprj[7]
port 749 nsew signal input
rlabel metal2 s 146574 -400 146630 60 8 la_oen_mprj[80]
port 750 nsew signal input
rlabel metal2 s 147034 -400 147090 60 8 la_oen_mprj[81]
port 751 nsew signal input
rlabel metal2 s 147402 -400 147458 60 8 la_oen_mprj[82]
port 752 nsew signal input
rlabel metal2 s 147862 -400 147918 60 8 la_oen_mprj[83]
port 753 nsew signal input
rlabel metal2 s 148322 -400 148378 60 8 la_oen_mprj[84]
port 754 nsew signal input
rlabel metal2 s 148782 -400 148838 60 8 la_oen_mprj[85]
port 755 nsew signal input
rlabel metal2 s 149150 -400 149206 60 8 la_oen_mprj[86]
port 756 nsew signal input
rlabel metal2 s 149610 -400 149666 60 8 la_oen_mprj[87]
port 757 nsew signal input
rlabel metal2 s 150070 -400 150126 60 8 la_oen_mprj[88]
port 758 nsew signal input
rlabel metal2 s 150530 -400 150586 60 8 la_oen_mprj[89]
port 759 nsew signal input
rlabel metal2 s 115202 -400 115258 60 8 la_oen_mprj[8]
port 760 nsew signal input
rlabel metal2 s 150898 -400 150954 60 8 la_oen_mprj[90]
port 761 nsew signal input
rlabel metal2 s 151358 -400 151414 60 8 la_oen_mprj[91]
port 762 nsew signal input
rlabel metal2 s 151818 -400 151874 60 8 la_oen_mprj[92]
port 763 nsew signal input
rlabel metal2 s 152186 -400 152242 60 8 la_oen_mprj[93]
port 764 nsew signal input
rlabel metal2 s 152646 -400 152702 60 8 la_oen_mprj[94]
port 765 nsew signal input
rlabel metal2 s 153106 -400 153162 60 8 la_oen_mprj[95]
port 766 nsew signal input
rlabel metal2 s 153566 -400 153622 60 8 la_oen_mprj[96]
port 767 nsew signal input
rlabel metal2 s 153934 -400 153990 60 8 la_oen_mprj[97]
port 768 nsew signal input
rlabel metal2 s 154394 -400 154450 60 8 la_oen_mprj[98]
port 769 nsew signal input
rlabel metal2 s 154854 -400 154910 60 8 la_oen_mprj[99]
port 770 nsew signal input
rlabel metal2 s 115662 -400 115718 60 8 la_oen_mprj[9]
port 771 nsew signal input
rlabel metal2 s 168746 -400 168802 60 8 mprj_adr_o_core[0]
port 772 nsew signal input
rlabel metal2 s 179234 -400 179290 60 8 mprj_adr_o_core[10]
port 773 nsew signal input
rlabel metal2 s 180154 -400 180210 60 8 mprj_adr_o_core[11]
port 774 nsew signal input
rlabel metal2 s 180982 -400 181038 60 8 mprj_adr_o_core[12]
port 775 nsew signal input
rlabel metal2 s 181902 -400 181958 60 8 mprj_adr_o_core[13]
port 776 nsew signal input
rlabel metal2 s 182730 -400 182786 60 8 mprj_adr_o_core[14]
port 777 nsew signal input
rlabel metal2 s 183650 -400 183706 60 8 mprj_adr_o_core[15]
port 778 nsew signal input
rlabel metal2 s 184478 -400 184534 60 8 mprj_adr_o_core[16]
port 779 nsew signal input
rlabel metal2 s 185306 -400 185362 60 8 mprj_adr_o_core[17]
port 780 nsew signal input
rlabel metal2 s 186226 -400 186282 60 8 mprj_adr_o_core[18]
port 781 nsew signal input
rlabel metal2 s 187054 -400 187110 60 8 mprj_adr_o_core[19]
port 782 nsew signal input
rlabel metal2 s 170126 -400 170182 60 8 mprj_adr_o_core[1]
port 783 nsew signal input
rlabel metal2 s 187974 -400 188030 60 8 mprj_adr_o_core[20]
port 784 nsew signal input
rlabel metal2 s 188802 -400 188858 60 8 mprj_adr_o_core[21]
port 785 nsew signal input
rlabel metal2 s 189722 -400 189778 60 8 mprj_adr_o_core[22]
port 786 nsew signal input
rlabel metal2 s 190550 -400 190606 60 8 mprj_adr_o_core[23]
port 787 nsew signal input
rlabel metal2 s 191470 -400 191526 60 8 mprj_adr_o_core[24]
port 788 nsew signal input
rlabel metal2 s 192298 -400 192354 60 8 mprj_adr_o_core[25]
port 789 nsew signal input
rlabel metal2 s 193218 -400 193274 60 8 mprj_adr_o_core[26]
port 790 nsew signal input
rlabel metal2 s 194046 -400 194102 60 8 mprj_adr_o_core[27]
port 791 nsew signal input
rlabel metal2 s 194966 -400 195022 60 8 mprj_adr_o_core[28]
port 792 nsew signal input
rlabel metal2 s 195794 -400 195850 60 8 mprj_adr_o_core[29]
port 793 nsew signal input
rlabel metal2 s 171414 -400 171470 60 8 mprj_adr_o_core[2]
port 794 nsew signal input
rlabel metal2 s 196714 -400 196770 60 8 mprj_adr_o_core[30]
port 795 nsew signal input
rlabel metal2 s 197542 -400 197598 60 8 mprj_adr_o_core[31]
port 796 nsew signal input
rlabel metal2 s 172702 -400 172758 60 8 mprj_adr_o_core[3]
port 797 nsew signal input
rlabel metal2 s 173990 -400 174046 60 8 mprj_adr_o_core[4]
port 798 nsew signal input
rlabel metal2 s 174910 -400 174966 60 8 mprj_adr_o_core[5]
port 799 nsew signal input
rlabel metal2 s 175738 -400 175794 60 8 mprj_adr_o_core[6]
port 800 nsew signal input
rlabel metal2 s 176658 -400 176714 60 8 mprj_adr_o_core[7]
port 801 nsew signal input
rlabel metal2 s 177486 -400 177542 60 8 mprj_adr_o_core[8]
port 802 nsew signal input
rlabel metal2 s 178406 -400 178462 60 8 mprj_adr_o_core[9]
port 803 nsew signal input
rlabel metal2 s 170494 17940 170550 18400 6 mprj_adr_o_user[0]
port 804 nsew signal output
rlabel metal2 s 180982 17940 181038 18400 6 mprj_adr_o_user[10]
port 805 nsew signal output
rlabel metal2 s 181902 17940 181958 18400 6 mprj_adr_o_user[11]
port 806 nsew signal output
rlabel metal2 s 182730 17940 182786 18400 6 mprj_adr_o_user[12]
port 807 nsew signal output
rlabel metal2 s 183650 17940 183706 18400 6 mprj_adr_o_user[13]
port 808 nsew signal output
rlabel metal2 s 184478 17940 184534 18400 6 mprj_adr_o_user[14]
port 809 nsew signal output
rlabel metal2 s 185306 17940 185362 18400 6 mprj_adr_o_user[15]
port 810 nsew signal output
rlabel metal2 s 186226 17940 186282 18400 6 mprj_adr_o_user[16]
port 811 nsew signal output
rlabel metal2 s 187054 17940 187110 18400 6 mprj_adr_o_user[17]
port 812 nsew signal output
rlabel metal2 s 187974 17940 188030 18400 6 mprj_adr_o_user[18]
port 813 nsew signal output
rlabel metal2 s 188802 17940 188858 18400 6 mprj_adr_o_user[19]
port 814 nsew signal output
rlabel metal2 s 171874 17940 171930 18400 6 mprj_adr_o_user[1]
port 815 nsew signal output
rlabel metal2 s 189722 17940 189778 18400 6 mprj_adr_o_user[20]
port 816 nsew signal output
rlabel metal2 s 190550 17940 190606 18400 6 mprj_adr_o_user[21]
port 817 nsew signal output
rlabel metal2 s 191470 17940 191526 18400 6 mprj_adr_o_user[22]
port 818 nsew signal output
rlabel metal2 s 192298 17940 192354 18400 6 mprj_adr_o_user[23]
port 819 nsew signal output
rlabel metal2 s 193218 17940 193274 18400 6 mprj_adr_o_user[24]
port 820 nsew signal output
rlabel metal2 s 194046 17940 194102 18400 6 mprj_adr_o_user[25]
port 821 nsew signal output
rlabel metal2 s 194966 17940 195022 18400 6 mprj_adr_o_user[26]
port 822 nsew signal output
rlabel metal2 s 195794 17940 195850 18400 6 mprj_adr_o_user[27]
port 823 nsew signal output
rlabel metal2 s 196714 17940 196770 18400 6 mprj_adr_o_user[28]
port 824 nsew signal output
rlabel metal2 s 197542 17940 197598 18400 6 mprj_adr_o_user[29]
port 825 nsew signal output
rlabel metal2 s 173162 17940 173218 18400 6 mprj_adr_o_user[2]
port 826 nsew signal output
rlabel metal2 s 198462 17940 198518 18400 6 mprj_adr_o_user[30]
port 827 nsew signal output
rlabel metal2 s 199290 17940 199346 18400 6 mprj_adr_o_user[31]
port 828 nsew signal output
rlabel metal2 s 174450 17940 174506 18400 6 mprj_adr_o_user[3]
port 829 nsew signal output
rlabel metal2 s 175738 17940 175794 18400 6 mprj_adr_o_user[4]
port 830 nsew signal output
rlabel metal2 s 176658 17940 176714 18400 6 mprj_adr_o_user[5]
port 831 nsew signal output
rlabel metal2 s 177486 17940 177542 18400 6 mprj_adr_o_user[6]
port 832 nsew signal output
rlabel metal2 s 178406 17940 178462 18400 6 mprj_adr_o_user[7]
port 833 nsew signal output
rlabel metal2 s 179234 17940 179290 18400 6 mprj_adr_o_user[8]
port 834 nsew signal output
rlabel metal2 s 180154 17940 180210 18400 6 mprj_adr_o_user[9]
port 835 nsew signal output
rlabel metal2 s 167458 -400 167514 60 8 mprj_cyc_o_core
port 836 nsew signal input
rlabel metal2 s 169206 17940 169262 18400 6 mprj_cyc_o_user
port 837 nsew signal output
rlabel metal2 s 169206 -400 169262 60 8 mprj_dat_o_core[0]
port 838 nsew signal input
rlabel metal2 s 179694 -400 179750 60 8 mprj_dat_o_core[10]
port 839 nsew signal input
rlabel metal2 s 180522 -400 180578 60 8 mprj_dat_o_core[11]
port 840 nsew signal input
rlabel metal2 s 181442 -400 181498 60 8 mprj_dat_o_core[12]
port 841 nsew signal input
rlabel metal2 s 182270 -400 182326 60 8 mprj_dat_o_core[13]
port 842 nsew signal input
rlabel metal2 s 183190 -400 183246 60 8 mprj_dat_o_core[14]
port 843 nsew signal input
rlabel metal2 s 184018 -400 184074 60 8 mprj_dat_o_core[15]
port 844 nsew signal input
rlabel metal2 s 184938 -400 184994 60 8 mprj_dat_o_core[16]
port 845 nsew signal input
rlabel metal2 s 185766 -400 185822 60 8 mprj_dat_o_core[17]
port 846 nsew signal input
rlabel metal2 s 186686 -400 186742 60 8 mprj_dat_o_core[18]
port 847 nsew signal input
rlabel metal2 s 187514 -400 187570 60 8 mprj_dat_o_core[19]
port 848 nsew signal input
rlabel metal2 s 170494 -400 170550 60 8 mprj_dat_o_core[1]
port 849 nsew signal input
rlabel metal2 s 188434 -400 188490 60 8 mprj_dat_o_core[20]
port 850 nsew signal input
rlabel metal2 s 189262 -400 189318 60 8 mprj_dat_o_core[21]
port 851 nsew signal input
rlabel metal2 s 190182 -400 190238 60 8 mprj_dat_o_core[22]
port 852 nsew signal input
rlabel metal2 s 191010 -400 191066 60 8 mprj_dat_o_core[23]
port 853 nsew signal input
rlabel metal2 s 191930 -400 191986 60 8 mprj_dat_o_core[24]
port 854 nsew signal input
rlabel metal2 s 192758 -400 192814 60 8 mprj_dat_o_core[25]
port 855 nsew signal input
rlabel metal2 s 193586 -400 193642 60 8 mprj_dat_o_core[26]
port 856 nsew signal input
rlabel metal2 s 194506 -400 194562 60 8 mprj_dat_o_core[27]
port 857 nsew signal input
rlabel metal2 s 195334 -400 195390 60 8 mprj_dat_o_core[28]
port 858 nsew signal input
rlabel metal2 s 196254 -400 196310 60 8 mprj_dat_o_core[29]
port 859 nsew signal input
rlabel metal2 s 171874 -400 171930 60 8 mprj_dat_o_core[2]
port 860 nsew signal input
rlabel metal2 s 197082 -400 197138 60 8 mprj_dat_o_core[30]
port 861 nsew signal input
rlabel metal2 s 198002 -400 198058 60 8 mprj_dat_o_core[31]
port 862 nsew signal input
rlabel metal2 s 173162 -400 173218 60 8 mprj_dat_o_core[3]
port 863 nsew signal input
rlabel metal2 s 174450 -400 174506 60 8 mprj_dat_o_core[4]
port 864 nsew signal input
rlabel metal2 s 175370 -400 175426 60 8 mprj_dat_o_core[5]
port 865 nsew signal input
rlabel metal2 s 176198 -400 176254 60 8 mprj_dat_o_core[6]
port 866 nsew signal input
rlabel metal2 s 177026 -400 177082 60 8 mprj_dat_o_core[7]
port 867 nsew signal input
rlabel metal2 s 177946 -400 178002 60 8 mprj_dat_o_core[8]
port 868 nsew signal input
rlabel metal2 s 178774 -400 178830 60 8 mprj_dat_o_core[9]
port 869 nsew signal input
rlabel metal2 s 170954 17940 171010 18400 6 mprj_dat_o_user[0]
port 870 nsew signal output
rlabel metal2 s 181442 17940 181498 18400 6 mprj_dat_o_user[10]
port 871 nsew signal output
rlabel metal2 s 182270 17940 182326 18400 6 mprj_dat_o_user[11]
port 872 nsew signal output
rlabel metal2 s 183190 17940 183246 18400 6 mprj_dat_o_user[12]
port 873 nsew signal output
rlabel metal2 s 184018 17940 184074 18400 6 mprj_dat_o_user[13]
port 874 nsew signal output
rlabel metal2 s 184938 17940 184994 18400 6 mprj_dat_o_user[14]
port 875 nsew signal output
rlabel metal2 s 185766 17940 185822 18400 6 mprj_dat_o_user[15]
port 876 nsew signal output
rlabel metal2 s 186686 17940 186742 18400 6 mprj_dat_o_user[16]
port 877 nsew signal output
rlabel metal2 s 187514 17940 187570 18400 6 mprj_dat_o_user[17]
port 878 nsew signal output
rlabel metal2 s 188434 17940 188490 18400 6 mprj_dat_o_user[18]
port 879 nsew signal output
rlabel metal2 s 189262 17940 189318 18400 6 mprj_dat_o_user[19]
port 880 nsew signal output
rlabel metal2 s 172242 17940 172298 18400 6 mprj_dat_o_user[1]
port 881 nsew signal output
rlabel metal2 s 190182 17940 190238 18400 6 mprj_dat_o_user[20]
port 882 nsew signal output
rlabel metal2 s 191010 17940 191066 18400 6 mprj_dat_o_user[21]
port 883 nsew signal output
rlabel metal2 s 191930 17940 191986 18400 6 mprj_dat_o_user[22]
port 884 nsew signal output
rlabel metal2 s 192758 17940 192814 18400 6 mprj_dat_o_user[23]
port 885 nsew signal output
rlabel metal2 s 193586 17940 193642 18400 6 mprj_dat_o_user[24]
port 886 nsew signal output
rlabel metal2 s 194506 17940 194562 18400 6 mprj_dat_o_user[25]
port 887 nsew signal output
rlabel metal2 s 195334 17940 195390 18400 6 mprj_dat_o_user[26]
port 888 nsew signal output
rlabel metal2 s 196254 17940 196310 18400 6 mprj_dat_o_user[27]
port 889 nsew signal output
rlabel metal2 s 197082 17940 197138 18400 6 mprj_dat_o_user[28]
port 890 nsew signal output
rlabel metal2 s 198002 17940 198058 18400 6 mprj_dat_o_user[29]
port 891 nsew signal output
rlabel metal2 s 173622 17940 173678 18400 6 mprj_dat_o_user[2]
port 892 nsew signal output
rlabel metal2 s 198830 17940 198886 18400 6 mprj_dat_o_user[30]
port 893 nsew signal output
rlabel metal2 s 199750 17940 199806 18400 6 mprj_dat_o_user[31]
port 894 nsew signal output
rlabel metal2 s 174910 17940 174966 18400 6 mprj_dat_o_user[3]
port 895 nsew signal output
rlabel metal2 s 176198 17940 176254 18400 6 mprj_dat_o_user[4]
port 896 nsew signal output
rlabel metal2 s 177026 17940 177082 18400 6 mprj_dat_o_user[5]
port 897 nsew signal output
rlabel metal2 s 177946 17940 178002 18400 6 mprj_dat_o_user[6]
port 898 nsew signal output
rlabel metal2 s 178774 17940 178830 18400 6 mprj_dat_o_user[7]
port 899 nsew signal output
rlabel metal2 s 179694 17940 179750 18400 6 mprj_dat_o_user[8]
port 900 nsew signal output
rlabel metal2 s 180522 17940 180578 18400 6 mprj_dat_o_user[9]
port 901 nsew signal output
rlabel metal2 s 169666 -400 169722 60 8 mprj_sel_o_core[0]
port 902 nsew signal input
rlabel metal2 s 170954 -400 171010 60 8 mprj_sel_o_core[1]
port 903 nsew signal input
rlabel metal2 s 172242 -400 172298 60 8 mprj_sel_o_core[2]
port 904 nsew signal input
rlabel metal2 s 173622 -400 173678 60 8 mprj_sel_o_core[3]
port 905 nsew signal input
rlabel metal2 s 171414 17940 171470 18400 6 mprj_sel_o_user[0]
port 906 nsew signal output
rlabel metal2 s 172702 17940 172758 18400 6 mprj_sel_o_user[1]
port 907 nsew signal output
rlabel metal2 s 173990 17940 174046 18400 6 mprj_sel_o_user[2]
port 908 nsew signal output
rlabel metal2 s 175370 17940 175426 18400 6 mprj_sel_o_user[3]
port 909 nsew signal output
rlabel metal2 s 167918 -400 167974 60 8 mprj_stb_o_core
port 910 nsew signal input
rlabel metal2 s 169666 17940 169722 18400 6 mprj_stb_o_user
port 911 nsew signal output
rlabel metal2 s 168378 -400 168434 60 8 mprj_we_o_core
port 912 nsew signal input
rlabel metal2 s 170126 17940 170182 18400 6 mprj_we_o_user
port 913 nsew signal output
rlabel metal2 s 198462 -400 198518 60 8 user1_vcc_powergood
port 914 nsew signal output
rlabel metal2 s 198830 -400 198886 60 8 user1_vdd_powergood
port 915 nsew signal output
rlabel metal2 s 199290 -400 199346 60 8 user2_vcc_powergood
port 916 nsew signal output
rlabel metal2 s 199750 -400 199806 60 8 user2_vdd_powergood
port 917 nsew signal output
rlabel metal2 s 202 17940 258 18400 6 user_clock
port 918 nsew signal output
rlabel metal2 s 570 17940 626 18400 6 user_clock2
port 919 nsew signal output
rlabel metal2 s 1030 17940 1086 18400 6 user_reset
port 920 nsew signal output
rlabel metal2 s 1490 17940 1546 18400 6 user_resetn
port 921 nsew signal output
rlabel metal4 s 200122 -402 200302 18354 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 184014 -666 184194 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 154014 -666 154194 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 124014 -666 124194 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 94014 -666 94194 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 64014 -666 64194 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 34014 -666 34194 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 4014 -666 4194 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 184014 17940 184194 18618 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 154014 17940 154194 18618 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 124014 17940 124194 18618 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 94014 17940 94194 18618 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 64014 17940 64194 18618 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 34014 17940 34194 18618 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 4014 17940 4194 18618 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s -386 -402 -206 18354 4 vccd
port 922 nsew power bidirectional
rlabel via3 s 200220 -384 200284 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 200140 -384 200204 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 184112 -384 184176 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 184032 -384 184096 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 154112 -384 154176 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 154032 -384 154096 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 124112 -384 124176 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 124032 -384 124096 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 94112 -384 94176 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 94032 -384 94096 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 64112 -384 64176 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 64032 -384 64096 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 34112 -384 34176 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 34032 -384 34096 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 4112 -384 4176 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 4032 -384 4096 -320 8 vccd
port 922 nsew power bidirectional
rlabel via3 s -288 -384 -224 -320 2 vccd
port 922 nsew power bidirectional
rlabel via3 s -368 -384 -304 -320 2 vccd
port 922 nsew power bidirectional
rlabel via3 s 200220 -304 200284 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 200140 -304 200204 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 184112 -304 184176 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 184032 -304 184096 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 154112 -304 154176 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 154032 -304 154096 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 124112 -304 124176 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 124032 -304 124096 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 94112 -304 94176 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 94032 -304 94096 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 64112 -304 64176 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 64032 -304 64096 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 34112 -304 34176 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 34032 -304 34096 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 4112 -304 4176 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 4032 -304 4096 -240 8 vccd
port 922 nsew power bidirectional
rlabel via3 s -288 -304 -224 -240 2 vccd
port 922 nsew power bidirectional
rlabel via3 s -368 -304 -304 -240 2 vccd
port 922 nsew power bidirectional
rlabel via3 s 200220 18192 200284 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 200140 18192 200204 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 184112 18192 184176 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 184032 18192 184096 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 154112 18192 154176 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 154032 18192 154096 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 124112 18192 124176 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 124032 18192 124096 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 94112 18192 94176 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 94032 18192 94096 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 64112 18192 64176 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 64032 18192 64096 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 34112 18192 34176 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 34032 18192 34096 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 4112 18192 4176 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 4032 18192 4096 18256 6 vccd
port 922 nsew power bidirectional
rlabel via3 s -288 18192 -224 18256 4 vccd
port 922 nsew power bidirectional
rlabel via3 s -368 18192 -304 18256 4 vccd
port 922 nsew power bidirectional
rlabel via3 s 200220 18272 200284 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 200140 18272 200204 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 184112 18272 184176 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 184032 18272 184096 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 154112 18272 154176 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 154032 18272 154096 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 124112 18272 124176 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 124032 18272 124096 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 94112 18272 94176 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 94032 18272 94096 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 64112 18272 64176 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 64032 18272 64096 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 34112 18272 34176 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 34032 18272 34096 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 4112 18272 4176 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 4032 18272 4096 18336 6 vccd
port 922 nsew power bidirectional
rlabel via3 s -288 18272 -224 18336 4 vccd
port 922 nsew power bidirectional
rlabel via3 s -368 18272 -304 18336 4 vccd
port 922 nsew power bidirectional
rlabel metal3 s -386 -402 200302 -222 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s -386 18174 200302 18354 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 200386 -666 200566 18618 6 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 169014 -666 169194 60 8 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 139014 -666 139194 60 8 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 109014 -666 109194 60 8 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 79014 -666 79194 60 8 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 49014 -666 49194 60 8 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 19014 -666 19194 60 8 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 169014 17940 169194 18618 6 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 139014 17940 139194 18618 6 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 109014 17940 109194 18618 6 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 79014 17940 79194 18618 6 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 49014 17940 49194 18618 6 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 19014 17940 19194 18618 6 vssd
port 923 nsew ground bidirectional
rlabel metal4 s -650 -666 -470 18618 4 vssd
port 923 nsew ground bidirectional
rlabel via3 s 200484 -648 200548 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 200404 -648 200468 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 169112 -648 169176 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 169032 -648 169096 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 139112 -648 139176 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 139032 -648 139096 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 109112 -648 109176 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 109032 -648 109096 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 79112 -648 79176 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 79032 -648 79096 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 49112 -648 49176 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 49032 -648 49096 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 19112 -648 19176 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 19032 -648 19096 -584 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s -552 -648 -488 -584 2 vssd
port 923 nsew ground bidirectional
rlabel via3 s -632 -648 -568 -584 2 vssd
port 923 nsew ground bidirectional
rlabel via3 s 200484 -568 200548 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 200404 -568 200468 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 169112 -568 169176 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 169032 -568 169096 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 139112 -568 139176 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 139032 -568 139096 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 109112 -568 109176 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 109032 -568 109096 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 79112 -568 79176 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 79032 -568 79096 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 49112 -568 49176 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 49032 -568 49096 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 19112 -568 19176 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s 19032 -568 19096 -504 8 vssd
port 923 nsew ground bidirectional
rlabel via3 s -552 -568 -488 -504 2 vssd
port 923 nsew ground bidirectional
rlabel via3 s -632 -568 -568 -504 2 vssd
port 923 nsew ground bidirectional
rlabel via3 s 200484 18456 200548 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 200404 18456 200468 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 169112 18456 169176 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 169032 18456 169096 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 139112 18456 139176 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 139032 18456 139096 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 109112 18456 109176 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 109032 18456 109096 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 79112 18456 79176 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 79032 18456 79096 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 49112 18456 49176 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 49032 18456 49096 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 19112 18456 19176 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 19032 18456 19096 18520 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s -552 18456 -488 18520 4 vssd
port 923 nsew ground bidirectional
rlabel via3 s -632 18456 -568 18520 4 vssd
port 923 nsew ground bidirectional
rlabel via3 s 200484 18536 200548 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 200404 18536 200468 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 169112 18536 169176 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 169032 18536 169096 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 139112 18536 139176 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 139032 18536 139096 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 109112 18536 109176 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 109032 18536 109096 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 79112 18536 79176 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 79032 18536 79096 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 49112 18536 49176 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 49032 18536 49096 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 19112 18536 19176 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s 19032 18536 19096 18600 6 vssd
port 923 nsew ground bidirectional
rlabel via3 s -552 18536 -488 18600 4 vssd
port 923 nsew ground bidirectional
rlabel via3 s -632 18536 -568 18600 4 vssd
port 923 nsew ground bidirectional
rlabel metal3 s -650 -666 200566 -486 8 vssd
port 923 nsew ground bidirectional
rlabel metal3 s -650 18438 200566 18618 6 vssd
port 923 nsew ground bidirectional
rlabel metal4 s 200650 -930 200830 18882 6 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 184834 -1194 185014 60 8 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 154834 -1194 155014 60 8 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 124834 -1194 125014 60 8 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 94834 -1194 95014 60 8 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 64834 -1194 65014 60 8 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 34834 -1194 35014 60 8 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 4834 -1194 5014 60 8 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 184834 17940 185014 19146 6 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 154834 17940 155014 19146 6 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 124834 17940 125014 19146 6 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 94834 17940 95014 19146 6 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 64834 17940 65014 19146 6 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 34834 17940 35014 19146 6 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 4834 17940 5014 19146 6 vccd1
port 924 nsew power bidirectional
rlabel metal4 s -914 -930 -734 18882 4 vccd1
port 924 nsew power bidirectional
rlabel via3 s 200748 -912 200812 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 200668 -912 200732 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 184932 -912 184996 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 184852 -912 184916 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 154932 -912 154996 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 154852 -912 154916 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 124932 -912 124996 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 124852 -912 124916 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 94932 -912 94996 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 94852 -912 94916 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 64932 -912 64996 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 64852 -912 64916 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 34932 -912 34996 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 34852 -912 34916 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 4932 -912 4996 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 4852 -912 4916 -848 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s -816 -912 -752 -848 2 vccd1
port 924 nsew power bidirectional
rlabel via3 s -896 -912 -832 -848 2 vccd1
port 924 nsew power bidirectional
rlabel via3 s 200748 -832 200812 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 200668 -832 200732 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 184932 -832 184996 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 184852 -832 184916 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 154932 -832 154996 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 154852 -832 154916 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 124932 -832 124996 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 124852 -832 124916 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 94932 -832 94996 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 94852 -832 94916 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 64932 -832 64996 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 64852 -832 64916 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 34932 -832 34996 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 34852 -832 34916 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 4932 -832 4996 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s 4852 -832 4916 -768 8 vccd1
port 924 nsew power bidirectional
rlabel via3 s -816 -832 -752 -768 2 vccd1
port 924 nsew power bidirectional
rlabel via3 s -896 -832 -832 -768 2 vccd1
port 924 nsew power bidirectional
rlabel via3 s 200748 18720 200812 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 200668 18720 200732 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 184932 18720 184996 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 184852 18720 184916 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 154932 18720 154996 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 154852 18720 154916 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 124932 18720 124996 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 124852 18720 124916 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 94932 18720 94996 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 94852 18720 94916 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 64932 18720 64996 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 64852 18720 64916 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 34932 18720 34996 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 34852 18720 34916 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 4932 18720 4996 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 4852 18720 4916 18784 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s -816 18720 -752 18784 4 vccd1
port 924 nsew power bidirectional
rlabel via3 s -896 18720 -832 18784 4 vccd1
port 924 nsew power bidirectional
rlabel via3 s 200748 18800 200812 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 200668 18800 200732 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 184932 18800 184996 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 184852 18800 184916 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 154932 18800 154996 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 154852 18800 154916 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 124932 18800 124996 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 124852 18800 124916 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 94932 18800 94996 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 94852 18800 94916 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 64932 18800 64996 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 64852 18800 64916 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 34932 18800 34996 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 34852 18800 34916 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 4932 18800 4996 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s 4852 18800 4916 18864 6 vccd1
port 924 nsew power bidirectional
rlabel via3 s -816 18800 -752 18864 4 vccd1
port 924 nsew power bidirectional
rlabel via3 s -896 18800 -832 18864 4 vccd1
port 924 nsew power bidirectional
rlabel metal3 s -914 -930 200830 -750 8 vccd1
port 924 nsew power bidirectional
rlabel metal3 s -914 18702 200830 18882 6 vccd1
port 924 nsew power bidirectional
rlabel metal4 s 200914 -1194 201094 19146 6 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 169834 -1194 170014 60 8 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 139834 -1194 140014 60 8 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 109834 -1194 110014 60 8 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 79834 -1194 80014 60 8 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 49834 -1194 50014 60 8 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 19834 -1194 20014 60 8 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 169834 17940 170014 19146 6 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 139834 17940 140014 19146 6 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 109834 17940 110014 19146 6 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 79834 17940 80014 19146 6 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 49834 17940 50014 19146 6 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 19834 17940 20014 19146 6 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s -1178 -1194 -998 19146 4 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 201012 -1176 201076 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 200932 -1176 200996 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 169932 -1176 169996 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 169852 -1176 169916 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 139932 -1176 139996 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 139852 -1176 139916 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 109932 -1176 109996 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 109852 -1176 109916 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 79932 -1176 79996 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 79852 -1176 79916 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 49932 -1176 49996 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 49852 -1176 49916 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 19932 -1176 19996 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 19852 -1176 19916 -1112 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s -1080 -1176 -1016 -1112 2 vssd1
port 925 nsew ground bidirectional
rlabel via3 s -1160 -1176 -1096 -1112 2 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 201012 -1096 201076 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 200932 -1096 200996 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 169932 -1096 169996 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 169852 -1096 169916 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 139932 -1096 139996 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 139852 -1096 139916 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 109932 -1096 109996 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 109852 -1096 109916 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 79932 -1096 79996 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 79852 -1096 79916 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 49932 -1096 49996 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 49852 -1096 49916 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 19932 -1096 19996 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 19852 -1096 19916 -1032 8 vssd1
port 925 nsew ground bidirectional
rlabel via3 s -1080 -1096 -1016 -1032 2 vssd1
port 925 nsew ground bidirectional
rlabel via3 s -1160 -1096 -1096 -1032 2 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 201012 18984 201076 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 200932 18984 200996 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 169932 18984 169996 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 169852 18984 169916 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 139932 18984 139996 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 139852 18984 139916 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 109932 18984 109996 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 109852 18984 109916 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 79932 18984 79996 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 79852 18984 79916 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 49932 18984 49996 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 49852 18984 49916 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 19932 18984 19996 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 19852 18984 19916 19048 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s -1080 18984 -1016 19048 4 vssd1
port 925 nsew ground bidirectional
rlabel via3 s -1160 18984 -1096 19048 4 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 201012 19064 201076 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 200932 19064 200996 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 169932 19064 169996 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 169852 19064 169916 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 139932 19064 139996 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 139852 19064 139916 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 109932 19064 109996 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 109852 19064 109916 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 79932 19064 79996 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 79852 19064 79916 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 49932 19064 49996 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 49852 19064 49916 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 19932 19064 19996 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s 19852 19064 19916 19128 6 vssd1
port 925 nsew ground bidirectional
rlabel via3 s -1080 19064 -1016 19128 4 vssd1
port 925 nsew ground bidirectional
rlabel via3 s -1160 19064 -1096 19128 4 vssd1
port 925 nsew ground bidirectional
rlabel metal3 s -1178 -1194 201094 -1014 8 vssd1
port 925 nsew ground bidirectional
rlabel metal3 s -1178 18966 201094 19146 6 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 201178 -1458 201358 19410 6 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 185654 -1722 185834 60 8 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 155654 -1722 155834 60 8 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 125654 -1722 125834 60 8 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 95654 -1722 95834 60 8 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 65654 -1722 65834 60 8 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 35654 -1722 35834 60 8 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 5654 -1722 5834 60 8 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 185654 17940 185834 19674 6 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 155654 17940 155834 19674 6 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 125654 17940 125834 19674 6 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 95654 17940 95834 19674 6 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 65654 17940 65834 19674 6 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 35654 17940 35834 19674 6 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 5654 17940 5834 19674 6 vccd2
port 926 nsew power bidirectional
rlabel metal4 s -1442 -1458 -1262 19410 4 vccd2
port 926 nsew power bidirectional
rlabel via3 s 201276 -1440 201340 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 201196 -1440 201260 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 185752 -1440 185816 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 185672 -1440 185736 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 155752 -1440 155816 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 155672 -1440 155736 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 125752 -1440 125816 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 125672 -1440 125736 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 95752 -1440 95816 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 95672 -1440 95736 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 65752 -1440 65816 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 65672 -1440 65736 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 35752 -1440 35816 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 35672 -1440 35736 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 5752 -1440 5816 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 5672 -1440 5736 -1376 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s -1344 -1440 -1280 -1376 2 vccd2
port 926 nsew power bidirectional
rlabel via3 s -1424 -1440 -1360 -1376 2 vccd2
port 926 nsew power bidirectional
rlabel via3 s 201276 -1360 201340 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 201196 -1360 201260 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 185752 -1360 185816 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 185672 -1360 185736 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 155752 -1360 155816 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 155672 -1360 155736 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 125752 -1360 125816 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 125672 -1360 125736 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 95752 -1360 95816 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 95672 -1360 95736 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 65752 -1360 65816 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 65672 -1360 65736 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 35752 -1360 35816 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 35672 -1360 35736 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 5752 -1360 5816 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s 5672 -1360 5736 -1296 8 vccd2
port 926 nsew power bidirectional
rlabel via3 s -1344 -1360 -1280 -1296 2 vccd2
port 926 nsew power bidirectional
rlabel via3 s -1424 -1360 -1360 -1296 2 vccd2
port 926 nsew power bidirectional
rlabel via3 s 201276 19248 201340 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 201196 19248 201260 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 185752 19248 185816 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 185672 19248 185736 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 155752 19248 155816 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 155672 19248 155736 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 125752 19248 125816 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 125672 19248 125736 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 95752 19248 95816 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 95672 19248 95736 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 65752 19248 65816 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 65672 19248 65736 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 35752 19248 35816 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 35672 19248 35736 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 5752 19248 5816 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 5672 19248 5736 19312 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s -1344 19248 -1280 19312 4 vccd2
port 926 nsew power bidirectional
rlabel via3 s -1424 19248 -1360 19312 4 vccd2
port 926 nsew power bidirectional
rlabel via3 s 201276 19328 201340 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 201196 19328 201260 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 185752 19328 185816 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 185672 19328 185736 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 155752 19328 155816 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 155672 19328 155736 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 125752 19328 125816 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 125672 19328 125736 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 95752 19328 95816 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 95672 19328 95736 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 65752 19328 65816 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 65672 19328 65736 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 35752 19328 35816 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 35672 19328 35736 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 5752 19328 5816 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s 5672 19328 5736 19392 6 vccd2
port 926 nsew power bidirectional
rlabel via3 s -1344 19328 -1280 19392 4 vccd2
port 926 nsew power bidirectional
rlabel via3 s -1424 19328 -1360 19392 4 vccd2
port 926 nsew power bidirectional
rlabel metal3 s -1442 -1458 201358 -1278 8 vccd2
port 926 nsew power bidirectional
rlabel metal3 s -1442 19230 201358 19410 6 vccd2
port 926 nsew power bidirectional
rlabel metal4 s 201442 -1722 201622 19674 6 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 170654 -1722 170834 60 8 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 140654 -1722 140834 60 8 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 110654 -1722 110834 60 8 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 80654 -1722 80834 60 8 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 50654 -1722 50834 60 8 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 20654 -1722 20834 60 8 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 170654 17940 170834 19674 6 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 140654 17940 140834 19674 6 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 110654 17940 110834 19674 6 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 80654 17940 80834 19674 6 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 50654 17940 50834 19674 6 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 20654 17940 20834 19674 6 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s -1706 -1722 -1526 19674 4 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 201540 -1704 201604 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 201460 -1704 201524 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 170752 -1704 170816 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 170672 -1704 170736 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 140752 -1704 140816 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 140672 -1704 140736 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 110752 -1704 110816 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 110672 -1704 110736 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 80752 -1704 80816 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 80672 -1704 80736 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 50752 -1704 50816 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 50672 -1704 50736 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 20752 -1704 20816 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 20672 -1704 20736 -1640 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s -1608 -1704 -1544 -1640 2 vssd2
port 927 nsew ground bidirectional
rlabel via3 s -1688 -1704 -1624 -1640 2 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 201540 -1624 201604 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 201460 -1624 201524 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 170752 -1624 170816 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 170672 -1624 170736 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 140752 -1624 140816 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 140672 -1624 140736 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 110752 -1624 110816 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 110672 -1624 110736 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 80752 -1624 80816 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 80672 -1624 80736 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 50752 -1624 50816 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 50672 -1624 50736 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 20752 -1624 20816 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 20672 -1624 20736 -1560 8 vssd2
port 927 nsew ground bidirectional
rlabel via3 s -1608 -1624 -1544 -1560 2 vssd2
port 927 nsew ground bidirectional
rlabel via3 s -1688 -1624 -1624 -1560 2 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 201540 19512 201604 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 201460 19512 201524 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 170752 19512 170816 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 170672 19512 170736 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 140752 19512 140816 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 140672 19512 140736 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 110752 19512 110816 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 110672 19512 110736 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 80752 19512 80816 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 80672 19512 80736 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 50752 19512 50816 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 50672 19512 50736 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 20752 19512 20816 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 20672 19512 20736 19576 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s -1608 19512 -1544 19576 4 vssd2
port 927 nsew ground bidirectional
rlabel via3 s -1688 19512 -1624 19576 4 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 201540 19592 201604 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 201460 19592 201524 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 170752 19592 170816 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 170672 19592 170736 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 140752 19592 140816 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 140672 19592 140736 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 110752 19592 110816 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 110672 19592 110736 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 80752 19592 80816 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 80672 19592 80736 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 50752 19592 50816 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 50672 19592 50736 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 20752 19592 20816 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s 20672 19592 20736 19656 6 vssd2
port 927 nsew ground bidirectional
rlabel via3 s -1608 19592 -1544 19656 4 vssd2
port 927 nsew ground bidirectional
rlabel via3 s -1688 19592 -1624 19656 4 vssd2
port 927 nsew ground bidirectional
rlabel metal3 s -1706 -1722 201622 -1542 8 vssd2
port 927 nsew ground bidirectional
rlabel metal3 s -1706 19494 201622 19674 6 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 201706 -1986 201886 19938 6 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 186474 -2250 186654 60 8 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 156474 -2250 156654 60 8 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 126474 -2250 126654 60 8 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 96474 -2250 96654 60 8 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 66474 -2250 66654 60 8 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 36474 -2250 36654 60 8 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 6474 -2250 6654 60 8 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 186474 17940 186654 20202 6 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 156474 17940 156654 20202 6 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 126474 17940 126654 20202 6 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 96474 17940 96654 20202 6 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 66474 17940 66654 20202 6 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 36474 17940 36654 20202 6 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 6474 17940 6654 20202 6 vdda1
port 928 nsew power bidirectional
rlabel metal4 s -1970 -1986 -1790 19938 4 vdda1
port 928 nsew power bidirectional
rlabel via3 s 201804 -1968 201868 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 201724 -1968 201788 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 186572 -1968 186636 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 186492 -1968 186556 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 156572 -1968 156636 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 156492 -1968 156556 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 126572 -1968 126636 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 126492 -1968 126556 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 96572 -1968 96636 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 96492 -1968 96556 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 66572 -1968 66636 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 66492 -1968 66556 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 36572 -1968 36636 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 36492 -1968 36556 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 6572 -1968 6636 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 6492 -1968 6556 -1904 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s -1872 -1968 -1808 -1904 2 vdda1
port 928 nsew power bidirectional
rlabel via3 s -1952 -1968 -1888 -1904 2 vdda1
port 928 nsew power bidirectional
rlabel via3 s 201804 -1888 201868 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 201724 -1888 201788 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 186572 -1888 186636 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 186492 -1888 186556 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 156572 -1888 156636 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 156492 -1888 156556 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 126572 -1888 126636 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 126492 -1888 126556 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 96572 -1888 96636 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 96492 -1888 96556 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 66572 -1888 66636 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 66492 -1888 66556 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 36572 -1888 36636 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 36492 -1888 36556 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 6572 -1888 6636 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s 6492 -1888 6556 -1824 8 vdda1
port 928 nsew power bidirectional
rlabel via3 s -1872 -1888 -1808 -1824 2 vdda1
port 928 nsew power bidirectional
rlabel via3 s -1952 -1888 -1888 -1824 2 vdda1
port 928 nsew power bidirectional
rlabel via3 s 201804 19776 201868 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 201724 19776 201788 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 186572 19776 186636 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 186492 19776 186556 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 156572 19776 156636 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 156492 19776 156556 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 126572 19776 126636 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 126492 19776 126556 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 96572 19776 96636 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 96492 19776 96556 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 66572 19776 66636 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 66492 19776 66556 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 36572 19776 36636 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 36492 19776 36556 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 6572 19776 6636 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 6492 19776 6556 19840 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s -1872 19776 -1808 19840 4 vdda1
port 928 nsew power bidirectional
rlabel via3 s -1952 19776 -1888 19840 4 vdda1
port 928 nsew power bidirectional
rlabel via3 s 201804 19856 201868 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 201724 19856 201788 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 186572 19856 186636 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 186492 19856 186556 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 156572 19856 156636 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 156492 19856 156556 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 126572 19856 126636 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 126492 19856 126556 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 96572 19856 96636 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 96492 19856 96556 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 66572 19856 66636 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 66492 19856 66556 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 36572 19856 36636 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 36492 19856 36556 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 6572 19856 6636 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s 6492 19856 6556 19920 6 vdda1
port 928 nsew power bidirectional
rlabel via3 s -1872 19856 -1808 19920 4 vdda1
port 928 nsew power bidirectional
rlabel via3 s -1952 19856 -1888 19920 4 vdda1
port 928 nsew power bidirectional
rlabel metal3 s -1970 -1986 201886 -1806 8 vdda1
port 928 nsew power bidirectional
rlabel metal3 s -1970 19758 201886 19938 6 vdda1
port 928 nsew power bidirectional
rlabel metal4 s 201970 -2250 202150 20202 6 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 171474 -2250 171654 60 8 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 141474 -2250 141654 60 8 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 111474 -2250 111654 60 8 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 81474 -2250 81654 60 8 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 51474 -2250 51654 60 8 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 21474 -2250 21654 60 8 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 171474 17940 171654 20202 6 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 141474 17940 141654 20202 6 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 111474 17940 111654 20202 6 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 81474 17940 81654 20202 6 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 51474 17940 51654 20202 6 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 21474 17940 21654 20202 6 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s -2234 -2250 -2054 20202 4 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 202068 -2232 202132 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 201988 -2232 202052 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 171572 -2232 171636 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 171492 -2232 171556 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 141572 -2232 141636 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 141492 -2232 141556 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 111572 -2232 111636 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 111492 -2232 111556 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 81572 -2232 81636 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 81492 -2232 81556 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 51572 -2232 51636 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 51492 -2232 51556 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 21572 -2232 21636 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 21492 -2232 21556 -2168 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s -2136 -2232 -2072 -2168 2 vssa1
port 929 nsew ground bidirectional
rlabel via3 s -2216 -2232 -2152 -2168 2 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 202068 -2152 202132 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 201988 -2152 202052 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 171572 -2152 171636 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 171492 -2152 171556 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 141572 -2152 141636 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 141492 -2152 141556 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 111572 -2152 111636 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 111492 -2152 111556 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 81572 -2152 81636 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 81492 -2152 81556 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 51572 -2152 51636 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 51492 -2152 51556 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 21572 -2152 21636 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 21492 -2152 21556 -2088 8 vssa1
port 929 nsew ground bidirectional
rlabel via3 s -2136 -2152 -2072 -2088 2 vssa1
port 929 nsew ground bidirectional
rlabel via3 s -2216 -2152 -2152 -2088 2 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 202068 20040 202132 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 201988 20040 202052 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 171572 20040 171636 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 171492 20040 171556 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 141572 20040 141636 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 141492 20040 141556 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 111572 20040 111636 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 111492 20040 111556 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 81572 20040 81636 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 81492 20040 81556 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 51572 20040 51636 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 51492 20040 51556 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 21572 20040 21636 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 21492 20040 21556 20104 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s -2136 20040 -2072 20104 4 vssa1
port 929 nsew ground bidirectional
rlabel via3 s -2216 20040 -2152 20104 4 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 202068 20120 202132 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 201988 20120 202052 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 171572 20120 171636 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 171492 20120 171556 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 141572 20120 141636 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 141492 20120 141556 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 111572 20120 111636 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 111492 20120 111556 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 81572 20120 81636 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 81492 20120 81556 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 51572 20120 51636 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 51492 20120 51556 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 21572 20120 21636 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s 21492 20120 21556 20184 6 vssa1
port 929 nsew ground bidirectional
rlabel via3 s -2136 20120 -2072 20184 4 vssa1
port 929 nsew ground bidirectional
rlabel via3 s -2216 20120 -2152 20184 4 vssa1
port 929 nsew ground bidirectional
rlabel metal3 s -2234 -2250 202150 -2070 8 vssa1
port 929 nsew ground bidirectional
rlabel metal3 s -2234 20022 202150 20202 6 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 202234 -2514 202414 20466 6 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 187294 -2778 187474 60 8 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 157294 -2778 157474 60 8 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 127294 -2778 127474 60 8 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 97294 -2778 97474 60 8 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 67294 -2778 67474 60 8 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 37294 -2778 37474 60 8 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 7294 -2778 7474 60 8 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 187294 17940 187474 20730 6 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 157294 17940 157474 20730 6 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 127294 17940 127474 20730 6 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 97294 17940 97474 20730 6 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 67294 17940 67474 20730 6 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 37294 17940 37474 20730 6 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 7294 17940 7474 20730 6 vdda2
port 930 nsew power bidirectional
rlabel metal4 s -2498 -2514 -2318 20466 4 vdda2
port 930 nsew power bidirectional
rlabel via3 s 202332 -2496 202396 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 202252 -2496 202316 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 187392 -2496 187456 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 187312 -2496 187376 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 157392 -2496 157456 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 157312 -2496 157376 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 127392 -2496 127456 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 127312 -2496 127376 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 97392 -2496 97456 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 97312 -2496 97376 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 67392 -2496 67456 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 67312 -2496 67376 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 37392 -2496 37456 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 37312 -2496 37376 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 7392 -2496 7456 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 7312 -2496 7376 -2432 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s -2400 -2496 -2336 -2432 2 vdda2
port 930 nsew power bidirectional
rlabel via3 s -2480 -2496 -2416 -2432 2 vdda2
port 930 nsew power bidirectional
rlabel via3 s 202332 -2416 202396 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 202252 -2416 202316 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 187392 -2416 187456 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 187312 -2416 187376 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 157392 -2416 157456 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 157312 -2416 157376 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 127392 -2416 127456 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 127312 -2416 127376 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 97392 -2416 97456 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 97312 -2416 97376 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 67392 -2416 67456 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 67312 -2416 67376 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 37392 -2416 37456 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 37312 -2416 37376 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 7392 -2416 7456 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s 7312 -2416 7376 -2352 8 vdda2
port 930 nsew power bidirectional
rlabel via3 s -2400 -2416 -2336 -2352 2 vdda2
port 930 nsew power bidirectional
rlabel via3 s -2480 -2416 -2416 -2352 2 vdda2
port 930 nsew power bidirectional
rlabel via3 s 202332 20304 202396 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 202252 20304 202316 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 187392 20304 187456 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 187312 20304 187376 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 157392 20304 157456 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 157312 20304 157376 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 127392 20304 127456 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 127312 20304 127376 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 97392 20304 97456 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 97312 20304 97376 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 67392 20304 67456 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 67312 20304 67376 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 37392 20304 37456 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 37312 20304 37376 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 7392 20304 7456 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 7312 20304 7376 20368 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s -2400 20304 -2336 20368 4 vdda2
port 930 nsew power bidirectional
rlabel via3 s -2480 20304 -2416 20368 4 vdda2
port 930 nsew power bidirectional
rlabel via3 s 202332 20384 202396 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 202252 20384 202316 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 187392 20384 187456 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 187312 20384 187376 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 157392 20384 157456 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 157312 20384 157376 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 127392 20384 127456 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 127312 20384 127376 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 97392 20384 97456 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 97312 20384 97376 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 67392 20384 67456 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 67312 20384 67376 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 37392 20384 37456 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 37312 20384 37376 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 7392 20384 7456 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s 7312 20384 7376 20448 6 vdda2
port 930 nsew power bidirectional
rlabel via3 s -2400 20384 -2336 20448 4 vdda2
port 930 nsew power bidirectional
rlabel via3 s -2480 20384 -2416 20448 4 vdda2
port 930 nsew power bidirectional
rlabel metal3 s -2498 -2514 202414 -2334 8 vdda2
port 930 nsew power bidirectional
rlabel metal3 s -2498 20286 202414 20466 6 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 202498 -2778 202678 20730 6 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 172294 -2778 172474 60 8 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 142294 -2778 142474 60 8 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 112294 -2778 112474 60 8 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 82294 -2778 82474 60 8 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 52294 -2778 52474 60 8 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 22294 -2778 22474 60 8 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 172294 17940 172474 20730 6 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 142294 17940 142474 20730 6 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 112294 17940 112474 20730 6 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 82294 17940 82474 20730 6 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 52294 17940 52474 20730 6 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 22294 17940 22474 20730 6 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s -2762 -2778 -2582 20730 4 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 202596 -2760 202660 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 202516 -2760 202580 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 172392 -2760 172456 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 172312 -2760 172376 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 142392 -2760 142456 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 142312 -2760 142376 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 112392 -2760 112456 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 112312 -2760 112376 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 82392 -2760 82456 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 82312 -2760 82376 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 52392 -2760 52456 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 52312 -2760 52376 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 22392 -2760 22456 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 22312 -2760 22376 -2696 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s -2664 -2760 -2600 -2696 2 vssa2
port 931 nsew ground bidirectional
rlabel via3 s -2744 -2760 -2680 -2696 2 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 202596 -2680 202660 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 202516 -2680 202580 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 172392 -2680 172456 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 172312 -2680 172376 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 142392 -2680 142456 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 142312 -2680 142376 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 112392 -2680 112456 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 112312 -2680 112376 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 82392 -2680 82456 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 82312 -2680 82376 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 52392 -2680 52456 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 52312 -2680 52376 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 22392 -2680 22456 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 22312 -2680 22376 -2616 8 vssa2
port 931 nsew ground bidirectional
rlabel via3 s -2664 -2680 -2600 -2616 2 vssa2
port 931 nsew ground bidirectional
rlabel via3 s -2744 -2680 -2680 -2616 2 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 202596 20568 202660 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 202516 20568 202580 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 172392 20568 172456 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 172312 20568 172376 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 142392 20568 142456 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 142312 20568 142376 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 112392 20568 112456 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 112312 20568 112376 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 82392 20568 82456 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 82312 20568 82376 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 52392 20568 52456 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 52312 20568 52376 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 22392 20568 22456 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 22312 20568 22376 20632 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s -2664 20568 -2600 20632 4 vssa2
port 931 nsew ground bidirectional
rlabel via3 s -2744 20568 -2680 20632 4 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 202596 20648 202660 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 202516 20648 202580 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 172392 20648 172456 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 172312 20648 172376 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 142392 20648 142456 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 142312 20648 142376 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 112392 20648 112456 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 112312 20648 112376 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 82392 20648 82456 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 82312 20648 82376 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 52392 20648 52456 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 52312 20648 52376 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 22392 20648 22456 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s 22312 20648 22376 20712 6 vssa2
port 931 nsew ground bidirectional
rlabel via3 s -2664 20648 -2600 20712 4 vssa2
port 931 nsew ground bidirectional
rlabel via3 s -2744 20648 -2680 20712 4 vssa2
port 931 nsew ground bidirectional
rlabel metal3 s -2762 -2778 202678 -2598 8 vssa2
port 931 nsew ground bidirectional
rlabel metal3 s -2762 20550 202678 20730 6 vssa2
port 931 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 200000 18000
string LEFview TRUE
<< end >>
