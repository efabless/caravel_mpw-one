magic
tech sky130A
magscale 1 2
timestamp 1624759901
<< error_p >>
rect 13273 237181 17273 237186
rect 12953 236861 17593 236866
rect 625657 236228 629657 236246
rect 625337 235908 629977 235926
<< metal3 >>
rect 537138 958512 541918 958985
rect 537138 956582 537238 958512
rect 541806 956582 541918 958512
rect 537138 956486 541918 956582
rect 547117 958490 551897 958978
rect 547117 956560 547188 958490
rect 551756 956560 551897 958490
rect 547117 956479 551897 956560
rect 781 888076 17286 888232
rect 781 883570 1793 888076
rect 17130 883570 17286 888076
rect 781 883443 17286 883570
rect 620598 883639 639620 883792
rect 620598 879190 620797 883639
rect 638082 879190 639620 883639
rect 620598 878992 639620 879190
rect 889 878028 17274 878192
rect 889 873522 1744 878028
rect 17081 873522 17274 878028
rect 889 873392 17274 873522
rect 620598 873616 639538 873741
rect 620598 869167 620810 873616
rect 638095 869167 639538 873616
rect 620598 868952 639538 869167
rect 1313 803652 5324 803750
rect 1313 799066 4359 803652
rect 5171 799066 5324 803652
rect 1313 798970 5324 799066
rect 633613 794462 639114 794593
rect 1294 793675 5299 793771
rect 1294 789089 4351 793675
rect 5163 789089 5299 793675
rect 633613 789897 633781 794462
rect 635118 789897 639114 794462
rect 633613 789813 639114 789897
rect 1294 788991 5299 789089
rect 633613 784517 639083 784614
rect 633613 779952 633749 784517
rect 635086 779952 639083 784517
rect 633613 779834 639083 779952
rect 630630 479910 639074 479993
rect 630630 475283 630713 479910
rect 632588 475283 639074 479910
rect 630630 475213 639074 475283
rect 630612 469932 639056 470014
rect 630612 465305 630706 469932
rect 632581 465305 639056 469932
rect 630612 465234 639056 465305
rect 1282 459103 7279 459135
rect 1282 454442 6326 459103
rect 7225 454442 7279 459103
rect 1282 454370 7279 454442
rect 1311 449139 7308 449171
rect 1311 444435 6315 449139
rect 7201 444435 7308 449139
rect 1311 444392 7308 444435
rect 625608 435779 639543 435992
rect 625608 431386 625855 435779
rect 638381 431386 639543 435779
rect 625608 431192 639543 431386
rect 625608 425749 639630 425941
rect 625608 421357 625811 425749
rect 638601 421357 639630 425749
rect 625608 421152 639630 421357
rect 904 416868 12379 417032
rect 904 412396 5639 416868
rect 12132 412396 12379 416868
rect 904 412243 12379 412396
rect 890 406832 12365 406992
rect 890 402360 5697 406832
rect 12190 402360 12365 406832
rect 890 402192 12365 402360
rect 633606 391672 639149 391793
rect 633606 387094 633737 391672
rect 635564 387094 639149 391672
rect 633606 387013 639149 387094
rect 633579 381734 639122 381814
rect 633579 377156 633726 381734
rect 635553 377156 639122 381734
rect 633579 377034 639122 377156
rect 1333 86219 13326 86350
rect 1333 81681 10344 86219
rect 13143 81681 13326 86219
rect 1333 81570 13326 81681
rect 1333 76201 13326 76371
rect 1333 71741 10357 76201
rect 13169 71741 13326 76201
rect 1333 71591 13326 71741
rect 770 44026 9140 44232
rect 770 39587 1813 44026
rect 8962 39587 9140 44026
rect 770 39443 9140 39587
rect 583 34000 9140 34192
rect 583 29539 1559 34000
rect 8951 29539 9140 34000
rect 583 29392 9140 29539
rect 202699 15152 207488 15425
rect 202699 9725 202830 15152
rect 207269 9725 207488 15152
rect 107896 9117 108610 9119
rect 104677 9102 108616 9117
rect 104677 8664 104698 9102
rect 105042 8664 108616 9102
rect 104677 8643 108616 8664
rect 104883 8641 108616 8643
rect 107896 3755 108610 8641
rect 107896 1861 107928 3755
rect 108561 1861 108610 3755
rect 107896 1818 108610 1861
rect 202699 620 207488 9725
rect 212739 15120 217539 15425
rect 212739 9693 212909 15120
rect 217348 9693 217539 15120
rect 212739 599 217539 9693
rect 530581 6582 535361 6705
rect 530581 2784 530645 6582
rect 535200 2784 535361 6582
rect 530581 1218 535361 2784
rect 540560 6573 545340 6714
rect 540560 2775 540643 6573
rect 545198 2775 545340 6573
rect 540560 1227 545340 2775
<< via3 >>
rect 537238 956582 541806 958512
rect 547188 956560 551756 958490
rect 1793 883570 17130 888076
rect 620797 879190 638082 883639
rect 1744 873522 17081 878028
rect 620810 869167 638095 873616
rect 4359 799066 5171 803652
rect 4351 789089 5163 793675
rect 633781 789897 635118 794462
rect 633749 779952 635086 784517
rect 630713 475283 632588 479910
rect 630706 465305 632581 469932
rect 6326 454442 7225 459103
rect 6315 444435 7201 449139
rect 625855 431386 638381 435779
rect 625811 421357 638601 425749
rect 5639 412396 12132 416868
rect 5697 402360 12190 406832
rect 633737 387094 635564 391672
rect 633726 377156 635553 381734
rect 10344 81681 13143 86219
rect 10357 71741 13169 76201
rect 1813 39587 8962 44026
rect 1559 29539 8951 34000
rect 202830 9725 207269 15152
rect 104698 8664 105042 9102
rect 107928 1861 108561 3755
rect 212909 9693 217348 15120
rect 530645 2784 535200 6582
rect 540643 2775 545198 6573
<< metal4 >>
rect 537142 958512 541910 958586
rect 537142 956582 537238 958512
rect 541806 956582 541910 958512
rect 537142 956220 541910 956582
rect 537142 953456 537238 956220
rect 541828 953456 541910 956220
rect 537142 953337 541910 953456
rect 547106 958490 551874 958572
rect 547106 956560 547188 958490
rect 551756 956560 551874 958490
rect 547106 956205 551874 956560
rect 547106 953441 547180 956205
rect 551770 953441 551874 956205
rect 547106 953323 551874 953441
rect 1648 888076 17286 888256
rect 1648 883570 1793 888076
rect 17130 883570 17286 888076
rect 1648 883473 17286 883570
rect 620660 883639 638402 883817
rect 620660 879190 620797 883639
rect 638082 879190 638402 883639
rect 620660 879028 638402 879190
rect 1612 878028 17250 878185
rect 1612 873522 1744 878028
rect 17081 878016 17250 878028
rect 17165 873619 17250 878016
rect 17081 873522 17250 873619
rect 1612 873402 17250 873522
rect 620598 873616 638332 873741
rect 620598 869167 620810 873616
rect 638095 869167 638332 873616
rect 620598 868952 638332 869167
rect 4270 803652 5272 803759
rect 4270 799066 4359 803652
rect 5171 799066 5272 803652
rect 4270 798985 5272 799066
rect 633661 794462 635232 794563
rect 4269 793675 5271 793760
rect 4269 789089 4351 793675
rect 5163 789089 5271 793675
rect 633661 789897 633781 794462
rect 635118 789897 635232 794462
rect 633661 789817 635232 789897
rect 4269 788986 5271 789089
rect 633673 784517 635244 784599
rect 633673 779952 633749 784517
rect 635086 779952 635244 784517
rect 633673 779853 635244 779952
rect 630652 479910 632660 479992
rect 630652 475283 630713 479910
rect 632588 475283 632660 479910
rect 630652 475222 632660 475283
rect 630648 469932 632656 470000
rect 630648 465305 630706 469932
rect 632581 465305 632656 469932
rect 630648 465230 632656 465305
rect 6245 459103 7322 459189
rect 6245 454442 6326 459103
rect 7225 454442 7322 459103
rect 6245 454364 7322 454442
rect 6220 449139 7297 449200
rect 6220 444435 6315 449139
rect 7201 444435 7297 449139
rect 6220 444375 7297 444435
rect 625608 435866 638675 435998
rect 625608 431326 625815 435866
rect 629491 435779 638675 435866
rect 638381 431386 638675 435779
rect 629491 431326 638675 431386
rect 625608 431192 638675 431326
rect 625608 425749 638807 425935
rect 625608 421357 625811 425749
rect 638601 421357 638807 425749
rect 625608 421152 638807 421357
rect 5551 416912 12278 417071
rect 5551 416868 8417 416912
rect 5551 412396 5639 416868
rect 12175 412440 12278 416912
rect 12132 412396 12278 412440
rect 5551 412250 12278 412396
rect 5551 406832 12278 407006
rect 5551 402360 5697 406832
rect 12190 402360 12278 406832
rect 5551 402185 12278 402360
rect 633661 391672 635651 391772
rect 633661 387094 633737 391672
rect 635564 387094 635651 391672
rect 633661 386987 635651 387094
rect 633639 381734 635651 381821
rect 633639 377156 633726 381734
rect 635553 377156 635651 381734
rect 633639 377052 635651 377156
rect 620641 242438 624668 242587
rect 8286 240968 12286 241061
rect 6237 238811 7262 238942
rect 6237 233558 6344 238811
rect 7160 233558 7262 238811
rect 6237 231502 7262 233558
rect 6237 227791 6355 231502
rect 7149 227791 7262 231502
rect 6237 227659 7262 227791
rect 8286 234855 8378 240968
rect 12145 234855 12286 240968
rect 8286 231501 12286 234855
rect 8286 227903 8423 231501
rect 12144 227903 12286 231501
rect 8286 227701 12286 227903
rect 13282 240911 17282 241061
rect 13282 237313 13396 240911
rect 17117 237313 17282 240911
rect 13282 231468 17282 237313
rect 13282 227870 13419 231468
rect 17140 227870 17282 231468
rect 620641 239279 620804 242438
rect 624519 239279 624668 242438
rect 620641 233434 624668 239279
rect 620641 230071 620817 233434
rect 624505 230071 624668 233434
rect 620641 229841 624668 230071
rect 625658 242425 629685 242587
rect 625658 236341 625807 242425
rect 629455 236341 629685 242425
rect 625658 233407 629685 236341
rect 625658 230044 625848 233407
rect 629536 230044 629685 233407
rect 625658 229841 629685 230044
rect 630635 242425 632682 242547
rect 630635 235468 630784 242425
rect 632547 235468 632682 242425
rect 630635 233461 632682 235468
rect 630635 230058 630865 233461
rect 632506 230058 632682 233461
rect 630635 229868 632682 230058
rect 13282 227701 17282 227870
rect 159182 225528 159543 225563
rect 159182 224103 159217 225528
rect 159507 224103 159543 225528
rect 159182 224066 159543 224103
rect 189282 225528 189643 225563
rect 189282 224103 189317 225528
rect 189607 224103 189643 225528
rect 189282 224066 189643 224103
rect 219382 225528 219743 225563
rect 219382 224103 219417 225528
rect 219707 224103 219743 225528
rect 219382 224066 219743 224103
rect 249482 225528 249843 225563
rect 249482 224103 249517 225528
rect 249807 224103 249843 225528
rect 249482 224066 249843 224103
rect 279582 225528 279943 225563
rect 279582 224103 279617 225528
rect 279907 224103 279943 225528
rect 279582 224066 279943 224103
rect 309682 225528 310043 225563
rect 309682 224103 309717 225528
rect 310007 224103 310043 225528
rect 309682 224066 310043 224103
rect 339782 225528 340143 225563
rect 339782 224103 339817 225528
rect 340107 224103 340143 225528
rect 339782 224066 340143 224103
rect 369882 225528 370243 225563
rect 369882 224103 369917 225528
rect 370207 224103 370243 225528
rect 369882 224066 370243 224103
rect 174229 223017 174620 223066
rect 174229 221605 174274 223017
rect 174572 221605 174620 223017
rect 174229 221563 174620 221605
rect 204329 223017 204720 223066
rect 204329 221605 204374 223017
rect 204672 221605 204720 223017
rect 204329 221563 204720 221605
rect 234429 223017 234820 223066
rect 234429 221605 234474 223017
rect 234772 221605 234820 223017
rect 234429 221563 234820 221605
rect 264529 223017 264920 223066
rect 264529 221605 264574 223017
rect 264872 221605 264920 223017
rect 264529 221563 264920 221605
rect 294629 223017 295020 223066
rect 294629 221605 294674 223017
rect 294972 221605 295020 223017
rect 294629 221563 295020 221605
rect 324729 223017 325120 223066
rect 324729 221605 324774 223017
rect 325072 221605 325120 223017
rect 324729 221563 325120 221605
rect 354829 223017 355220 223066
rect 354829 221605 354874 223017
rect 355172 221605 355220 223017
rect 354829 221563 355220 221605
rect 159984 220516 160416 220561
rect 159984 219105 160027 220516
rect 160382 219105 160416 220516
rect 159984 219067 160416 219105
rect 190084 220516 190516 220561
rect 190084 219105 190127 220516
rect 190482 219105 190516 220516
rect 190084 219067 190516 219105
rect 220184 220516 220616 220561
rect 220184 219105 220227 220516
rect 220582 219105 220616 220516
rect 220184 219067 220616 219105
rect 250224 220516 250576 220561
rect 250224 219105 250267 220516
rect 250542 219105 250576 220516
rect 250224 219067 250576 219105
rect 280384 220516 280816 220561
rect 280384 219105 280427 220516
rect 280782 219105 280816 220516
rect 280384 219067 280816 219105
rect 310484 220516 310916 220561
rect 310484 219105 310527 220516
rect 310882 219105 310916 220516
rect 310484 219067 310916 219105
rect 340584 220516 341016 220561
rect 340584 219105 340627 220516
rect 340982 219105 341016 220516
rect 340584 219067 341016 219105
rect 370684 220516 371116 220561
rect 370684 219105 370727 220516
rect 371082 219105 371116 220516
rect 370684 219067 371116 219105
rect 175882 218030 176215 218067
rect 175882 216608 175919 218030
rect 176178 216608 176215 218030
rect 175882 216567 176215 216608
rect 205982 218030 206315 218067
rect 205982 216608 206019 218030
rect 206278 216608 206315 218030
rect 205982 216567 206315 216608
rect 236082 218030 236415 218067
rect 236082 216608 236119 218030
rect 236378 216608 236415 218030
rect 236082 216567 236415 216608
rect 266182 218030 266515 218067
rect 266182 216608 266219 218030
rect 266478 216608 266515 218030
rect 266182 216567 266515 216608
rect 296282 218030 296615 218067
rect 296282 216608 296319 218030
rect 296578 216608 296615 218030
rect 296282 216567 296615 216608
rect 326382 218030 326715 218067
rect 326382 216608 326419 218030
rect 326678 216608 326715 218030
rect 326382 216567 326715 216608
rect 356482 218030 356815 218067
rect 356482 216608 356519 218030
rect 356778 216608 356815 218030
rect 356482 216567 356815 216608
rect 158364 215526 158733 215566
rect 158364 214096 158407 215526
rect 158695 214096 158733 215526
rect 158364 214066 158733 214096
rect 188464 215526 188833 215566
rect 188464 214096 188507 215526
rect 188795 214096 188833 215526
rect 188464 214066 188833 214096
rect 218564 215526 218933 215566
rect 218564 214096 218607 215526
rect 218895 214096 218933 215526
rect 218564 214066 218933 214096
rect 248754 215526 249113 215566
rect 248754 214096 248797 215526
rect 249075 214096 249113 215526
rect 248754 214066 249113 214096
rect 278764 215526 279083 215566
rect 278764 214096 278807 215526
rect 279045 214096 279083 215526
rect 278764 214066 279083 214096
rect 308864 215526 309233 215566
rect 308864 214096 308907 215526
rect 309195 214096 309233 215526
rect 308864 214066 309233 214096
rect 338964 215526 339333 215566
rect 338964 214096 339007 215526
rect 339295 214096 339333 215526
rect 338964 214066 339333 214096
rect 369064 215526 369433 215566
rect 369064 214096 369107 215526
rect 369395 214096 369433 215526
rect 369064 214066 369433 214096
rect 109921 213365 116936 213753
rect 109921 207012 110403 213365
rect 116528 207012 116936 213365
rect 109921 200162 116936 207012
rect 109921 199698 110021 200162
rect 116816 199698 116936 200162
rect 109921 197631 116936 199698
rect 109936 190162 116936 197631
rect 129936 213365 136936 213574
rect 129936 207012 130322 213365
rect 136447 207012 136936 213365
rect 173422 213029 173760 213061
rect 173422 211601 173451 213029
rect 173725 211601 173760 213029
rect 173422 211564 173760 211601
rect 203522 213029 203860 213061
rect 203522 211601 203551 213029
rect 203825 211601 203860 213029
rect 203522 211564 203860 211601
rect 233672 213029 234010 213061
rect 233672 211601 233701 213029
rect 233975 211601 234010 213029
rect 293822 213029 294160 213061
rect 233672 211564 234010 211601
rect 263662 212949 264000 212981
rect 263662 211601 263691 212949
rect 263965 211601 264000 212949
rect 263662 211564 264000 211601
rect 293822 211601 293851 213029
rect 294125 211601 294160 213029
rect 293822 211564 294160 211601
rect 323922 213029 324260 213061
rect 323922 211601 323951 213029
rect 324225 211601 324260 213029
rect 323922 211564 324260 211601
rect 354022 213029 354360 213061
rect 354022 211601 354051 213029
rect 354325 211601 354360 213029
rect 354022 211564 354360 211601
rect 160062 210533 160393 210565
rect 160062 209096 160095 210533
rect 160347 209096 160393 210533
rect 160062 209060 160393 209096
rect 190162 210533 190493 210565
rect 190162 209096 190195 210533
rect 190447 209096 190493 210533
rect 190162 209060 190493 209096
rect 220262 210533 220593 210565
rect 220262 209096 220295 210533
rect 220547 209096 220593 210533
rect 220262 209060 220593 209096
rect 250242 210533 250573 210565
rect 250242 209096 250275 210533
rect 250527 209096 250573 210533
rect 250242 209060 250573 209096
rect 280462 210533 280793 210565
rect 280462 209096 280495 210533
rect 280747 209096 280793 210533
rect 280462 209060 280793 209096
rect 310562 210533 310893 210565
rect 310562 209096 310595 210533
rect 310847 209096 310893 210533
rect 310562 209060 310893 209096
rect 340662 210533 340993 210565
rect 340662 209096 340695 210533
rect 340947 209096 340993 210533
rect 340662 209060 340993 209096
rect 370762 210533 371093 210565
rect 370762 209096 370795 210533
rect 371047 209096 371093 210533
rect 370762 209060 371093 209096
rect 109936 189698 110021 190162
rect 116816 189698 116936 190162
rect 109936 180162 116936 189698
rect 109936 179698 110021 180162
rect 116816 179698 116936 180162
rect 109936 170162 116936 179698
rect 109936 169698 110021 170162
rect 116816 169698 116936 170162
rect 109936 160162 116936 169698
rect 109936 159698 110021 160162
rect 116816 159698 116936 160162
rect 109936 150162 116936 159698
rect 109936 149698 110021 150162
rect 116816 149698 116936 150162
rect 109936 140162 116936 149698
rect 109936 139698 110021 140162
rect 116816 139698 116936 140162
rect 109936 130162 116936 139698
rect 109936 129698 110021 130162
rect 116816 129698 116936 130162
rect 109936 120162 116936 129698
rect 109936 119698 110021 120162
rect 116816 119698 116936 120162
rect 109936 110162 116936 119698
rect 109936 109698 110021 110162
rect 116816 109698 116936 110162
rect 109936 100162 116936 109698
rect 109936 99698 110021 100162
rect 116816 99698 116936 100162
rect 109936 90162 116936 99698
rect 109936 89698 110021 90162
rect 116816 89698 116936 90162
rect 10265 86219 13265 86428
rect 10265 81681 10344 86219
rect 13143 81681 13265 86219
rect 10265 76201 13265 81681
rect 10265 71741 10357 76201
rect 13169 71741 13265 76201
rect 1687 44026 9128 44216
rect 1687 39587 1813 44026
rect 8962 39587 9128 44026
rect 1687 39426 9128 39587
rect 1399 34000 9121 34185
rect 1399 29539 1559 34000
rect 8951 29539 9121 34000
rect 1399 29395 9121 29539
rect 10265 8084 13265 71741
rect 109936 80162 116936 89698
rect 109936 79698 110021 80162
rect 116816 79698 116936 80162
rect 109936 70162 116936 79698
rect 109936 69698 110021 70162
rect 116816 69698 116936 70162
rect 109936 60162 116936 69698
rect 109936 59698 110021 60162
rect 116816 59698 116936 60162
rect 109936 50162 116936 59698
rect 109936 49698 110021 50162
rect 116816 49698 116936 50162
rect 109936 40162 116936 49698
rect 109936 39698 110021 40162
rect 116816 39698 116936 40162
rect 109936 30162 116936 39698
rect 109936 29698 110021 30162
rect 116816 29698 116936 30162
rect 109936 20162 116936 29698
rect 119936 195145 126936 195210
rect 119936 194628 119991 195145
rect 126852 194628 126936 195145
rect 119936 188265 126936 194628
rect 119936 183580 120133 188265
rect 126688 183580 126936 188265
rect 119936 175168 126936 183580
rect 119936 174631 120020 175168
rect 126822 174631 126936 175168
rect 119936 165168 126936 174631
rect 119936 164631 120020 165168
rect 126822 164631 126936 165168
rect 119936 155168 126936 164631
rect 119936 154631 120020 155168
rect 126822 154631 126936 155168
rect 119936 145168 126936 154631
rect 119936 144631 120020 145168
rect 126822 144631 126936 145168
rect 119936 135168 126936 144631
rect 119936 134631 120020 135168
rect 126822 134631 126936 135168
rect 119936 125168 126936 134631
rect 119936 124631 120020 125168
rect 126822 124631 126936 125168
rect 119936 115168 126936 124631
rect 119936 114631 120020 115168
rect 126822 114631 126936 115168
rect 119936 105168 126936 114631
rect 119936 104631 120020 105168
rect 126822 104631 126936 105168
rect 119936 95168 126936 104631
rect 119936 94631 120020 95168
rect 126822 94631 126936 95168
rect 119936 85168 126936 94631
rect 119936 84631 120020 85168
rect 126822 84631 126936 85168
rect 119936 75168 126936 84631
rect 119936 74631 120020 75168
rect 126822 74631 126936 75168
rect 119936 65168 126936 74631
rect 119936 64631 120020 65168
rect 126822 64631 126936 65168
rect 119936 55168 126936 64631
rect 119936 54631 120020 55168
rect 126822 54631 126936 55168
rect 119936 45168 126936 54631
rect 119936 44631 120020 45168
rect 126822 44631 126936 45168
rect 119936 35168 126936 44631
rect 119936 34631 120020 35168
rect 126822 34631 126936 35168
rect 119936 26772 126936 34631
rect 119936 22141 120212 26772
rect 126733 22141 126936 26772
rect 119936 21906 126936 22141
rect 129936 176657 136936 207012
rect 175073 208037 175402 208065
rect 175073 206605 175100 208037
rect 175364 206605 175402 208037
rect 175073 206567 175402 206605
rect 205173 208037 205502 208065
rect 205173 206605 205200 208037
rect 205464 206605 205502 208037
rect 205173 206567 205502 206605
rect 235333 208037 235662 208065
rect 235333 206605 235360 208037
rect 235624 206605 235662 208037
rect 235333 206567 235662 206605
rect 265323 208037 265652 208065
rect 265323 206605 265350 208037
rect 265614 206605 265652 208037
rect 265323 206567 265652 206605
rect 295473 208037 295802 208065
rect 295473 206605 295500 208037
rect 295764 206605 295802 208037
rect 295473 206567 295802 206605
rect 325573 208037 325902 208065
rect 325573 206605 325600 208037
rect 325864 206605 325902 208037
rect 325573 206567 325902 206605
rect 355673 208037 356002 208065
rect 355673 206605 355700 208037
rect 355964 206605 356002 208037
rect 355673 206567 356002 206605
rect 157538 205533 157910 205564
rect 157538 204093 157566 205533
rect 157877 204093 157910 205533
rect 157538 204068 157910 204093
rect 187638 205533 188010 205564
rect 187638 204093 187666 205533
rect 187977 204093 188010 205533
rect 187638 204068 188010 204093
rect 217738 205533 218110 205564
rect 217738 204093 217766 205533
rect 218077 204093 218110 205533
rect 217738 204068 218110 204093
rect 247788 205533 248160 205564
rect 247788 204093 247816 205533
rect 248127 204093 248160 205533
rect 247788 204068 248160 204093
rect 278018 205533 278340 205564
rect 278018 204093 278046 205533
rect 278307 204093 278340 205533
rect 278018 204068 278340 204093
rect 308038 205533 308410 205564
rect 308038 204093 308066 205533
rect 308377 204093 308410 205533
rect 308038 204068 308410 204093
rect 338138 205533 338510 205564
rect 338138 204093 338166 205533
rect 338477 204093 338510 205533
rect 338138 204068 338510 204093
rect 368238 205533 368610 205564
rect 368238 204093 368266 205533
rect 368577 204093 368610 205533
rect 368238 204068 368610 204093
rect 172596 203026 172965 203066
rect 172596 201601 172628 203026
rect 172929 201601 172965 203026
rect 172596 201566 172965 201601
rect 202696 203026 203065 203066
rect 202696 201601 202728 203026
rect 203029 201601 203065 203026
rect 202696 201566 203065 201601
rect 232796 203026 233165 203066
rect 232796 201601 232828 203026
rect 233129 201601 233165 203026
rect 232796 201566 233165 201601
rect 262896 203026 263265 203066
rect 262896 201601 262928 203026
rect 263229 201601 263265 203026
rect 262896 201566 263265 201601
rect 292886 203026 293255 203066
rect 292886 201601 292918 203026
rect 293219 201601 293255 203026
rect 292886 201566 293255 201601
rect 323096 203026 323465 203066
rect 323096 201601 323128 203026
rect 323429 201601 323465 203026
rect 323096 201566 323465 201601
rect 353196 203026 353565 203066
rect 353196 201601 353228 203026
rect 353529 201601 353565 203026
rect 353196 201566 353565 201601
rect 387736 202845 394099 203087
rect 387736 201297 387985 202845
rect 393910 201297 394099 202845
rect 129936 176107 130009 176657
rect 136855 176107 136936 176657
rect 129936 150657 136936 176107
rect 129936 150107 130009 150657
rect 136855 150107 136936 150657
rect 129936 124657 136936 150107
rect 129936 124107 130009 124657
rect 136855 124107 136936 124657
rect 129936 98657 136936 124107
rect 129936 98107 130009 98657
rect 136855 98107 136936 98657
rect 129936 72657 136936 98107
rect 129936 72107 130009 72657
rect 136855 72107 136936 72657
rect 129936 46657 136936 72107
rect 129936 46107 130009 46657
rect 136855 46107 136936 46657
rect 129936 29832 136936 46107
rect 129936 29243 129997 29832
rect 136890 29243 136936 29832
rect 109936 19698 110021 20162
rect 116816 19698 116936 20162
rect 103995 16262 104641 16287
rect 103995 15523 104025 16262
rect 104608 15523 104641 16262
rect 103995 15490 104641 15523
rect 103999 8961 104179 15490
rect 109936 14272 116936 19698
rect 105009 13315 105775 13367
rect 105009 12252 105051 13315
rect 105711 12252 105775 13315
rect 105009 12187 105775 12252
rect 105299 10514 105479 12187
rect 109936 9641 110144 14272
rect 116665 9641 116936 14272
rect 109936 9338 116936 9641
rect 129936 14174 136936 29243
rect 138936 188234 145936 188621
rect 138936 183549 139135 188234
rect 145690 183549 145936 188234
rect 138936 163654 145936 183549
rect 387736 188204 394099 201297
rect 608559 195168 613559 195344
rect 608559 190557 608763 195168
rect 613356 190557 613559 195168
rect 387736 183649 388000 188204
rect 393895 183649 394099 188204
rect 387736 183011 394099 183649
rect 602559 188229 607559 188383
rect 602559 183618 602772 188229
rect 607365 183618 607559 188229
rect 138936 163065 138995 163654
rect 145878 163065 145936 163654
rect 138936 137654 145936 163065
rect 138936 137065 138995 137654
rect 145878 137065 145936 137654
rect 138936 111654 145936 137065
rect 138936 111065 138995 111654
rect 145878 111065 145936 111654
rect 138936 85654 145936 111065
rect 138936 85065 138995 85654
rect 145878 85065 145936 85654
rect 138936 59654 145936 85065
rect 138936 59065 138995 59654
rect 145878 59065 145936 59654
rect 138936 33654 145936 59065
rect 138936 33065 138995 33654
rect 145878 33065 145936 33654
rect 138936 26804 145936 33065
rect 138936 22173 139167 26804
rect 145688 22173 145936 26804
rect 138936 21906 145936 22173
rect 602559 163571 607559 183618
rect 602559 163148 602628 163571
rect 607445 163148 607559 163571
rect 602559 137571 607559 163148
rect 602559 137148 602628 137571
rect 607445 137148 607559 137571
rect 602559 111571 607559 137148
rect 602559 111148 602628 111571
rect 607445 111148 607559 111571
rect 602559 85571 607559 111148
rect 602559 85148 602628 85571
rect 607445 85148 607559 85571
rect 602559 59571 607559 85148
rect 602559 59148 602628 59571
rect 607445 59148 607559 59571
rect 602559 46757 607559 59148
rect 602559 46284 602636 46757
rect 607470 46284 607559 46757
rect 602559 45120 607559 46284
rect 602559 44647 602600 45120
rect 607434 44647 607559 45120
rect 602559 33615 607559 44647
rect 602559 33085 602623 33615
rect 607495 33085 607559 33615
rect 602559 18529 607559 33085
rect 129936 9543 130166 14174
rect 136687 9543 136936 14174
rect 129936 9207 136936 9543
rect 202686 15232 207477 15441
rect 202686 10634 202782 15232
rect 207285 10634 207477 15232
rect 202686 9725 202830 10634
rect 207269 9725 207477 10634
rect 202686 9501 207477 9725
rect 212765 15200 217556 15393
rect 212765 10602 212877 15200
rect 217380 10602 217556 15200
rect 602559 14168 602693 18529
rect 607423 14168 607559 18529
rect 608559 176601 613559 190557
rect 608559 176153 608613 176601
rect 613500 176153 613559 176601
rect 608559 150601 613559 176153
rect 608559 150153 608613 150601
rect 613500 150153 613559 150601
rect 608559 124601 613559 150153
rect 608559 124153 608613 124601
rect 613500 124153 613559 124601
rect 608559 98601 613559 124153
rect 608559 98153 608613 98601
rect 613500 98153 613559 98601
rect 608559 72601 613559 98153
rect 608559 72153 608613 72601
rect 613500 72153 613559 72601
rect 608559 65265 613559 72153
rect 614123 75734 615417 75779
rect 614123 74690 614156 75734
rect 615367 74690 615417 75734
rect 614123 66919 615417 74690
rect 614123 66521 616130 66919
rect 614173 66519 616130 66521
rect 608559 64636 608612 65265
rect 613504 64636 613559 65265
rect 608559 47558 613559 64636
rect 614106 65891 615647 66209
rect 622876 66145 626729 66212
rect 614106 63098 615400 65891
rect 622870 65883 626729 66145
rect 622870 65118 624708 65883
rect 622870 64798 622897 65118
rect 624672 64798 624708 65118
rect 622870 64757 624708 64798
rect 614106 61750 614165 63098
rect 615335 61750 615400 63098
rect 614106 61685 615400 61750
rect 608559 47085 608618 47558
rect 613452 47085 613559 47558
rect 608559 45911 613559 47085
rect 608559 45438 608633 45911
rect 613467 45438 613559 45911
rect 608559 44256 613559 45438
rect 608559 43861 608607 44256
rect 613498 43861 613559 44256
rect 608559 20655 613559 43861
rect 608559 16294 608661 20655
rect 613391 16294 613559 20655
rect 608559 16161 613559 16294
rect 602559 14061 607559 14168
rect 222286 11866 631506 11878
rect 222231 11854 631506 11866
rect 212765 9693 212909 10602
rect 217348 9693 217556 10602
rect 212765 9453 217556 9693
rect 222053 11787 631506 11854
rect 104677 9102 105059 9117
rect 104677 8664 104698 9102
rect 105042 8664 105059 9102
rect 104677 8643 105059 8664
rect 106179 8084 106359 8902
rect 222053 8084 628597 11787
rect 10265 7973 628597 8084
rect 631428 7973 631506 11787
rect 10265 7878 631506 7973
rect 10265 4775 225362 7878
rect 229032 6588 635531 6686
rect 229032 6582 632642 6588
rect 10265 3815 106953 4775
rect 229032 3803 530645 6582
rect 107864 3755 530645 3803
rect 107864 1861 107928 3755
rect 108561 2784 530645 3755
rect 535200 6573 632642 6582
rect 535200 2784 540643 6573
rect 108561 2775 540643 2784
rect 545198 2815 632642 6573
rect 635402 2815 635531 6588
rect 545198 2775 635531 2815
rect 108561 2686 635531 2775
rect 108561 1861 231437 2686
rect 107864 1803 231437 1861
<< via4 >>
rect 537238 953456 541828 956220
rect 547180 953441 551770 956205
rect 13382 883618 17116 888015
rect 620860 879253 624447 883577
rect 13431 873619 17081 878016
rect 17081 873619 17165 878016
rect 620810 869167 624397 873491
rect 4359 799066 5171 803652
rect 4351 789089 5163 793675
rect 633781 789897 635118 794462
rect 633749 779952 635086 784517
rect 630713 475283 632588 479910
rect 630706 465305 632581 469932
rect 6326 454442 7225 459103
rect 6315 444435 7201 449139
rect 625815 435779 629491 435866
rect 625815 431386 625855 435779
rect 625855 431386 629491 435779
rect 625815 431326 629491 431386
rect 625811 421357 629472 425749
rect 8417 416868 12175 416912
rect 8417 412440 12132 416868
rect 12132 412440 12175 416868
rect 8374 402360 12132 406832
rect 633737 387094 635564 391672
rect 633726 377156 635553 381734
rect 6344 233558 7160 238811
rect 6355 227791 7149 231502
rect 8378 234855 12145 240968
rect 8423 227903 12144 231501
rect 13396 237313 17117 240911
rect 13419 227870 17140 231468
rect 620804 239279 624519 242438
rect 620817 230071 624505 233434
rect 625807 236341 629455 242425
rect 625848 230044 629536 233407
rect 630784 235468 632547 242425
rect 630865 230058 632506 233461
rect 159217 224103 159507 225528
rect 189317 224103 189607 225528
rect 219417 224103 219707 225528
rect 249517 224103 249807 225528
rect 279617 224103 279907 225528
rect 309717 224103 310007 225528
rect 339817 224103 340107 225528
rect 369917 224103 370207 225528
rect 174274 221605 174572 223017
rect 204374 221605 204672 223017
rect 234474 221605 234772 223017
rect 264574 221605 264872 223017
rect 294674 221605 294972 223017
rect 324774 221605 325072 223017
rect 354874 221605 355172 223017
rect 160027 219105 160382 220516
rect 190127 219105 190482 220516
rect 220227 219105 220582 220516
rect 250267 219105 250542 220516
rect 280427 219105 280782 220516
rect 310527 219105 310882 220516
rect 340627 219105 340982 220516
rect 370727 219105 371082 220516
rect 175919 216608 176178 218030
rect 206019 216608 206278 218030
rect 236119 216608 236378 218030
rect 266219 216608 266478 218030
rect 296319 216608 296578 218030
rect 326419 216608 326678 218030
rect 356519 216608 356778 218030
rect 158407 214096 158695 215526
rect 188507 214096 188795 215526
rect 218607 214096 218895 215526
rect 248797 214096 249075 215526
rect 278807 214096 279045 215526
rect 308907 214096 309195 215526
rect 339007 214096 339295 215526
rect 369107 214096 369395 215526
rect 110403 207012 116528 213365
rect 110021 199698 116816 200162
rect 130322 207012 136447 213365
rect 173451 211601 173725 213029
rect 203551 211601 203825 213029
rect 233701 211601 233975 213029
rect 263691 211601 263965 212949
rect 293851 211601 294125 213029
rect 323951 211601 324225 213029
rect 354051 211601 354325 213029
rect 160095 209096 160347 210533
rect 190195 209096 190447 210533
rect 220295 209096 220547 210533
rect 250275 209096 250527 210533
rect 280495 209096 280747 210533
rect 310595 209096 310847 210533
rect 340695 209096 340947 210533
rect 370795 209096 371047 210533
rect 110021 189698 116816 190162
rect 110021 179698 116816 180162
rect 110021 169698 116816 170162
rect 110021 159698 116816 160162
rect 110021 149698 116816 150162
rect 110021 139698 116816 140162
rect 110021 129698 116816 130162
rect 110021 119698 116816 120162
rect 110021 109698 116816 110162
rect 110021 99698 116816 100162
rect 110021 89698 116816 90162
rect 4302 39598 8940 43927
rect 4280 30314 8918 33967
rect 4280 29638 8917 30314
rect 110021 79698 116816 80162
rect 110021 69698 116816 70162
rect 110021 59698 116816 60162
rect 110021 49698 116816 50162
rect 110021 39698 116816 40162
rect 110021 29698 116816 30162
rect 119991 194628 126852 195145
rect 120133 183580 126688 188265
rect 120020 174631 126822 175168
rect 120020 164631 126822 165168
rect 120020 154631 126822 155168
rect 120020 144631 126822 145168
rect 120020 134631 126822 135168
rect 120020 124631 126822 125168
rect 120020 114631 126822 115168
rect 120020 104631 126822 105168
rect 120020 94631 126822 95168
rect 120020 84631 126822 85168
rect 120020 74631 126822 75168
rect 120020 64631 126822 65168
rect 120020 54631 126822 55168
rect 120020 44631 126822 45168
rect 120020 34631 126822 35168
rect 120212 22141 126733 26772
rect 175100 206605 175364 208037
rect 205200 206605 205464 208037
rect 235360 206605 235624 208037
rect 265350 206605 265614 208037
rect 295500 206605 295764 208037
rect 325600 206605 325864 208037
rect 355700 206605 355964 208037
rect 157566 204093 157877 205533
rect 187666 204093 187977 205533
rect 217766 204093 218077 205533
rect 247816 204093 248127 205533
rect 278046 204093 278307 205533
rect 308066 204093 308377 205533
rect 338166 204093 338477 205533
rect 368266 204093 368577 205533
rect 172628 201601 172929 203026
rect 202728 201601 203029 203026
rect 232828 201601 233129 203026
rect 262928 201601 263229 203026
rect 292918 201601 293219 203026
rect 323128 201601 323429 203026
rect 353228 201601 353529 203026
rect 387985 201297 393910 202845
rect 130009 176107 136855 176657
rect 130009 150107 136855 150657
rect 130009 124107 136855 124657
rect 130009 98107 136855 98657
rect 130009 72107 136855 72657
rect 130009 46107 136855 46657
rect 129997 29243 136890 29832
rect 110021 19698 116816 20162
rect 104025 15523 104608 16262
rect 105051 12252 105711 13315
rect 110144 9641 116665 14272
rect 139135 183549 145690 188234
rect 608763 190557 613356 195168
rect 388000 183649 393895 188204
rect 602772 183618 607365 188229
rect 138995 163065 145878 163654
rect 138995 137065 145878 137654
rect 138995 111065 145878 111654
rect 138995 85065 145878 85654
rect 138995 59065 145878 59654
rect 138995 33065 145878 33654
rect 139167 22173 145688 26804
rect 602628 163148 607445 163571
rect 602628 137148 607445 137571
rect 602628 111148 607445 111571
rect 602628 85148 607445 85571
rect 602628 59148 607445 59571
rect 602636 46284 607470 46757
rect 602600 44647 607434 45120
rect 602623 33085 607495 33615
rect 130166 9543 136687 14174
rect 202782 15152 207285 15232
rect 202782 10634 202830 15152
rect 202830 10634 207269 15152
rect 207269 10634 207285 15152
rect 212877 15120 217380 15200
rect 212877 10602 212909 15120
rect 212909 10602 217348 15120
rect 217348 10602 217380 15120
rect 602693 14168 607423 18529
rect 608613 176153 613500 176601
rect 608613 150153 613500 150601
rect 608613 124153 613500 124601
rect 608613 98153 613500 98601
rect 608613 72153 613500 72601
rect 614156 74690 615367 75734
rect 608612 64636 613504 65265
rect 622897 64798 624672 65118
rect 614165 61750 615335 63098
rect 608618 47085 613452 47558
rect 608633 45438 613467 45911
rect 608607 43861 613498 44256
rect 608661 16294 613391 20655
rect 628597 7973 631428 11787
rect 632642 2815 635402 6588
<< metal5 >>
rect 633657 956325 635657 956329
rect 537099 956220 635657 956325
rect 537099 953456 537238 956220
rect 541828 956205 635657 956220
rect 541828 953456 547180 956205
rect 537099 953441 547180 953456
rect 551770 953441 635657 956205
rect 537099 953325 635657 953441
rect 4273 950850 18820 951450
rect 4273 803652 5273 950850
rect 4273 799066 4359 803652
rect 5171 799066 5273 803652
rect 4273 793675 5273 799066
rect 4273 789089 4351 793675
rect 5163 789089 5273 793675
rect 4273 233106 5273 789089
rect 6273 949910 19792 950510
rect 6273 459103 7273 949910
rect 633657 949570 635657 953325
rect 616645 948970 635657 949570
rect 615787 948030 632657 948630
rect 6273 454442 6326 459103
rect 7225 454442 7273 459103
rect 6273 449139 7273 454442
rect 6273 444435 6315 449139
rect 7201 444435 7273 449139
rect 6273 238811 7273 444435
rect 6273 233558 6344 238811
rect 7160 234046 7273 238811
rect 8273 947090 22611 947690
rect 8273 416912 12273 947090
rect 8273 412440 8417 416912
rect 12175 412440 12273 416912
rect 8273 406832 12273 412440
rect 8273 402360 8374 406832
rect 12132 402360 12273 406832
rect 8273 240968 12273 402360
rect 8273 234855 8378 240968
rect 12145 236866 12273 240968
rect 13273 946150 23511 946750
rect 13273 888015 17273 946150
rect 625657 945810 629657 945814
rect 612964 945210 629657 945810
rect 612016 944847 624648 944870
rect 612016 944270 624657 944847
rect 13273 883618 13382 888015
rect 17116 883618 17273 888015
rect 13273 878016 17273 883618
rect 13273 873619 13431 878016
rect 17165 873619 17273 878016
rect 13273 240911 17273 873619
rect 13273 237313 13396 240911
rect 17117 237806 17273 240911
rect 620657 883577 624657 944270
rect 620657 879253 620860 883577
rect 624447 879253 624657 883577
rect 620657 873491 624657 879253
rect 620657 869167 620810 873491
rect 624397 869167 624657 873491
rect 620657 242438 624657 869167
rect 620657 239686 620804 242438
rect 611967 239279 620804 239686
rect 624519 239279 624657 242438
rect 611967 239093 624657 239279
rect 625657 435866 629657 945210
rect 625657 431326 625815 435866
rect 629491 431326 629657 435866
rect 625657 425749 629657 431326
rect 625657 421357 625811 425749
rect 629472 421357 629657 425749
rect 625657 242425 629657 421357
rect 611967 239086 624610 239093
rect 625657 238746 625807 242425
rect 612951 238146 625807 238746
rect 17117 237313 23509 237806
rect 13273 237206 23509 237313
rect 13273 237181 17273 237206
rect 12145 236266 22611 236866
rect 625657 236341 625807 238146
rect 629455 238746 629657 242425
rect 630657 479910 632657 948030
rect 630657 475283 630713 479910
rect 632588 475283 632657 479910
rect 630657 469932 632657 475283
rect 630657 465305 630706 469932
rect 632581 465305 632657 469932
rect 630657 242425 632657 465305
rect 629455 238146 629686 238746
rect 629455 236341 629657 238146
rect 12145 234855 12273 236266
rect 625657 236228 629657 236341
rect 630657 235926 630784 242425
rect 615700 235468 630784 235926
rect 632547 235468 632657 242425
rect 615700 235326 632657 235468
rect 630657 235323 632657 235326
rect 633657 794462 635657 948970
rect 633657 789897 633781 794462
rect 635118 789897 635657 794462
rect 633657 784517 635657 789897
rect 633657 779952 633749 784517
rect 635086 779952 635657 784517
rect 633657 391672 635657 779952
rect 633657 387094 633737 391672
rect 635564 387094 635657 391672
rect 633657 381734 635657 387094
rect 633657 377156 633726 381734
rect 635553 377156 635657 381734
rect 630657 235315 632621 235323
rect 633657 234986 635657 377156
rect 8273 234697 12273 234855
rect 616560 234386 635657 234986
rect 7160 233558 19774 234046
rect 6273 233446 19774 233558
rect 6273 233435 7273 233446
rect 620657 233434 624657 233624
rect 4273 232506 18789 233106
rect 4273 217854 5273 232506
rect 6273 231502 7273 231631
rect 6273 227791 6355 231502
rect 7149 227791 7273 231502
rect 6273 220854 7273 227791
rect 8273 231501 12273 231631
rect 8273 227903 8423 231501
rect 12144 227903 12273 231501
rect 8273 224854 12273 227903
rect 13273 231468 17273 231631
rect 13273 227870 13419 231468
rect 17140 229854 17273 231468
rect 620657 230071 620817 233434
rect 624505 230071 624657 233434
rect 17140 227870 144995 229854
rect 13273 226854 144995 227870
rect 620657 227074 624657 230071
rect 143495 225564 144995 226854
rect 143495 225528 372157 225564
rect 8273 223064 141281 224854
rect 143495 224103 159217 225528
rect 159507 224103 189317 225528
rect 189607 224103 219417 225528
rect 219707 224103 249517 225528
rect 249807 224103 279617 225528
rect 279907 224103 309717 225528
rect 310007 224103 339817 225528
rect 340107 224103 369917 225528
rect 370207 224103 372157 225528
rect 143495 224064 372157 224103
rect 383256 223074 624657 227074
rect 625657 233407 629657 233624
rect 625657 230044 625848 233407
rect 629536 230044 629657 233407
rect 8273 223017 372157 223064
rect 8273 221854 174274 223017
rect 139781 221605 174274 221854
rect 174572 221605 204374 223017
rect 204672 221605 234474 223017
rect 234772 221605 264574 223017
rect 264872 221605 294674 223017
rect 294972 221605 324774 223017
rect 325072 221605 354874 223017
rect 355172 221605 372157 223017
rect 139781 221564 372157 221605
rect 6273 220564 137328 220854
rect 6273 220516 372157 220564
rect 6273 219105 160027 220516
rect 160382 219105 190127 220516
rect 190482 219105 220227 220516
rect 220582 219105 250267 220516
rect 250542 219105 280427 220516
rect 280782 219105 310527 220516
rect 310882 219105 340627 220516
rect 340982 219105 370727 220516
rect 371082 219105 372157 220516
rect 6273 219064 372157 219105
rect 6273 218854 137328 219064
rect 138364 218030 357099 218064
rect 138364 217854 175919 218030
rect 4273 216608 175919 217854
rect 176178 216608 206019 218030
rect 206278 216608 236119 218030
rect 236378 216608 266219 218030
rect 266478 216608 296319 218030
rect 296578 216608 326419 218030
rect 326678 216608 356519 218030
rect 356778 216608 357099 218030
rect 4273 216564 357099 216608
rect 4273 215854 140993 216564
rect 383256 215564 387256 223074
rect 625657 221074 629657 230044
rect 158192 215526 387256 215564
rect 158192 214096 158407 215526
rect 158695 214096 188507 215526
rect 188795 214096 218607 215526
rect 218895 214096 248797 215526
rect 249075 214096 278807 215526
rect 279045 214096 308907 215526
rect 309195 214096 339007 215526
rect 339295 214096 369107 215526
rect 369395 214096 387256 215526
rect 158192 214064 387256 214096
rect 389353 217074 629657 221074
rect 630657 233461 632657 233624
rect 630657 230058 630865 233461
rect 632506 230058 632657 233461
rect 5106 213365 145906 213604
rect 5106 207012 110403 213365
rect 116528 207012 130322 213365
rect 136447 207012 145906 213365
rect 389353 213064 393353 217074
rect 630657 213074 632657 230058
rect 173291 213029 393353 213064
rect 173291 211601 173451 213029
rect 173725 211601 203551 213029
rect 203825 211601 233701 213029
rect 233975 212949 293851 213029
rect 233975 211601 263691 212949
rect 263965 211601 293851 212949
rect 294125 211601 323951 213029
rect 324225 211601 354051 213029
rect 354325 211601 393353 213029
rect 173291 211564 393353 211601
rect 395119 210564 632657 213074
rect 159813 210533 632657 210564
rect 159813 209096 160095 210533
rect 160347 209096 190195 210533
rect 190447 209096 220295 210533
rect 220547 209096 250275 210533
rect 250527 209096 280495 210533
rect 280747 209096 310595 210533
rect 310847 209096 340695 210533
rect 340947 209096 370795 210533
rect 371047 210074 632657 210533
rect 371047 209096 398119 210074
rect 159813 209064 398119 209096
rect 633657 209074 635657 234386
rect 401055 208064 635657 209074
rect 5106 206604 145906 207012
rect 5106 200066 10106 206604
rect 138906 205564 145906 206604
rect 174811 208037 635657 208064
rect 174811 206605 175100 208037
rect 175364 206605 205200 208037
rect 205464 206605 235360 208037
rect 235624 206605 265350 208037
rect 265614 206605 295500 208037
rect 295764 206605 325600 208037
rect 325864 206605 355700 208037
rect 355964 206605 635657 208037
rect 174811 206564 635657 206605
rect 401055 206074 635657 206564
rect 138906 205533 368771 205564
rect 138906 204093 157566 205533
rect 157877 204093 187666 205533
rect 187977 204093 217766 205533
rect 218077 204093 247816 205533
rect 248127 204093 278046 205533
rect 278307 204093 308066 205533
rect 308377 204093 338166 205533
rect 338477 204093 368266 205533
rect 368577 204093 368771 205533
rect 138906 204064 368771 204093
rect 109924 200162 116943 200253
rect 109924 200066 110021 200162
rect 5106 199746 14895 200066
rect 104047 199746 110021 200066
rect 5106 190066 10106 199746
rect 109924 199698 110021 199746
rect 116816 200066 116943 200162
rect 116816 199746 116961 200066
rect 116816 199698 116943 199746
rect 109924 199612 116943 199698
rect 138906 195370 145906 204064
rect 172379 203026 394268 203064
rect 172379 201601 172628 203026
rect 172929 201601 202728 203026
rect 203029 201601 232828 203026
rect 233129 201601 262928 203026
rect 263229 201601 292918 203026
rect 293219 201601 323128 203026
rect 323429 201601 353228 203026
rect 353529 202845 394268 203026
rect 353529 201601 387985 202845
rect 172379 201564 387985 201601
rect 387723 201297 387985 201564
rect 393910 201297 394268 202845
rect 387723 201064 394268 201297
rect 387741 201053 394235 201064
rect 119933 195145 126973 195272
rect 119933 195066 119991 195145
rect 104047 194746 119991 195066
rect 119933 194628 119991 194746
rect 126852 195066 126973 195145
rect 138906 195168 613563 195370
rect 126852 194746 126975 195066
rect 126852 194628 126973 194746
rect 119933 194559 126973 194628
rect 138906 190557 608763 195168
rect 613356 190557 613563 195168
rect 138906 190370 613563 190557
rect 138906 190347 145906 190370
rect 109924 190162 116943 190253
rect 109924 190066 110021 190162
rect 5106 189746 14884 190066
rect 104047 189746 110021 190066
rect 5106 180066 10106 189746
rect 109924 189698 110021 189746
rect 116816 189698 116943 190162
rect 109924 189612 116943 189698
rect 119975 188265 607566 188370
rect 119975 185066 120133 188265
rect 104047 184746 120133 185066
rect 119975 183580 120133 184746
rect 126688 188234 607566 188265
rect 126688 183580 139135 188234
rect 119975 183549 139135 183580
rect 145690 188229 607566 188234
rect 145690 188204 602772 188229
rect 145690 183649 388000 188204
rect 393895 183649 602772 188204
rect 145690 183618 602772 183649
rect 607365 183618 607566 188229
rect 145690 183549 607566 183618
rect 119975 183370 607566 183549
rect 109924 180162 116943 180253
rect 109924 180066 110021 180162
rect 5106 179746 14884 180066
rect 104047 179746 110021 180066
rect 5106 170066 10106 179746
rect 109924 179698 110021 179746
rect 116816 179698 116943 180162
rect 109924 179612 116943 179698
rect 129802 176657 136933 176729
rect 129802 176107 130009 176657
rect 136855 176512 136933 176657
rect 608556 176601 613582 176652
rect 608556 176512 608613 176601
rect 136855 176192 153297 176512
rect 600378 176192 608613 176512
rect 136855 176107 136933 176192
rect 129802 176012 136933 176107
rect 608556 176153 608613 176192
rect 613500 176512 613582 176601
rect 613500 176192 613584 176512
rect 613500 176153 613582 176192
rect 608556 176088 613582 176153
rect 119938 175168 126930 175245
rect 119938 175066 120020 175168
rect 104047 174746 120020 175066
rect 119938 174631 120020 174746
rect 126822 175066 126930 175168
rect 126822 174746 126933 175066
rect 126822 174631 126930 174746
rect 119938 174555 126930 174631
rect 109924 170162 116943 170253
rect 109924 170066 110021 170162
rect 5106 169746 14884 170066
rect 104005 169746 110021 170066
rect 5106 160066 10106 169746
rect 109924 169698 110021 169746
rect 116816 169698 116943 170162
rect 109924 169612 116943 169698
rect 119938 165168 126930 165245
rect 119938 165066 120020 165168
rect 104047 164746 120020 165066
rect 119938 164631 120020 164746
rect 126822 165066 126930 165168
rect 126822 164746 126968 165066
rect 126822 164631 126930 164746
rect 119938 164555 126930 164631
rect 138925 163654 145941 163717
rect 138925 163065 138995 163654
rect 145878 163512 145941 163654
rect 602550 163571 607549 163646
rect 602550 163512 602628 163571
rect 145878 163192 153297 163512
rect 600421 163192 602628 163512
rect 145878 163065 145941 163192
rect 602550 163148 602628 163192
rect 607445 163512 607549 163571
rect 607445 163192 607587 163512
rect 607445 163148 607549 163192
rect 602550 163065 607549 163148
rect 138925 163012 145941 163065
rect 109924 160162 116943 160253
rect 109924 160066 110021 160162
rect 5106 159746 14884 160066
rect 104047 159746 110021 160066
rect 5106 150066 10106 159746
rect 109924 159698 110021 159746
rect 116816 159698 116943 160162
rect 109924 159612 116943 159698
rect 119938 155168 126930 155245
rect 119938 155066 120020 155168
rect 104006 154746 120020 155066
rect 119938 154631 120020 154746
rect 126822 155066 126930 155168
rect 126822 154746 126947 155066
rect 126822 154631 126930 154746
rect 119938 154555 126930 154631
rect 129802 150657 136933 150729
rect 109924 150162 116943 150253
rect 109924 150066 110021 150162
rect 5106 149746 14884 150066
rect 104047 149746 110021 150066
rect 5106 140066 10106 149746
rect 109924 149698 110021 149746
rect 116816 150066 116943 150162
rect 129802 150107 130009 150657
rect 136855 150512 136933 150657
rect 608556 150601 613582 150652
rect 608556 150512 608613 150601
rect 136855 150192 153297 150512
rect 600420 150192 608613 150512
rect 136855 150107 136933 150192
rect 116816 149746 116951 150066
rect 129802 150012 136933 150107
rect 608556 150153 608613 150192
rect 613500 150512 613582 150601
rect 613500 150192 613584 150512
rect 613500 150153 613582 150192
rect 608556 150088 613582 150153
rect 116816 149698 116943 149746
rect 109924 149612 116943 149698
rect 119938 145168 126930 145245
rect 119938 145066 120020 145168
rect 104017 144746 120020 145066
rect 119938 144631 120020 144746
rect 126822 145066 126930 145168
rect 126822 144746 126958 145066
rect 126822 144631 126930 144746
rect 119938 144555 126930 144631
rect 109924 140162 116943 140253
rect 109924 140066 110021 140162
rect 5106 139746 14884 140066
rect 104047 139746 110021 140066
rect 5106 130066 10106 139746
rect 109924 139698 110021 139746
rect 116816 139698 116943 140162
rect 109924 139612 116943 139698
rect 138925 137654 145941 137717
rect 138925 137065 138995 137654
rect 145878 137512 145941 137654
rect 602550 137571 607549 137646
rect 602550 137512 602628 137571
rect 145878 137192 153327 137512
rect 600392 137192 602628 137512
rect 145878 137065 145941 137192
rect 602550 137148 602628 137192
rect 607445 137512 607549 137571
rect 607445 137192 607573 137512
rect 607445 137148 607549 137192
rect 602550 137065 607549 137148
rect 138925 137012 145941 137065
rect 119938 135168 126930 135245
rect 119938 135066 120020 135168
rect 104047 134746 120020 135066
rect 119938 134631 120020 134746
rect 126822 135066 126930 135168
rect 126822 134746 126937 135066
rect 126822 134631 126930 134746
rect 119938 134555 126930 134631
rect 109924 130162 116943 130253
rect 109924 130066 110021 130162
rect 5106 129746 14884 130066
rect 104047 129746 110021 130066
rect 5106 120066 10106 129746
rect 109924 129698 110021 129746
rect 116816 130066 116943 130162
rect 116816 129746 116951 130066
rect 116816 129698 116943 129746
rect 109924 129612 116943 129698
rect 119938 125168 126930 125245
rect 119938 125066 120020 125168
rect 104047 124746 120020 125066
rect 119938 124631 120020 124746
rect 126822 125066 126930 125168
rect 126822 124746 126979 125066
rect 126822 124631 126930 124746
rect 119938 124555 126930 124631
rect 129802 124657 136933 124729
rect 129802 124107 130009 124657
rect 136855 124512 136933 124657
rect 608556 124601 613582 124652
rect 608556 124512 608613 124601
rect 136855 124192 153297 124512
rect 600421 124192 608613 124512
rect 136855 124107 136933 124192
rect 129802 124012 136933 124107
rect 608556 124153 608613 124192
rect 613500 124512 613582 124601
rect 613500 124192 613612 124512
rect 613500 124153 613582 124192
rect 608556 124088 613582 124153
rect 109924 120162 116943 120253
rect 109924 120066 110021 120162
rect 5106 119746 14884 120066
rect 104047 119746 110021 120066
rect 5106 110066 10106 119746
rect 109924 119698 110021 119746
rect 116816 119698 116943 120162
rect 109924 119612 116943 119698
rect 119938 115168 126930 115245
rect 119938 115066 120020 115168
rect 104047 114746 120020 115066
rect 119938 114631 120020 114746
rect 126822 115066 126930 115168
rect 126822 114746 126958 115066
rect 126822 114631 126930 114746
rect 119938 114555 126930 114631
rect 138925 111654 145941 111717
rect 138925 111512 138995 111654
rect 138912 111192 138995 111512
rect 138925 111065 138995 111192
rect 145878 111512 145941 111654
rect 602550 111571 607549 111646
rect 602550 111512 602628 111571
rect 145878 111192 153297 111512
rect 600421 111192 602628 111512
rect 145878 111065 145941 111192
rect 602550 111148 602628 111192
rect 607445 111148 607549 111571
rect 602550 111065 607549 111148
rect 138925 111012 145941 111065
rect 109924 110162 116943 110253
rect 109924 110066 110021 110162
rect 5106 109746 14884 110066
rect 104047 109746 110021 110066
rect 5106 100066 10106 109746
rect 109924 109698 110021 109746
rect 116816 110066 116943 110162
rect 116816 109746 116972 110066
rect 116816 109698 116943 109746
rect 109924 109612 116943 109698
rect 119938 105168 126930 105245
rect 119938 105066 120020 105168
rect 104047 104746 120020 105066
rect 119938 104631 120020 104746
rect 126822 105066 126930 105168
rect 126822 104746 126947 105066
rect 126822 104631 126930 104746
rect 119938 104555 126930 104631
rect 109924 100162 116943 100253
rect 109924 100066 110021 100162
rect 5106 99746 14884 100066
rect 104047 99746 110021 100066
rect 5106 98794 10106 99746
rect 109924 99698 110021 99746
rect 116816 99698 116943 100162
rect 109924 99612 116943 99698
rect 4106 93783 10106 98794
rect 129802 98657 136933 98729
rect 129802 98107 130009 98657
rect 136855 98512 136933 98657
rect 608556 98601 613582 98652
rect 608556 98512 608613 98601
rect 136855 98192 153344 98512
rect 600421 98192 608613 98512
rect 136855 98107 136933 98192
rect 129802 98012 136933 98107
rect 608556 98153 608613 98192
rect 613500 98512 613582 98601
rect 613500 98192 613584 98512
rect 613500 98153 613582 98192
rect 608556 98088 613582 98153
rect 119938 95168 126930 95245
rect 119938 95066 120020 95168
rect 103996 94746 120020 95066
rect 119938 94631 120020 94746
rect 126822 95066 126930 95168
rect 126822 94746 126958 95066
rect 126822 94631 126930 94746
rect 119938 94555 126930 94631
rect 4106 90066 9106 93783
rect 109924 90162 116943 90253
rect 109924 90066 110021 90162
rect 4106 89746 14884 90066
rect 104047 89746 110021 90066
rect 4106 80066 9106 89746
rect 109924 89698 110021 89746
rect 116816 90066 116943 90162
rect 116816 89746 116983 90066
rect 116816 89698 116943 89746
rect 109924 89612 116943 89698
rect 138925 85654 145941 85717
rect 138925 85512 138995 85654
rect 119938 85168 126930 85245
rect 138878 85192 138995 85512
rect 119938 85066 120020 85168
rect 104047 84746 120020 85066
rect 119938 84631 120020 84746
rect 126822 85066 126930 85168
rect 126822 84746 126958 85066
rect 138925 85065 138995 85192
rect 145878 85512 145941 85654
rect 602550 85571 607549 85646
rect 602550 85512 602628 85571
rect 145878 85192 153327 85512
rect 600421 85192 602628 85512
rect 145878 85065 145941 85192
rect 602550 85148 602628 85192
rect 607445 85512 607549 85571
rect 607445 85192 607593 85512
rect 607445 85148 607549 85192
rect 602550 85065 607549 85148
rect 138925 85012 145941 85065
rect 126822 84631 126930 84746
rect 119938 84555 126930 84631
rect 109924 80162 116943 80253
rect 109924 80066 110021 80162
rect 4106 79746 14854 80066
rect 104047 79746 110021 80066
rect 4106 70066 9106 79746
rect 109924 79698 110021 79746
rect 116816 79698 116943 80162
rect 109924 79612 116943 79698
rect 628513 75779 631513 75781
rect 614103 75734 635513 75779
rect 119938 75168 126930 75245
rect 119938 75066 120020 75168
rect 104047 74746 120020 75066
rect 119938 74631 120020 74746
rect 126822 75066 126930 75168
rect 126822 74746 126958 75066
rect 126822 74631 126930 74746
rect 614103 74690 614156 75734
rect 615367 74690 635513 75734
rect 614103 74653 635513 74690
rect 628513 74650 631513 74653
rect 119938 74555 126930 74631
rect 129802 72657 136933 72729
rect 129802 72107 130009 72657
rect 136855 72512 136933 72657
rect 608556 72601 613582 72652
rect 608556 72512 608613 72601
rect 136855 72192 153297 72512
rect 600395 72192 608613 72512
rect 136855 72107 136933 72192
rect 129802 72012 136933 72107
rect 608556 72153 608613 72192
rect 613500 72512 613582 72601
rect 613500 72192 613584 72512
rect 613500 72153 613582 72192
rect 608556 72088 613582 72153
rect 109924 70162 116943 70253
rect 109924 70066 110021 70162
rect 4106 69746 14854 70066
rect 104047 69746 110021 70066
rect 4106 60066 9106 69746
rect 109924 69698 110021 69746
rect 116816 69698 116943 70162
rect 109924 69612 116943 69698
rect 608537 65265 613556 65312
rect 119938 65168 126930 65245
rect 119938 65066 120020 65168
rect 104027 64746 120020 65066
rect 119938 64631 120020 64746
rect 126822 65066 126930 65168
rect 126822 64746 126947 65066
rect 126822 64631 126930 64746
rect 119938 64555 126930 64631
rect 608537 64636 608612 65265
rect 613504 65160 613556 65265
rect 613504 65118 624709 65160
rect 613504 64798 622897 65118
rect 624672 64798 624709 65118
rect 613504 64760 624709 64798
rect 613504 64636 613556 64760
rect 608537 64599 613556 64636
rect 614106 63098 631513 63171
rect 614106 61750 614165 63098
rect 615335 61750 631513 63098
rect 614106 61685 631513 61750
rect 109924 60162 116943 60253
rect 109924 60066 110021 60162
rect 4106 59746 14854 60066
rect 104047 59746 110021 60066
rect 4106 50066 9106 59746
rect 109924 59698 110021 59746
rect 116816 60066 116943 60162
rect 116816 59746 116983 60066
rect 116816 59698 116943 59746
rect 109924 59612 116943 59698
rect 138925 59654 145941 59717
rect 138925 59065 138995 59654
rect 145878 59512 145941 59654
rect 602550 59571 607549 59646
rect 602550 59512 602628 59571
rect 145878 59192 153302 59512
rect 600406 59192 602628 59512
rect 145878 59065 145941 59192
rect 602550 59148 602628 59192
rect 607445 59148 607549 59571
rect 602550 59065 607549 59148
rect 138925 59012 145941 59065
rect 119938 55168 126930 55245
rect 119938 55066 120020 55168
rect 104047 54746 120020 55066
rect 119938 54631 120020 54746
rect 126822 55066 126930 55168
rect 126822 54746 126979 55066
rect 126822 54631 126930 54746
rect 119938 54555 126930 54631
rect 109924 50162 116943 50253
rect 109924 50066 110021 50162
rect 4106 49746 14854 50066
rect 103996 49746 110021 50066
rect 4106 43927 9106 49746
rect 109924 49698 110021 49746
rect 116816 49698 116943 50162
rect 109924 49612 116943 49698
rect 608557 47558 613537 47628
rect 608557 47498 608618 47558
rect 601533 47418 608618 47498
rect 601528 47178 608618 47418
rect 129802 46657 136933 46729
rect 129802 46107 130009 46657
rect 136855 46512 136933 46657
rect 601528 46512 601848 47178
rect 608557 47085 608618 47178
rect 613452 47498 613537 47558
rect 613452 47178 619487 47498
rect 613452 47085 613537 47178
rect 608557 47039 613537 47085
rect 136855 46192 153355 46512
rect 600421 46192 601848 46512
rect 602565 46757 607545 46812
rect 602565 46284 602636 46757
rect 607470 46682 607545 46757
rect 607470 46362 619530 46682
rect 607470 46284 607545 46362
rect 602565 46223 607545 46284
rect 136855 46107 136933 46192
rect 129802 46012 136933 46107
rect 608567 45911 613547 45972
rect 608567 45438 608633 45911
rect 613467 45866 613547 45911
rect 613467 45546 619512 45866
rect 613467 45438 613547 45546
rect 608567 45383 613547 45438
rect 119938 45168 126930 45245
rect 119938 45066 120020 45168
rect 103967 44746 120020 45066
rect 119938 44631 120020 44746
rect 126822 45066 126930 45168
rect 602560 45120 607540 45171
rect 126822 44746 126933 45066
rect 126822 44631 126930 44746
rect 119938 44555 126930 44631
rect 602560 44647 602600 45120
rect 607434 45050 607540 45120
rect 607434 44730 619487 45050
rect 607434 44647 607540 44730
rect 602560 44582 607540 44647
rect 608552 44256 613571 44314
rect 608552 44234 608607 44256
rect 4106 39598 4302 43927
rect 8940 40066 9106 43927
rect 608551 43914 608607 44234
rect 608552 43861 608607 43914
rect 613498 44234 613571 44256
rect 613498 43914 619487 44234
rect 613498 43861 613571 43914
rect 608552 43813 613571 43861
rect 109924 40162 116943 40253
rect 109924 40066 110021 40162
rect 8940 39746 14854 40066
rect 103764 39746 110021 40066
rect 8940 39598 9106 39746
rect 109924 39698 110021 39746
rect 116816 40066 116943 40162
rect 116816 39746 116988 40066
rect 116816 39698 116943 39746
rect 109924 39612 116943 39698
rect 4106 33967 9106 39598
rect 119938 35168 126930 35245
rect 119938 35066 120020 35168
rect 103906 34746 120020 35066
rect 119938 34631 120020 34746
rect 126822 35066 126930 35168
rect 126822 34746 126933 35066
rect 126822 34631 126930 34746
rect 119938 34555 126930 34631
rect 4106 29638 4280 33967
rect 8918 30314 9106 33967
rect 138925 33654 145941 33717
rect 138925 33065 138995 33654
rect 145878 33512 145941 33654
rect 602565 33615 607553 33681
rect 602565 33512 602623 33615
rect 145878 33192 153446 33512
rect 600415 33192 602623 33512
rect 145878 33065 145941 33192
rect 138925 33012 145941 33065
rect 602565 33085 602623 33192
rect 607495 33512 607553 33615
rect 607495 33192 607560 33512
rect 607495 33085 607553 33192
rect 602565 33039 607553 33085
rect 8917 30066 9106 30314
rect 109924 30162 116943 30253
rect 109924 30066 110021 30162
rect 8917 29746 14854 30066
rect 104047 29746 110021 30066
rect 8917 29638 9106 29746
rect 4106 20066 9106 29638
rect 109924 29698 110021 29746
rect 116816 29698 116943 30162
rect 109924 29612 116943 29698
rect 129908 29832 136938 29895
rect 129908 29243 129997 29832
rect 136890 29708 136938 29832
rect 136890 29388 149780 29708
rect 136890 29243 136938 29388
rect 129908 29189 136938 29243
rect 119814 26804 145999 26947
rect 119814 26772 139167 26804
rect 119814 25066 120212 26772
rect 103886 24746 120212 25066
rect 119814 22141 120212 24746
rect 126733 22173 139167 26772
rect 145688 22173 145999 26804
rect 126733 22141 145999 22173
rect 119814 21947 145999 22141
rect 109924 20162 116943 20253
rect 109924 20066 110021 20162
rect 4106 19746 14854 20066
rect 104021 19746 110021 20066
rect 4106 14415 9106 19746
rect 109924 19698 110021 19746
rect 116816 19698 116943 20162
rect 109924 19612 116943 19698
rect 140999 16289 145999 21947
rect 149460 20512 149780 29388
rect 608551 20655 613551 20812
rect 608551 20512 608661 20655
rect 149460 20192 153471 20512
rect 600421 20192 608661 20512
rect 104033 16287 145999 16289
rect 103984 16262 145999 16287
rect 103984 15523 104025 16262
rect 104608 15523 145999 16262
rect 103984 15490 145999 15523
rect 104033 15489 145999 15490
rect 140999 15415 145999 15489
rect 602560 18529 607560 18653
rect 602560 15415 602693 18529
rect 140999 15232 602693 15415
rect 131993 14415 136993 14418
rect 4106 14272 136993 14415
rect 4106 13315 110144 14272
rect 4106 12252 105051 13315
rect 105711 12252 110144 13315
rect 4106 9641 110144 12252
rect 116665 14174 136993 14272
rect 116665 9641 130166 14174
rect 4106 9543 130166 9641
rect 136687 9543 136993 14174
rect 140999 10634 202782 15232
rect 207285 15200 602693 15232
rect 207285 10634 212877 15200
rect 140999 10602 212877 10634
rect 217380 14168 602693 15200
rect 607423 14168 607560 18529
rect 217380 10602 607560 14168
rect 140999 10415 607560 10602
rect 608551 16294 608661 20192
rect 613391 16294 613551 20655
rect 4106 9415 136993 9543
rect 131993 8415 136993 9415
rect 608551 8415 613551 16294
rect 131993 3415 613551 8415
rect 628513 11787 631513 61685
rect 628513 7973 628597 11787
rect 631428 7973 631513 11787
rect 628513 7887 631513 7973
rect 632513 6588 635513 74653
rect 632513 2815 632642 6588
rect 635402 2815 635513 6588
rect 632513 2669 635513 2815
<< labels >>
flabel metal5 145438 217320 145438 217320 0 FreeSans 8000 0 0 0 VSSA2
flabel metal5 144640 219774 144640 219774 0 FreeSans 8000 0 0 0 VDDA2
flabel metal5 144395 222474 144395 222474 0 FreeSans 8000 0 0 0 VSSD2
flabel metal5 146359 224867 146359 224867 0 FreeSans 8000 0 0 0 VCCD2
flabel metal5 147893 204740 147893 204740 0 FreeSans 8000 0 0 0 VCCD
flabel metal5 379355 202224 379355 202224 0 FreeSans 8000 0 0 0 VSSD
flabel metal5 379539 207256 379539 207256 0 FreeSans 8000 0 0 0 VSSA1
flabel metal5 379232 209895 379232 209895 0 FreeSans 8000 0 0 0 VDDA1
flabel metal5 378925 212288 378925 212288 0 FreeSans 8000 0 0 0 VSSD1
flabel metal5 378557 214804 378557 214804 0 FreeSans 8000 0 0 0 VCCD1
<< end >>
