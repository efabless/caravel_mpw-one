VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel
  CLASS BLOCK ;
  FOREIGN caravel ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.010 BY 5188.010 ;
  OBS
      LAYER li1 ;
        RECT 0.225 0.225 3587.785 5187.715 ;
      LAYER met1 ;
        RECT 0.000 0.000 3588.010 5188.010 ;
      LAYER met2 ;
        RECT 0.000 0.000 3588.010 5188.010 ;
      LAYER met3 ;
        RECT 0.000 0.000 3588.010 5188.010 ;
      LAYER met4 ;
        RECT 0.000 0.000 3588.010 5188.010 ;
      LAYER met5 ;
        RECT 0.000 0.000 3588.010 5188.010 ;
  END
END caravel
END LIBRARY

