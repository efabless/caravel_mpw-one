magic
tech sky130A
magscale 1 2
timestamp 1606421840
<< error_p >>
rect -7050 799 -6992 805
rect -6932 799 -6874 805
rect -6814 799 -6756 805
rect -6696 799 -6638 805
rect -6578 799 -6520 805
rect -6460 799 -6402 805
rect -6342 799 -6284 805
rect -6224 799 -6166 805
rect -6106 799 -6048 805
rect -5988 799 -5930 805
rect -5870 799 -5812 805
rect -5752 799 -5694 805
rect -5634 799 -5576 805
rect -5516 799 -5458 805
rect -5398 799 -5340 805
rect -5280 799 -5222 805
rect -5162 799 -5104 805
rect -5044 799 -4986 805
rect -4926 799 -4868 805
rect -4808 799 -4750 805
rect -4690 799 -4632 805
rect -4572 799 -4514 805
rect -4454 799 -4396 805
rect -4336 799 -4278 805
rect -4218 799 -4160 805
rect -4100 799 -4042 805
rect -3982 799 -3924 805
rect -3864 799 -3806 805
rect -3746 799 -3688 805
rect -3628 799 -3570 805
rect -3510 799 -3452 805
rect -3392 799 -3334 805
rect -3274 799 -3216 805
rect -3156 799 -3098 805
rect -3038 799 -2980 805
rect -2920 799 -2862 805
rect -2802 799 -2744 805
rect -2684 799 -2626 805
rect -2566 799 -2508 805
rect -2448 799 -2390 805
rect -2330 799 -2272 805
rect -2212 799 -2154 805
rect -2094 799 -2036 805
rect -1976 799 -1918 805
rect -1858 799 -1800 805
rect -1740 799 -1682 805
rect -1622 799 -1564 805
rect -1504 799 -1446 805
rect -1386 799 -1328 805
rect -1268 799 -1210 805
rect -1150 799 -1092 805
rect -1032 799 -974 805
rect -914 799 -856 805
rect -796 799 -738 805
rect -678 799 -620 805
rect -560 799 -502 805
rect -442 799 -384 805
rect -324 799 -266 805
rect -206 799 -148 805
rect -88 799 -30 805
rect 30 799 88 805
rect 148 799 206 805
rect 266 799 324 805
rect 384 799 442 805
rect 502 799 560 805
rect 620 799 678 805
rect 738 799 796 805
rect 856 799 914 805
rect 974 799 1032 805
rect 1092 799 1150 805
rect 1210 799 1268 805
rect 1328 799 1386 805
rect 1446 799 1504 805
rect 1564 799 1622 805
rect 1682 799 1740 805
rect 1800 799 1858 805
rect 1918 799 1976 805
rect 2036 799 2094 805
rect 2154 799 2212 805
rect 2272 799 2330 805
rect 2390 799 2448 805
rect 2508 799 2566 805
rect 2626 799 2684 805
rect 2744 799 2802 805
rect 2862 799 2920 805
rect 2980 799 3038 805
rect 3098 799 3156 805
rect 3216 799 3274 805
rect 3334 799 3392 805
rect 3452 799 3510 805
rect 3570 799 3628 805
rect 3688 799 3746 805
rect 3806 799 3864 805
rect 3924 799 3982 805
rect 4042 799 4100 805
rect 4160 799 4218 805
rect 4278 799 4336 805
rect 4396 799 4454 805
rect 4514 799 4572 805
rect 4632 799 4690 805
rect 4750 799 4808 805
rect 4868 799 4926 805
rect 4986 799 5044 805
rect 5104 799 5162 805
rect 5222 799 5280 805
rect 5340 799 5398 805
rect 5458 799 5516 805
rect 5576 799 5634 805
rect 5694 799 5752 805
rect 5812 799 5870 805
rect 5930 799 5988 805
rect 6048 799 6106 805
rect 6166 799 6224 805
rect 6284 799 6342 805
rect 6402 799 6460 805
rect 6520 799 6578 805
rect 6638 799 6696 805
rect 6756 799 6814 805
rect 6874 799 6932 805
rect 6992 799 7050 805
rect -7050 765 -7038 799
rect -6932 765 -6920 799
rect -6814 765 -6802 799
rect -6696 765 -6684 799
rect -6578 765 -6566 799
rect -6460 765 -6448 799
rect -6342 765 -6330 799
rect -6224 765 -6212 799
rect -6106 765 -6094 799
rect -5988 765 -5976 799
rect -5870 765 -5858 799
rect -5752 765 -5740 799
rect -5634 765 -5622 799
rect -5516 765 -5504 799
rect -5398 765 -5386 799
rect -5280 765 -5268 799
rect -5162 765 -5150 799
rect -5044 765 -5032 799
rect -4926 765 -4914 799
rect -4808 765 -4796 799
rect -4690 765 -4678 799
rect -4572 765 -4560 799
rect -4454 765 -4442 799
rect -4336 765 -4324 799
rect -4218 765 -4206 799
rect -4100 765 -4088 799
rect -3982 765 -3970 799
rect -3864 765 -3852 799
rect -3746 765 -3734 799
rect -3628 765 -3616 799
rect -3510 765 -3498 799
rect -3392 765 -3380 799
rect -3274 765 -3262 799
rect -3156 765 -3144 799
rect -3038 765 -3026 799
rect -2920 765 -2908 799
rect -2802 765 -2790 799
rect -2684 765 -2672 799
rect -2566 765 -2554 799
rect -2448 765 -2436 799
rect -2330 765 -2318 799
rect -2212 765 -2200 799
rect -2094 765 -2082 799
rect -1976 765 -1964 799
rect -1858 765 -1846 799
rect -1740 765 -1728 799
rect -1622 765 -1610 799
rect -1504 765 -1492 799
rect -1386 765 -1374 799
rect -1268 765 -1256 799
rect -1150 765 -1138 799
rect -1032 765 -1020 799
rect -914 765 -902 799
rect -796 765 -784 799
rect -678 765 -666 799
rect -560 765 -548 799
rect -442 765 -430 799
rect -324 765 -312 799
rect -206 765 -194 799
rect -88 765 -76 799
rect 30 765 42 799
rect 148 765 160 799
rect 266 765 278 799
rect 384 765 396 799
rect 502 765 514 799
rect 620 765 632 799
rect 738 765 750 799
rect 856 765 868 799
rect 974 765 986 799
rect 1092 765 1104 799
rect 1210 765 1222 799
rect 1328 765 1340 799
rect 1446 765 1458 799
rect 1564 765 1576 799
rect 1682 765 1694 799
rect 1800 765 1812 799
rect 1918 765 1930 799
rect 2036 765 2048 799
rect 2154 765 2166 799
rect 2272 765 2284 799
rect 2390 765 2402 799
rect 2508 765 2520 799
rect 2626 765 2638 799
rect 2744 765 2756 799
rect 2862 765 2874 799
rect 2980 765 2992 799
rect 3098 765 3110 799
rect 3216 765 3228 799
rect 3334 765 3346 799
rect 3452 765 3464 799
rect 3570 765 3582 799
rect 3688 765 3700 799
rect 3806 765 3818 799
rect 3924 765 3936 799
rect 4042 765 4054 799
rect 4160 765 4172 799
rect 4278 765 4290 799
rect 4396 765 4408 799
rect 4514 765 4526 799
rect 4632 765 4644 799
rect 4750 765 4762 799
rect 4868 765 4880 799
rect 4986 765 4998 799
rect 5104 765 5116 799
rect 5222 765 5234 799
rect 5340 765 5352 799
rect 5458 765 5470 799
rect 5576 765 5588 799
rect 5694 765 5706 799
rect 5812 765 5824 799
rect 5930 765 5942 799
rect 6048 765 6060 799
rect 6166 765 6178 799
rect 6284 765 6296 799
rect 6402 765 6414 799
rect 6520 765 6532 799
rect 6638 765 6650 799
rect 6756 765 6768 799
rect 6874 765 6886 799
rect 6992 765 7004 799
rect -7050 759 -6992 765
rect -6932 759 -6874 765
rect -6814 759 -6756 765
rect -6696 759 -6638 765
rect -6578 759 -6520 765
rect -6460 759 -6402 765
rect -6342 759 -6284 765
rect -6224 759 -6166 765
rect -6106 759 -6048 765
rect -5988 759 -5930 765
rect -5870 759 -5812 765
rect -5752 759 -5694 765
rect -5634 759 -5576 765
rect -5516 759 -5458 765
rect -5398 759 -5340 765
rect -5280 759 -5222 765
rect -5162 759 -5104 765
rect -5044 759 -4986 765
rect -4926 759 -4868 765
rect -4808 759 -4750 765
rect -4690 759 -4632 765
rect -4572 759 -4514 765
rect -4454 759 -4396 765
rect -4336 759 -4278 765
rect -4218 759 -4160 765
rect -4100 759 -4042 765
rect -3982 759 -3924 765
rect -3864 759 -3806 765
rect -3746 759 -3688 765
rect -3628 759 -3570 765
rect -3510 759 -3452 765
rect -3392 759 -3334 765
rect -3274 759 -3216 765
rect -3156 759 -3098 765
rect -3038 759 -2980 765
rect -2920 759 -2862 765
rect -2802 759 -2744 765
rect -2684 759 -2626 765
rect -2566 759 -2508 765
rect -2448 759 -2390 765
rect -2330 759 -2272 765
rect -2212 759 -2154 765
rect -2094 759 -2036 765
rect -1976 759 -1918 765
rect -1858 759 -1800 765
rect -1740 759 -1682 765
rect -1622 759 -1564 765
rect -1504 759 -1446 765
rect -1386 759 -1328 765
rect -1268 759 -1210 765
rect -1150 759 -1092 765
rect -1032 759 -974 765
rect -914 759 -856 765
rect -796 759 -738 765
rect -678 759 -620 765
rect -560 759 -502 765
rect -442 759 -384 765
rect -324 759 -266 765
rect -206 759 -148 765
rect -88 759 -30 765
rect 30 759 88 765
rect 148 759 206 765
rect 266 759 324 765
rect 384 759 442 765
rect 502 759 560 765
rect 620 759 678 765
rect 738 759 796 765
rect 856 759 914 765
rect 974 759 1032 765
rect 1092 759 1150 765
rect 1210 759 1268 765
rect 1328 759 1386 765
rect 1446 759 1504 765
rect 1564 759 1622 765
rect 1682 759 1740 765
rect 1800 759 1858 765
rect 1918 759 1976 765
rect 2036 759 2094 765
rect 2154 759 2212 765
rect 2272 759 2330 765
rect 2390 759 2448 765
rect 2508 759 2566 765
rect 2626 759 2684 765
rect 2744 759 2802 765
rect 2862 759 2920 765
rect 2980 759 3038 765
rect 3098 759 3156 765
rect 3216 759 3274 765
rect 3334 759 3392 765
rect 3452 759 3510 765
rect 3570 759 3628 765
rect 3688 759 3746 765
rect 3806 759 3864 765
rect 3924 759 3982 765
rect 4042 759 4100 765
rect 4160 759 4218 765
rect 4278 759 4336 765
rect 4396 759 4454 765
rect 4514 759 4572 765
rect 4632 759 4690 765
rect 4750 759 4808 765
rect 4868 759 4926 765
rect 4986 759 5044 765
rect 5104 759 5162 765
rect 5222 759 5280 765
rect 5340 759 5398 765
rect 5458 759 5516 765
rect 5576 759 5634 765
rect 5694 759 5752 765
rect 5812 759 5870 765
rect 5930 759 5988 765
rect 6048 759 6106 765
rect 6166 759 6224 765
rect 6284 759 6342 765
rect 6402 759 6460 765
rect 6520 759 6578 765
rect 6638 759 6696 765
rect 6756 759 6814 765
rect 6874 759 6932 765
rect 6992 759 7050 765
rect -7050 71 -6992 77
rect -6932 71 -6874 77
rect -6814 71 -6756 77
rect -6696 71 -6638 77
rect -6578 71 -6520 77
rect -6460 71 -6402 77
rect -6342 71 -6284 77
rect -6224 71 -6166 77
rect -6106 71 -6048 77
rect -5988 71 -5930 77
rect -5870 71 -5812 77
rect -5752 71 -5694 77
rect -5634 71 -5576 77
rect -5516 71 -5458 77
rect -5398 71 -5340 77
rect -5280 71 -5222 77
rect -5162 71 -5104 77
rect -5044 71 -4986 77
rect -4926 71 -4868 77
rect -4808 71 -4750 77
rect -4690 71 -4632 77
rect -4572 71 -4514 77
rect -4454 71 -4396 77
rect -4336 71 -4278 77
rect -4218 71 -4160 77
rect -4100 71 -4042 77
rect -3982 71 -3924 77
rect -3864 71 -3806 77
rect -3746 71 -3688 77
rect -3628 71 -3570 77
rect -3510 71 -3452 77
rect -3392 71 -3334 77
rect -3274 71 -3216 77
rect -3156 71 -3098 77
rect -3038 71 -2980 77
rect -2920 71 -2862 77
rect -2802 71 -2744 77
rect -2684 71 -2626 77
rect -2566 71 -2508 77
rect -2448 71 -2390 77
rect -2330 71 -2272 77
rect -2212 71 -2154 77
rect -2094 71 -2036 77
rect -1976 71 -1918 77
rect -1858 71 -1800 77
rect -1740 71 -1682 77
rect -1622 71 -1564 77
rect -1504 71 -1446 77
rect -1386 71 -1328 77
rect -1268 71 -1210 77
rect -1150 71 -1092 77
rect -1032 71 -974 77
rect -914 71 -856 77
rect -796 71 -738 77
rect -678 71 -620 77
rect -560 71 -502 77
rect -442 71 -384 77
rect -324 71 -266 77
rect -206 71 -148 77
rect -88 71 -30 77
rect 30 71 88 77
rect 148 71 206 77
rect 266 71 324 77
rect 384 71 442 77
rect 502 71 560 77
rect 620 71 678 77
rect 738 71 796 77
rect 856 71 914 77
rect 974 71 1032 77
rect 1092 71 1150 77
rect 1210 71 1268 77
rect 1328 71 1386 77
rect 1446 71 1504 77
rect 1564 71 1622 77
rect 1682 71 1740 77
rect 1800 71 1858 77
rect 1918 71 1976 77
rect 2036 71 2094 77
rect 2154 71 2212 77
rect 2272 71 2330 77
rect 2390 71 2448 77
rect 2508 71 2566 77
rect 2626 71 2684 77
rect 2744 71 2802 77
rect 2862 71 2920 77
rect 2980 71 3038 77
rect 3098 71 3156 77
rect 3216 71 3274 77
rect 3334 71 3392 77
rect 3452 71 3510 77
rect 3570 71 3628 77
rect 3688 71 3746 77
rect 3806 71 3864 77
rect 3924 71 3982 77
rect 4042 71 4100 77
rect 4160 71 4218 77
rect 4278 71 4336 77
rect 4396 71 4454 77
rect 4514 71 4572 77
rect 4632 71 4690 77
rect 4750 71 4808 77
rect 4868 71 4926 77
rect 4986 71 5044 77
rect 5104 71 5162 77
rect 5222 71 5280 77
rect 5340 71 5398 77
rect 5458 71 5516 77
rect 5576 71 5634 77
rect 5694 71 5752 77
rect 5812 71 5870 77
rect 5930 71 5988 77
rect 6048 71 6106 77
rect 6166 71 6224 77
rect 6284 71 6342 77
rect 6402 71 6460 77
rect 6520 71 6578 77
rect 6638 71 6696 77
rect 6756 71 6814 77
rect 6874 71 6932 77
rect 6992 71 7050 77
rect -7050 37 -7038 71
rect -6932 37 -6920 71
rect -6814 37 -6802 71
rect -6696 37 -6684 71
rect -6578 37 -6566 71
rect -6460 37 -6448 71
rect -6342 37 -6330 71
rect -6224 37 -6212 71
rect -6106 37 -6094 71
rect -5988 37 -5976 71
rect -5870 37 -5858 71
rect -5752 37 -5740 71
rect -5634 37 -5622 71
rect -5516 37 -5504 71
rect -5398 37 -5386 71
rect -5280 37 -5268 71
rect -5162 37 -5150 71
rect -5044 37 -5032 71
rect -4926 37 -4914 71
rect -4808 37 -4796 71
rect -4690 37 -4678 71
rect -4572 37 -4560 71
rect -4454 37 -4442 71
rect -4336 37 -4324 71
rect -4218 37 -4206 71
rect -4100 37 -4088 71
rect -3982 37 -3970 71
rect -3864 37 -3852 71
rect -3746 37 -3734 71
rect -3628 37 -3616 71
rect -3510 37 -3498 71
rect -3392 37 -3380 71
rect -3274 37 -3262 71
rect -3156 37 -3144 71
rect -3038 37 -3026 71
rect -2920 37 -2908 71
rect -2802 37 -2790 71
rect -2684 37 -2672 71
rect -2566 37 -2554 71
rect -2448 37 -2436 71
rect -2330 37 -2318 71
rect -2212 37 -2200 71
rect -2094 37 -2082 71
rect -1976 37 -1964 71
rect -1858 37 -1846 71
rect -1740 37 -1728 71
rect -1622 37 -1610 71
rect -1504 37 -1492 71
rect -1386 37 -1374 71
rect -1268 37 -1256 71
rect -1150 37 -1138 71
rect -1032 37 -1020 71
rect -914 37 -902 71
rect -796 37 -784 71
rect -678 37 -666 71
rect -560 37 -548 71
rect -442 37 -430 71
rect -324 37 -312 71
rect -206 37 -194 71
rect -88 37 -76 71
rect 30 37 42 71
rect 148 37 160 71
rect 266 37 278 71
rect 384 37 396 71
rect 502 37 514 71
rect 620 37 632 71
rect 738 37 750 71
rect 856 37 868 71
rect 974 37 986 71
rect 1092 37 1104 71
rect 1210 37 1222 71
rect 1328 37 1340 71
rect 1446 37 1458 71
rect 1564 37 1576 71
rect 1682 37 1694 71
rect 1800 37 1812 71
rect 1918 37 1930 71
rect 2036 37 2048 71
rect 2154 37 2166 71
rect 2272 37 2284 71
rect 2390 37 2402 71
rect 2508 37 2520 71
rect 2626 37 2638 71
rect 2744 37 2756 71
rect 2862 37 2874 71
rect 2980 37 2992 71
rect 3098 37 3110 71
rect 3216 37 3228 71
rect 3334 37 3346 71
rect 3452 37 3464 71
rect 3570 37 3582 71
rect 3688 37 3700 71
rect 3806 37 3818 71
rect 3924 37 3936 71
rect 4042 37 4054 71
rect 4160 37 4172 71
rect 4278 37 4290 71
rect 4396 37 4408 71
rect 4514 37 4526 71
rect 4632 37 4644 71
rect 4750 37 4762 71
rect 4868 37 4880 71
rect 4986 37 4998 71
rect 5104 37 5116 71
rect 5222 37 5234 71
rect 5340 37 5352 71
rect 5458 37 5470 71
rect 5576 37 5588 71
rect 5694 37 5706 71
rect 5812 37 5824 71
rect 5930 37 5942 71
rect 6048 37 6060 71
rect 6166 37 6178 71
rect 6284 37 6296 71
rect 6402 37 6414 71
rect 6520 37 6532 71
rect 6638 37 6650 71
rect 6756 37 6768 71
rect 6874 37 6886 71
rect 6992 37 7004 71
rect -7050 31 -6992 37
rect -6932 31 -6874 37
rect -6814 31 -6756 37
rect -6696 31 -6638 37
rect -6578 31 -6520 37
rect -6460 31 -6402 37
rect -6342 31 -6284 37
rect -6224 31 -6166 37
rect -6106 31 -6048 37
rect -5988 31 -5930 37
rect -5870 31 -5812 37
rect -5752 31 -5694 37
rect -5634 31 -5576 37
rect -5516 31 -5458 37
rect -5398 31 -5340 37
rect -5280 31 -5222 37
rect -5162 31 -5104 37
rect -5044 31 -4986 37
rect -4926 31 -4868 37
rect -4808 31 -4750 37
rect -4690 31 -4632 37
rect -4572 31 -4514 37
rect -4454 31 -4396 37
rect -4336 31 -4278 37
rect -4218 31 -4160 37
rect -4100 31 -4042 37
rect -3982 31 -3924 37
rect -3864 31 -3806 37
rect -3746 31 -3688 37
rect -3628 31 -3570 37
rect -3510 31 -3452 37
rect -3392 31 -3334 37
rect -3274 31 -3216 37
rect -3156 31 -3098 37
rect -3038 31 -2980 37
rect -2920 31 -2862 37
rect -2802 31 -2744 37
rect -2684 31 -2626 37
rect -2566 31 -2508 37
rect -2448 31 -2390 37
rect -2330 31 -2272 37
rect -2212 31 -2154 37
rect -2094 31 -2036 37
rect -1976 31 -1918 37
rect -1858 31 -1800 37
rect -1740 31 -1682 37
rect -1622 31 -1564 37
rect -1504 31 -1446 37
rect -1386 31 -1328 37
rect -1268 31 -1210 37
rect -1150 31 -1092 37
rect -1032 31 -974 37
rect -914 31 -856 37
rect -796 31 -738 37
rect -678 31 -620 37
rect -560 31 -502 37
rect -442 31 -384 37
rect -324 31 -266 37
rect -206 31 -148 37
rect -88 31 -30 37
rect 30 31 88 37
rect 148 31 206 37
rect 266 31 324 37
rect 384 31 442 37
rect 502 31 560 37
rect 620 31 678 37
rect 738 31 796 37
rect 856 31 914 37
rect 974 31 1032 37
rect 1092 31 1150 37
rect 1210 31 1268 37
rect 1328 31 1386 37
rect 1446 31 1504 37
rect 1564 31 1622 37
rect 1682 31 1740 37
rect 1800 31 1858 37
rect 1918 31 1976 37
rect 2036 31 2094 37
rect 2154 31 2212 37
rect 2272 31 2330 37
rect 2390 31 2448 37
rect 2508 31 2566 37
rect 2626 31 2684 37
rect 2744 31 2802 37
rect 2862 31 2920 37
rect 2980 31 3038 37
rect 3098 31 3156 37
rect 3216 31 3274 37
rect 3334 31 3392 37
rect 3452 31 3510 37
rect 3570 31 3628 37
rect 3688 31 3746 37
rect 3806 31 3864 37
rect 3924 31 3982 37
rect 4042 31 4100 37
rect 4160 31 4218 37
rect 4278 31 4336 37
rect 4396 31 4454 37
rect 4514 31 4572 37
rect 4632 31 4690 37
rect 4750 31 4808 37
rect 4868 31 4926 37
rect 4986 31 5044 37
rect 5104 31 5162 37
rect 5222 31 5280 37
rect 5340 31 5398 37
rect 5458 31 5516 37
rect 5576 31 5634 37
rect 5694 31 5752 37
rect 5812 31 5870 37
rect 5930 31 5988 37
rect 6048 31 6106 37
rect 6166 31 6224 37
rect 6284 31 6342 37
rect 6402 31 6460 37
rect 6520 31 6578 37
rect 6638 31 6696 37
rect 6756 31 6814 37
rect 6874 31 6932 37
rect 6992 31 7050 37
rect -7050 -37 -6992 -31
rect -6932 -37 -6874 -31
rect -6814 -37 -6756 -31
rect -6696 -37 -6638 -31
rect -6578 -37 -6520 -31
rect -6460 -37 -6402 -31
rect -6342 -37 -6284 -31
rect -6224 -37 -6166 -31
rect -6106 -37 -6048 -31
rect -5988 -37 -5930 -31
rect -5870 -37 -5812 -31
rect -5752 -37 -5694 -31
rect -5634 -37 -5576 -31
rect -5516 -37 -5458 -31
rect -5398 -37 -5340 -31
rect -5280 -37 -5222 -31
rect -5162 -37 -5104 -31
rect -5044 -37 -4986 -31
rect -4926 -37 -4868 -31
rect -4808 -37 -4750 -31
rect -4690 -37 -4632 -31
rect -4572 -37 -4514 -31
rect -4454 -37 -4396 -31
rect -4336 -37 -4278 -31
rect -4218 -37 -4160 -31
rect -4100 -37 -4042 -31
rect -3982 -37 -3924 -31
rect -3864 -37 -3806 -31
rect -3746 -37 -3688 -31
rect -3628 -37 -3570 -31
rect -3510 -37 -3452 -31
rect -3392 -37 -3334 -31
rect -3274 -37 -3216 -31
rect -3156 -37 -3098 -31
rect -3038 -37 -2980 -31
rect -2920 -37 -2862 -31
rect -2802 -37 -2744 -31
rect -2684 -37 -2626 -31
rect -2566 -37 -2508 -31
rect -2448 -37 -2390 -31
rect -2330 -37 -2272 -31
rect -2212 -37 -2154 -31
rect -2094 -37 -2036 -31
rect -1976 -37 -1918 -31
rect -1858 -37 -1800 -31
rect -1740 -37 -1682 -31
rect -1622 -37 -1564 -31
rect -1504 -37 -1446 -31
rect -1386 -37 -1328 -31
rect -1268 -37 -1210 -31
rect -1150 -37 -1092 -31
rect -1032 -37 -974 -31
rect -914 -37 -856 -31
rect -796 -37 -738 -31
rect -678 -37 -620 -31
rect -560 -37 -502 -31
rect -442 -37 -384 -31
rect -324 -37 -266 -31
rect -206 -37 -148 -31
rect -88 -37 -30 -31
rect 30 -37 88 -31
rect 148 -37 206 -31
rect 266 -37 324 -31
rect 384 -37 442 -31
rect 502 -37 560 -31
rect 620 -37 678 -31
rect 738 -37 796 -31
rect 856 -37 914 -31
rect 974 -37 1032 -31
rect 1092 -37 1150 -31
rect 1210 -37 1268 -31
rect 1328 -37 1386 -31
rect 1446 -37 1504 -31
rect 1564 -37 1622 -31
rect 1682 -37 1740 -31
rect 1800 -37 1858 -31
rect 1918 -37 1976 -31
rect 2036 -37 2094 -31
rect 2154 -37 2212 -31
rect 2272 -37 2330 -31
rect 2390 -37 2448 -31
rect 2508 -37 2566 -31
rect 2626 -37 2684 -31
rect 2744 -37 2802 -31
rect 2862 -37 2920 -31
rect 2980 -37 3038 -31
rect 3098 -37 3156 -31
rect 3216 -37 3274 -31
rect 3334 -37 3392 -31
rect 3452 -37 3510 -31
rect 3570 -37 3628 -31
rect 3688 -37 3746 -31
rect 3806 -37 3864 -31
rect 3924 -37 3982 -31
rect 4042 -37 4100 -31
rect 4160 -37 4218 -31
rect 4278 -37 4336 -31
rect 4396 -37 4454 -31
rect 4514 -37 4572 -31
rect 4632 -37 4690 -31
rect 4750 -37 4808 -31
rect 4868 -37 4926 -31
rect 4986 -37 5044 -31
rect 5104 -37 5162 -31
rect 5222 -37 5280 -31
rect 5340 -37 5398 -31
rect 5458 -37 5516 -31
rect 5576 -37 5634 -31
rect 5694 -37 5752 -31
rect 5812 -37 5870 -31
rect 5930 -37 5988 -31
rect 6048 -37 6106 -31
rect 6166 -37 6224 -31
rect 6284 -37 6342 -31
rect 6402 -37 6460 -31
rect 6520 -37 6578 -31
rect 6638 -37 6696 -31
rect 6756 -37 6814 -31
rect 6874 -37 6932 -31
rect 6992 -37 7050 -31
rect -7050 -71 -7038 -37
rect -6932 -71 -6920 -37
rect -6814 -71 -6802 -37
rect -6696 -71 -6684 -37
rect -6578 -71 -6566 -37
rect -6460 -71 -6448 -37
rect -6342 -71 -6330 -37
rect -6224 -71 -6212 -37
rect -6106 -71 -6094 -37
rect -5988 -71 -5976 -37
rect -5870 -71 -5858 -37
rect -5752 -71 -5740 -37
rect -5634 -71 -5622 -37
rect -5516 -71 -5504 -37
rect -5398 -71 -5386 -37
rect -5280 -71 -5268 -37
rect -5162 -71 -5150 -37
rect -5044 -71 -5032 -37
rect -4926 -71 -4914 -37
rect -4808 -71 -4796 -37
rect -4690 -71 -4678 -37
rect -4572 -71 -4560 -37
rect -4454 -71 -4442 -37
rect -4336 -71 -4324 -37
rect -4218 -71 -4206 -37
rect -4100 -71 -4088 -37
rect -3982 -71 -3970 -37
rect -3864 -71 -3852 -37
rect -3746 -71 -3734 -37
rect -3628 -71 -3616 -37
rect -3510 -71 -3498 -37
rect -3392 -71 -3380 -37
rect -3274 -71 -3262 -37
rect -3156 -71 -3144 -37
rect -3038 -71 -3026 -37
rect -2920 -71 -2908 -37
rect -2802 -71 -2790 -37
rect -2684 -71 -2672 -37
rect -2566 -71 -2554 -37
rect -2448 -71 -2436 -37
rect -2330 -71 -2318 -37
rect -2212 -71 -2200 -37
rect -2094 -71 -2082 -37
rect -1976 -71 -1964 -37
rect -1858 -71 -1846 -37
rect -1740 -71 -1728 -37
rect -1622 -71 -1610 -37
rect -1504 -71 -1492 -37
rect -1386 -71 -1374 -37
rect -1268 -71 -1256 -37
rect -1150 -71 -1138 -37
rect -1032 -71 -1020 -37
rect -914 -71 -902 -37
rect -796 -71 -784 -37
rect -678 -71 -666 -37
rect -560 -71 -548 -37
rect -442 -71 -430 -37
rect -324 -71 -312 -37
rect -206 -71 -194 -37
rect -88 -71 -76 -37
rect 30 -71 42 -37
rect 148 -71 160 -37
rect 266 -71 278 -37
rect 384 -71 396 -37
rect 502 -71 514 -37
rect 620 -71 632 -37
rect 738 -71 750 -37
rect 856 -71 868 -37
rect 974 -71 986 -37
rect 1092 -71 1104 -37
rect 1210 -71 1222 -37
rect 1328 -71 1340 -37
rect 1446 -71 1458 -37
rect 1564 -71 1576 -37
rect 1682 -71 1694 -37
rect 1800 -71 1812 -37
rect 1918 -71 1930 -37
rect 2036 -71 2048 -37
rect 2154 -71 2166 -37
rect 2272 -71 2284 -37
rect 2390 -71 2402 -37
rect 2508 -71 2520 -37
rect 2626 -71 2638 -37
rect 2744 -71 2756 -37
rect 2862 -71 2874 -37
rect 2980 -71 2992 -37
rect 3098 -71 3110 -37
rect 3216 -71 3228 -37
rect 3334 -71 3346 -37
rect 3452 -71 3464 -37
rect 3570 -71 3582 -37
rect 3688 -71 3700 -37
rect 3806 -71 3818 -37
rect 3924 -71 3936 -37
rect 4042 -71 4054 -37
rect 4160 -71 4172 -37
rect 4278 -71 4290 -37
rect 4396 -71 4408 -37
rect 4514 -71 4526 -37
rect 4632 -71 4644 -37
rect 4750 -71 4762 -37
rect 4868 -71 4880 -37
rect 4986 -71 4998 -37
rect 5104 -71 5116 -37
rect 5222 -71 5234 -37
rect 5340 -71 5352 -37
rect 5458 -71 5470 -37
rect 5576 -71 5588 -37
rect 5694 -71 5706 -37
rect 5812 -71 5824 -37
rect 5930 -71 5942 -37
rect 6048 -71 6060 -37
rect 6166 -71 6178 -37
rect 6284 -71 6296 -37
rect 6402 -71 6414 -37
rect 6520 -71 6532 -37
rect 6638 -71 6650 -37
rect 6756 -71 6768 -37
rect 6874 -71 6886 -37
rect 6992 -71 7004 -37
rect -7050 -77 -6992 -71
rect -6932 -77 -6874 -71
rect -6814 -77 -6756 -71
rect -6696 -77 -6638 -71
rect -6578 -77 -6520 -71
rect -6460 -77 -6402 -71
rect -6342 -77 -6284 -71
rect -6224 -77 -6166 -71
rect -6106 -77 -6048 -71
rect -5988 -77 -5930 -71
rect -5870 -77 -5812 -71
rect -5752 -77 -5694 -71
rect -5634 -77 -5576 -71
rect -5516 -77 -5458 -71
rect -5398 -77 -5340 -71
rect -5280 -77 -5222 -71
rect -5162 -77 -5104 -71
rect -5044 -77 -4986 -71
rect -4926 -77 -4868 -71
rect -4808 -77 -4750 -71
rect -4690 -77 -4632 -71
rect -4572 -77 -4514 -71
rect -4454 -77 -4396 -71
rect -4336 -77 -4278 -71
rect -4218 -77 -4160 -71
rect -4100 -77 -4042 -71
rect -3982 -77 -3924 -71
rect -3864 -77 -3806 -71
rect -3746 -77 -3688 -71
rect -3628 -77 -3570 -71
rect -3510 -77 -3452 -71
rect -3392 -77 -3334 -71
rect -3274 -77 -3216 -71
rect -3156 -77 -3098 -71
rect -3038 -77 -2980 -71
rect -2920 -77 -2862 -71
rect -2802 -77 -2744 -71
rect -2684 -77 -2626 -71
rect -2566 -77 -2508 -71
rect -2448 -77 -2390 -71
rect -2330 -77 -2272 -71
rect -2212 -77 -2154 -71
rect -2094 -77 -2036 -71
rect -1976 -77 -1918 -71
rect -1858 -77 -1800 -71
rect -1740 -77 -1682 -71
rect -1622 -77 -1564 -71
rect -1504 -77 -1446 -71
rect -1386 -77 -1328 -71
rect -1268 -77 -1210 -71
rect -1150 -77 -1092 -71
rect -1032 -77 -974 -71
rect -914 -77 -856 -71
rect -796 -77 -738 -71
rect -678 -77 -620 -71
rect -560 -77 -502 -71
rect -442 -77 -384 -71
rect -324 -77 -266 -71
rect -206 -77 -148 -71
rect -88 -77 -30 -71
rect 30 -77 88 -71
rect 148 -77 206 -71
rect 266 -77 324 -71
rect 384 -77 442 -71
rect 502 -77 560 -71
rect 620 -77 678 -71
rect 738 -77 796 -71
rect 856 -77 914 -71
rect 974 -77 1032 -71
rect 1092 -77 1150 -71
rect 1210 -77 1268 -71
rect 1328 -77 1386 -71
rect 1446 -77 1504 -71
rect 1564 -77 1622 -71
rect 1682 -77 1740 -71
rect 1800 -77 1858 -71
rect 1918 -77 1976 -71
rect 2036 -77 2094 -71
rect 2154 -77 2212 -71
rect 2272 -77 2330 -71
rect 2390 -77 2448 -71
rect 2508 -77 2566 -71
rect 2626 -77 2684 -71
rect 2744 -77 2802 -71
rect 2862 -77 2920 -71
rect 2980 -77 3038 -71
rect 3098 -77 3156 -71
rect 3216 -77 3274 -71
rect 3334 -77 3392 -71
rect 3452 -77 3510 -71
rect 3570 -77 3628 -71
rect 3688 -77 3746 -71
rect 3806 -77 3864 -71
rect 3924 -77 3982 -71
rect 4042 -77 4100 -71
rect 4160 -77 4218 -71
rect 4278 -77 4336 -71
rect 4396 -77 4454 -71
rect 4514 -77 4572 -71
rect 4632 -77 4690 -71
rect 4750 -77 4808 -71
rect 4868 -77 4926 -71
rect 4986 -77 5044 -71
rect 5104 -77 5162 -71
rect 5222 -77 5280 -71
rect 5340 -77 5398 -71
rect 5458 -77 5516 -71
rect 5576 -77 5634 -71
rect 5694 -77 5752 -71
rect 5812 -77 5870 -71
rect 5930 -77 5988 -71
rect 6048 -77 6106 -71
rect 6166 -77 6224 -71
rect 6284 -77 6342 -71
rect 6402 -77 6460 -71
rect 6520 -77 6578 -71
rect 6638 -77 6696 -71
rect 6756 -77 6814 -71
rect 6874 -77 6932 -71
rect 6992 -77 7050 -71
rect -7050 -765 -6992 -759
rect -6932 -765 -6874 -759
rect -6814 -765 -6756 -759
rect -6696 -765 -6638 -759
rect -6578 -765 -6520 -759
rect -6460 -765 -6402 -759
rect -6342 -765 -6284 -759
rect -6224 -765 -6166 -759
rect -6106 -765 -6048 -759
rect -5988 -765 -5930 -759
rect -5870 -765 -5812 -759
rect -5752 -765 -5694 -759
rect -5634 -765 -5576 -759
rect -5516 -765 -5458 -759
rect -5398 -765 -5340 -759
rect -5280 -765 -5222 -759
rect -5162 -765 -5104 -759
rect -5044 -765 -4986 -759
rect -4926 -765 -4868 -759
rect -4808 -765 -4750 -759
rect -4690 -765 -4632 -759
rect -4572 -765 -4514 -759
rect -4454 -765 -4396 -759
rect -4336 -765 -4278 -759
rect -4218 -765 -4160 -759
rect -4100 -765 -4042 -759
rect -3982 -765 -3924 -759
rect -3864 -765 -3806 -759
rect -3746 -765 -3688 -759
rect -3628 -765 -3570 -759
rect -3510 -765 -3452 -759
rect -3392 -765 -3334 -759
rect -3274 -765 -3216 -759
rect -3156 -765 -3098 -759
rect -3038 -765 -2980 -759
rect -2920 -765 -2862 -759
rect -2802 -765 -2744 -759
rect -2684 -765 -2626 -759
rect -2566 -765 -2508 -759
rect -2448 -765 -2390 -759
rect -2330 -765 -2272 -759
rect -2212 -765 -2154 -759
rect -2094 -765 -2036 -759
rect -1976 -765 -1918 -759
rect -1858 -765 -1800 -759
rect -1740 -765 -1682 -759
rect -1622 -765 -1564 -759
rect -1504 -765 -1446 -759
rect -1386 -765 -1328 -759
rect -1268 -765 -1210 -759
rect -1150 -765 -1092 -759
rect -1032 -765 -974 -759
rect -914 -765 -856 -759
rect -796 -765 -738 -759
rect -678 -765 -620 -759
rect -560 -765 -502 -759
rect -442 -765 -384 -759
rect -324 -765 -266 -759
rect -206 -765 -148 -759
rect -88 -765 -30 -759
rect 30 -765 88 -759
rect 148 -765 206 -759
rect 266 -765 324 -759
rect 384 -765 442 -759
rect 502 -765 560 -759
rect 620 -765 678 -759
rect 738 -765 796 -759
rect 856 -765 914 -759
rect 974 -765 1032 -759
rect 1092 -765 1150 -759
rect 1210 -765 1268 -759
rect 1328 -765 1386 -759
rect 1446 -765 1504 -759
rect 1564 -765 1622 -759
rect 1682 -765 1740 -759
rect 1800 -765 1858 -759
rect 1918 -765 1976 -759
rect 2036 -765 2094 -759
rect 2154 -765 2212 -759
rect 2272 -765 2330 -759
rect 2390 -765 2448 -759
rect 2508 -765 2566 -759
rect 2626 -765 2684 -759
rect 2744 -765 2802 -759
rect 2862 -765 2920 -759
rect 2980 -765 3038 -759
rect 3098 -765 3156 -759
rect 3216 -765 3274 -759
rect 3334 -765 3392 -759
rect 3452 -765 3510 -759
rect 3570 -765 3628 -759
rect 3688 -765 3746 -759
rect 3806 -765 3864 -759
rect 3924 -765 3982 -759
rect 4042 -765 4100 -759
rect 4160 -765 4218 -759
rect 4278 -765 4336 -759
rect 4396 -765 4454 -759
rect 4514 -765 4572 -759
rect 4632 -765 4690 -759
rect 4750 -765 4808 -759
rect 4868 -765 4926 -759
rect 4986 -765 5044 -759
rect 5104 -765 5162 -759
rect 5222 -765 5280 -759
rect 5340 -765 5398 -759
rect 5458 -765 5516 -759
rect 5576 -765 5634 -759
rect 5694 -765 5752 -759
rect 5812 -765 5870 -759
rect 5930 -765 5988 -759
rect 6048 -765 6106 -759
rect 6166 -765 6224 -759
rect 6284 -765 6342 -759
rect 6402 -765 6460 -759
rect 6520 -765 6578 -759
rect 6638 -765 6696 -759
rect 6756 -765 6814 -759
rect 6874 -765 6932 -759
rect 6992 -765 7050 -759
rect -7050 -799 -7038 -765
rect -6932 -799 -6920 -765
rect -6814 -799 -6802 -765
rect -6696 -799 -6684 -765
rect -6578 -799 -6566 -765
rect -6460 -799 -6448 -765
rect -6342 -799 -6330 -765
rect -6224 -799 -6212 -765
rect -6106 -799 -6094 -765
rect -5988 -799 -5976 -765
rect -5870 -799 -5858 -765
rect -5752 -799 -5740 -765
rect -5634 -799 -5622 -765
rect -5516 -799 -5504 -765
rect -5398 -799 -5386 -765
rect -5280 -799 -5268 -765
rect -5162 -799 -5150 -765
rect -5044 -799 -5032 -765
rect -4926 -799 -4914 -765
rect -4808 -799 -4796 -765
rect -4690 -799 -4678 -765
rect -4572 -799 -4560 -765
rect -4454 -799 -4442 -765
rect -4336 -799 -4324 -765
rect -4218 -799 -4206 -765
rect -4100 -799 -4088 -765
rect -3982 -799 -3970 -765
rect -3864 -799 -3852 -765
rect -3746 -799 -3734 -765
rect -3628 -799 -3616 -765
rect -3510 -799 -3498 -765
rect -3392 -799 -3380 -765
rect -3274 -799 -3262 -765
rect -3156 -799 -3144 -765
rect -3038 -799 -3026 -765
rect -2920 -799 -2908 -765
rect -2802 -799 -2790 -765
rect -2684 -799 -2672 -765
rect -2566 -799 -2554 -765
rect -2448 -799 -2436 -765
rect -2330 -799 -2318 -765
rect -2212 -799 -2200 -765
rect -2094 -799 -2082 -765
rect -1976 -799 -1964 -765
rect -1858 -799 -1846 -765
rect -1740 -799 -1728 -765
rect -1622 -799 -1610 -765
rect -1504 -799 -1492 -765
rect -1386 -799 -1374 -765
rect -1268 -799 -1256 -765
rect -1150 -799 -1138 -765
rect -1032 -799 -1020 -765
rect -914 -799 -902 -765
rect -796 -799 -784 -765
rect -678 -799 -666 -765
rect -560 -799 -548 -765
rect -442 -799 -430 -765
rect -324 -799 -312 -765
rect -206 -799 -194 -765
rect -88 -799 -76 -765
rect 30 -799 42 -765
rect 148 -799 160 -765
rect 266 -799 278 -765
rect 384 -799 396 -765
rect 502 -799 514 -765
rect 620 -799 632 -765
rect 738 -799 750 -765
rect 856 -799 868 -765
rect 974 -799 986 -765
rect 1092 -799 1104 -765
rect 1210 -799 1222 -765
rect 1328 -799 1340 -765
rect 1446 -799 1458 -765
rect 1564 -799 1576 -765
rect 1682 -799 1694 -765
rect 1800 -799 1812 -765
rect 1918 -799 1930 -765
rect 2036 -799 2048 -765
rect 2154 -799 2166 -765
rect 2272 -799 2284 -765
rect 2390 -799 2402 -765
rect 2508 -799 2520 -765
rect 2626 -799 2638 -765
rect 2744 -799 2756 -765
rect 2862 -799 2874 -765
rect 2980 -799 2992 -765
rect 3098 -799 3110 -765
rect 3216 -799 3228 -765
rect 3334 -799 3346 -765
rect 3452 -799 3464 -765
rect 3570 -799 3582 -765
rect 3688 -799 3700 -765
rect 3806 -799 3818 -765
rect 3924 -799 3936 -765
rect 4042 -799 4054 -765
rect 4160 -799 4172 -765
rect 4278 -799 4290 -765
rect 4396 -799 4408 -765
rect 4514 -799 4526 -765
rect 4632 -799 4644 -765
rect 4750 -799 4762 -765
rect 4868 -799 4880 -765
rect 4986 -799 4998 -765
rect 5104 -799 5116 -765
rect 5222 -799 5234 -765
rect 5340 -799 5352 -765
rect 5458 -799 5470 -765
rect 5576 -799 5588 -765
rect 5694 -799 5706 -765
rect 5812 -799 5824 -765
rect 5930 -799 5942 -765
rect 6048 -799 6060 -765
rect 6166 -799 6178 -765
rect 6284 -799 6296 -765
rect 6402 -799 6414 -765
rect 6520 -799 6532 -765
rect 6638 -799 6650 -765
rect 6756 -799 6768 -765
rect 6874 -799 6886 -765
rect 6992 -799 7004 -765
rect -7050 -805 -6992 -799
rect -6932 -805 -6874 -799
rect -6814 -805 -6756 -799
rect -6696 -805 -6638 -799
rect -6578 -805 -6520 -799
rect -6460 -805 -6402 -799
rect -6342 -805 -6284 -799
rect -6224 -805 -6166 -799
rect -6106 -805 -6048 -799
rect -5988 -805 -5930 -799
rect -5870 -805 -5812 -799
rect -5752 -805 -5694 -799
rect -5634 -805 -5576 -799
rect -5516 -805 -5458 -799
rect -5398 -805 -5340 -799
rect -5280 -805 -5222 -799
rect -5162 -805 -5104 -799
rect -5044 -805 -4986 -799
rect -4926 -805 -4868 -799
rect -4808 -805 -4750 -799
rect -4690 -805 -4632 -799
rect -4572 -805 -4514 -799
rect -4454 -805 -4396 -799
rect -4336 -805 -4278 -799
rect -4218 -805 -4160 -799
rect -4100 -805 -4042 -799
rect -3982 -805 -3924 -799
rect -3864 -805 -3806 -799
rect -3746 -805 -3688 -799
rect -3628 -805 -3570 -799
rect -3510 -805 -3452 -799
rect -3392 -805 -3334 -799
rect -3274 -805 -3216 -799
rect -3156 -805 -3098 -799
rect -3038 -805 -2980 -799
rect -2920 -805 -2862 -799
rect -2802 -805 -2744 -799
rect -2684 -805 -2626 -799
rect -2566 -805 -2508 -799
rect -2448 -805 -2390 -799
rect -2330 -805 -2272 -799
rect -2212 -805 -2154 -799
rect -2094 -805 -2036 -799
rect -1976 -805 -1918 -799
rect -1858 -805 -1800 -799
rect -1740 -805 -1682 -799
rect -1622 -805 -1564 -799
rect -1504 -805 -1446 -799
rect -1386 -805 -1328 -799
rect -1268 -805 -1210 -799
rect -1150 -805 -1092 -799
rect -1032 -805 -974 -799
rect -914 -805 -856 -799
rect -796 -805 -738 -799
rect -678 -805 -620 -799
rect -560 -805 -502 -799
rect -442 -805 -384 -799
rect -324 -805 -266 -799
rect -206 -805 -148 -799
rect -88 -805 -30 -799
rect 30 -805 88 -799
rect 148 -805 206 -799
rect 266 -805 324 -799
rect 384 -805 442 -799
rect 502 -805 560 -799
rect 620 -805 678 -799
rect 738 -805 796 -799
rect 856 -805 914 -799
rect 974 -805 1032 -799
rect 1092 -805 1150 -799
rect 1210 -805 1268 -799
rect 1328 -805 1386 -799
rect 1446 -805 1504 -799
rect 1564 -805 1622 -799
rect 1682 -805 1740 -799
rect 1800 -805 1858 -799
rect 1918 -805 1976 -799
rect 2036 -805 2094 -799
rect 2154 -805 2212 -799
rect 2272 -805 2330 -799
rect 2390 -805 2448 -799
rect 2508 -805 2566 -799
rect 2626 -805 2684 -799
rect 2744 -805 2802 -799
rect 2862 -805 2920 -799
rect 2980 -805 3038 -799
rect 3098 -805 3156 -799
rect 3216 -805 3274 -799
rect 3334 -805 3392 -799
rect 3452 -805 3510 -799
rect 3570 -805 3628 -799
rect 3688 -805 3746 -799
rect 3806 -805 3864 -799
rect 3924 -805 3982 -799
rect 4042 -805 4100 -799
rect 4160 -805 4218 -799
rect 4278 -805 4336 -799
rect 4396 -805 4454 -799
rect 4514 -805 4572 -799
rect 4632 -805 4690 -799
rect 4750 -805 4808 -799
rect 4868 -805 4926 -799
rect 4986 -805 5044 -799
rect 5104 -805 5162 -799
rect 5222 -805 5280 -799
rect 5340 -805 5398 -799
rect 5458 -805 5516 -799
rect 5576 -805 5634 -799
rect 5694 -805 5752 -799
rect 5812 -805 5870 -799
rect 5930 -805 5988 -799
rect 6048 -805 6106 -799
rect 6166 -805 6224 -799
rect 6284 -805 6342 -799
rect 6402 -805 6460 -799
rect 6520 -805 6578 -799
rect 6638 -805 6696 -799
rect 6756 -805 6814 -799
rect 6874 -805 6932 -799
rect 6992 -805 7050 -799
<< nwell >>
rect -7247 -937 7247 937
<< pmos >>
rect -7051 118 -6991 718
rect -6933 118 -6873 718
rect -6815 118 -6755 718
rect -6697 118 -6637 718
rect -6579 118 -6519 718
rect -6461 118 -6401 718
rect -6343 118 -6283 718
rect -6225 118 -6165 718
rect -6107 118 -6047 718
rect -5989 118 -5929 718
rect -5871 118 -5811 718
rect -5753 118 -5693 718
rect -5635 118 -5575 718
rect -5517 118 -5457 718
rect -5399 118 -5339 718
rect -5281 118 -5221 718
rect -5163 118 -5103 718
rect -5045 118 -4985 718
rect -4927 118 -4867 718
rect -4809 118 -4749 718
rect -4691 118 -4631 718
rect -4573 118 -4513 718
rect -4455 118 -4395 718
rect -4337 118 -4277 718
rect -4219 118 -4159 718
rect -4101 118 -4041 718
rect -3983 118 -3923 718
rect -3865 118 -3805 718
rect -3747 118 -3687 718
rect -3629 118 -3569 718
rect -3511 118 -3451 718
rect -3393 118 -3333 718
rect -3275 118 -3215 718
rect -3157 118 -3097 718
rect -3039 118 -2979 718
rect -2921 118 -2861 718
rect -2803 118 -2743 718
rect -2685 118 -2625 718
rect -2567 118 -2507 718
rect -2449 118 -2389 718
rect -2331 118 -2271 718
rect -2213 118 -2153 718
rect -2095 118 -2035 718
rect -1977 118 -1917 718
rect -1859 118 -1799 718
rect -1741 118 -1681 718
rect -1623 118 -1563 718
rect -1505 118 -1445 718
rect -1387 118 -1327 718
rect -1269 118 -1209 718
rect -1151 118 -1091 718
rect -1033 118 -973 718
rect -915 118 -855 718
rect -797 118 -737 718
rect -679 118 -619 718
rect -561 118 -501 718
rect -443 118 -383 718
rect -325 118 -265 718
rect -207 118 -147 718
rect -89 118 -29 718
rect 29 118 89 718
rect 147 118 207 718
rect 265 118 325 718
rect 383 118 443 718
rect 501 118 561 718
rect 619 118 679 718
rect 737 118 797 718
rect 855 118 915 718
rect 973 118 1033 718
rect 1091 118 1151 718
rect 1209 118 1269 718
rect 1327 118 1387 718
rect 1445 118 1505 718
rect 1563 118 1623 718
rect 1681 118 1741 718
rect 1799 118 1859 718
rect 1917 118 1977 718
rect 2035 118 2095 718
rect 2153 118 2213 718
rect 2271 118 2331 718
rect 2389 118 2449 718
rect 2507 118 2567 718
rect 2625 118 2685 718
rect 2743 118 2803 718
rect 2861 118 2921 718
rect 2979 118 3039 718
rect 3097 118 3157 718
rect 3215 118 3275 718
rect 3333 118 3393 718
rect 3451 118 3511 718
rect 3569 118 3629 718
rect 3687 118 3747 718
rect 3805 118 3865 718
rect 3923 118 3983 718
rect 4041 118 4101 718
rect 4159 118 4219 718
rect 4277 118 4337 718
rect 4395 118 4455 718
rect 4513 118 4573 718
rect 4631 118 4691 718
rect 4749 118 4809 718
rect 4867 118 4927 718
rect 4985 118 5045 718
rect 5103 118 5163 718
rect 5221 118 5281 718
rect 5339 118 5399 718
rect 5457 118 5517 718
rect 5575 118 5635 718
rect 5693 118 5753 718
rect 5811 118 5871 718
rect 5929 118 5989 718
rect 6047 118 6107 718
rect 6165 118 6225 718
rect 6283 118 6343 718
rect 6401 118 6461 718
rect 6519 118 6579 718
rect 6637 118 6697 718
rect 6755 118 6815 718
rect 6873 118 6933 718
rect 6991 118 7051 718
rect -7051 -718 -6991 -118
rect -6933 -718 -6873 -118
rect -6815 -718 -6755 -118
rect -6697 -718 -6637 -118
rect -6579 -718 -6519 -118
rect -6461 -718 -6401 -118
rect -6343 -718 -6283 -118
rect -6225 -718 -6165 -118
rect -6107 -718 -6047 -118
rect -5989 -718 -5929 -118
rect -5871 -718 -5811 -118
rect -5753 -718 -5693 -118
rect -5635 -718 -5575 -118
rect -5517 -718 -5457 -118
rect -5399 -718 -5339 -118
rect -5281 -718 -5221 -118
rect -5163 -718 -5103 -118
rect -5045 -718 -4985 -118
rect -4927 -718 -4867 -118
rect -4809 -718 -4749 -118
rect -4691 -718 -4631 -118
rect -4573 -718 -4513 -118
rect -4455 -718 -4395 -118
rect -4337 -718 -4277 -118
rect -4219 -718 -4159 -118
rect -4101 -718 -4041 -118
rect -3983 -718 -3923 -118
rect -3865 -718 -3805 -118
rect -3747 -718 -3687 -118
rect -3629 -718 -3569 -118
rect -3511 -718 -3451 -118
rect -3393 -718 -3333 -118
rect -3275 -718 -3215 -118
rect -3157 -718 -3097 -118
rect -3039 -718 -2979 -118
rect -2921 -718 -2861 -118
rect -2803 -718 -2743 -118
rect -2685 -718 -2625 -118
rect -2567 -718 -2507 -118
rect -2449 -718 -2389 -118
rect -2331 -718 -2271 -118
rect -2213 -718 -2153 -118
rect -2095 -718 -2035 -118
rect -1977 -718 -1917 -118
rect -1859 -718 -1799 -118
rect -1741 -718 -1681 -118
rect -1623 -718 -1563 -118
rect -1505 -718 -1445 -118
rect -1387 -718 -1327 -118
rect -1269 -718 -1209 -118
rect -1151 -718 -1091 -118
rect -1033 -718 -973 -118
rect -915 -718 -855 -118
rect -797 -718 -737 -118
rect -679 -718 -619 -118
rect -561 -718 -501 -118
rect -443 -718 -383 -118
rect -325 -718 -265 -118
rect -207 -718 -147 -118
rect -89 -718 -29 -118
rect 29 -718 89 -118
rect 147 -718 207 -118
rect 265 -718 325 -118
rect 383 -718 443 -118
rect 501 -718 561 -118
rect 619 -718 679 -118
rect 737 -718 797 -118
rect 855 -718 915 -118
rect 973 -718 1033 -118
rect 1091 -718 1151 -118
rect 1209 -718 1269 -118
rect 1327 -718 1387 -118
rect 1445 -718 1505 -118
rect 1563 -718 1623 -118
rect 1681 -718 1741 -118
rect 1799 -718 1859 -118
rect 1917 -718 1977 -118
rect 2035 -718 2095 -118
rect 2153 -718 2213 -118
rect 2271 -718 2331 -118
rect 2389 -718 2449 -118
rect 2507 -718 2567 -118
rect 2625 -718 2685 -118
rect 2743 -718 2803 -118
rect 2861 -718 2921 -118
rect 2979 -718 3039 -118
rect 3097 -718 3157 -118
rect 3215 -718 3275 -118
rect 3333 -718 3393 -118
rect 3451 -718 3511 -118
rect 3569 -718 3629 -118
rect 3687 -718 3747 -118
rect 3805 -718 3865 -118
rect 3923 -718 3983 -118
rect 4041 -718 4101 -118
rect 4159 -718 4219 -118
rect 4277 -718 4337 -118
rect 4395 -718 4455 -118
rect 4513 -718 4573 -118
rect 4631 -718 4691 -118
rect 4749 -718 4809 -118
rect 4867 -718 4927 -118
rect 4985 -718 5045 -118
rect 5103 -718 5163 -118
rect 5221 -718 5281 -118
rect 5339 -718 5399 -118
rect 5457 -718 5517 -118
rect 5575 -718 5635 -118
rect 5693 -718 5753 -118
rect 5811 -718 5871 -118
rect 5929 -718 5989 -118
rect 6047 -718 6107 -118
rect 6165 -718 6225 -118
rect 6283 -718 6343 -118
rect 6401 -718 6461 -118
rect 6519 -718 6579 -118
rect 6637 -718 6697 -118
rect 6755 -718 6815 -118
rect 6873 -718 6933 -118
rect 6991 -718 7051 -118
<< pdiff >>
rect -7109 706 -7051 718
rect -7109 130 -7097 706
rect -7063 130 -7051 706
rect -7109 118 -7051 130
rect -6991 706 -6933 718
rect -6991 130 -6979 706
rect -6945 130 -6933 706
rect -6991 118 -6933 130
rect -6873 706 -6815 718
rect -6873 130 -6861 706
rect -6827 130 -6815 706
rect -6873 118 -6815 130
rect -6755 706 -6697 718
rect -6755 130 -6743 706
rect -6709 130 -6697 706
rect -6755 118 -6697 130
rect -6637 706 -6579 718
rect -6637 130 -6625 706
rect -6591 130 -6579 706
rect -6637 118 -6579 130
rect -6519 706 -6461 718
rect -6519 130 -6507 706
rect -6473 130 -6461 706
rect -6519 118 -6461 130
rect -6401 706 -6343 718
rect -6401 130 -6389 706
rect -6355 130 -6343 706
rect -6401 118 -6343 130
rect -6283 706 -6225 718
rect -6283 130 -6271 706
rect -6237 130 -6225 706
rect -6283 118 -6225 130
rect -6165 706 -6107 718
rect -6165 130 -6153 706
rect -6119 130 -6107 706
rect -6165 118 -6107 130
rect -6047 706 -5989 718
rect -6047 130 -6035 706
rect -6001 130 -5989 706
rect -6047 118 -5989 130
rect -5929 706 -5871 718
rect -5929 130 -5917 706
rect -5883 130 -5871 706
rect -5929 118 -5871 130
rect -5811 706 -5753 718
rect -5811 130 -5799 706
rect -5765 130 -5753 706
rect -5811 118 -5753 130
rect -5693 706 -5635 718
rect -5693 130 -5681 706
rect -5647 130 -5635 706
rect -5693 118 -5635 130
rect -5575 706 -5517 718
rect -5575 130 -5563 706
rect -5529 130 -5517 706
rect -5575 118 -5517 130
rect -5457 706 -5399 718
rect -5457 130 -5445 706
rect -5411 130 -5399 706
rect -5457 118 -5399 130
rect -5339 706 -5281 718
rect -5339 130 -5327 706
rect -5293 130 -5281 706
rect -5339 118 -5281 130
rect -5221 706 -5163 718
rect -5221 130 -5209 706
rect -5175 130 -5163 706
rect -5221 118 -5163 130
rect -5103 706 -5045 718
rect -5103 130 -5091 706
rect -5057 130 -5045 706
rect -5103 118 -5045 130
rect -4985 706 -4927 718
rect -4985 130 -4973 706
rect -4939 130 -4927 706
rect -4985 118 -4927 130
rect -4867 706 -4809 718
rect -4867 130 -4855 706
rect -4821 130 -4809 706
rect -4867 118 -4809 130
rect -4749 706 -4691 718
rect -4749 130 -4737 706
rect -4703 130 -4691 706
rect -4749 118 -4691 130
rect -4631 706 -4573 718
rect -4631 130 -4619 706
rect -4585 130 -4573 706
rect -4631 118 -4573 130
rect -4513 706 -4455 718
rect -4513 130 -4501 706
rect -4467 130 -4455 706
rect -4513 118 -4455 130
rect -4395 706 -4337 718
rect -4395 130 -4383 706
rect -4349 130 -4337 706
rect -4395 118 -4337 130
rect -4277 706 -4219 718
rect -4277 130 -4265 706
rect -4231 130 -4219 706
rect -4277 118 -4219 130
rect -4159 706 -4101 718
rect -4159 130 -4147 706
rect -4113 130 -4101 706
rect -4159 118 -4101 130
rect -4041 706 -3983 718
rect -4041 130 -4029 706
rect -3995 130 -3983 706
rect -4041 118 -3983 130
rect -3923 706 -3865 718
rect -3923 130 -3911 706
rect -3877 130 -3865 706
rect -3923 118 -3865 130
rect -3805 706 -3747 718
rect -3805 130 -3793 706
rect -3759 130 -3747 706
rect -3805 118 -3747 130
rect -3687 706 -3629 718
rect -3687 130 -3675 706
rect -3641 130 -3629 706
rect -3687 118 -3629 130
rect -3569 706 -3511 718
rect -3569 130 -3557 706
rect -3523 130 -3511 706
rect -3569 118 -3511 130
rect -3451 706 -3393 718
rect -3451 130 -3439 706
rect -3405 130 -3393 706
rect -3451 118 -3393 130
rect -3333 706 -3275 718
rect -3333 130 -3321 706
rect -3287 130 -3275 706
rect -3333 118 -3275 130
rect -3215 706 -3157 718
rect -3215 130 -3203 706
rect -3169 130 -3157 706
rect -3215 118 -3157 130
rect -3097 706 -3039 718
rect -3097 130 -3085 706
rect -3051 130 -3039 706
rect -3097 118 -3039 130
rect -2979 706 -2921 718
rect -2979 130 -2967 706
rect -2933 130 -2921 706
rect -2979 118 -2921 130
rect -2861 706 -2803 718
rect -2861 130 -2849 706
rect -2815 130 -2803 706
rect -2861 118 -2803 130
rect -2743 706 -2685 718
rect -2743 130 -2731 706
rect -2697 130 -2685 706
rect -2743 118 -2685 130
rect -2625 706 -2567 718
rect -2625 130 -2613 706
rect -2579 130 -2567 706
rect -2625 118 -2567 130
rect -2507 706 -2449 718
rect -2507 130 -2495 706
rect -2461 130 -2449 706
rect -2507 118 -2449 130
rect -2389 706 -2331 718
rect -2389 130 -2377 706
rect -2343 130 -2331 706
rect -2389 118 -2331 130
rect -2271 706 -2213 718
rect -2271 130 -2259 706
rect -2225 130 -2213 706
rect -2271 118 -2213 130
rect -2153 706 -2095 718
rect -2153 130 -2141 706
rect -2107 130 -2095 706
rect -2153 118 -2095 130
rect -2035 706 -1977 718
rect -2035 130 -2023 706
rect -1989 130 -1977 706
rect -2035 118 -1977 130
rect -1917 706 -1859 718
rect -1917 130 -1905 706
rect -1871 130 -1859 706
rect -1917 118 -1859 130
rect -1799 706 -1741 718
rect -1799 130 -1787 706
rect -1753 130 -1741 706
rect -1799 118 -1741 130
rect -1681 706 -1623 718
rect -1681 130 -1669 706
rect -1635 130 -1623 706
rect -1681 118 -1623 130
rect -1563 706 -1505 718
rect -1563 130 -1551 706
rect -1517 130 -1505 706
rect -1563 118 -1505 130
rect -1445 706 -1387 718
rect -1445 130 -1433 706
rect -1399 130 -1387 706
rect -1445 118 -1387 130
rect -1327 706 -1269 718
rect -1327 130 -1315 706
rect -1281 130 -1269 706
rect -1327 118 -1269 130
rect -1209 706 -1151 718
rect -1209 130 -1197 706
rect -1163 130 -1151 706
rect -1209 118 -1151 130
rect -1091 706 -1033 718
rect -1091 130 -1079 706
rect -1045 130 -1033 706
rect -1091 118 -1033 130
rect -973 706 -915 718
rect -973 130 -961 706
rect -927 130 -915 706
rect -973 118 -915 130
rect -855 706 -797 718
rect -855 130 -843 706
rect -809 130 -797 706
rect -855 118 -797 130
rect -737 706 -679 718
rect -737 130 -725 706
rect -691 130 -679 706
rect -737 118 -679 130
rect -619 706 -561 718
rect -619 130 -607 706
rect -573 130 -561 706
rect -619 118 -561 130
rect -501 706 -443 718
rect -501 130 -489 706
rect -455 130 -443 706
rect -501 118 -443 130
rect -383 706 -325 718
rect -383 130 -371 706
rect -337 130 -325 706
rect -383 118 -325 130
rect -265 706 -207 718
rect -265 130 -253 706
rect -219 130 -207 706
rect -265 118 -207 130
rect -147 706 -89 718
rect -147 130 -135 706
rect -101 130 -89 706
rect -147 118 -89 130
rect -29 706 29 718
rect -29 130 -17 706
rect 17 130 29 706
rect -29 118 29 130
rect 89 706 147 718
rect 89 130 101 706
rect 135 130 147 706
rect 89 118 147 130
rect 207 706 265 718
rect 207 130 219 706
rect 253 130 265 706
rect 207 118 265 130
rect 325 706 383 718
rect 325 130 337 706
rect 371 130 383 706
rect 325 118 383 130
rect 443 706 501 718
rect 443 130 455 706
rect 489 130 501 706
rect 443 118 501 130
rect 561 706 619 718
rect 561 130 573 706
rect 607 130 619 706
rect 561 118 619 130
rect 679 706 737 718
rect 679 130 691 706
rect 725 130 737 706
rect 679 118 737 130
rect 797 706 855 718
rect 797 130 809 706
rect 843 130 855 706
rect 797 118 855 130
rect 915 706 973 718
rect 915 130 927 706
rect 961 130 973 706
rect 915 118 973 130
rect 1033 706 1091 718
rect 1033 130 1045 706
rect 1079 130 1091 706
rect 1033 118 1091 130
rect 1151 706 1209 718
rect 1151 130 1163 706
rect 1197 130 1209 706
rect 1151 118 1209 130
rect 1269 706 1327 718
rect 1269 130 1281 706
rect 1315 130 1327 706
rect 1269 118 1327 130
rect 1387 706 1445 718
rect 1387 130 1399 706
rect 1433 130 1445 706
rect 1387 118 1445 130
rect 1505 706 1563 718
rect 1505 130 1517 706
rect 1551 130 1563 706
rect 1505 118 1563 130
rect 1623 706 1681 718
rect 1623 130 1635 706
rect 1669 130 1681 706
rect 1623 118 1681 130
rect 1741 706 1799 718
rect 1741 130 1753 706
rect 1787 130 1799 706
rect 1741 118 1799 130
rect 1859 706 1917 718
rect 1859 130 1871 706
rect 1905 130 1917 706
rect 1859 118 1917 130
rect 1977 706 2035 718
rect 1977 130 1989 706
rect 2023 130 2035 706
rect 1977 118 2035 130
rect 2095 706 2153 718
rect 2095 130 2107 706
rect 2141 130 2153 706
rect 2095 118 2153 130
rect 2213 706 2271 718
rect 2213 130 2225 706
rect 2259 130 2271 706
rect 2213 118 2271 130
rect 2331 706 2389 718
rect 2331 130 2343 706
rect 2377 130 2389 706
rect 2331 118 2389 130
rect 2449 706 2507 718
rect 2449 130 2461 706
rect 2495 130 2507 706
rect 2449 118 2507 130
rect 2567 706 2625 718
rect 2567 130 2579 706
rect 2613 130 2625 706
rect 2567 118 2625 130
rect 2685 706 2743 718
rect 2685 130 2697 706
rect 2731 130 2743 706
rect 2685 118 2743 130
rect 2803 706 2861 718
rect 2803 130 2815 706
rect 2849 130 2861 706
rect 2803 118 2861 130
rect 2921 706 2979 718
rect 2921 130 2933 706
rect 2967 130 2979 706
rect 2921 118 2979 130
rect 3039 706 3097 718
rect 3039 130 3051 706
rect 3085 130 3097 706
rect 3039 118 3097 130
rect 3157 706 3215 718
rect 3157 130 3169 706
rect 3203 130 3215 706
rect 3157 118 3215 130
rect 3275 706 3333 718
rect 3275 130 3287 706
rect 3321 130 3333 706
rect 3275 118 3333 130
rect 3393 706 3451 718
rect 3393 130 3405 706
rect 3439 130 3451 706
rect 3393 118 3451 130
rect 3511 706 3569 718
rect 3511 130 3523 706
rect 3557 130 3569 706
rect 3511 118 3569 130
rect 3629 706 3687 718
rect 3629 130 3641 706
rect 3675 130 3687 706
rect 3629 118 3687 130
rect 3747 706 3805 718
rect 3747 130 3759 706
rect 3793 130 3805 706
rect 3747 118 3805 130
rect 3865 706 3923 718
rect 3865 130 3877 706
rect 3911 130 3923 706
rect 3865 118 3923 130
rect 3983 706 4041 718
rect 3983 130 3995 706
rect 4029 130 4041 706
rect 3983 118 4041 130
rect 4101 706 4159 718
rect 4101 130 4113 706
rect 4147 130 4159 706
rect 4101 118 4159 130
rect 4219 706 4277 718
rect 4219 130 4231 706
rect 4265 130 4277 706
rect 4219 118 4277 130
rect 4337 706 4395 718
rect 4337 130 4349 706
rect 4383 130 4395 706
rect 4337 118 4395 130
rect 4455 706 4513 718
rect 4455 130 4467 706
rect 4501 130 4513 706
rect 4455 118 4513 130
rect 4573 706 4631 718
rect 4573 130 4585 706
rect 4619 130 4631 706
rect 4573 118 4631 130
rect 4691 706 4749 718
rect 4691 130 4703 706
rect 4737 130 4749 706
rect 4691 118 4749 130
rect 4809 706 4867 718
rect 4809 130 4821 706
rect 4855 130 4867 706
rect 4809 118 4867 130
rect 4927 706 4985 718
rect 4927 130 4939 706
rect 4973 130 4985 706
rect 4927 118 4985 130
rect 5045 706 5103 718
rect 5045 130 5057 706
rect 5091 130 5103 706
rect 5045 118 5103 130
rect 5163 706 5221 718
rect 5163 130 5175 706
rect 5209 130 5221 706
rect 5163 118 5221 130
rect 5281 706 5339 718
rect 5281 130 5293 706
rect 5327 130 5339 706
rect 5281 118 5339 130
rect 5399 706 5457 718
rect 5399 130 5411 706
rect 5445 130 5457 706
rect 5399 118 5457 130
rect 5517 706 5575 718
rect 5517 130 5529 706
rect 5563 130 5575 706
rect 5517 118 5575 130
rect 5635 706 5693 718
rect 5635 130 5647 706
rect 5681 130 5693 706
rect 5635 118 5693 130
rect 5753 706 5811 718
rect 5753 130 5765 706
rect 5799 130 5811 706
rect 5753 118 5811 130
rect 5871 706 5929 718
rect 5871 130 5883 706
rect 5917 130 5929 706
rect 5871 118 5929 130
rect 5989 706 6047 718
rect 5989 130 6001 706
rect 6035 130 6047 706
rect 5989 118 6047 130
rect 6107 706 6165 718
rect 6107 130 6119 706
rect 6153 130 6165 706
rect 6107 118 6165 130
rect 6225 706 6283 718
rect 6225 130 6237 706
rect 6271 130 6283 706
rect 6225 118 6283 130
rect 6343 706 6401 718
rect 6343 130 6355 706
rect 6389 130 6401 706
rect 6343 118 6401 130
rect 6461 706 6519 718
rect 6461 130 6473 706
rect 6507 130 6519 706
rect 6461 118 6519 130
rect 6579 706 6637 718
rect 6579 130 6591 706
rect 6625 130 6637 706
rect 6579 118 6637 130
rect 6697 706 6755 718
rect 6697 130 6709 706
rect 6743 130 6755 706
rect 6697 118 6755 130
rect 6815 706 6873 718
rect 6815 130 6827 706
rect 6861 130 6873 706
rect 6815 118 6873 130
rect 6933 706 6991 718
rect 6933 130 6945 706
rect 6979 130 6991 706
rect 6933 118 6991 130
rect 7051 706 7109 718
rect 7051 130 7063 706
rect 7097 130 7109 706
rect 7051 118 7109 130
rect -7109 -130 -7051 -118
rect -7109 -706 -7097 -130
rect -7063 -706 -7051 -130
rect -7109 -718 -7051 -706
rect -6991 -130 -6933 -118
rect -6991 -706 -6979 -130
rect -6945 -706 -6933 -130
rect -6991 -718 -6933 -706
rect -6873 -130 -6815 -118
rect -6873 -706 -6861 -130
rect -6827 -706 -6815 -130
rect -6873 -718 -6815 -706
rect -6755 -130 -6697 -118
rect -6755 -706 -6743 -130
rect -6709 -706 -6697 -130
rect -6755 -718 -6697 -706
rect -6637 -130 -6579 -118
rect -6637 -706 -6625 -130
rect -6591 -706 -6579 -130
rect -6637 -718 -6579 -706
rect -6519 -130 -6461 -118
rect -6519 -706 -6507 -130
rect -6473 -706 -6461 -130
rect -6519 -718 -6461 -706
rect -6401 -130 -6343 -118
rect -6401 -706 -6389 -130
rect -6355 -706 -6343 -130
rect -6401 -718 -6343 -706
rect -6283 -130 -6225 -118
rect -6283 -706 -6271 -130
rect -6237 -706 -6225 -130
rect -6283 -718 -6225 -706
rect -6165 -130 -6107 -118
rect -6165 -706 -6153 -130
rect -6119 -706 -6107 -130
rect -6165 -718 -6107 -706
rect -6047 -130 -5989 -118
rect -6047 -706 -6035 -130
rect -6001 -706 -5989 -130
rect -6047 -718 -5989 -706
rect -5929 -130 -5871 -118
rect -5929 -706 -5917 -130
rect -5883 -706 -5871 -130
rect -5929 -718 -5871 -706
rect -5811 -130 -5753 -118
rect -5811 -706 -5799 -130
rect -5765 -706 -5753 -130
rect -5811 -718 -5753 -706
rect -5693 -130 -5635 -118
rect -5693 -706 -5681 -130
rect -5647 -706 -5635 -130
rect -5693 -718 -5635 -706
rect -5575 -130 -5517 -118
rect -5575 -706 -5563 -130
rect -5529 -706 -5517 -130
rect -5575 -718 -5517 -706
rect -5457 -130 -5399 -118
rect -5457 -706 -5445 -130
rect -5411 -706 -5399 -130
rect -5457 -718 -5399 -706
rect -5339 -130 -5281 -118
rect -5339 -706 -5327 -130
rect -5293 -706 -5281 -130
rect -5339 -718 -5281 -706
rect -5221 -130 -5163 -118
rect -5221 -706 -5209 -130
rect -5175 -706 -5163 -130
rect -5221 -718 -5163 -706
rect -5103 -130 -5045 -118
rect -5103 -706 -5091 -130
rect -5057 -706 -5045 -130
rect -5103 -718 -5045 -706
rect -4985 -130 -4927 -118
rect -4985 -706 -4973 -130
rect -4939 -706 -4927 -130
rect -4985 -718 -4927 -706
rect -4867 -130 -4809 -118
rect -4867 -706 -4855 -130
rect -4821 -706 -4809 -130
rect -4867 -718 -4809 -706
rect -4749 -130 -4691 -118
rect -4749 -706 -4737 -130
rect -4703 -706 -4691 -130
rect -4749 -718 -4691 -706
rect -4631 -130 -4573 -118
rect -4631 -706 -4619 -130
rect -4585 -706 -4573 -130
rect -4631 -718 -4573 -706
rect -4513 -130 -4455 -118
rect -4513 -706 -4501 -130
rect -4467 -706 -4455 -130
rect -4513 -718 -4455 -706
rect -4395 -130 -4337 -118
rect -4395 -706 -4383 -130
rect -4349 -706 -4337 -130
rect -4395 -718 -4337 -706
rect -4277 -130 -4219 -118
rect -4277 -706 -4265 -130
rect -4231 -706 -4219 -130
rect -4277 -718 -4219 -706
rect -4159 -130 -4101 -118
rect -4159 -706 -4147 -130
rect -4113 -706 -4101 -130
rect -4159 -718 -4101 -706
rect -4041 -130 -3983 -118
rect -4041 -706 -4029 -130
rect -3995 -706 -3983 -130
rect -4041 -718 -3983 -706
rect -3923 -130 -3865 -118
rect -3923 -706 -3911 -130
rect -3877 -706 -3865 -130
rect -3923 -718 -3865 -706
rect -3805 -130 -3747 -118
rect -3805 -706 -3793 -130
rect -3759 -706 -3747 -130
rect -3805 -718 -3747 -706
rect -3687 -130 -3629 -118
rect -3687 -706 -3675 -130
rect -3641 -706 -3629 -130
rect -3687 -718 -3629 -706
rect -3569 -130 -3511 -118
rect -3569 -706 -3557 -130
rect -3523 -706 -3511 -130
rect -3569 -718 -3511 -706
rect -3451 -130 -3393 -118
rect -3451 -706 -3439 -130
rect -3405 -706 -3393 -130
rect -3451 -718 -3393 -706
rect -3333 -130 -3275 -118
rect -3333 -706 -3321 -130
rect -3287 -706 -3275 -130
rect -3333 -718 -3275 -706
rect -3215 -130 -3157 -118
rect -3215 -706 -3203 -130
rect -3169 -706 -3157 -130
rect -3215 -718 -3157 -706
rect -3097 -130 -3039 -118
rect -3097 -706 -3085 -130
rect -3051 -706 -3039 -130
rect -3097 -718 -3039 -706
rect -2979 -130 -2921 -118
rect -2979 -706 -2967 -130
rect -2933 -706 -2921 -130
rect -2979 -718 -2921 -706
rect -2861 -130 -2803 -118
rect -2861 -706 -2849 -130
rect -2815 -706 -2803 -130
rect -2861 -718 -2803 -706
rect -2743 -130 -2685 -118
rect -2743 -706 -2731 -130
rect -2697 -706 -2685 -130
rect -2743 -718 -2685 -706
rect -2625 -130 -2567 -118
rect -2625 -706 -2613 -130
rect -2579 -706 -2567 -130
rect -2625 -718 -2567 -706
rect -2507 -130 -2449 -118
rect -2507 -706 -2495 -130
rect -2461 -706 -2449 -130
rect -2507 -718 -2449 -706
rect -2389 -130 -2331 -118
rect -2389 -706 -2377 -130
rect -2343 -706 -2331 -130
rect -2389 -718 -2331 -706
rect -2271 -130 -2213 -118
rect -2271 -706 -2259 -130
rect -2225 -706 -2213 -130
rect -2271 -718 -2213 -706
rect -2153 -130 -2095 -118
rect -2153 -706 -2141 -130
rect -2107 -706 -2095 -130
rect -2153 -718 -2095 -706
rect -2035 -130 -1977 -118
rect -2035 -706 -2023 -130
rect -1989 -706 -1977 -130
rect -2035 -718 -1977 -706
rect -1917 -130 -1859 -118
rect -1917 -706 -1905 -130
rect -1871 -706 -1859 -130
rect -1917 -718 -1859 -706
rect -1799 -130 -1741 -118
rect -1799 -706 -1787 -130
rect -1753 -706 -1741 -130
rect -1799 -718 -1741 -706
rect -1681 -130 -1623 -118
rect -1681 -706 -1669 -130
rect -1635 -706 -1623 -130
rect -1681 -718 -1623 -706
rect -1563 -130 -1505 -118
rect -1563 -706 -1551 -130
rect -1517 -706 -1505 -130
rect -1563 -718 -1505 -706
rect -1445 -130 -1387 -118
rect -1445 -706 -1433 -130
rect -1399 -706 -1387 -130
rect -1445 -718 -1387 -706
rect -1327 -130 -1269 -118
rect -1327 -706 -1315 -130
rect -1281 -706 -1269 -130
rect -1327 -718 -1269 -706
rect -1209 -130 -1151 -118
rect -1209 -706 -1197 -130
rect -1163 -706 -1151 -130
rect -1209 -718 -1151 -706
rect -1091 -130 -1033 -118
rect -1091 -706 -1079 -130
rect -1045 -706 -1033 -130
rect -1091 -718 -1033 -706
rect -973 -130 -915 -118
rect -973 -706 -961 -130
rect -927 -706 -915 -130
rect -973 -718 -915 -706
rect -855 -130 -797 -118
rect -855 -706 -843 -130
rect -809 -706 -797 -130
rect -855 -718 -797 -706
rect -737 -130 -679 -118
rect -737 -706 -725 -130
rect -691 -706 -679 -130
rect -737 -718 -679 -706
rect -619 -130 -561 -118
rect -619 -706 -607 -130
rect -573 -706 -561 -130
rect -619 -718 -561 -706
rect -501 -130 -443 -118
rect -501 -706 -489 -130
rect -455 -706 -443 -130
rect -501 -718 -443 -706
rect -383 -130 -325 -118
rect -383 -706 -371 -130
rect -337 -706 -325 -130
rect -383 -718 -325 -706
rect -265 -130 -207 -118
rect -265 -706 -253 -130
rect -219 -706 -207 -130
rect -265 -718 -207 -706
rect -147 -130 -89 -118
rect -147 -706 -135 -130
rect -101 -706 -89 -130
rect -147 -718 -89 -706
rect -29 -130 29 -118
rect -29 -706 -17 -130
rect 17 -706 29 -130
rect -29 -718 29 -706
rect 89 -130 147 -118
rect 89 -706 101 -130
rect 135 -706 147 -130
rect 89 -718 147 -706
rect 207 -130 265 -118
rect 207 -706 219 -130
rect 253 -706 265 -130
rect 207 -718 265 -706
rect 325 -130 383 -118
rect 325 -706 337 -130
rect 371 -706 383 -130
rect 325 -718 383 -706
rect 443 -130 501 -118
rect 443 -706 455 -130
rect 489 -706 501 -130
rect 443 -718 501 -706
rect 561 -130 619 -118
rect 561 -706 573 -130
rect 607 -706 619 -130
rect 561 -718 619 -706
rect 679 -130 737 -118
rect 679 -706 691 -130
rect 725 -706 737 -130
rect 679 -718 737 -706
rect 797 -130 855 -118
rect 797 -706 809 -130
rect 843 -706 855 -130
rect 797 -718 855 -706
rect 915 -130 973 -118
rect 915 -706 927 -130
rect 961 -706 973 -130
rect 915 -718 973 -706
rect 1033 -130 1091 -118
rect 1033 -706 1045 -130
rect 1079 -706 1091 -130
rect 1033 -718 1091 -706
rect 1151 -130 1209 -118
rect 1151 -706 1163 -130
rect 1197 -706 1209 -130
rect 1151 -718 1209 -706
rect 1269 -130 1327 -118
rect 1269 -706 1281 -130
rect 1315 -706 1327 -130
rect 1269 -718 1327 -706
rect 1387 -130 1445 -118
rect 1387 -706 1399 -130
rect 1433 -706 1445 -130
rect 1387 -718 1445 -706
rect 1505 -130 1563 -118
rect 1505 -706 1517 -130
rect 1551 -706 1563 -130
rect 1505 -718 1563 -706
rect 1623 -130 1681 -118
rect 1623 -706 1635 -130
rect 1669 -706 1681 -130
rect 1623 -718 1681 -706
rect 1741 -130 1799 -118
rect 1741 -706 1753 -130
rect 1787 -706 1799 -130
rect 1741 -718 1799 -706
rect 1859 -130 1917 -118
rect 1859 -706 1871 -130
rect 1905 -706 1917 -130
rect 1859 -718 1917 -706
rect 1977 -130 2035 -118
rect 1977 -706 1989 -130
rect 2023 -706 2035 -130
rect 1977 -718 2035 -706
rect 2095 -130 2153 -118
rect 2095 -706 2107 -130
rect 2141 -706 2153 -130
rect 2095 -718 2153 -706
rect 2213 -130 2271 -118
rect 2213 -706 2225 -130
rect 2259 -706 2271 -130
rect 2213 -718 2271 -706
rect 2331 -130 2389 -118
rect 2331 -706 2343 -130
rect 2377 -706 2389 -130
rect 2331 -718 2389 -706
rect 2449 -130 2507 -118
rect 2449 -706 2461 -130
rect 2495 -706 2507 -130
rect 2449 -718 2507 -706
rect 2567 -130 2625 -118
rect 2567 -706 2579 -130
rect 2613 -706 2625 -130
rect 2567 -718 2625 -706
rect 2685 -130 2743 -118
rect 2685 -706 2697 -130
rect 2731 -706 2743 -130
rect 2685 -718 2743 -706
rect 2803 -130 2861 -118
rect 2803 -706 2815 -130
rect 2849 -706 2861 -130
rect 2803 -718 2861 -706
rect 2921 -130 2979 -118
rect 2921 -706 2933 -130
rect 2967 -706 2979 -130
rect 2921 -718 2979 -706
rect 3039 -130 3097 -118
rect 3039 -706 3051 -130
rect 3085 -706 3097 -130
rect 3039 -718 3097 -706
rect 3157 -130 3215 -118
rect 3157 -706 3169 -130
rect 3203 -706 3215 -130
rect 3157 -718 3215 -706
rect 3275 -130 3333 -118
rect 3275 -706 3287 -130
rect 3321 -706 3333 -130
rect 3275 -718 3333 -706
rect 3393 -130 3451 -118
rect 3393 -706 3405 -130
rect 3439 -706 3451 -130
rect 3393 -718 3451 -706
rect 3511 -130 3569 -118
rect 3511 -706 3523 -130
rect 3557 -706 3569 -130
rect 3511 -718 3569 -706
rect 3629 -130 3687 -118
rect 3629 -706 3641 -130
rect 3675 -706 3687 -130
rect 3629 -718 3687 -706
rect 3747 -130 3805 -118
rect 3747 -706 3759 -130
rect 3793 -706 3805 -130
rect 3747 -718 3805 -706
rect 3865 -130 3923 -118
rect 3865 -706 3877 -130
rect 3911 -706 3923 -130
rect 3865 -718 3923 -706
rect 3983 -130 4041 -118
rect 3983 -706 3995 -130
rect 4029 -706 4041 -130
rect 3983 -718 4041 -706
rect 4101 -130 4159 -118
rect 4101 -706 4113 -130
rect 4147 -706 4159 -130
rect 4101 -718 4159 -706
rect 4219 -130 4277 -118
rect 4219 -706 4231 -130
rect 4265 -706 4277 -130
rect 4219 -718 4277 -706
rect 4337 -130 4395 -118
rect 4337 -706 4349 -130
rect 4383 -706 4395 -130
rect 4337 -718 4395 -706
rect 4455 -130 4513 -118
rect 4455 -706 4467 -130
rect 4501 -706 4513 -130
rect 4455 -718 4513 -706
rect 4573 -130 4631 -118
rect 4573 -706 4585 -130
rect 4619 -706 4631 -130
rect 4573 -718 4631 -706
rect 4691 -130 4749 -118
rect 4691 -706 4703 -130
rect 4737 -706 4749 -130
rect 4691 -718 4749 -706
rect 4809 -130 4867 -118
rect 4809 -706 4821 -130
rect 4855 -706 4867 -130
rect 4809 -718 4867 -706
rect 4927 -130 4985 -118
rect 4927 -706 4939 -130
rect 4973 -706 4985 -130
rect 4927 -718 4985 -706
rect 5045 -130 5103 -118
rect 5045 -706 5057 -130
rect 5091 -706 5103 -130
rect 5045 -718 5103 -706
rect 5163 -130 5221 -118
rect 5163 -706 5175 -130
rect 5209 -706 5221 -130
rect 5163 -718 5221 -706
rect 5281 -130 5339 -118
rect 5281 -706 5293 -130
rect 5327 -706 5339 -130
rect 5281 -718 5339 -706
rect 5399 -130 5457 -118
rect 5399 -706 5411 -130
rect 5445 -706 5457 -130
rect 5399 -718 5457 -706
rect 5517 -130 5575 -118
rect 5517 -706 5529 -130
rect 5563 -706 5575 -130
rect 5517 -718 5575 -706
rect 5635 -130 5693 -118
rect 5635 -706 5647 -130
rect 5681 -706 5693 -130
rect 5635 -718 5693 -706
rect 5753 -130 5811 -118
rect 5753 -706 5765 -130
rect 5799 -706 5811 -130
rect 5753 -718 5811 -706
rect 5871 -130 5929 -118
rect 5871 -706 5883 -130
rect 5917 -706 5929 -130
rect 5871 -718 5929 -706
rect 5989 -130 6047 -118
rect 5989 -706 6001 -130
rect 6035 -706 6047 -130
rect 5989 -718 6047 -706
rect 6107 -130 6165 -118
rect 6107 -706 6119 -130
rect 6153 -706 6165 -130
rect 6107 -718 6165 -706
rect 6225 -130 6283 -118
rect 6225 -706 6237 -130
rect 6271 -706 6283 -130
rect 6225 -718 6283 -706
rect 6343 -130 6401 -118
rect 6343 -706 6355 -130
rect 6389 -706 6401 -130
rect 6343 -718 6401 -706
rect 6461 -130 6519 -118
rect 6461 -706 6473 -130
rect 6507 -706 6519 -130
rect 6461 -718 6519 -706
rect 6579 -130 6637 -118
rect 6579 -706 6591 -130
rect 6625 -706 6637 -130
rect 6579 -718 6637 -706
rect 6697 -130 6755 -118
rect 6697 -706 6709 -130
rect 6743 -706 6755 -130
rect 6697 -718 6755 -706
rect 6815 -130 6873 -118
rect 6815 -706 6827 -130
rect 6861 -706 6873 -130
rect 6815 -718 6873 -706
rect 6933 -130 6991 -118
rect 6933 -706 6945 -130
rect 6979 -706 6991 -130
rect 6933 -718 6991 -706
rect 7051 -130 7109 -118
rect 7051 -706 7063 -130
rect 7097 -706 7109 -130
rect 7051 -718 7109 -706
<< pdiffc >>
rect -7097 130 -7063 706
rect -6979 130 -6945 706
rect -6861 130 -6827 706
rect -6743 130 -6709 706
rect -6625 130 -6591 706
rect -6507 130 -6473 706
rect -6389 130 -6355 706
rect -6271 130 -6237 706
rect -6153 130 -6119 706
rect -6035 130 -6001 706
rect -5917 130 -5883 706
rect -5799 130 -5765 706
rect -5681 130 -5647 706
rect -5563 130 -5529 706
rect -5445 130 -5411 706
rect -5327 130 -5293 706
rect -5209 130 -5175 706
rect -5091 130 -5057 706
rect -4973 130 -4939 706
rect -4855 130 -4821 706
rect -4737 130 -4703 706
rect -4619 130 -4585 706
rect -4501 130 -4467 706
rect -4383 130 -4349 706
rect -4265 130 -4231 706
rect -4147 130 -4113 706
rect -4029 130 -3995 706
rect -3911 130 -3877 706
rect -3793 130 -3759 706
rect -3675 130 -3641 706
rect -3557 130 -3523 706
rect -3439 130 -3405 706
rect -3321 130 -3287 706
rect -3203 130 -3169 706
rect -3085 130 -3051 706
rect -2967 130 -2933 706
rect -2849 130 -2815 706
rect -2731 130 -2697 706
rect -2613 130 -2579 706
rect -2495 130 -2461 706
rect -2377 130 -2343 706
rect -2259 130 -2225 706
rect -2141 130 -2107 706
rect -2023 130 -1989 706
rect -1905 130 -1871 706
rect -1787 130 -1753 706
rect -1669 130 -1635 706
rect -1551 130 -1517 706
rect -1433 130 -1399 706
rect -1315 130 -1281 706
rect -1197 130 -1163 706
rect -1079 130 -1045 706
rect -961 130 -927 706
rect -843 130 -809 706
rect -725 130 -691 706
rect -607 130 -573 706
rect -489 130 -455 706
rect -371 130 -337 706
rect -253 130 -219 706
rect -135 130 -101 706
rect -17 130 17 706
rect 101 130 135 706
rect 219 130 253 706
rect 337 130 371 706
rect 455 130 489 706
rect 573 130 607 706
rect 691 130 725 706
rect 809 130 843 706
rect 927 130 961 706
rect 1045 130 1079 706
rect 1163 130 1197 706
rect 1281 130 1315 706
rect 1399 130 1433 706
rect 1517 130 1551 706
rect 1635 130 1669 706
rect 1753 130 1787 706
rect 1871 130 1905 706
rect 1989 130 2023 706
rect 2107 130 2141 706
rect 2225 130 2259 706
rect 2343 130 2377 706
rect 2461 130 2495 706
rect 2579 130 2613 706
rect 2697 130 2731 706
rect 2815 130 2849 706
rect 2933 130 2967 706
rect 3051 130 3085 706
rect 3169 130 3203 706
rect 3287 130 3321 706
rect 3405 130 3439 706
rect 3523 130 3557 706
rect 3641 130 3675 706
rect 3759 130 3793 706
rect 3877 130 3911 706
rect 3995 130 4029 706
rect 4113 130 4147 706
rect 4231 130 4265 706
rect 4349 130 4383 706
rect 4467 130 4501 706
rect 4585 130 4619 706
rect 4703 130 4737 706
rect 4821 130 4855 706
rect 4939 130 4973 706
rect 5057 130 5091 706
rect 5175 130 5209 706
rect 5293 130 5327 706
rect 5411 130 5445 706
rect 5529 130 5563 706
rect 5647 130 5681 706
rect 5765 130 5799 706
rect 5883 130 5917 706
rect 6001 130 6035 706
rect 6119 130 6153 706
rect 6237 130 6271 706
rect 6355 130 6389 706
rect 6473 130 6507 706
rect 6591 130 6625 706
rect 6709 130 6743 706
rect 6827 130 6861 706
rect 6945 130 6979 706
rect 7063 130 7097 706
rect -7097 -706 -7063 -130
rect -6979 -706 -6945 -130
rect -6861 -706 -6827 -130
rect -6743 -706 -6709 -130
rect -6625 -706 -6591 -130
rect -6507 -706 -6473 -130
rect -6389 -706 -6355 -130
rect -6271 -706 -6237 -130
rect -6153 -706 -6119 -130
rect -6035 -706 -6001 -130
rect -5917 -706 -5883 -130
rect -5799 -706 -5765 -130
rect -5681 -706 -5647 -130
rect -5563 -706 -5529 -130
rect -5445 -706 -5411 -130
rect -5327 -706 -5293 -130
rect -5209 -706 -5175 -130
rect -5091 -706 -5057 -130
rect -4973 -706 -4939 -130
rect -4855 -706 -4821 -130
rect -4737 -706 -4703 -130
rect -4619 -706 -4585 -130
rect -4501 -706 -4467 -130
rect -4383 -706 -4349 -130
rect -4265 -706 -4231 -130
rect -4147 -706 -4113 -130
rect -4029 -706 -3995 -130
rect -3911 -706 -3877 -130
rect -3793 -706 -3759 -130
rect -3675 -706 -3641 -130
rect -3557 -706 -3523 -130
rect -3439 -706 -3405 -130
rect -3321 -706 -3287 -130
rect -3203 -706 -3169 -130
rect -3085 -706 -3051 -130
rect -2967 -706 -2933 -130
rect -2849 -706 -2815 -130
rect -2731 -706 -2697 -130
rect -2613 -706 -2579 -130
rect -2495 -706 -2461 -130
rect -2377 -706 -2343 -130
rect -2259 -706 -2225 -130
rect -2141 -706 -2107 -130
rect -2023 -706 -1989 -130
rect -1905 -706 -1871 -130
rect -1787 -706 -1753 -130
rect -1669 -706 -1635 -130
rect -1551 -706 -1517 -130
rect -1433 -706 -1399 -130
rect -1315 -706 -1281 -130
rect -1197 -706 -1163 -130
rect -1079 -706 -1045 -130
rect -961 -706 -927 -130
rect -843 -706 -809 -130
rect -725 -706 -691 -130
rect -607 -706 -573 -130
rect -489 -706 -455 -130
rect -371 -706 -337 -130
rect -253 -706 -219 -130
rect -135 -706 -101 -130
rect -17 -706 17 -130
rect 101 -706 135 -130
rect 219 -706 253 -130
rect 337 -706 371 -130
rect 455 -706 489 -130
rect 573 -706 607 -130
rect 691 -706 725 -130
rect 809 -706 843 -130
rect 927 -706 961 -130
rect 1045 -706 1079 -130
rect 1163 -706 1197 -130
rect 1281 -706 1315 -130
rect 1399 -706 1433 -130
rect 1517 -706 1551 -130
rect 1635 -706 1669 -130
rect 1753 -706 1787 -130
rect 1871 -706 1905 -130
rect 1989 -706 2023 -130
rect 2107 -706 2141 -130
rect 2225 -706 2259 -130
rect 2343 -706 2377 -130
rect 2461 -706 2495 -130
rect 2579 -706 2613 -130
rect 2697 -706 2731 -130
rect 2815 -706 2849 -130
rect 2933 -706 2967 -130
rect 3051 -706 3085 -130
rect 3169 -706 3203 -130
rect 3287 -706 3321 -130
rect 3405 -706 3439 -130
rect 3523 -706 3557 -130
rect 3641 -706 3675 -130
rect 3759 -706 3793 -130
rect 3877 -706 3911 -130
rect 3995 -706 4029 -130
rect 4113 -706 4147 -130
rect 4231 -706 4265 -130
rect 4349 -706 4383 -130
rect 4467 -706 4501 -130
rect 4585 -706 4619 -130
rect 4703 -706 4737 -130
rect 4821 -706 4855 -130
rect 4939 -706 4973 -130
rect 5057 -706 5091 -130
rect 5175 -706 5209 -130
rect 5293 -706 5327 -130
rect 5411 -706 5445 -130
rect 5529 -706 5563 -130
rect 5647 -706 5681 -130
rect 5765 -706 5799 -130
rect 5883 -706 5917 -130
rect 6001 -706 6035 -130
rect 6119 -706 6153 -130
rect 6237 -706 6271 -130
rect 6355 -706 6389 -130
rect 6473 -706 6507 -130
rect 6591 -706 6625 -130
rect 6709 -706 6743 -130
rect 6827 -706 6861 -130
rect 6945 -706 6979 -130
rect 7063 -706 7097 -130
<< nsubdiff >>
rect -7211 867 -7115 901
rect 7115 867 7211 901
rect -7211 805 -7177 867
rect 7177 805 7211 867
rect -7211 -867 -7177 -805
rect 7177 -867 7211 -805
rect -7211 -901 -7115 -867
rect 7115 -901 7211 -867
<< nsubdiffcont >>
rect -7115 867 7115 901
rect -7211 -805 -7177 805
rect 7177 -805 7211 805
rect -7115 -901 7115 -867
<< poly >>
rect -7054 799 -6988 815
rect -7054 765 -7038 799
rect -7004 765 -6988 799
rect -7054 749 -6988 765
rect -6936 799 -6870 815
rect -6936 765 -6920 799
rect -6886 765 -6870 799
rect -6936 749 -6870 765
rect -6818 799 -6752 815
rect -6818 765 -6802 799
rect -6768 765 -6752 799
rect -6818 749 -6752 765
rect -6700 799 -6634 815
rect -6700 765 -6684 799
rect -6650 765 -6634 799
rect -6700 749 -6634 765
rect -6582 799 -6516 815
rect -6582 765 -6566 799
rect -6532 765 -6516 799
rect -6582 749 -6516 765
rect -6464 799 -6398 815
rect -6464 765 -6448 799
rect -6414 765 -6398 799
rect -6464 749 -6398 765
rect -6346 799 -6280 815
rect -6346 765 -6330 799
rect -6296 765 -6280 799
rect -6346 749 -6280 765
rect -6228 799 -6162 815
rect -6228 765 -6212 799
rect -6178 765 -6162 799
rect -6228 749 -6162 765
rect -6110 799 -6044 815
rect -6110 765 -6094 799
rect -6060 765 -6044 799
rect -6110 749 -6044 765
rect -5992 799 -5926 815
rect -5992 765 -5976 799
rect -5942 765 -5926 799
rect -5992 749 -5926 765
rect -5874 799 -5808 815
rect -5874 765 -5858 799
rect -5824 765 -5808 799
rect -5874 749 -5808 765
rect -5756 799 -5690 815
rect -5756 765 -5740 799
rect -5706 765 -5690 799
rect -5756 749 -5690 765
rect -5638 799 -5572 815
rect -5638 765 -5622 799
rect -5588 765 -5572 799
rect -5638 749 -5572 765
rect -5520 799 -5454 815
rect -5520 765 -5504 799
rect -5470 765 -5454 799
rect -5520 749 -5454 765
rect -5402 799 -5336 815
rect -5402 765 -5386 799
rect -5352 765 -5336 799
rect -5402 749 -5336 765
rect -5284 799 -5218 815
rect -5284 765 -5268 799
rect -5234 765 -5218 799
rect -5284 749 -5218 765
rect -5166 799 -5100 815
rect -5166 765 -5150 799
rect -5116 765 -5100 799
rect -5166 749 -5100 765
rect -5048 799 -4982 815
rect -5048 765 -5032 799
rect -4998 765 -4982 799
rect -5048 749 -4982 765
rect -4930 799 -4864 815
rect -4930 765 -4914 799
rect -4880 765 -4864 799
rect -4930 749 -4864 765
rect -4812 799 -4746 815
rect -4812 765 -4796 799
rect -4762 765 -4746 799
rect -4812 749 -4746 765
rect -4694 799 -4628 815
rect -4694 765 -4678 799
rect -4644 765 -4628 799
rect -4694 749 -4628 765
rect -4576 799 -4510 815
rect -4576 765 -4560 799
rect -4526 765 -4510 799
rect -4576 749 -4510 765
rect -4458 799 -4392 815
rect -4458 765 -4442 799
rect -4408 765 -4392 799
rect -4458 749 -4392 765
rect -4340 799 -4274 815
rect -4340 765 -4324 799
rect -4290 765 -4274 799
rect -4340 749 -4274 765
rect -4222 799 -4156 815
rect -4222 765 -4206 799
rect -4172 765 -4156 799
rect -4222 749 -4156 765
rect -4104 799 -4038 815
rect -4104 765 -4088 799
rect -4054 765 -4038 799
rect -4104 749 -4038 765
rect -3986 799 -3920 815
rect -3986 765 -3970 799
rect -3936 765 -3920 799
rect -3986 749 -3920 765
rect -3868 799 -3802 815
rect -3868 765 -3852 799
rect -3818 765 -3802 799
rect -3868 749 -3802 765
rect -3750 799 -3684 815
rect -3750 765 -3734 799
rect -3700 765 -3684 799
rect -3750 749 -3684 765
rect -3632 799 -3566 815
rect -3632 765 -3616 799
rect -3582 765 -3566 799
rect -3632 749 -3566 765
rect -3514 799 -3448 815
rect -3514 765 -3498 799
rect -3464 765 -3448 799
rect -3514 749 -3448 765
rect -3396 799 -3330 815
rect -3396 765 -3380 799
rect -3346 765 -3330 799
rect -3396 749 -3330 765
rect -3278 799 -3212 815
rect -3278 765 -3262 799
rect -3228 765 -3212 799
rect -3278 749 -3212 765
rect -3160 799 -3094 815
rect -3160 765 -3144 799
rect -3110 765 -3094 799
rect -3160 749 -3094 765
rect -3042 799 -2976 815
rect -3042 765 -3026 799
rect -2992 765 -2976 799
rect -3042 749 -2976 765
rect -2924 799 -2858 815
rect -2924 765 -2908 799
rect -2874 765 -2858 799
rect -2924 749 -2858 765
rect -2806 799 -2740 815
rect -2806 765 -2790 799
rect -2756 765 -2740 799
rect -2806 749 -2740 765
rect -2688 799 -2622 815
rect -2688 765 -2672 799
rect -2638 765 -2622 799
rect -2688 749 -2622 765
rect -2570 799 -2504 815
rect -2570 765 -2554 799
rect -2520 765 -2504 799
rect -2570 749 -2504 765
rect -2452 799 -2386 815
rect -2452 765 -2436 799
rect -2402 765 -2386 799
rect -2452 749 -2386 765
rect -2334 799 -2268 815
rect -2334 765 -2318 799
rect -2284 765 -2268 799
rect -2334 749 -2268 765
rect -2216 799 -2150 815
rect -2216 765 -2200 799
rect -2166 765 -2150 799
rect -2216 749 -2150 765
rect -2098 799 -2032 815
rect -2098 765 -2082 799
rect -2048 765 -2032 799
rect -2098 749 -2032 765
rect -1980 799 -1914 815
rect -1980 765 -1964 799
rect -1930 765 -1914 799
rect -1980 749 -1914 765
rect -1862 799 -1796 815
rect -1862 765 -1846 799
rect -1812 765 -1796 799
rect -1862 749 -1796 765
rect -1744 799 -1678 815
rect -1744 765 -1728 799
rect -1694 765 -1678 799
rect -1744 749 -1678 765
rect -1626 799 -1560 815
rect -1626 765 -1610 799
rect -1576 765 -1560 799
rect -1626 749 -1560 765
rect -1508 799 -1442 815
rect -1508 765 -1492 799
rect -1458 765 -1442 799
rect -1508 749 -1442 765
rect -1390 799 -1324 815
rect -1390 765 -1374 799
rect -1340 765 -1324 799
rect -1390 749 -1324 765
rect -1272 799 -1206 815
rect -1272 765 -1256 799
rect -1222 765 -1206 799
rect -1272 749 -1206 765
rect -1154 799 -1088 815
rect -1154 765 -1138 799
rect -1104 765 -1088 799
rect -1154 749 -1088 765
rect -1036 799 -970 815
rect -1036 765 -1020 799
rect -986 765 -970 799
rect -1036 749 -970 765
rect -918 799 -852 815
rect -918 765 -902 799
rect -868 765 -852 799
rect -918 749 -852 765
rect -800 799 -734 815
rect -800 765 -784 799
rect -750 765 -734 799
rect -800 749 -734 765
rect -682 799 -616 815
rect -682 765 -666 799
rect -632 765 -616 799
rect -682 749 -616 765
rect -564 799 -498 815
rect -564 765 -548 799
rect -514 765 -498 799
rect -564 749 -498 765
rect -446 799 -380 815
rect -446 765 -430 799
rect -396 765 -380 799
rect -446 749 -380 765
rect -328 799 -262 815
rect -328 765 -312 799
rect -278 765 -262 799
rect -328 749 -262 765
rect -210 799 -144 815
rect -210 765 -194 799
rect -160 765 -144 799
rect -210 749 -144 765
rect -92 799 -26 815
rect -92 765 -76 799
rect -42 765 -26 799
rect -92 749 -26 765
rect 26 799 92 815
rect 26 765 42 799
rect 76 765 92 799
rect 26 749 92 765
rect 144 799 210 815
rect 144 765 160 799
rect 194 765 210 799
rect 144 749 210 765
rect 262 799 328 815
rect 262 765 278 799
rect 312 765 328 799
rect 262 749 328 765
rect 380 799 446 815
rect 380 765 396 799
rect 430 765 446 799
rect 380 749 446 765
rect 498 799 564 815
rect 498 765 514 799
rect 548 765 564 799
rect 498 749 564 765
rect 616 799 682 815
rect 616 765 632 799
rect 666 765 682 799
rect 616 749 682 765
rect 734 799 800 815
rect 734 765 750 799
rect 784 765 800 799
rect 734 749 800 765
rect 852 799 918 815
rect 852 765 868 799
rect 902 765 918 799
rect 852 749 918 765
rect 970 799 1036 815
rect 970 765 986 799
rect 1020 765 1036 799
rect 970 749 1036 765
rect 1088 799 1154 815
rect 1088 765 1104 799
rect 1138 765 1154 799
rect 1088 749 1154 765
rect 1206 799 1272 815
rect 1206 765 1222 799
rect 1256 765 1272 799
rect 1206 749 1272 765
rect 1324 799 1390 815
rect 1324 765 1340 799
rect 1374 765 1390 799
rect 1324 749 1390 765
rect 1442 799 1508 815
rect 1442 765 1458 799
rect 1492 765 1508 799
rect 1442 749 1508 765
rect 1560 799 1626 815
rect 1560 765 1576 799
rect 1610 765 1626 799
rect 1560 749 1626 765
rect 1678 799 1744 815
rect 1678 765 1694 799
rect 1728 765 1744 799
rect 1678 749 1744 765
rect 1796 799 1862 815
rect 1796 765 1812 799
rect 1846 765 1862 799
rect 1796 749 1862 765
rect 1914 799 1980 815
rect 1914 765 1930 799
rect 1964 765 1980 799
rect 1914 749 1980 765
rect 2032 799 2098 815
rect 2032 765 2048 799
rect 2082 765 2098 799
rect 2032 749 2098 765
rect 2150 799 2216 815
rect 2150 765 2166 799
rect 2200 765 2216 799
rect 2150 749 2216 765
rect 2268 799 2334 815
rect 2268 765 2284 799
rect 2318 765 2334 799
rect 2268 749 2334 765
rect 2386 799 2452 815
rect 2386 765 2402 799
rect 2436 765 2452 799
rect 2386 749 2452 765
rect 2504 799 2570 815
rect 2504 765 2520 799
rect 2554 765 2570 799
rect 2504 749 2570 765
rect 2622 799 2688 815
rect 2622 765 2638 799
rect 2672 765 2688 799
rect 2622 749 2688 765
rect 2740 799 2806 815
rect 2740 765 2756 799
rect 2790 765 2806 799
rect 2740 749 2806 765
rect 2858 799 2924 815
rect 2858 765 2874 799
rect 2908 765 2924 799
rect 2858 749 2924 765
rect 2976 799 3042 815
rect 2976 765 2992 799
rect 3026 765 3042 799
rect 2976 749 3042 765
rect 3094 799 3160 815
rect 3094 765 3110 799
rect 3144 765 3160 799
rect 3094 749 3160 765
rect 3212 799 3278 815
rect 3212 765 3228 799
rect 3262 765 3278 799
rect 3212 749 3278 765
rect 3330 799 3396 815
rect 3330 765 3346 799
rect 3380 765 3396 799
rect 3330 749 3396 765
rect 3448 799 3514 815
rect 3448 765 3464 799
rect 3498 765 3514 799
rect 3448 749 3514 765
rect 3566 799 3632 815
rect 3566 765 3582 799
rect 3616 765 3632 799
rect 3566 749 3632 765
rect 3684 799 3750 815
rect 3684 765 3700 799
rect 3734 765 3750 799
rect 3684 749 3750 765
rect 3802 799 3868 815
rect 3802 765 3818 799
rect 3852 765 3868 799
rect 3802 749 3868 765
rect 3920 799 3986 815
rect 3920 765 3936 799
rect 3970 765 3986 799
rect 3920 749 3986 765
rect 4038 799 4104 815
rect 4038 765 4054 799
rect 4088 765 4104 799
rect 4038 749 4104 765
rect 4156 799 4222 815
rect 4156 765 4172 799
rect 4206 765 4222 799
rect 4156 749 4222 765
rect 4274 799 4340 815
rect 4274 765 4290 799
rect 4324 765 4340 799
rect 4274 749 4340 765
rect 4392 799 4458 815
rect 4392 765 4408 799
rect 4442 765 4458 799
rect 4392 749 4458 765
rect 4510 799 4576 815
rect 4510 765 4526 799
rect 4560 765 4576 799
rect 4510 749 4576 765
rect 4628 799 4694 815
rect 4628 765 4644 799
rect 4678 765 4694 799
rect 4628 749 4694 765
rect 4746 799 4812 815
rect 4746 765 4762 799
rect 4796 765 4812 799
rect 4746 749 4812 765
rect 4864 799 4930 815
rect 4864 765 4880 799
rect 4914 765 4930 799
rect 4864 749 4930 765
rect 4982 799 5048 815
rect 4982 765 4998 799
rect 5032 765 5048 799
rect 4982 749 5048 765
rect 5100 799 5166 815
rect 5100 765 5116 799
rect 5150 765 5166 799
rect 5100 749 5166 765
rect 5218 799 5284 815
rect 5218 765 5234 799
rect 5268 765 5284 799
rect 5218 749 5284 765
rect 5336 799 5402 815
rect 5336 765 5352 799
rect 5386 765 5402 799
rect 5336 749 5402 765
rect 5454 799 5520 815
rect 5454 765 5470 799
rect 5504 765 5520 799
rect 5454 749 5520 765
rect 5572 799 5638 815
rect 5572 765 5588 799
rect 5622 765 5638 799
rect 5572 749 5638 765
rect 5690 799 5756 815
rect 5690 765 5706 799
rect 5740 765 5756 799
rect 5690 749 5756 765
rect 5808 799 5874 815
rect 5808 765 5824 799
rect 5858 765 5874 799
rect 5808 749 5874 765
rect 5926 799 5992 815
rect 5926 765 5942 799
rect 5976 765 5992 799
rect 5926 749 5992 765
rect 6044 799 6110 815
rect 6044 765 6060 799
rect 6094 765 6110 799
rect 6044 749 6110 765
rect 6162 799 6228 815
rect 6162 765 6178 799
rect 6212 765 6228 799
rect 6162 749 6228 765
rect 6280 799 6346 815
rect 6280 765 6296 799
rect 6330 765 6346 799
rect 6280 749 6346 765
rect 6398 799 6464 815
rect 6398 765 6414 799
rect 6448 765 6464 799
rect 6398 749 6464 765
rect 6516 799 6582 815
rect 6516 765 6532 799
rect 6566 765 6582 799
rect 6516 749 6582 765
rect 6634 799 6700 815
rect 6634 765 6650 799
rect 6684 765 6700 799
rect 6634 749 6700 765
rect 6752 799 6818 815
rect 6752 765 6768 799
rect 6802 765 6818 799
rect 6752 749 6818 765
rect 6870 799 6936 815
rect 6870 765 6886 799
rect 6920 765 6936 799
rect 6870 749 6936 765
rect 6988 799 7054 815
rect 6988 765 7004 799
rect 7038 765 7054 799
rect 6988 749 7054 765
rect -7051 718 -6991 749
rect -6933 718 -6873 749
rect -6815 718 -6755 749
rect -6697 718 -6637 749
rect -6579 718 -6519 749
rect -6461 718 -6401 749
rect -6343 718 -6283 749
rect -6225 718 -6165 749
rect -6107 718 -6047 749
rect -5989 718 -5929 749
rect -5871 718 -5811 749
rect -5753 718 -5693 749
rect -5635 718 -5575 749
rect -5517 718 -5457 749
rect -5399 718 -5339 749
rect -5281 718 -5221 749
rect -5163 718 -5103 749
rect -5045 718 -4985 749
rect -4927 718 -4867 749
rect -4809 718 -4749 749
rect -4691 718 -4631 749
rect -4573 718 -4513 749
rect -4455 718 -4395 749
rect -4337 718 -4277 749
rect -4219 718 -4159 749
rect -4101 718 -4041 749
rect -3983 718 -3923 749
rect -3865 718 -3805 749
rect -3747 718 -3687 749
rect -3629 718 -3569 749
rect -3511 718 -3451 749
rect -3393 718 -3333 749
rect -3275 718 -3215 749
rect -3157 718 -3097 749
rect -3039 718 -2979 749
rect -2921 718 -2861 749
rect -2803 718 -2743 749
rect -2685 718 -2625 749
rect -2567 718 -2507 749
rect -2449 718 -2389 749
rect -2331 718 -2271 749
rect -2213 718 -2153 749
rect -2095 718 -2035 749
rect -1977 718 -1917 749
rect -1859 718 -1799 749
rect -1741 718 -1681 749
rect -1623 718 -1563 749
rect -1505 718 -1445 749
rect -1387 718 -1327 749
rect -1269 718 -1209 749
rect -1151 718 -1091 749
rect -1033 718 -973 749
rect -915 718 -855 749
rect -797 718 -737 749
rect -679 718 -619 749
rect -561 718 -501 749
rect -443 718 -383 749
rect -325 718 -265 749
rect -207 718 -147 749
rect -89 718 -29 749
rect 29 718 89 749
rect 147 718 207 749
rect 265 718 325 749
rect 383 718 443 749
rect 501 718 561 749
rect 619 718 679 749
rect 737 718 797 749
rect 855 718 915 749
rect 973 718 1033 749
rect 1091 718 1151 749
rect 1209 718 1269 749
rect 1327 718 1387 749
rect 1445 718 1505 749
rect 1563 718 1623 749
rect 1681 718 1741 749
rect 1799 718 1859 749
rect 1917 718 1977 749
rect 2035 718 2095 749
rect 2153 718 2213 749
rect 2271 718 2331 749
rect 2389 718 2449 749
rect 2507 718 2567 749
rect 2625 718 2685 749
rect 2743 718 2803 749
rect 2861 718 2921 749
rect 2979 718 3039 749
rect 3097 718 3157 749
rect 3215 718 3275 749
rect 3333 718 3393 749
rect 3451 718 3511 749
rect 3569 718 3629 749
rect 3687 718 3747 749
rect 3805 718 3865 749
rect 3923 718 3983 749
rect 4041 718 4101 749
rect 4159 718 4219 749
rect 4277 718 4337 749
rect 4395 718 4455 749
rect 4513 718 4573 749
rect 4631 718 4691 749
rect 4749 718 4809 749
rect 4867 718 4927 749
rect 4985 718 5045 749
rect 5103 718 5163 749
rect 5221 718 5281 749
rect 5339 718 5399 749
rect 5457 718 5517 749
rect 5575 718 5635 749
rect 5693 718 5753 749
rect 5811 718 5871 749
rect 5929 718 5989 749
rect 6047 718 6107 749
rect 6165 718 6225 749
rect 6283 718 6343 749
rect 6401 718 6461 749
rect 6519 718 6579 749
rect 6637 718 6697 749
rect 6755 718 6815 749
rect 6873 718 6933 749
rect 6991 718 7051 749
rect -7051 87 -6991 118
rect -6933 87 -6873 118
rect -6815 87 -6755 118
rect -6697 87 -6637 118
rect -6579 87 -6519 118
rect -6461 87 -6401 118
rect -6343 87 -6283 118
rect -6225 87 -6165 118
rect -6107 87 -6047 118
rect -5989 87 -5929 118
rect -5871 87 -5811 118
rect -5753 87 -5693 118
rect -5635 87 -5575 118
rect -5517 87 -5457 118
rect -5399 87 -5339 118
rect -5281 87 -5221 118
rect -5163 87 -5103 118
rect -5045 87 -4985 118
rect -4927 87 -4867 118
rect -4809 87 -4749 118
rect -4691 87 -4631 118
rect -4573 87 -4513 118
rect -4455 87 -4395 118
rect -4337 87 -4277 118
rect -4219 87 -4159 118
rect -4101 87 -4041 118
rect -3983 87 -3923 118
rect -3865 87 -3805 118
rect -3747 87 -3687 118
rect -3629 87 -3569 118
rect -3511 87 -3451 118
rect -3393 87 -3333 118
rect -3275 87 -3215 118
rect -3157 87 -3097 118
rect -3039 87 -2979 118
rect -2921 87 -2861 118
rect -2803 87 -2743 118
rect -2685 87 -2625 118
rect -2567 87 -2507 118
rect -2449 87 -2389 118
rect -2331 87 -2271 118
rect -2213 87 -2153 118
rect -2095 87 -2035 118
rect -1977 87 -1917 118
rect -1859 87 -1799 118
rect -1741 87 -1681 118
rect -1623 87 -1563 118
rect -1505 87 -1445 118
rect -1387 87 -1327 118
rect -1269 87 -1209 118
rect -1151 87 -1091 118
rect -1033 87 -973 118
rect -915 87 -855 118
rect -797 87 -737 118
rect -679 87 -619 118
rect -561 87 -501 118
rect -443 87 -383 118
rect -325 87 -265 118
rect -207 87 -147 118
rect -89 87 -29 118
rect 29 87 89 118
rect 147 87 207 118
rect 265 87 325 118
rect 383 87 443 118
rect 501 87 561 118
rect 619 87 679 118
rect 737 87 797 118
rect 855 87 915 118
rect 973 87 1033 118
rect 1091 87 1151 118
rect 1209 87 1269 118
rect 1327 87 1387 118
rect 1445 87 1505 118
rect 1563 87 1623 118
rect 1681 87 1741 118
rect 1799 87 1859 118
rect 1917 87 1977 118
rect 2035 87 2095 118
rect 2153 87 2213 118
rect 2271 87 2331 118
rect 2389 87 2449 118
rect 2507 87 2567 118
rect 2625 87 2685 118
rect 2743 87 2803 118
rect 2861 87 2921 118
rect 2979 87 3039 118
rect 3097 87 3157 118
rect 3215 87 3275 118
rect 3333 87 3393 118
rect 3451 87 3511 118
rect 3569 87 3629 118
rect 3687 87 3747 118
rect 3805 87 3865 118
rect 3923 87 3983 118
rect 4041 87 4101 118
rect 4159 87 4219 118
rect 4277 87 4337 118
rect 4395 87 4455 118
rect 4513 87 4573 118
rect 4631 87 4691 118
rect 4749 87 4809 118
rect 4867 87 4927 118
rect 4985 87 5045 118
rect 5103 87 5163 118
rect 5221 87 5281 118
rect 5339 87 5399 118
rect 5457 87 5517 118
rect 5575 87 5635 118
rect 5693 87 5753 118
rect 5811 87 5871 118
rect 5929 87 5989 118
rect 6047 87 6107 118
rect 6165 87 6225 118
rect 6283 87 6343 118
rect 6401 87 6461 118
rect 6519 87 6579 118
rect 6637 87 6697 118
rect 6755 87 6815 118
rect 6873 87 6933 118
rect 6991 87 7051 118
rect -7054 71 -6988 87
rect -7054 37 -7038 71
rect -7004 37 -6988 71
rect -7054 21 -6988 37
rect -6936 71 -6870 87
rect -6936 37 -6920 71
rect -6886 37 -6870 71
rect -6936 21 -6870 37
rect -6818 71 -6752 87
rect -6818 37 -6802 71
rect -6768 37 -6752 71
rect -6818 21 -6752 37
rect -6700 71 -6634 87
rect -6700 37 -6684 71
rect -6650 37 -6634 71
rect -6700 21 -6634 37
rect -6582 71 -6516 87
rect -6582 37 -6566 71
rect -6532 37 -6516 71
rect -6582 21 -6516 37
rect -6464 71 -6398 87
rect -6464 37 -6448 71
rect -6414 37 -6398 71
rect -6464 21 -6398 37
rect -6346 71 -6280 87
rect -6346 37 -6330 71
rect -6296 37 -6280 71
rect -6346 21 -6280 37
rect -6228 71 -6162 87
rect -6228 37 -6212 71
rect -6178 37 -6162 71
rect -6228 21 -6162 37
rect -6110 71 -6044 87
rect -6110 37 -6094 71
rect -6060 37 -6044 71
rect -6110 21 -6044 37
rect -5992 71 -5926 87
rect -5992 37 -5976 71
rect -5942 37 -5926 71
rect -5992 21 -5926 37
rect -5874 71 -5808 87
rect -5874 37 -5858 71
rect -5824 37 -5808 71
rect -5874 21 -5808 37
rect -5756 71 -5690 87
rect -5756 37 -5740 71
rect -5706 37 -5690 71
rect -5756 21 -5690 37
rect -5638 71 -5572 87
rect -5638 37 -5622 71
rect -5588 37 -5572 71
rect -5638 21 -5572 37
rect -5520 71 -5454 87
rect -5520 37 -5504 71
rect -5470 37 -5454 71
rect -5520 21 -5454 37
rect -5402 71 -5336 87
rect -5402 37 -5386 71
rect -5352 37 -5336 71
rect -5402 21 -5336 37
rect -5284 71 -5218 87
rect -5284 37 -5268 71
rect -5234 37 -5218 71
rect -5284 21 -5218 37
rect -5166 71 -5100 87
rect -5166 37 -5150 71
rect -5116 37 -5100 71
rect -5166 21 -5100 37
rect -5048 71 -4982 87
rect -5048 37 -5032 71
rect -4998 37 -4982 71
rect -5048 21 -4982 37
rect -4930 71 -4864 87
rect -4930 37 -4914 71
rect -4880 37 -4864 71
rect -4930 21 -4864 37
rect -4812 71 -4746 87
rect -4812 37 -4796 71
rect -4762 37 -4746 71
rect -4812 21 -4746 37
rect -4694 71 -4628 87
rect -4694 37 -4678 71
rect -4644 37 -4628 71
rect -4694 21 -4628 37
rect -4576 71 -4510 87
rect -4576 37 -4560 71
rect -4526 37 -4510 71
rect -4576 21 -4510 37
rect -4458 71 -4392 87
rect -4458 37 -4442 71
rect -4408 37 -4392 71
rect -4458 21 -4392 37
rect -4340 71 -4274 87
rect -4340 37 -4324 71
rect -4290 37 -4274 71
rect -4340 21 -4274 37
rect -4222 71 -4156 87
rect -4222 37 -4206 71
rect -4172 37 -4156 71
rect -4222 21 -4156 37
rect -4104 71 -4038 87
rect -4104 37 -4088 71
rect -4054 37 -4038 71
rect -4104 21 -4038 37
rect -3986 71 -3920 87
rect -3986 37 -3970 71
rect -3936 37 -3920 71
rect -3986 21 -3920 37
rect -3868 71 -3802 87
rect -3868 37 -3852 71
rect -3818 37 -3802 71
rect -3868 21 -3802 37
rect -3750 71 -3684 87
rect -3750 37 -3734 71
rect -3700 37 -3684 71
rect -3750 21 -3684 37
rect -3632 71 -3566 87
rect -3632 37 -3616 71
rect -3582 37 -3566 71
rect -3632 21 -3566 37
rect -3514 71 -3448 87
rect -3514 37 -3498 71
rect -3464 37 -3448 71
rect -3514 21 -3448 37
rect -3396 71 -3330 87
rect -3396 37 -3380 71
rect -3346 37 -3330 71
rect -3396 21 -3330 37
rect -3278 71 -3212 87
rect -3278 37 -3262 71
rect -3228 37 -3212 71
rect -3278 21 -3212 37
rect -3160 71 -3094 87
rect -3160 37 -3144 71
rect -3110 37 -3094 71
rect -3160 21 -3094 37
rect -3042 71 -2976 87
rect -3042 37 -3026 71
rect -2992 37 -2976 71
rect -3042 21 -2976 37
rect -2924 71 -2858 87
rect -2924 37 -2908 71
rect -2874 37 -2858 71
rect -2924 21 -2858 37
rect -2806 71 -2740 87
rect -2806 37 -2790 71
rect -2756 37 -2740 71
rect -2806 21 -2740 37
rect -2688 71 -2622 87
rect -2688 37 -2672 71
rect -2638 37 -2622 71
rect -2688 21 -2622 37
rect -2570 71 -2504 87
rect -2570 37 -2554 71
rect -2520 37 -2504 71
rect -2570 21 -2504 37
rect -2452 71 -2386 87
rect -2452 37 -2436 71
rect -2402 37 -2386 71
rect -2452 21 -2386 37
rect -2334 71 -2268 87
rect -2334 37 -2318 71
rect -2284 37 -2268 71
rect -2334 21 -2268 37
rect -2216 71 -2150 87
rect -2216 37 -2200 71
rect -2166 37 -2150 71
rect -2216 21 -2150 37
rect -2098 71 -2032 87
rect -2098 37 -2082 71
rect -2048 37 -2032 71
rect -2098 21 -2032 37
rect -1980 71 -1914 87
rect -1980 37 -1964 71
rect -1930 37 -1914 71
rect -1980 21 -1914 37
rect -1862 71 -1796 87
rect -1862 37 -1846 71
rect -1812 37 -1796 71
rect -1862 21 -1796 37
rect -1744 71 -1678 87
rect -1744 37 -1728 71
rect -1694 37 -1678 71
rect -1744 21 -1678 37
rect -1626 71 -1560 87
rect -1626 37 -1610 71
rect -1576 37 -1560 71
rect -1626 21 -1560 37
rect -1508 71 -1442 87
rect -1508 37 -1492 71
rect -1458 37 -1442 71
rect -1508 21 -1442 37
rect -1390 71 -1324 87
rect -1390 37 -1374 71
rect -1340 37 -1324 71
rect -1390 21 -1324 37
rect -1272 71 -1206 87
rect -1272 37 -1256 71
rect -1222 37 -1206 71
rect -1272 21 -1206 37
rect -1154 71 -1088 87
rect -1154 37 -1138 71
rect -1104 37 -1088 71
rect -1154 21 -1088 37
rect -1036 71 -970 87
rect -1036 37 -1020 71
rect -986 37 -970 71
rect -1036 21 -970 37
rect -918 71 -852 87
rect -918 37 -902 71
rect -868 37 -852 71
rect -918 21 -852 37
rect -800 71 -734 87
rect -800 37 -784 71
rect -750 37 -734 71
rect -800 21 -734 37
rect -682 71 -616 87
rect -682 37 -666 71
rect -632 37 -616 71
rect -682 21 -616 37
rect -564 71 -498 87
rect -564 37 -548 71
rect -514 37 -498 71
rect -564 21 -498 37
rect -446 71 -380 87
rect -446 37 -430 71
rect -396 37 -380 71
rect -446 21 -380 37
rect -328 71 -262 87
rect -328 37 -312 71
rect -278 37 -262 71
rect -328 21 -262 37
rect -210 71 -144 87
rect -210 37 -194 71
rect -160 37 -144 71
rect -210 21 -144 37
rect -92 71 -26 87
rect -92 37 -76 71
rect -42 37 -26 71
rect -92 21 -26 37
rect 26 71 92 87
rect 26 37 42 71
rect 76 37 92 71
rect 26 21 92 37
rect 144 71 210 87
rect 144 37 160 71
rect 194 37 210 71
rect 144 21 210 37
rect 262 71 328 87
rect 262 37 278 71
rect 312 37 328 71
rect 262 21 328 37
rect 380 71 446 87
rect 380 37 396 71
rect 430 37 446 71
rect 380 21 446 37
rect 498 71 564 87
rect 498 37 514 71
rect 548 37 564 71
rect 498 21 564 37
rect 616 71 682 87
rect 616 37 632 71
rect 666 37 682 71
rect 616 21 682 37
rect 734 71 800 87
rect 734 37 750 71
rect 784 37 800 71
rect 734 21 800 37
rect 852 71 918 87
rect 852 37 868 71
rect 902 37 918 71
rect 852 21 918 37
rect 970 71 1036 87
rect 970 37 986 71
rect 1020 37 1036 71
rect 970 21 1036 37
rect 1088 71 1154 87
rect 1088 37 1104 71
rect 1138 37 1154 71
rect 1088 21 1154 37
rect 1206 71 1272 87
rect 1206 37 1222 71
rect 1256 37 1272 71
rect 1206 21 1272 37
rect 1324 71 1390 87
rect 1324 37 1340 71
rect 1374 37 1390 71
rect 1324 21 1390 37
rect 1442 71 1508 87
rect 1442 37 1458 71
rect 1492 37 1508 71
rect 1442 21 1508 37
rect 1560 71 1626 87
rect 1560 37 1576 71
rect 1610 37 1626 71
rect 1560 21 1626 37
rect 1678 71 1744 87
rect 1678 37 1694 71
rect 1728 37 1744 71
rect 1678 21 1744 37
rect 1796 71 1862 87
rect 1796 37 1812 71
rect 1846 37 1862 71
rect 1796 21 1862 37
rect 1914 71 1980 87
rect 1914 37 1930 71
rect 1964 37 1980 71
rect 1914 21 1980 37
rect 2032 71 2098 87
rect 2032 37 2048 71
rect 2082 37 2098 71
rect 2032 21 2098 37
rect 2150 71 2216 87
rect 2150 37 2166 71
rect 2200 37 2216 71
rect 2150 21 2216 37
rect 2268 71 2334 87
rect 2268 37 2284 71
rect 2318 37 2334 71
rect 2268 21 2334 37
rect 2386 71 2452 87
rect 2386 37 2402 71
rect 2436 37 2452 71
rect 2386 21 2452 37
rect 2504 71 2570 87
rect 2504 37 2520 71
rect 2554 37 2570 71
rect 2504 21 2570 37
rect 2622 71 2688 87
rect 2622 37 2638 71
rect 2672 37 2688 71
rect 2622 21 2688 37
rect 2740 71 2806 87
rect 2740 37 2756 71
rect 2790 37 2806 71
rect 2740 21 2806 37
rect 2858 71 2924 87
rect 2858 37 2874 71
rect 2908 37 2924 71
rect 2858 21 2924 37
rect 2976 71 3042 87
rect 2976 37 2992 71
rect 3026 37 3042 71
rect 2976 21 3042 37
rect 3094 71 3160 87
rect 3094 37 3110 71
rect 3144 37 3160 71
rect 3094 21 3160 37
rect 3212 71 3278 87
rect 3212 37 3228 71
rect 3262 37 3278 71
rect 3212 21 3278 37
rect 3330 71 3396 87
rect 3330 37 3346 71
rect 3380 37 3396 71
rect 3330 21 3396 37
rect 3448 71 3514 87
rect 3448 37 3464 71
rect 3498 37 3514 71
rect 3448 21 3514 37
rect 3566 71 3632 87
rect 3566 37 3582 71
rect 3616 37 3632 71
rect 3566 21 3632 37
rect 3684 71 3750 87
rect 3684 37 3700 71
rect 3734 37 3750 71
rect 3684 21 3750 37
rect 3802 71 3868 87
rect 3802 37 3818 71
rect 3852 37 3868 71
rect 3802 21 3868 37
rect 3920 71 3986 87
rect 3920 37 3936 71
rect 3970 37 3986 71
rect 3920 21 3986 37
rect 4038 71 4104 87
rect 4038 37 4054 71
rect 4088 37 4104 71
rect 4038 21 4104 37
rect 4156 71 4222 87
rect 4156 37 4172 71
rect 4206 37 4222 71
rect 4156 21 4222 37
rect 4274 71 4340 87
rect 4274 37 4290 71
rect 4324 37 4340 71
rect 4274 21 4340 37
rect 4392 71 4458 87
rect 4392 37 4408 71
rect 4442 37 4458 71
rect 4392 21 4458 37
rect 4510 71 4576 87
rect 4510 37 4526 71
rect 4560 37 4576 71
rect 4510 21 4576 37
rect 4628 71 4694 87
rect 4628 37 4644 71
rect 4678 37 4694 71
rect 4628 21 4694 37
rect 4746 71 4812 87
rect 4746 37 4762 71
rect 4796 37 4812 71
rect 4746 21 4812 37
rect 4864 71 4930 87
rect 4864 37 4880 71
rect 4914 37 4930 71
rect 4864 21 4930 37
rect 4982 71 5048 87
rect 4982 37 4998 71
rect 5032 37 5048 71
rect 4982 21 5048 37
rect 5100 71 5166 87
rect 5100 37 5116 71
rect 5150 37 5166 71
rect 5100 21 5166 37
rect 5218 71 5284 87
rect 5218 37 5234 71
rect 5268 37 5284 71
rect 5218 21 5284 37
rect 5336 71 5402 87
rect 5336 37 5352 71
rect 5386 37 5402 71
rect 5336 21 5402 37
rect 5454 71 5520 87
rect 5454 37 5470 71
rect 5504 37 5520 71
rect 5454 21 5520 37
rect 5572 71 5638 87
rect 5572 37 5588 71
rect 5622 37 5638 71
rect 5572 21 5638 37
rect 5690 71 5756 87
rect 5690 37 5706 71
rect 5740 37 5756 71
rect 5690 21 5756 37
rect 5808 71 5874 87
rect 5808 37 5824 71
rect 5858 37 5874 71
rect 5808 21 5874 37
rect 5926 71 5992 87
rect 5926 37 5942 71
rect 5976 37 5992 71
rect 5926 21 5992 37
rect 6044 71 6110 87
rect 6044 37 6060 71
rect 6094 37 6110 71
rect 6044 21 6110 37
rect 6162 71 6228 87
rect 6162 37 6178 71
rect 6212 37 6228 71
rect 6162 21 6228 37
rect 6280 71 6346 87
rect 6280 37 6296 71
rect 6330 37 6346 71
rect 6280 21 6346 37
rect 6398 71 6464 87
rect 6398 37 6414 71
rect 6448 37 6464 71
rect 6398 21 6464 37
rect 6516 71 6582 87
rect 6516 37 6532 71
rect 6566 37 6582 71
rect 6516 21 6582 37
rect 6634 71 6700 87
rect 6634 37 6650 71
rect 6684 37 6700 71
rect 6634 21 6700 37
rect 6752 71 6818 87
rect 6752 37 6768 71
rect 6802 37 6818 71
rect 6752 21 6818 37
rect 6870 71 6936 87
rect 6870 37 6886 71
rect 6920 37 6936 71
rect 6870 21 6936 37
rect 6988 71 7054 87
rect 6988 37 7004 71
rect 7038 37 7054 71
rect 6988 21 7054 37
rect -7054 -37 -6988 -21
rect -7054 -71 -7038 -37
rect -7004 -71 -6988 -37
rect -7054 -87 -6988 -71
rect -6936 -37 -6870 -21
rect -6936 -71 -6920 -37
rect -6886 -71 -6870 -37
rect -6936 -87 -6870 -71
rect -6818 -37 -6752 -21
rect -6818 -71 -6802 -37
rect -6768 -71 -6752 -37
rect -6818 -87 -6752 -71
rect -6700 -37 -6634 -21
rect -6700 -71 -6684 -37
rect -6650 -71 -6634 -37
rect -6700 -87 -6634 -71
rect -6582 -37 -6516 -21
rect -6582 -71 -6566 -37
rect -6532 -71 -6516 -37
rect -6582 -87 -6516 -71
rect -6464 -37 -6398 -21
rect -6464 -71 -6448 -37
rect -6414 -71 -6398 -37
rect -6464 -87 -6398 -71
rect -6346 -37 -6280 -21
rect -6346 -71 -6330 -37
rect -6296 -71 -6280 -37
rect -6346 -87 -6280 -71
rect -6228 -37 -6162 -21
rect -6228 -71 -6212 -37
rect -6178 -71 -6162 -37
rect -6228 -87 -6162 -71
rect -6110 -37 -6044 -21
rect -6110 -71 -6094 -37
rect -6060 -71 -6044 -37
rect -6110 -87 -6044 -71
rect -5992 -37 -5926 -21
rect -5992 -71 -5976 -37
rect -5942 -71 -5926 -37
rect -5992 -87 -5926 -71
rect -5874 -37 -5808 -21
rect -5874 -71 -5858 -37
rect -5824 -71 -5808 -37
rect -5874 -87 -5808 -71
rect -5756 -37 -5690 -21
rect -5756 -71 -5740 -37
rect -5706 -71 -5690 -37
rect -5756 -87 -5690 -71
rect -5638 -37 -5572 -21
rect -5638 -71 -5622 -37
rect -5588 -71 -5572 -37
rect -5638 -87 -5572 -71
rect -5520 -37 -5454 -21
rect -5520 -71 -5504 -37
rect -5470 -71 -5454 -37
rect -5520 -87 -5454 -71
rect -5402 -37 -5336 -21
rect -5402 -71 -5386 -37
rect -5352 -71 -5336 -37
rect -5402 -87 -5336 -71
rect -5284 -37 -5218 -21
rect -5284 -71 -5268 -37
rect -5234 -71 -5218 -37
rect -5284 -87 -5218 -71
rect -5166 -37 -5100 -21
rect -5166 -71 -5150 -37
rect -5116 -71 -5100 -37
rect -5166 -87 -5100 -71
rect -5048 -37 -4982 -21
rect -5048 -71 -5032 -37
rect -4998 -71 -4982 -37
rect -5048 -87 -4982 -71
rect -4930 -37 -4864 -21
rect -4930 -71 -4914 -37
rect -4880 -71 -4864 -37
rect -4930 -87 -4864 -71
rect -4812 -37 -4746 -21
rect -4812 -71 -4796 -37
rect -4762 -71 -4746 -37
rect -4812 -87 -4746 -71
rect -4694 -37 -4628 -21
rect -4694 -71 -4678 -37
rect -4644 -71 -4628 -37
rect -4694 -87 -4628 -71
rect -4576 -37 -4510 -21
rect -4576 -71 -4560 -37
rect -4526 -71 -4510 -37
rect -4576 -87 -4510 -71
rect -4458 -37 -4392 -21
rect -4458 -71 -4442 -37
rect -4408 -71 -4392 -37
rect -4458 -87 -4392 -71
rect -4340 -37 -4274 -21
rect -4340 -71 -4324 -37
rect -4290 -71 -4274 -37
rect -4340 -87 -4274 -71
rect -4222 -37 -4156 -21
rect -4222 -71 -4206 -37
rect -4172 -71 -4156 -37
rect -4222 -87 -4156 -71
rect -4104 -37 -4038 -21
rect -4104 -71 -4088 -37
rect -4054 -71 -4038 -37
rect -4104 -87 -4038 -71
rect -3986 -37 -3920 -21
rect -3986 -71 -3970 -37
rect -3936 -71 -3920 -37
rect -3986 -87 -3920 -71
rect -3868 -37 -3802 -21
rect -3868 -71 -3852 -37
rect -3818 -71 -3802 -37
rect -3868 -87 -3802 -71
rect -3750 -37 -3684 -21
rect -3750 -71 -3734 -37
rect -3700 -71 -3684 -37
rect -3750 -87 -3684 -71
rect -3632 -37 -3566 -21
rect -3632 -71 -3616 -37
rect -3582 -71 -3566 -37
rect -3632 -87 -3566 -71
rect -3514 -37 -3448 -21
rect -3514 -71 -3498 -37
rect -3464 -71 -3448 -37
rect -3514 -87 -3448 -71
rect -3396 -37 -3330 -21
rect -3396 -71 -3380 -37
rect -3346 -71 -3330 -37
rect -3396 -87 -3330 -71
rect -3278 -37 -3212 -21
rect -3278 -71 -3262 -37
rect -3228 -71 -3212 -37
rect -3278 -87 -3212 -71
rect -3160 -37 -3094 -21
rect -3160 -71 -3144 -37
rect -3110 -71 -3094 -37
rect -3160 -87 -3094 -71
rect -3042 -37 -2976 -21
rect -3042 -71 -3026 -37
rect -2992 -71 -2976 -37
rect -3042 -87 -2976 -71
rect -2924 -37 -2858 -21
rect -2924 -71 -2908 -37
rect -2874 -71 -2858 -37
rect -2924 -87 -2858 -71
rect -2806 -37 -2740 -21
rect -2806 -71 -2790 -37
rect -2756 -71 -2740 -37
rect -2806 -87 -2740 -71
rect -2688 -37 -2622 -21
rect -2688 -71 -2672 -37
rect -2638 -71 -2622 -37
rect -2688 -87 -2622 -71
rect -2570 -37 -2504 -21
rect -2570 -71 -2554 -37
rect -2520 -71 -2504 -37
rect -2570 -87 -2504 -71
rect -2452 -37 -2386 -21
rect -2452 -71 -2436 -37
rect -2402 -71 -2386 -37
rect -2452 -87 -2386 -71
rect -2334 -37 -2268 -21
rect -2334 -71 -2318 -37
rect -2284 -71 -2268 -37
rect -2334 -87 -2268 -71
rect -2216 -37 -2150 -21
rect -2216 -71 -2200 -37
rect -2166 -71 -2150 -37
rect -2216 -87 -2150 -71
rect -2098 -37 -2032 -21
rect -2098 -71 -2082 -37
rect -2048 -71 -2032 -37
rect -2098 -87 -2032 -71
rect -1980 -37 -1914 -21
rect -1980 -71 -1964 -37
rect -1930 -71 -1914 -37
rect -1980 -87 -1914 -71
rect -1862 -37 -1796 -21
rect -1862 -71 -1846 -37
rect -1812 -71 -1796 -37
rect -1862 -87 -1796 -71
rect -1744 -37 -1678 -21
rect -1744 -71 -1728 -37
rect -1694 -71 -1678 -37
rect -1744 -87 -1678 -71
rect -1626 -37 -1560 -21
rect -1626 -71 -1610 -37
rect -1576 -71 -1560 -37
rect -1626 -87 -1560 -71
rect -1508 -37 -1442 -21
rect -1508 -71 -1492 -37
rect -1458 -71 -1442 -37
rect -1508 -87 -1442 -71
rect -1390 -37 -1324 -21
rect -1390 -71 -1374 -37
rect -1340 -71 -1324 -37
rect -1390 -87 -1324 -71
rect -1272 -37 -1206 -21
rect -1272 -71 -1256 -37
rect -1222 -71 -1206 -37
rect -1272 -87 -1206 -71
rect -1154 -37 -1088 -21
rect -1154 -71 -1138 -37
rect -1104 -71 -1088 -37
rect -1154 -87 -1088 -71
rect -1036 -37 -970 -21
rect -1036 -71 -1020 -37
rect -986 -71 -970 -37
rect -1036 -87 -970 -71
rect -918 -37 -852 -21
rect -918 -71 -902 -37
rect -868 -71 -852 -37
rect -918 -87 -852 -71
rect -800 -37 -734 -21
rect -800 -71 -784 -37
rect -750 -71 -734 -37
rect -800 -87 -734 -71
rect -682 -37 -616 -21
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -682 -87 -616 -71
rect -564 -37 -498 -21
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -564 -87 -498 -71
rect -446 -37 -380 -21
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -446 -87 -380 -71
rect -328 -37 -262 -21
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -328 -87 -262 -71
rect -210 -37 -144 -21
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -210 -87 -144 -71
rect -92 -37 -26 -21
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect -92 -87 -26 -71
rect 26 -37 92 -21
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 26 -87 92 -71
rect 144 -37 210 -21
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 144 -87 210 -71
rect 262 -37 328 -21
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 262 -87 328 -71
rect 380 -37 446 -21
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 380 -87 446 -71
rect 498 -37 564 -21
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 498 -87 564 -71
rect 616 -37 682 -21
rect 616 -71 632 -37
rect 666 -71 682 -37
rect 616 -87 682 -71
rect 734 -37 800 -21
rect 734 -71 750 -37
rect 784 -71 800 -37
rect 734 -87 800 -71
rect 852 -37 918 -21
rect 852 -71 868 -37
rect 902 -71 918 -37
rect 852 -87 918 -71
rect 970 -37 1036 -21
rect 970 -71 986 -37
rect 1020 -71 1036 -37
rect 970 -87 1036 -71
rect 1088 -37 1154 -21
rect 1088 -71 1104 -37
rect 1138 -71 1154 -37
rect 1088 -87 1154 -71
rect 1206 -37 1272 -21
rect 1206 -71 1222 -37
rect 1256 -71 1272 -37
rect 1206 -87 1272 -71
rect 1324 -37 1390 -21
rect 1324 -71 1340 -37
rect 1374 -71 1390 -37
rect 1324 -87 1390 -71
rect 1442 -37 1508 -21
rect 1442 -71 1458 -37
rect 1492 -71 1508 -37
rect 1442 -87 1508 -71
rect 1560 -37 1626 -21
rect 1560 -71 1576 -37
rect 1610 -71 1626 -37
rect 1560 -87 1626 -71
rect 1678 -37 1744 -21
rect 1678 -71 1694 -37
rect 1728 -71 1744 -37
rect 1678 -87 1744 -71
rect 1796 -37 1862 -21
rect 1796 -71 1812 -37
rect 1846 -71 1862 -37
rect 1796 -87 1862 -71
rect 1914 -37 1980 -21
rect 1914 -71 1930 -37
rect 1964 -71 1980 -37
rect 1914 -87 1980 -71
rect 2032 -37 2098 -21
rect 2032 -71 2048 -37
rect 2082 -71 2098 -37
rect 2032 -87 2098 -71
rect 2150 -37 2216 -21
rect 2150 -71 2166 -37
rect 2200 -71 2216 -37
rect 2150 -87 2216 -71
rect 2268 -37 2334 -21
rect 2268 -71 2284 -37
rect 2318 -71 2334 -37
rect 2268 -87 2334 -71
rect 2386 -37 2452 -21
rect 2386 -71 2402 -37
rect 2436 -71 2452 -37
rect 2386 -87 2452 -71
rect 2504 -37 2570 -21
rect 2504 -71 2520 -37
rect 2554 -71 2570 -37
rect 2504 -87 2570 -71
rect 2622 -37 2688 -21
rect 2622 -71 2638 -37
rect 2672 -71 2688 -37
rect 2622 -87 2688 -71
rect 2740 -37 2806 -21
rect 2740 -71 2756 -37
rect 2790 -71 2806 -37
rect 2740 -87 2806 -71
rect 2858 -37 2924 -21
rect 2858 -71 2874 -37
rect 2908 -71 2924 -37
rect 2858 -87 2924 -71
rect 2976 -37 3042 -21
rect 2976 -71 2992 -37
rect 3026 -71 3042 -37
rect 2976 -87 3042 -71
rect 3094 -37 3160 -21
rect 3094 -71 3110 -37
rect 3144 -71 3160 -37
rect 3094 -87 3160 -71
rect 3212 -37 3278 -21
rect 3212 -71 3228 -37
rect 3262 -71 3278 -37
rect 3212 -87 3278 -71
rect 3330 -37 3396 -21
rect 3330 -71 3346 -37
rect 3380 -71 3396 -37
rect 3330 -87 3396 -71
rect 3448 -37 3514 -21
rect 3448 -71 3464 -37
rect 3498 -71 3514 -37
rect 3448 -87 3514 -71
rect 3566 -37 3632 -21
rect 3566 -71 3582 -37
rect 3616 -71 3632 -37
rect 3566 -87 3632 -71
rect 3684 -37 3750 -21
rect 3684 -71 3700 -37
rect 3734 -71 3750 -37
rect 3684 -87 3750 -71
rect 3802 -37 3868 -21
rect 3802 -71 3818 -37
rect 3852 -71 3868 -37
rect 3802 -87 3868 -71
rect 3920 -37 3986 -21
rect 3920 -71 3936 -37
rect 3970 -71 3986 -37
rect 3920 -87 3986 -71
rect 4038 -37 4104 -21
rect 4038 -71 4054 -37
rect 4088 -71 4104 -37
rect 4038 -87 4104 -71
rect 4156 -37 4222 -21
rect 4156 -71 4172 -37
rect 4206 -71 4222 -37
rect 4156 -87 4222 -71
rect 4274 -37 4340 -21
rect 4274 -71 4290 -37
rect 4324 -71 4340 -37
rect 4274 -87 4340 -71
rect 4392 -37 4458 -21
rect 4392 -71 4408 -37
rect 4442 -71 4458 -37
rect 4392 -87 4458 -71
rect 4510 -37 4576 -21
rect 4510 -71 4526 -37
rect 4560 -71 4576 -37
rect 4510 -87 4576 -71
rect 4628 -37 4694 -21
rect 4628 -71 4644 -37
rect 4678 -71 4694 -37
rect 4628 -87 4694 -71
rect 4746 -37 4812 -21
rect 4746 -71 4762 -37
rect 4796 -71 4812 -37
rect 4746 -87 4812 -71
rect 4864 -37 4930 -21
rect 4864 -71 4880 -37
rect 4914 -71 4930 -37
rect 4864 -87 4930 -71
rect 4982 -37 5048 -21
rect 4982 -71 4998 -37
rect 5032 -71 5048 -37
rect 4982 -87 5048 -71
rect 5100 -37 5166 -21
rect 5100 -71 5116 -37
rect 5150 -71 5166 -37
rect 5100 -87 5166 -71
rect 5218 -37 5284 -21
rect 5218 -71 5234 -37
rect 5268 -71 5284 -37
rect 5218 -87 5284 -71
rect 5336 -37 5402 -21
rect 5336 -71 5352 -37
rect 5386 -71 5402 -37
rect 5336 -87 5402 -71
rect 5454 -37 5520 -21
rect 5454 -71 5470 -37
rect 5504 -71 5520 -37
rect 5454 -87 5520 -71
rect 5572 -37 5638 -21
rect 5572 -71 5588 -37
rect 5622 -71 5638 -37
rect 5572 -87 5638 -71
rect 5690 -37 5756 -21
rect 5690 -71 5706 -37
rect 5740 -71 5756 -37
rect 5690 -87 5756 -71
rect 5808 -37 5874 -21
rect 5808 -71 5824 -37
rect 5858 -71 5874 -37
rect 5808 -87 5874 -71
rect 5926 -37 5992 -21
rect 5926 -71 5942 -37
rect 5976 -71 5992 -37
rect 5926 -87 5992 -71
rect 6044 -37 6110 -21
rect 6044 -71 6060 -37
rect 6094 -71 6110 -37
rect 6044 -87 6110 -71
rect 6162 -37 6228 -21
rect 6162 -71 6178 -37
rect 6212 -71 6228 -37
rect 6162 -87 6228 -71
rect 6280 -37 6346 -21
rect 6280 -71 6296 -37
rect 6330 -71 6346 -37
rect 6280 -87 6346 -71
rect 6398 -37 6464 -21
rect 6398 -71 6414 -37
rect 6448 -71 6464 -37
rect 6398 -87 6464 -71
rect 6516 -37 6582 -21
rect 6516 -71 6532 -37
rect 6566 -71 6582 -37
rect 6516 -87 6582 -71
rect 6634 -37 6700 -21
rect 6634 -71 6650 -37
rect 6684 -71 6700 -37
rect 6634 -87 6700 -71
rect 6752 -37 6818 -21
rect 6752 -71 6768 -37
rect 6802 -71 6818 -37
rect 6752 -87 6818 -71
rect 6870 -37 6936 -21
rect 6870 -71 6886 -37
rect 6920 -71 6936 -37
rect 6870 -87 6936 -71
rect 6988 -37 7054 -21
rect 6988 -71 7004 -37
rect 7038 -71 7054 -37
rect 6988 -87 7054 -71
rect -7051 -118 -6991 -87
rect -6933 -118 -6873 -87
rect -6815 -118 -6755 -87
rect -6697 -118 -6637 -87
rect -6579 -118 -6519 -87
rect -6461 -118 -6401 -87
rect -6343 -118 -6283 -87
rect -6225 -118 -6165 -87
rect -6107 -118 -6047 -87
rect -5989 -118 -5929 -87
rect -5871 -118 -5811 -87
rect -5753 -118 -5693 -87
rect -5635 -118 -5575 -87
rect -5517 -118 -5457 -87
rect -5399 -118 -5339 -87
rect -5281 -118 -5221 -87
rect -5163 -118 -5103 -87
rect -5045 -118 -4985 -87
rect -4927 -118 -4867 -87
rect -4809 -118 -4749 -87
rect -4691 -118 -4631 -87
rect -4573 -118 -4513 -87
rect -4455 -118 -4395 -87
rect -4337 -118 -4277 -87
rect -4219 -118 -4159 -87
rect -4101 -118 -4041 -87
rect -3983 -118 -3923 -87
rect -3865 -118 -3805 -87
rect -3747 -118 -3687 -87
rect -3629 -118 -3569 -87
rect -3511 -118 -3451 -87
rect -3393 -118 -3333 -87
rect -3275 -118 -3215 -87
rect -3157 -118 -3097 -87
rect -3039 -118 -2979 -87
rect -2921 -118 -2861 -87
rect -2803 -118 -2743 -87
rect -2685 -118 -2625 -87
rect -2567 -118 -2507 -87
rect -2449 -118 -2389 -87
rect -2331 -118 -2271 -87
rect -2213 -118 -2153 -87
rect -2095 -118 -2035 -87
rect -1977 -118 -1917 -87
rect -1859 -118 -1799 -87
rect -1741 -118 -1681 -87
rect -1623 -118 -1563 -87
rect -1505 -118 -1445 -87
rect -1387 -118 -1327 -87
rect -1269 -118 -1209 -87
rect -1151 -118 -1091 -87
rect -1033 -118 -973 -87
rect -915 -118 -855 -87
rect -797 -118 -737 -87
rect -679 -118 -619 -87
rect -561 -118 -501 -87
rect -443 -118 -383 -87
rect -325 -118 -265 -87
rect -207 -118 -147 -87
rect -89 -118 -29 -87
rect 29 -118 89 -87
rect 147 -118 207 -87
rect 265 -118 325 -87
rect 383 -118 443 -87
rect 501 -118 561 -87
rect 619 -118 679 -87
rect 737 -118 797 -87
rect 855 -118 915 -87
rect 973 -118 1033 -87
rect 1091 -118 1151 -87
rect 1209 -118 1269 -87
rect 1327 -118 1387 -87
rect 1445 -118 1505 -87
rect 1563 -118 1623 -87
rect 1681 -118 1741 -87
rect 1799 -118 1859 -87
rect 1917 -118 1977 -87
rect 2035 -118 2095 -87
rect 2153 -118 2213 -87
rect 2271 -118 2331 -87
rect 2389 -118 2449 -87
rect 2507 -118 2567 -87
rect 2625 -118 2685 -87
rect 2743 -118 2803 -87
rect 2861 -118 2921 -87
rect 2979 -118 3039 -87
rect 3097 -118 3157 -87
rect 3215 -118 3275 -87
rect 3333 -118 3393 -87
rect 3451 -118 3511 -87
rect 3569 -118 3629 -87
rect 3687 -118 3747 -87
rect 3805 -118 3865 -87
rect 3923 -118 3983 -87
rect 4041 -118 4101 -87
rect 4159 -118 4219 -87
rect 4277 -118 4337 -87
rect 4395 -118 4455 -87
rect 4513 -118 4573 -87
rect 4631 -118 4691 -87
rect 4749 -118 4809 -87
rect 4867 -118 4927 -87
rect 4985 -118 5045 -87
rect 5103 -118 5163 -87
rect 5221 -118 5281 -87
rect 5339 -118 5399 -87
rect 5457 -118 5517 -87
rect 5575 -118 5635 -87
rect 5693 -118 5753 -87
rect 5811 -118 5871 -87
rect 5929 -118 5989 -87
rect 6047 -118 6107 -87
rect 6165 -118 6225 -87
rect 6283 -118 6343 -87
rect 6401 -118 6461 -87
rect 6519 -118 6579 -87
rect 6637 -118 6697 -87
rect 6755 -118 6815 -87
rect 6873 -118 6933 -87
rect 6991 -118 7051 -87
rect -7051 -749 -6991 -718
rect -6933 -749 -6873 -718
rect -6815 -749 -6755 -718
rect -6697 -749 -6637 -718
rect -6579 -749 -6519 -718
rect -6461 -749 -6401 -718
rect -6343 -749 -6283 -718
rect -6225 -749 -6165 -718
rect -6107 -749 -6047 -718
rect -5989 -749 -5929 -718
rect -5871 -749 -5811 -718
rect -5753 -749 -5693 -718
rect -5635 -749 -5575 -718
rect -5517 -749 -5457 -718
rect -5399 -749 -5339 -718
rect -5281 -749 -5221 -718
rect -5163 -749 -5103 -718
rect -5045 -749 -4985 -718
rect -4927 -749 -4867 -718
rect -4809 -749 -4749 -718
rect -4691 -749 -4631 -718
rect -4573 -749 -4513 -718
rect -4455 -749 -4395 -718
rect -4337 -749 -4277 -718
rect -4219 -749 -4159 -718
rect -4101 -749 -4041 -718
rect -3983 -749 -3923 -718
rect -3865 -749 -3805 -718
rect -3747 -749 -3687 -718
rect -3629 -749 -3569 -718
rect -3511 -749 -3451 -718
rect -3393 -749 -3333 -718
rect -3275 -749 -3215 -718
rect -3157 -749 -3097 -718
rect -3039 -749 -2979 -718
rect -2921 -749 -2861 -718
rect -2803 -749 -2743 -718
rect -2685 -749 -2625 -718
rect -2567 -749 -2507 -718
rect -2449 -749 -2389 -718
rect -2331 -749 -2271 -718
rect -2213 -749 -2153 -718
rect -2095 -749 -2035 -718
rect -1977 -749 -1917 -718
rect -1859 -749 -1799 -718
rect -1741 -749 -1681 -718
rect -1623 -749 -1563 -718
rect -1505 -749 -1445 -718
rect -1387 -749 -1327 -718
rect -1269 -749 -1209 -718
rect -1151 -749 -1091 -718
rect -1033 -749 -973 -718
rect -915 -749 -855 -718
rect -797 -749 -737 -718
rect -679 -749 -619 -718
rect -561 -749 -501 -718
rect -443 -749 -383 -718
rect -325 -749 -265 -718
rect -207 -749 -147 -718
rect -89 -749 -29 -718
rect 29 -749 89 -718
rect 147 -749 207 -718
rect 265 -749 325 -718
rect 383 -749 443 -718
rect 501 -749 561 -718
rect 619 -749 679 -718
rect 737 -749 797 -718
rect 855 -749 915 -718
rect 973 -749 1033 -718
rect 1091 -749 1151 -718
rect 1209 -749 1269 -718
rect 1327 -749 1387 -718
rect 1445 -749 1505 -718
rect 1563 -749 1623 -718
rect 1681 -749 1741 -718
rect 1799 -749 1859 -718
rect 1917 -749 1977 -718
rect 2035 -749 2095 -718
rect 2153 -749 2213 -718
rect 2271 -749 2331 -718
rect 2389 -749 2449 -718
rect 2507 -749 2567 -718
rect 2625 -749 2685 -718
rect 2743 -749 2803 -718
rect 2861 -749 2921 -718
rect 2979 -749 3039 -718
rect 3097 -749 3157 -718
rect 3215 -749 3275 -718
rect 3333 -749 3393 -718
rect 3451 -749 3511 -718
rect 3569 -749 3629 -718
rect 3687 -749 3747 -718
rect 3805 -749 3865 -718
rect 3923 -749 3983 -718
rect 4041 -749 4101 -718
rect 4159 -749 4219 -718
rect 4277 -749 4337 -718
rect 4395 -749 4455 -718
rect 4513 -749 4573 -718
rect 4631 -749 4691 -718
rect 4749 -749 4809 -718
rect 4867 -749 4927 -718
rect 4985 -749 5045 -718
rect 5103 -749 5163 -718
rect 5221 -749 5281 -718
rect 5339 -749 5399 -718
rect 5457 -749 5517 -718
rect 5575 -749 5635 -718
rect 5693 -749 5753 -718
rect 5811 -749 5871 -718
rect 5929 -749 5989 -718
rect 6047 -749 6107 -718
rect 6165 -749 6225 -718
rect 6283 -749 6343 -718
rect 6401 -749 6461 -718
rect 6519 -749 6579 -718
rect 6637 -749 6697 -718
rect 6755 -749 6815 -718
rect 6873 -749 6933 -718
rect 6991 -749 7051 -718
rect -7054 -765 -6988 -749
rect -7054 -799 -7038 -765
rect -7004 -799 -6988 -765
rect -7054 -815 -6988 -799
rect -6936 -765 -6870 -749
rect -6936 -799 -6920 -765
rect -6886 -799 -6870 -765
rect -6936 -815 -6870 -799
rect -6818 -765 -6752 -749
rect -6818 -799 -6802 -765
rect -6768 -799 -6752 -765
rect -6818 -815 -6752 -799
rect -6700 -765 -6634 -749
rect -6700 -799 -6684 -765
rect -6650 -799 -6634 -765
rect -6700 -815 -6634 -799
rect -6582 -765 -6516 -749
rect -6582 -799 -6566 -765
rect -6532 -799 -6516 -765
rect -6582 -815 -6516 -799
rect -6464 -765 -6398 -749
rect -6464 -799 -6448 -765
rect -6414 -799 -6398 -765
rect -6464 -815 -6398 -799
rect -6346 -765 -6280 -749
rect -6346 -799 -6330 -765
rect -6296 -799 -6280 -765
rect -6346 -815 -6280 -799
rect -6228 -765 -6162 -749
rect -6228 -799 -6212 -765
rect -6178 -799 -6162 -765
rect -6228 -815 -6162 -799
rect -6110 -765 -6044 -749
rect -6110 -799 -6094 -765
rect -6060 -799 -6044 -765
rect -6110 -815 -6044 -799
rect -5992 -765 -5926 -749
rect -5992 -799 -5976 -765
rect -5942 -799 -5926 -765
rect -5992 -815 -5926 -799
rect -5874 -765 -5808 -749
rect -5874 -799 -5858 -765
rect -5824 -799 -5808 -765
rect -5874 -815 -5808 -799
rect -5756 -765 -5690 -749
rect -5756 -799 -5740 -765
rect -5706 -799 -5690 -765
rect -5756 -815 -5690 -799
rect -5638 -765 -5572 -749
rect -5638 -799 -5622 -765
rect -5588 -799 -5572 -765
rect -5638 -815 -5572 -799
rect -5520 -765 -5454 -749
rect -5520 -799 -5504 -765
rect -5470 -799 -5454 -765
rect -5520 -815 -5454 -799
rect -5402 -765 -5336 -749
rect -5402 -799 -5386 -765
rect -5352 -799 -5336 -765
rect -5402 -815 -5336 -799
rect -5284 -765 -5218 -749
rect -5284 -799 -5268 -765
rect -5234 -799 -5218 -765
rect -5284 -815 -5218 -799
rect -5166 -765 -5100 -749
rect -5166 -799 -5150 -765
rect -5116 -799 -5100 -765
rect -5166 -815 -5100 -799
rect -5048 -765 -4982 -749
rect -5048 -799 -5032 -765
rect -4998 -799 -4982 -765
rect -5048 -815 -4982 -799
rect -4930 -765 -4864 -749
rect -4930 -799 -4914 -765
rect -4880 -799 -4864 -765
rect -4930 -815 -4864 -799
rect -4812 -765 -4746 -749
rect -4812 -799 -4796 -765
rect -4762 -799 -4746 -765
rect -4812 -815 -4746 -799
rect -4694 -765 -4628 -749
rect -4694 -799 -4678 -765
rect -4644 -799 -4628 -765
rect -4694 -815 -4628 -799
rect -4576 -765 -4510 -749
rect -4576 -799 -4560 -765
rect -4526 -799 -4510 -765
rect -4576 -815 -4510 -799
rect -4458 -765 -4392 -749
rect -4458 -799 -4442 -765
rect -4408 -799 -4392 -765
rect -4458 -815 -4392 -799
rect -4340 -765 -4274 -749
rect -4340 -799 -4324 -765
rect -4290 -799 -4274 -765
rect -4340 -815 -4274 -799
rect -4222 -765 -4156 -749
rect -4222 -799 -4206 -765
rect -4172 -799 -4156 -765
rect -4222 -815 -4156 -799
rect -4104 -765 -4038 -749
rect -4104 -799 -4088 -765
rect -4054 -799 -4038 -765
rect -4104 -815 -4038 -799
rect -3986 -765 -3920 -749
rect -3986 -799 -3970 -765
rect -3936 -799 -3920 -765
rect -3986 -815 -3920 -799
rect -3868 -765 -3802 -749
rect -3868 -799 -3852 -765
rect -3818 -799 -3802 -765
rect -3868 -815 -3802 -799
rect -3750 -765 -3684 -749
rect -3750 -799 -3734 -765
rect -3700 -799 -3684 -765
rect -3750 -815 -3684 -799
rect -3632 -765 -3566 -749
rect -3632 -799 -3616 -765
rect -3582 -799 -3566 -765
rect -3632 -815 -3566 -799
rect -3514 -765 -3448 -749
rect -3514 -799 -3498 -765
rect -3464 -799 -3448 -765
rect -3514 -815 -3448 -799
rect -3396 -765 -3330 -749
rect -3396 -799 -3380 -765
rect -3346 -799 -3330 -765
rect -3396 -815 -3330 -799
rect -3278 -765 -3212 -749
rect -3278 -799 -3262 -765
rect -3228 -799 -3212 -765
rect -3278 -815 -3212 -799
rect -3160 -765 -3094 -749
rect -3160 -799 -3144 -765
rect -3110 -799 -3094 -765
rect -3160 -815 -3094 -799
rect -3042 -765 -2976 -749
rect -3042 -799 -3026 -765
rect -2992 -799 -2976 -765
rect -3042 -815 -2976 -799
rect -2924 -765 -2858 -749
rect -2924 -799 -2908 -765
rect -2874 -799 -2858 -765
rect -2924 -815 -2858 -799
rect -2806 -765 -2740 -749
rect -2806 -799 -2790 -765
rect -2756 -799 -2740 -765
rect -2806 -815 -2740 -799
rect -2688 -765 -2622 -749
rect -2688 -799 -2672 -765
rect -2638 -799 -2622 -765
rect -2688 -815 -2622 -799
rect -2570 -765 -2504 -749
rect -2570 -799 -2554 -765
rect -2520 -799 -2504 -765
rect -2570 -815 -2504 -799
rect -2452 -765 -2386 -749
rect -2452 -799 -2436 -765
rect -2402 -799 -2386 -765
rect -2452 -815 -2386 -799
rect -2334 -765 -2268 -749
rect -2334 -799 -2318 -765
rect -2284 -799 -2268 -765
rect -2334 -815 -2268 -799
rect -2216 -765 -2150 -749
rect -2216 -799 -2200 -765
rect -2166 -799 -2150 -765
rect -2216 -815 -2150 -799
rect -2098 -765 -2032 -749
rect -2098 -799 -2082 -765
rect -2048 -799 -2032 -765
rect -2098 -815 -2032 -799
rect -1980 -765 -1914 -749
rect -1980 -799 -1964 -765
rect -1930 -799 -1914 -765
rect -1980 -815 -1914 -799
rect -1862 -765 -1796 -749
rect -1862 -799 -1846 -765
rect -1812 -799 -1796 -765
rect -1862 -815 -1796 -799
rect -1744 -765 -1678 -749
rect -1744 -799 -1728 -765
rect -1694 -799 -1678 -765
rect -1744 -815 -1678 -799
rect -1626 -765 -1560 -749
rect -1626 -799 -1610 -765
rect -1576 -799 -1560 -765
rect -1626 -815 -1560 -799
rect -1508 -765 -1442 -749
rect -1508 -799 -1492 -765
rect -1458 -799 -1442 -765
rect -1508 -815 -1442 -799
rect -1390 -765 -1324 -749
rect -1390 -799 -1374 -765
rect -1340 -799 -1324 -765
rect -1390 -815 -1324 -799
rect -1272 -765 -1206 -749
rect -1272 -799 -1256 -765
rect -1222 -799 -1206 -765
rect -1272 -815 -1206 -799
rect -1154 -765 -1088 -749
rect -1154 -799 -1138 -765
rect -1104 -799 -1088 -765
rect -1154 -815 -1088 -799
rect -1036 -765 -970 -749
rect -1036 -799 -1020 -765
rect -986 -799 -970 -765
rect -1036 -815 -970 -799
rect -918 -765 -852 -749
rect -918 -799 -902 -765
rect -868 -799 -852 -765
rect -918 -815 -852 -799
rect -800 -765 -734 -749
rect -800 -799 -784 -765
rect -750 -799 -734 -765
rect -800 -815 -734 -799
rect -682 -765 -616 -749
rect -682 -799 -666 -765
rect -632 -799 -616 -765
rect -682 -815 -616 -799
rect -564 -765 -498 -749
rect -564 -799 -548 -765
rect -514 -799 -498 -765
rect -564 -815 -498 -799
rect -446 -765 -380 -749
rect -446 -799 -430 -765
rect -396 -799 -380 -765
rect -446 -815 -380 -799
rect -328 -765 -262 -749
rect -328 -799 -312 -765
rect -278 -799 -262 -765
rect -328 -815 -262 -799
rect -210 -765 -144 -749
rect -210 -799 -194 -765
rect -160 -799 -144 -765
rect -210 -815 -144 -799
rect -92 -765 -26 -749
rect -92 -799 -76 -765
rect -42 -799 -26 -765
rect -92 -815 -26 -799
rect 26 -765 92 -749
rect 26 -799 42 -765
rect 76 -799 92 -765
rect 26 -815 92 -799
rect 144 -765 210 -749
rect 144 -799 160 -765
rect 194 -799 210 -765
rect 144 -815 210 -799
rect 262 -765 328 -749
rect 262 -799 278 -765
rect 312 -799 328 -765
rect 262 -815 328 -799
rect 380 -765 446 -749
rect 380 -799 396 -765
rect 430 -799 446 -765
rect 380 -815 446 -799
rect 498 -765 564 -749
rect 498 -799 514 -765
rect 548 -799 564 -765
rect 498 -815 564 -799
rect 616 -765 682 -749
rect 616 -799 632 -765
rect 666 -799 682 -765
rect 616 -815 682 -799
rect 734 -765 800 -749
rect 734 -799 750 -765
rect 784 -799 800 -765
rect 734 -815 800 -799
rect 852 -765 918 -749
rect 852 -799 868 -765
rect 902 -799 918 -765
rect 852 -815 918 -799
rect 970 -765 1036 -749
rect 970 -799 986 -765
rect 1020 -799 1036 -765
rect 970 -815 1036 -799
rect 1088 -765 1154 -749
rect 1088 -799 1104 -765
rect 1138 -799 1154 -765
rect 1088 -815 1154 -799
rect 1206 -765 1272 -749
rect 1206 -799 1222 -765
rect 1256 -799 1272 -765
rect 1206 -815 1272 -799
rect 1324 -765 1390 -749
rect 1324 -799 1340 -765
rect 1374 -799 1390 -765
rect 1324 -815 1390 -799
rect 1442 -765 1508 -749
rect 1442 -799 1458 -765
rect 1492 -799 1508 -765
rect 1442 -815 1508 -799
rect 1560 -765 1626 -749
rect 1560 -799 1576 -765
rect 1610 -799 1626 -765
rect 1560 -815 1626 -799
rect 1678 -765 1744 -749
rect 1678 -799 1694 -765
rect 1728 -799 1744 -765
rect 1678 -815 1744 -799
rect 1796 -765 1862 -749
rect 1796 -799 1812 -765
rect 1846 -799 1862 -765
rect 1796 -815 1862 -799
rect 1914 -765 1980 -749
rect 1914 -799 1930 -765
rect 1964 -799 1980 -765
rect 1914 -815 1980 -799
rect 2032 -765 2098 -749
rect 2032 -799 2048 -765
rect 2082 -799 2098 -765
rect 2032 -815 2098 -799
rect 2150 -765 2216 -749
rect 2150 -799 2166 -765
rect 2200 -799 2216 -765
rect 2150 -815 2216 -799
rect 2268 -765 2334 -749
rect 2268 -799 2284 -765
rect 2318 -799 2334 -765
rect 2268 -815 2334 -799
rect 2386 -765 2452 -749
rect 2386 -799 2402 -765
rect 2436 -799 2452 -765
rect 2386 -815 2452 -799
rect 2504 -765 2570 -749
rect 2504 -799 2520 -765
rect 2554 -799 2570 -765
rect 2504 -815 2570 -799
rect 2622 -765 2688 -749
rect 2622 -799 2638 -765
rect 2672 -799 2688 -765
rect 2622 -815 2688 -799
rect 2740 -765 2806 -749
rect 2740 -799 2756 -765
rect 2790 -799 2806 -765
rect 2740 -815 2806 -799
rect 2858 -765 2924 -749
rect 2858 -799 2874 -765
rect 2908 -799 2924 -765
rect 2858 -815 2924 -799
rect 2976 -765 3042 -749
rect 2976 -799 2992 -765
rect 3026 -799 3042 -765
rect 2976 -815 3042 -799
rect 3094 -765 3160 -749
rect 3094 -799 3110 -765
rect 3144 -799 3160 -765
rect 3094 -815 3160 -799
rect 3212 -765 3278 -749
rect 3212 -799 3228 -765
rect 3262 -799 3278 -765
rect 3212 -815 3278 -799
rect 3330 -765 3396 -749
rect 3330 -799 3346 -765
rect 3380 -799 3396 -765
rect 3330 -815 3396 -799
rect 3448 -765 3514 -749
rect 3448 -799 3464 -765
rect 3498 -799 3514 -765
rect 3448 -815 3514 -799
rect 3566 -765 3632 -749
rect 3566 -799 3582 -765
rect 3616 -799 3632 -765
rect 3566 -815 3632 -799
rect 3684 -765 3750 -749
rect 3684 -799 3700 -765
rect 3734 -799 3750 -765
rect 3684 -815 3750 -799
rect 3802 -765 3868 -749
rect 3802 -799 3818 -765
rect 3852 -799 3868 -765
rect 3802 -815 3868 -799
rect 3920 -765 3986 -749
rect 3920 -799 3936 -765
rect 3970 -799 3986 -765
rect 3920 -815 3986 -799
rect 4038 -765 4104 -749
rect 4038 -799 4054 -765
rect 4088 -799 4104 -765
rect 4038 -815 4104 -799
rect 4156 -765 4222 -749
rect 4156 -799 4172 -765
rect 4206 -799 4222 -765
rect 4156 -815 4222 -799
rect 4274 -765 4340 -749
rect 4274 -799 4290 -765
rect 4324 -799 4340 -765
rect 4274 -815 4340 -799
rect 4392 -765 4458 -749
rect 4392 -799 4408 -765
rect 4442 -799 4458 -765
rect 4392 -815 4458 -799
rect 4510 -765 4576 -749
rect 4510 -799 4526 -765
rect 4560 -799 4576 -765
rect 4510 -815 4576 -799
rect 4628 -765 4694 -749
rect 4628 -799 4644 -765
rect 4678 -799 4694 -765
rect 4628 -815 4694 -799
rect 4746 -765 4812 -749
rect 4746 -799 4762 -765
rect 4796 -799 4812 -765
rect 4746 -815 4812 -799
rect 4864 -765 4930 -749
rect 4864 -799 4880 -765
rect 4914 -799 4930 -765
rect 4864 -815 4930 -799
rect 4982 -765 5048 -749
rect 4982 -799 4998 -765
rect 5032 -799 5048 -765
rect 4982 -815 5048 -799
rect 5100 -765 5166 -749
rect 5100 -799 5116 -765
rect 5150 -799 5166 -765
rect 5100 -815 5166 -799
rect 5218 -765 5284 -749
rect 5218 -799 5234 -765
rect 5268 -799 5284 -765
rect 5218 -815 5284 -799
rect 5336 -765 5402 -749
rect 5336 -799 5352 -765
rect 5386 -799 5402 -765
rect 5336 -815 5402 -799
rect 5454 -765 5520 -749
rect 5454 -799 5470 -765
rect 5504 -799 5520 -765
rect 5454 -815 5520 -799
rect 5572 -765 5638 -749
rect 5572 -799 5588 -765
rect 5622 -799 5638 -765
rect 5572 -815 5638 -799
rect 5690 -765 5756 -749
rect 5690 -799 5706 -765
rect 5740 -799 5756 -765
rect 5690 -815 5756 -799
rect 5808 -765 5874 -749
rect 5808 -799 5824 -765
rect 5858 -799 5874 -765
rect 5808 -815 5874 -799
rect 5926 -765 5992 -749
rect 5926 -799 5942 -765
rect 5976 -799 5992 -765
rect 5926 -815 5992 -799
rect 6044 -765 6110 -749
rect 6044 -799 6060 -765
rect 6094 -799 6110 -765
rect 6044 -815 6110 -799
rect 6162 -765 6228 -749
rect 6162 -799 6178 -765
rect 6212 -799 6228 -765
rect 6162 -815 6228 -799
rect 6280 -765 6346 -749
rect 6280 -799 6296 -765
rect 6330 -799 6346 -765
rect 6280 -815 6346 -799
rect 6398 -765 6464 -749
rect 6398 -799 6414 -765
rect 6448 -799 6464 -765
rect 6398 -815 6464 -799
rect 6516 -765 6582 -749
rect 6516 -799 6532 -765
rect 6566 -799 6582 -765
rect 6516 -815 6582 -799
rect 6634 -765 6700 -749
rect 6634 -799 6650 -765
rect 6684 -799 6700 -765
rect 6634 -815 6700 -799
rect 6752 -765 6818 -749
rect 6752 -799 6768 -765
rect 6802 -799 6818 -765
rect 6752 -815 6818 -799
rect 6870 -765 6936 -749
rect 6870 -799 6886 -765
rect 6920 -799 6936 -765
rect 6870 -815 6936 -799
rect 6988 -765 7054 -749
rect 6988 -799 7004 -765
rect 7038 -799 7054 -765
rect 6988 -815 7054 -799
<< polycont >>
rect -7038 765 -7004 799
rect -6920 765 -6886 799
rect -6802 765 -6768 799
rect -6684 765 -6650 799
rect -6566 765 -6532 799
rect -6448 765 -6414 799
rect -6330 765 -6296 799
rect -6212 765 -6178 799
rect -6094 765 -6060 799
rect -5976 765 -5942 799
rect -5858 765 -5824 799
rect -5740 765 -5706 799
rect -5622 765 -5588 799
rect -5504 765 -5470 799
rect -5386 765 -5352 799
rect -5268 765 -5234 799
rect -5150 765 -5116 799
rect -5032 765 -4998 799
rect -4914 765 -4880 799
rect -4796 765 -4762 799
rect -4678 765 -4644 799
rect -4560 765 -4526 799
rect -4442 765 -4408 799
rect -4324 765 -4290 799
rect -4206 765 -4172 799
rect -4088 765 -4054 799
rect -3970 765 -3936 799
rect -3852 765 -3818 799
rect -3734 765 -3700 799
rect -3616 765 -3582 799
rect -3498 765 -3464 799
rect -3380 765 -3346 799
rect -3262 765 -3228 799
rect -3144 765 -3110 799
rect -3026 765 -2992 799
rect -2908 765 -2874 799
rect -2790 765 -2756 799
rect -2672 765 -2638 799
rect -2554 765 -2520 799
rect -2436 765 -2402 799
rect -2318 765 -2284 799
rect -2200 765 -2166 799
rect -2082 765 -2048 799
rect -1964 765 -1930 799
rect -1846 765 -1812 799
rect -1728 765 -1694 799
rect -1610 765 -1576 799
rect -1492 765 -1458 799
rect -1374 765 -1340 799
rect -1256 765 -1222 799
rect -1138 765 -1104 799
rect -1020 765 -986 799
rect -902 765 -868 799
rect -784 765 -750 799
rect -666 765 -632 799
rect -548 765 -514 799
rect -430 765 -396 799
rect -312 765 -278 799
rect -194 765 -160 799
rect -76 765 -42 799
rect 42 765 76 799
rect 160 765 194 799
rect 278 765 312 799
rect 396 765 430 799
rect 514 765 548 799
rect 632 765 666 799
rect 750 765 784 799
rect 868 765 902 799
rect 986 765 1020 799
rect 1104 765 1138 799
rect 1222 765 1256 799
rect 1340 765 1374 799
rect 1458 765 1492 799
rect 1576 765 1610 799
rect 1694 765 1728 799
rect 1812 765 1846 799
rect 1930 765 1964 799
rect 2048 765 2082 799
rect 2166 765 2200 799
rect 2284 765 2318 799
rect 2402 765 2436 799
rect 2520 765 2554 799
rect 2638 765 2672 799
rect 2756 765 2790 799
rect 2874 765 2908 799
rect 2992 765 3026 799
rect 3110 765 3144 799
rect 3228 765 3262 799
rect 3346 765 3380 799
rect 3464 765 3498 799
rect 3582 765 3616 799
rect 3700 765 3734 799
rect 3818 765 3852 799
rect 3936 765 3970 799
rect 4054 765 4088 799
rect 4172 765 4206 799
rect 4290 765 4324 799
rect 4408 765 4442 799
rect 4526 765 4560 799
rect 4644 765 4678 799
rect 4762 765 4796 799
rect 4880 765 4914 799
rect 4998 765 5032 799
rect 5116 765 5150 799
rect 5234 765 5268 799
rect 5352 765 5386 799
rect 5470 765 5504 799
rect 5588 765 5622 799
rect 5706 765 5740 799
rect 5824 765 5858 799
rect 5942 765 5976 799
rect 6060 765 6094 799
rect 6178 765 6212 799
rect 6296 765 6330 799
rect 6414 765 6448 799
rect 6532 765 6566 799
rect 6650 765 6684 799
rect 6768 765 6802 799
rect 6886 765 6920 799
rect 7004 765 7038 799
rect -7038 37 -7004 71
rect -6920 37 -6886 71
rect -6802 37 -6768 71
rect -6684 37 -6650 71
rect -6566 37 -6532 71
rect -6448 37 -6414 71
rect -6330 37 -6296 71
rect -6212 37 -6178 71
rect -6094 37 -6060 71
rect -5976 37 -5942 71
rect -5858 37 -5824 71
rect -5740 37 -5706 71
rect -5622 37 -5588 71
rect -5504 37 -5470 71
rect -5386 37 -5352 71
rect -5268 37 -5234 71
rect -5150 37 -5116 71
rect -5032 37 -4998 71
rect -4914 37 -4880 71
rect -4796 37 -4762 71
rect -4678 37 -4644 71
rect -4560 37 -4526 71
rect -4442 37 -4408 71
rect -4324 37 -4290 71
rect -4206 37 -4172 71
rect -4088 37 -4054 71
rect -3970 37 -3936 71
rect -3852 37 -3818 71
rect -3734 37 -3700 71
rect -3616 37 -3582 71
rect -3498 37 -3464 71
rect -3380 37 -3346 71
rect -3262 37 -3228 71
rect -3144 37 -3110 71
rect -3026 37 -2992 71
rect -2908 37 -2874 71
rect -2790 37 -2756 71
rect -2672 37 -2638 71
rect -2554 37 -2520 71
rect -2436 37 -2402 71
rect -2318 37 -2284 71
rect -2200 37 -2166 71
rect -2082 37 -2048 71
rect -1964 37 -1930 71
rect -1846 37 -1812 71
rect -1728 37 -1694 71
rect -1610 37 -1576 71
rect -1492 37 -1458 71
rect -1374 37 -1340 71
rect -1256 37 -1222 71
rect -1138 37 -1104 71
rect -1020 37 -986 71
rect -902 37 -868 71
rect -784 37 -750 71
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect 750 37 784 71
rect 868 37 902 71
rect 986 37 1020 71
rect 1104 37 1138 71
rect 1222 37 1256 71
rect 1340 37 1374 71
rect 1458 37 1492 71
rect 1576 37 1610 71
rect 1694 37 1728 71
rect 1812 37 1846 71
rect 1930 37 1964 71
rect 2048 37 2082 71
rect 2166 37 2200 71
rect 2284 37 2318 71
rect 2402 37 2436 71
rect 2520 37 2554 71
rect 2638 37 2672 71
rect 2756 37 2790 71
rect 2874 37 2908 71
rect 2992 37 3026 71
rect 3110 37 3144 71
rect 3228 37 3262 71
rect 3346 37 3380 71
rect 3464 37 3498 71
rect 3582 37 3616 71
rect 3700 37 3734 71
rect 3818 37 3852 71
rect 3936 37 3970 71
rect 4054 37 4088 71
rect 4172 37 4206 71
rect 4290 37 4324 71
rect 4408 37 4442 71
rect 4526 37 4560 71
rect 4644 37 4678 71
rect 4762 37 4796 71
rect 4880 37 4914 71
rect 4998 37 5032 71
rect 5116 37 5150 71
rect 5234 37 5268 71
rect 5352 37 5386 71
rect 5470 37 5504 71
rect 5588 37 5622 71
rect 5706 37 5740 71
rect 5824 37 5858 71
rect 5942 37 5976 71
rect 6060 37 6094 71
rect 6178 37 6212 71
rect 6296 37 6330 71
rect 6414 37 6448 71
rect 6532 37 6566 71
rect 6650 37 6684 71
rect 6768 37 6802 71
rect 6886 37 6920 71
rect 7004 37 7038 71
rect -7038 -71 -7004 -37
rect -6920 -71 -6886 -37
rect -6802 -71 -6768 -37
rect -6684 -71 -6650 -37
rect -6566 -71 -6532 -37
rect -6448 -71 -6414 -37
rect -6330 -71 -6296 -37
rect -6212 -71 -6178 -37
rect -6094 -71 -6060 -37
rect -5976 -71 -5942 -37
rect -5858 -71 -5824 -37
rect -5740 -71 -5706 -37
rect -5622 -71 -5588 -37
rect -5504 -71 -5470 -37
rect -5386 -71 -5352 -37
rect -5268 -71 -5234 -37
rect -5150 -71 -5116 -37
rect -5032 -71 -4998 -37
rect -4914 -71 -4880 -37
rect -4796 -71 -4762 -37
rect -4678 -71 -4644 -37
rect -4560 -71 -4526 -37
rect -4442 -71 -4408 -37
rect -4324 -71 -4290 -37
rect -4206 -71 -4172 -37
rect -4088 -71 -4054 -37
rect -3970 -71 -3936 -37
rect -3852 -71 -3818 -37
rect -3734 -71 -3700 -37
rect -3616 -71 -3582 -37
rect -3498 -71 -3464 -37
rect -3380 -71 -3346 -37
rect -3262 -71 -3228 -37
rect -3144 -71 -3110 -37
rect -3026 -71 -2992 -37
rect -2908 -71 -2874 -37
rect -2790 -71 -2756 -37
rect -2672 -71 -2638 -37
rect -2554 -71 -2520 -37
rect -2436 -71 -2402 -37
rect -2318 -71 -2284 -37
rect -2200 -71 -2166 -37
rect -2082 -71 -2048 -37
rect -1964 -71 -1930 -37
rect -1846 -71 -1812 -37
rect -1728 -71 -1694 -37
rect -1610 -71 -1576 -37
rect -1492 -71 -1458 -37
rect -1374 -71 -1340 -37
rect -1256 -71 -1222 -37
rect -1138 -71 -1104 -37
rect -1020 -71 -986 -37
rect -902 -71 -868 -37
rect -784 -71 -750 -37
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect 750 -71 784 -37
rect 868 -71 902 -37
rect 986 -71 1020 -37
rect 1104 -71 1138 -37
rect 1222 -71 1256 -37
rect 1340 -71 1374 -37
rect 1458 -71 1492 -37
rect 1576 -71 1610 -37
rect 1694 -71 1728 -37
rect 1812 -71 1846 -37
rect 1930 -71 1964 -37
rect 2048 -71 2082 -37
rect 2166 -71 2200 -37
rect 2284 -71 2318 -37
rect 2402 -71 2436 -37
rect 2520 -71 2554 -37
rect 2638 -71 2672 -37
rect 2756 -71 2790 -37
rect 2874 -71 2908 -37
rect 2992 -71 3026 -37
rect 3110 -71 3144 -37
rect 3228 -71 3262 -37
rect 3346 -71 3380 -37
rect 3464 -71 3498 -37
rect 3582 -71 3616 -37
rect 3700 -71 3734 -37
rect 3818 -71 3852 -37
rect 3936 -71 3970 -37
rect 4054 -71 4088 -37
rect 4172 -71 4206 -37
rect 4290 -71 4324 -37
rect 4408 -71 4442 -37
rect 4526 -71 4560 -37
rect 4644 -71 4678 -37
rect 4762 -71 4796 -37
rect 4880 -71 4914 -37
rect 4998 -71 5032 -37
rect 5116 -71 5150 -37
rect 5234 -71 5268 -37
rect 5352 -71 5386 -37
rect 5470 -71 5504 -37
rect 5588 -71 5622 -37
rect 5706 -71 5740 -37
rect 5824 -71 5858 -37
rect 5942 -71 5976 -37
rect 6060 -71 6094 -37
rect 6178 -71 6212 -37
rect 6296 -71 6330 -37
rect 6414 -71 6448 -37
rect 6532 -71 6566 -37
rect 6650 -71 6684 -37
rect 6768 -71 6802 -37
rect 6886 -71 6920 -37
rect 7004 -71 7038 -37
rect -7038 -799 -7004 -765
rect -6920 -799 -6886 -765
rect -6802 -799 -6768 -765
rect -6684 -799 -6650 -765
rect -6566 -799 -6532 -765
rect -6448 -799 -6414 -765
rect -6330 -799 -6296 -765
rect -6212 -799 -6178 -765
rect -6094 -799 -6060 -765
rect -5976 -799 -5942 -765
rect -5858 -799 -5824 -765
rect -5740 -799 -5706 -765
rect -5622 -799 -5588 -765
rect -5504 -799 -5470 -765
rect -5386 -799 -5352 -765
rect -5268 -799 -5234 -765
rect -5150 -799 -5116 -765
rect -5032 -799 -4998 -765
rect -4914 -799 -4880 -765
rect -4796 -799 -4762 -765
rect -4678 -799 -4644 -765
rect -4560 -799 -4526 -765
rect -4442 -799 -4408 -765
rect -4324 -799 -4290 -765
rect -4206 -799 -4172 -765
rect -4088 -799 -4054 -765
rect -3970 -799 -3936 -765
rect -3852 -799 -3818 -765
rect -3734 -799 -3700 -765
rect -3616 -799 -3582 -765
rect -3498 -799 -3464 -765
rect -3380 -799 -3346 -765
rect -3262 -799 -3228 -765
rect -3144 -799 -3110 -765
rect -3026 -799 -2992 -765
rect -2908 -799 -2874 -765
rect -2790 -799 -2756 -765
rect -2672 -799 -2638 -765
rect -2554 -799 -2520 -765
rect -2436 -799 -2402 -765
rect -2318 -799 -2284 -765
rect -2200 -799 -2166 -765
rect -2082 -799 -2048 -765
rect -1964 -799 -1930 -765
rect -1846 -799 -1812 -765
rect -1728 -799 -1694 -765
rect -1610 -799 -1576 -765
rect -1492 -799 -1458 -765
rect -1374 -799 -1340 -765
rect -1256 -799 -1222 -765
rect -1138 -799 -1104 -765
rect -1020 -799 -986 -765
rect -902 -799 -868 -765
rect -784 -799 -750 -765
rect -666 -799 -632 -765
rect -548 -799 -514 -765
rect -430 -799 -396 -765
rect -312 -799 -278 -765
rect -194 -799 -160 -765
rect -76 -799 -42 -765
rect 42 -799 76 -765
rect 160 -799 194 -765
rect 278 -799 312 -765
rect 396 -799 430 -765
rect 514 -799 548 -765
rect 632 -799 666 -765
rect 750 -799 784 -765
rect 868 -799 902 -765
rect 986 -799 1020 -765
rect 1104 -799 1138 -765
rect 1222 -799 1256 -765
rect 1340 -799 1374 -765
rect 1458 -799 1492 -765
rect 1576 -799 1610 -765
rect 1694 -799 1728 -765
rect 1812 -799 1846 -765
rect 1930 -799 1964 -765
rect 2048 -799 2082 -765
rect 2166 -799 2200 -765
rect 2284 -799 2318 -765
rect 2402 -799 2436 -765
rect 2520 -799 2554 -765
rect 2638 -799 2672 -765
rect 2756 -799 2790 -765
rect 2874 -799 2908 -765
rect 2992 -799 3026 -765
rect 3110 -799 3144 -765
rect 3228 -799 3262 -765
rect 3346 -799 3380 -765
rect 3464 -799 3498 -765
rect 3582 -799 3616 -765
rect 3700 -799 3734 -765
rect 3818 -799 3852 -765
rect 3936 -799 3970 -765
rect 4054 -799 4088 -765
rect 4172 -799 4206 -765
rect 4290 -799 4324 -765
rect 4408 -799 4442 -765
rect 4526 -799 4560 -765
rect 4644 -799 4678 -765
rect 4762 -799 4796 -765
rect 4880 -799 4914 -765
rect 4998 -799 5032 -765
rect 5116 -799 5150 -765
rect 5234 -799 5268 -765
rect 5352 -799 5386 -765
rect 5470 -799 5504 -765
rect 5588 -799 5622 -765
rect 5706 -799 5740 -765
rect 5824 -799 5858 -765
rect 5942 -799 5976 -765
rect 6060 -799 6094 -765
rect 6178 -799 6212 -765
rect 6296 -799 6330 -765
rect 6414 -799 6448 -765
rect 6532 -799 6566 -765
rect 6650 -799 6684 -765
rect 6768 -799 6802 -765
rect 6886 -799 6920 -765
rect 7004 -799 7038 -765
<< locali >>
rect -7211 867 -7115 901
rect 7115 867 7211 901
rect -7211 805 -7177 867
rect 7177 805 7211 867
rect -7054 765 -7038 799
rect -7004 765 -6988 799
rect -6936 765 -6920 799
rect -6886 765 -6870 799
rect -6818 765 -6802 799
rect -6768 765 -6752 799
rect -6700 765 -6684 799
rect -6650 765 -6634 799
rect -6582 765 -6566 799
rect -6532 765 -6516 799
rect -6464 765 -6448 799
rect -6414 765 -6398 799
rect -6346 765 -6330 799
rect -6296 765 -6280 799
rect -6228 765 -6212 799
rect -6178 765 -6162 799
rect -6110 765 -6094 799
rect -6060 765 -6044 799
rect -5992 765 -5976 799
rect -5942 765 -5926 799
rect -5874 765 -5858 799
rect -5824 765 -5808 799
rect -5756 765 -5740 799
rect -5706 765 -5690 799
rect -5638 765 -5622 799
rect -5588 765 -5572 799
rect -5520 765 -5504 799
rect -5470 765 -5454 799
rect -5402 765 -5386 799
rect -5352 765 -5336 799
rect -5284 765 -5268 799
rect -5234 765 -5218 799
rect -5166 765 -5150 799
rect -5116 765 -5100 799
rect -5048 765 -5032 799
rect -4998 765 -4982 799
rect -4930 765 -4914 799
rect -4880 765 -4864 799
rect -4812 765 -4796 799
rect -4762 765 -4746 799
rect -4694 765 -4678 799
rect -4644 765 -4628 799
rect -4576 765 -4560 799
rect -4526 765 -4510 799
rect -4458 765 -4442 799
rect -4408 765 -4392 799
rect -4340 765 -4324 799
rect -4290 765 -4274 799
rect -4222 765 -4206 799
rect -4172 765 -4156 799
rect -4104 765 -4088 799
rect -4054 765 -4038 799
rect -3986 765 -3970 799
rect -3936 765 -3920 799
rect -3868 765 -3852 799
rect -3818 765 -3802 799
rect -3750 765 -3734 799
rect -3700 765 -3684 799
rect -3632 765 -3616 799
rect -3582 765 -3566 799
rect -3514 765 -3498 799
rect -3464 765 -3448 799
rect -3396 765 -3380 799
rect -3346 765 -3330 799
rect -3278 765 -3262 799
rect -3228 765 -3212 799
rect -3160 765 -3144 799
rect -3110 765 -3094 799
rect -3042 765 -3026 799
rect -2992 765 -2976 799
rect -2924 765 -2908 799
rect -2874 765 -2858 799
rect -2806 765 -2790 799
rect -2756 765 -2740 799
rect -2688 765 -2672 799
rect -2638 765 -2622 799
rect -2570 765 -2554 799
rect -2520 765 -2504 799
rect -2452 765 -2436 799
rect -2402 765 -2386 799
rect -2334 765 -2318 799
rect -2284 765 -2268 799
rect -2216 765 -2200 799
rect -2166 765 -2150 799
rect -2098 765 -2082 799
rect -2048 765 -2032 799
rect -1980 765 -1964 799
rect -1930 765 -1914 799
rect -1862 765 -1846 799
rect -1812 765 -1796 799
rect -1744 765 -1728 799
rect -1694 765 -1678 799
rect -1626 765 -1610 799
rect -1576 765 -1560 799
rect -1508 765 -1492 799
rect -1458 765 -1442 799
rect -1390 765 -1374 799
rect -1340 765 -1324 799
rect -1272 765 -1256 799
rect -1222 765 -1206 799
rect -1154 765 -1138 799
rect -1104 765 -1088 799
rect -1036 765 -1020 799
rect -986 765 -970 799
rect -918 765 -902 799
rect -868 765 -852 799
rect -800 765 -784 799
rect -750 765 -734 799
rect -682 765 -666 799
rect -632 765 -616 799
rect -564 765 -548 799
rect -514 765 -498 799
rect -446 765 -430 799
rect -396 765 -380 799
rect -328 765 -312 799
rect -278 765 -262 799
rect -210 765 -194 799
rect -160 765 -144 799
rect -92 765 -76 799
rect -42 765 -26 799
rect 26 765 42 799
rect 76 765 92 799
rect 144 765 160 799
rect 194 765 210 799
rect 262 765 278 799
rect 312 765 328 799
rect 380 765 396 799
rect 430 765 446 799
rect 498 765 514 799
rect 548 765 564 799
rect 616 765 632 799
rect 666 765 682 799
rect 734 765 750 799
rect 784 765 800 799
rect 852 765 868 799
rect 902 765 918 799
rect 970 765 986 799
rect 1020 765 1036 799
rect 1088 765 1104 799
rect 1138 765 1154 799
rect 1206 765 1222 799
rect 1256 765 1272 799
rect 1324 765 1340 799
rect 1374 765 1390 799
rect 1442 765 1458 799
rect 1492 765 1508 799
rect 1560 765 1576 799
rect 1610 765 1626 799
rect 1678 765 1694 799
rect 1728 765 1744 799
rect 1796 765 1812 799
rect 1846 765 1862 799
rect 1914 765 1930 799
rect 1964 765 1980 799
rect 2032 765 2048 799
rect 2082 765 2098 799
rect 2150 765 2166 799
rect 2200 765 2216 799
rect 2268 765 2284 799
rect 2318 765 2334 799
rect 2386 765 2402 799
rect 2436 765 2452 799
rect 2504 765 2520 799
rect 2554 765 2570 799
rect 2622 765 2638 799
rect 2672 765 2688 799
rect 2740 765 2756 799
rect 2790 765 2806 799
rect 2858 765 2874 799
rect 2908 765 2924 799
rect 2976 765 2992 799
rect 3026 765 3042 799
rect 3094 765 3110 799
rect 3144 765 3160 799
rect 3212 765 3228 799
rect 3262 765 3278 799
rect 3330 765 3346 799
rect 3380 765 3396 799
rect 3448 765 3464 799
rect 3498 765 3514 799
rect 3566 765 3582 799
rect 3616 765 3632 799
rect 3684 765 3700 799
rect 3734 765 3750 799
rect 3802 765 3818 799
rect 3852 765 3868 799
rect 3920 765 3936 799
rect 3970 765 3986 799
rect 4038 765 4054 799
rect 4088 765 4104 799
rect 4156 765 4172 799
rect 4206 765 4222 799
rect 4274 765 4290 799
rect 4324 765 4340 799
rect 4392 765 4408 799
rect 4442 765 4458 799
rect 4510 765 4526 799
rect 4560 765 4576 799
rect 4628 765 4644 799
rect 4678 765 4694 799
rect 4746 765 4762 799
rect 4796 765 4812 799
rect 4864 765 4880 799
rect 4914 765 4930 799
rect 4982 765 4998 799
rect 5032 765 5048 799
rect 5100 765 5116 799
rect 5150 765 5166 799
rect 5218 765 5234 799
rect 5268 765 5284 799
rect 5336 765 5352 799
rect 5386 765 5402 799
rect 5454 765 5470 799
rect 5504 765 5520 799
rect 5572 765 5588 799
rect 5622 765 5638 799
rect 5690 765 5706 799
rect 5740 765 5756 799
rect 5808 765 5824 799
rect 5858 765 5874 799
rect 5926 765 5942 799
rect 5976 765 5992 799
rect 6044 765 6060 799
rect 6094 765 6110 799
rect 6162 765 6178 799
rect 6212 765 6228 799
rect 6280 765 6296 799
rect 6330 765 6346 799
rect 6398 765 6414 799
rect 6448 765 6464 799
rect 6516 765 6532 799
rect 6566 765 6582 799
rect 6634 765 6650 799
rect 6684 765 6700 799
rect 6752 765 6768 799
rect 6802 765 6818 799
rect 6870 765 6886 799
rect 6920 765 6936 799
rect 6988 765 7004 799
rect 7038 765 7054 799
rect -7097 706 -7063 722
rect -7097 114 -7063 130
rect -6979 706 -6945 722
rect -6979 114 -6945 130
rect -6861 706 -6827 722
rect -6861 114 -6827 130
rect -6743 706 -6709 722
rect -6743 114 -6709 130
rect -6625 706 -6591 722
rect -6625 114 -6591 130
rect -6507 706 -6473 722
rect -6507 114 -6473 130
rect -6389 706 -6355 722
rect -6389 114 -6355 130
rect -6271 706 -6237 722
rect -6271 114 -6237 130
rect -6153 706 -6119 722
rect -6153 114 -6119 130
rect -6035 706 -6001 722
rect -6035 114 -6001 130
rect -5917 706 -5883 722
rect -5917 114 -5883 130
rect -5799 706 -5765 722
rect -5799 114 -5765 130
rect -5681 706 -5647 722
rect -5681 114 -5647 130
rect -5563 706 -5529 722
rect -5563 114 -5529 130
rect -5445 706 -5411 722
rect -5445 114 -5411 130
rect -5327 706 -5293 722
rect -5327 114 -5293 130
rect -5209 706 -5175 722
rect -5209 114 -5175 130
rect -5091 706 -5057 722
rect -5091 114 -5057 130
rect -4973 706 -4939 722
rect -4973 114 -4939 130
rect -4855 706 -4821 722
rect -4855 114 -4821 130
rect -4737 706 -4703 722
rect -4737 114 -4703 130
rect -4619 706 -4585 722
rect -4619 114 -4585 130
rect -4501 706 -4467 722
rect -4501 114 -4467 130
rect -4383 706 -4349 722
rect -4383 114 -4349 130
rect -4265 706 -4231 722
rect -4265 114 -4231 130
rect -4147 706 -4113 722
rect -4147 114 -4113 130
rect -4029 706 -3995 722
rect -4029 114 -3995 130
rect -3911 706 -3877 722
rect -3911 114 -3877 130
rect -3793 706 -3759 722
rect -3793 114 -3759 130
rect -3675 706 -3641 722
rect -3675 114 -3641 130
rect -3557 706 -3523 722
rect -3557 114 -3523 130
rect -3439 706 -3405 722
rect -3439 114 -3405 130
rect -3321 706 -3287 722
rect -3321 114 -3287 130
rect -3203 706 -3169 722
rect -3203 114 -3169 130
rect -3085 706 -3051 722
rect -3085 114 -3051 130
rect -2967 706 -2933 722
rect -2967 114 -2933 130
rect -2849 706 -2815 722
rect -2849 114 -2815 130
rect -2731 706 -2697 722
rect -2731 114 -2697 130
rect -2613 706 -2579 722
rect -2613 114 -2579 130
rect -2495 706 -2461 722
rect -2495 114 -2461 130
rect -2377 706 -2343 722
rect -2377 114 -2343 130
rect -2259 706 -2225 722
rect -2259 114 -2225 130
rect -2141 706 -2107 722
rect -2141 114 -2107 130
rect -2023 706 -1989 722
rect -2023 114 -1989 130
rect -1905 706 -1871 722
rect -1905 114 -1871 130
rect -1787 706 -1753 722
rect -1787 114 -1753 130
rect -1669 706 -1635 722
rect -1669 114 -1635 130
rect -1551 706 -1517 722
rect -1551 114 -1517 130
rect -1433 706 -1399 722
rect -1433 114 -1399 130
rect -1315 706 -1281 722
rect -1315 114 -1281 130
rect -1197 706 -1163 722
rect -1197 114 -1163 130
rect -1079 706 -1045 722
rect -1079 114 -1045 130
rect -961 706 -927 722
rect -961 114 -927 130
rect -843 706 -809 722
rect -843 114 -809 130
rect -725 706 -691 722
rect -725 114 -691 130
rect -607 706 -573 722
rect -607 114 -573 130
rect -489 706 -455 722
rect -489 114 -455 130
rect -371 706 -337 722
rect -371 114 -337 130
rect -253 706 -219 722
rect -253 114 -219 130
rect -135 706 -101 722
rect -135 114 -101 130
rect -17 706 17 722
rect -17 114 17 130
rect 101 706 135 722
rect 101 114 135 130
rect 219 706 253 722
rect 219 114 253 130
rect 337 706 371 722
rect 337 114 371 130
rect 455 706 489 722
rect 455 114 489 130
rect 573 706 607 722
rect 573 114 607 130
rect 691 706 725 722
rect 691 114 725 130
rect 809 706 843 722
rect 809 114 843 130
rect 927 706 961 722
rect 927 114 961 130
rect 1045 706 1079 722
rect 1045 114 1079 130
rect 1163 706 1197 722
rect 1163 114 1197 130
rect 1281 706 1315 722
rect 1281 114 1315 130
rect 1399 706 1433 722
rect 1399 114 1433 130
rect 1517 706 1551 722
rect 1517 114 1551 130
rect 1635 706 1669 722
rect 1635 114 1669 130
rect 1753 706 1787 722
rect 1753 114 1787 130
rect 1871 706 1905 722
rect 1871 114 1905 130
rect 1989 706 2023 722
rect 1989 114 2023 130
rect 2107 706 2141 722
rect 2107 114 2141 130
rect 2225 706 2259 722
rect 2225 114 2259 130
rect 2343 706 2377 722
rect 2343 114 2377 130
rect 2461 706 2495 722
rect 2461 114 2495 130
rect 2579 706 2613 722
rect 2579 114 2613 130
rect 2697 706 2731 722
rect 2697 114 2731 130
rect 2815 706 2849 722
rect 2815 114 2849 130
rect 2933 706 2967 722
rect 2933 114 2967 130
rect 3051 706 3085 722
rect 3051 114 3085 130
rect 3169 706 3203 722
rect 3169 114 3203 130
rect 3287 706 3321 722
rect 3287 114 3321 130
rect 3405 706 3439 722
rect 3405 114 3439 130
rect 3523 706 3557 722
rect 3523 114 3557 130
rect 3641 706 3675 722
rect 3641 114 3675 130
rect 3759 706 3793 722
rect 3759 114 3793 130
rect 3877 706 3911 722
rect 3877 114 3911 130
rect 3995 706 4029 722
rect 3995 114 4029 130
rect 4113 706 4147 722
rect 4113 114 4147 130
rect 4231 706 4265 722
rect 4231 114 4265 130
rect 4349 706 4383 722
rect 4349 114 4383 130
rect 4467 706 4501 722
rect 4467 114 4501 130
rect 4585 706 4619 722
rect 4585 114 4619 130
rect 4703 706 4737 722
rect 4703 114 4737 130
rect 4821 706 4855 722
rect 4821 114 4855 130
rect 4939 706 4973 722
rect 4939 114 4973 130
rect 5057 706 5091 722
rect 5057 114 5091 130
rect 5175 706 5209 722
rect 5175 114 5209 130
rect 5293 706 5327 722
rect 5293 114 5327 130
rect 5411 706 5445 722
rect 5411 114 5445 130
rect 5529 706 5563 722
rect 5529 114 5563 130
rect 5647 706 5681 722
rect 5647 114 5681 130
rect 5765 706 5799 722
rect 5765 114 5799 130
rect 5883 706 5917 722
rect 5883 114 5917 130
rect 6001 706 6035 722
rect 6001 114 6035 130
rect 6119 706 6153 722
rect 6119 114 6153 130
rect 6237 706 6271 722
rect 6237 114 6271 130
rect 6355 706 6389 722
rect 6355 114 6389 130
rect 6473 706 6507 722
rect 6473 114 6507 130
rect 6591 706 6625 722
rect 6591 114 6625 130
rect 6709 706 6743 722
rect 6709 114 6743 130
rect 6827 706 6861 722
rect 6827 114 6861 130
rect 6945 706 6979 722
rect 6945 114 6979 130
rect 7063 706 7097 722
rect 7063 114 7097 130
rect -7054 37 -7038 71
rect -7004 37 -6988 71
rect -6936 37 -6920 71
rect -6886 37 -6870 71
rect -6818 37 -6802 71
rect -6768 37 -6752 71
rect -6700 37 -6684 71
rect -6650 37 -6634 71
rect -6582 37 -6566 71
rect -6532 37 -6516 71
rect -6464 37 -6448 71
rect -6414 37 -6398 71
rect -6346 37 -6330 71
rect -6296 37 -6280 71
rect -6228 37 -6212 71
rect -6178 37 -6162 71
rect -6110 37 -6094 71
rect -6060 37 -6044 71
rect -5992 37 -5976 71
rect -5942 37 -5926 71
rect -5874 37 -5858 71
rect -5824 37 -5808 71
rect -5756 37 -5740 71
rect -5706 37 -5690 71
rect -5638 37 -5622 71
rect -5588 37 -5572 71
rect -5520 37 -5504 71
rect -5470 37 -5454 71
rect -5402 37 -5386 71
rect -5352 37 -5336 71
rect -5284 37 -5268 71
rect -5234 37 -5218 71
rect -5166 37 -5150 71
rect -5116 37 -5100 71
rect -5048 37 -5032 71
rect -4998 37 -4982 71
rect -4930 37 -4914 71
rect -4880 37 -4864 71
rect -4812 37 -4796 71
rect -4762 37 -4746 71
rect -4694 37 -4678 71
rect -4644 37 -4628 71
rect -4576 37 -4560 71
rect -4526 37 -4510 71
rect -4458 37 -4442 71
rect -4408 37 -4392 71
rect -4340 37 -4324 71
rect -4290 37 -4274 71
rect -4222 37 -4206 71
rect -4172 37 -4156 71
rect -4104 37 -4088 71
rect -4054 37 -4038 71
rect -3986 37 -3970 71
rect -3936 37 -3920 71
rect -3868 37 -3852 71
rect -3818 37 -3802 71
rect -3750 37 -3734 71
rect -3700 37 -3684 71
rect -3632 37 -3616 71
rect -3582 37 -3566 71
rect -3514 37 -3498 71
rect -3464 37 -3448 71
rect -3396 37 -3380 71
rect -3346 37 -3330 71
rect -3278 37 -3262 71
rect -3228 37 -3212 71
rect -3160 37 -3144 71
rect -3110 37 -3094 71
rect -3042 37 -3026 71
rect -2992 37 -2976 71
rect -2924 37 -2908 71
rect -2874 37 -2858 71
rect -2806 37 -2790 71
rect -2756 37 -2740 71
rect -2688 37 -2672 71
rect -2638 37 -2622 71
rect -2570 37 -2554 71
rect -2520 37 -2504 71
rect -2452 37 -2436 71
rect -2402 37 -2386 71
rect -2334 37 -2318 71
rect -2284 37 -2268 71
rect -2216 37 -2200 71
rect -2166 37 -2150 71
rect -2098 37 -2082 71
rect -2048 37 -2032 71
rect -1980 37 -1964 71
rect -1930 37 -1914 71
rect -1862 37 -1846 71
rect -1812 37 -1796 71
rect -1744 37 -1728 71
rect -1694 37 -1678 71
rect -1626 37 -1610 71
rect -1576 37 -1560 71
rect -1508 37 -1492 71
rect -1458 37 -1442 71
rect -1390 37 -1374 71
rect -1340 37 -1324 71
rect -1272 37 -1256 71
rect -1222 37 -1206 71
rect -1154 37 -1138 71
rect -1104 37 -1088 71
rect -1036 37 -1020 71
rect -986 37 -970 71
rect -918 37 -902 71
rect -868 37 -852 71
rect -800 37 -784 71
rect -750 37 -734 71
rect -682 37 -666 71
rect -632 37 -616 71
rect -564 37 -548 71
rect -514 37 -498 71
rect -446 37 -430 71
rect -396 37 -380 71
rect -328 37 -312 71
rect -278 37 -262 71
rect -210 37 -194 71
rect -160 37 -144 71
rect -92 37 -76 71
rect -42 37 -26 71
rect 26 37 42 71
rect 76 37 92 71
rect 144 37 160 71
rect 194 37 210 71
rect 262 37 278 71
rect 312 37 328 71
rect 380 37 396 71
rect 430 37 446 71
rect 498 37 514 71
rect 548 37 564 71
rect 616 37 632 71
rect 666 37 682 71
rect 734 37 750 71
rect 784 37 800 71
rect 852 37 868 71
rect 902 37 918 71
rect 970 37 986 71
rect 1020 37 1036 71
rect 1088 37 1104 71
rect 1138 37 1154 71
rect 1206 37 1222 71
rect 1256 37 1272 71
rect 1324 37 1340 71
rect 1374 37 1390 71
rect 1442 37 1458 71
rect 1492 37 1508 71
rect 1560 37 1576 71
rect 1610 37 1626 71
rect 1678 37 1694 71
rect 1728 37 1744 71
rect 1796 37 1812 71
rect 1846 37 1862 71
rect 1914 37 1930 71
rect 1964 37 1980 71
rect 2032 37 2048 71
rect 2082 37 2098 71
rect 2150 37 2166 71
rect 2200 37 2216 71
rect 2268 37 2284 71
rect 2318 37 2334 71
rect 2386 37 2402 71
rect 2436 37 2452 71
rect 2504 37 2520 71
rect 2554 37 2570 71
rect 2622 37 2638 71
rect 2672 37 2688 71
rect 2740 37 2756 71
rect 2790 37 2806 71
rect 2858 37 2874 71
rect 2908 37 2924 71
rect 2976 37 2992 71
rect 3026 37 3042 71
rect 3094 37 3110 71
rect 3144 37 3160 71
rect 3212 37 3228 71
rect 3262 37 3278 71
rect 3330 37 3346 71
rect 3380 37 3396 71
rect 3448 37 3464 71
rect 3498 37 3514 71
rect 3566 37 3582 71
rect 3616 37 3632 71
rect 3684 37 3700 71
rect 3734 37 3750 71
rect 3802 37 3818 71
rect 3852 37 3868 71
rect 3920 37 3936 71
rect 3970 37 3986 71
rect 4038 37 4054 71
rect 4088 37 4104 71
rect 4156 37 4172 71
rect 4206 37 4222 71
rect 4274 37 4290 71
rect 4324 37 4340 71
rect 4392 37 4408 71
rect 4442 37 4458 71
rect 4510 37 4526 71
rect 4560 37 4576 71
rect 4628 37 4644 71
rect 4678 37 4694 71
rect 4746 37 4762 71
rect 4796 37 4812 71
rect 4864 37 4880 71
rect 4914 37 4930 71
rect 4982 37 4998 71
rect 5032 37 5048 71
rect 5100 37 5116 71
rect 5150 37 5166 71
rect 5218 37 5234 71
rect 5268 37 5284 71
rect 5336 37 5352 71
rect 5386 37 5402 71
rect 5454 37 5470 71
rect 5504 37 5520 71
rect 5572 37 5588 71
rect 5622 37 5638 71
rect 5690 37 5706 71
rect 5740 37 5756 71
rect 5808 37 5824 71
rect 5858 37 5874 71
rect 5926 37 5942 71
rect 5976 37 5992 71
rect 6044 37 6060 71
rect 6094 37 6110 71
rect 6162 37 6178 71
rect 6212 37 6228 71
rect 6280 37 6296 71
rect 6330 37 6346 71
rect 6398 37 6414 71
rect 6448 37 6464 71
rect 6516 37 6532 71
rect 6566 37 6582 71
rect 6634 37 6650 71
rect 6684 37 6700 71
rect 6752 37 6768 71
rect 6802 37 6818 71
rect 6870 37 6886 71
rect 6920 37 6936 71
rect 6988 37 7004 71
rect 7038 37 7054 71
rect -7054 -71 -7038 -37
rect -7004 -71 -6988 -37
rect -6936 -71 -6920 -37
rect -6886 -71 -6870 -37
rect -6818 -71 -6802 -37
rect -6768 -71 -6752 -37
rect -6700 -71 -6684 -37
rect -6650 -71 -6634 -37
rect -6582 -71 -6566 -37
rect -6532 -71 -6516 -37
rect -6464 -71 -6448 -37
rect -6414 -71 -6398 -37
rect -6346 -71 -6330 -37
rect -6296 -71 -6280 -37
rect -6228 -71 -6212 -37
rect -6178 -71 -6162 -37
rect -6110 -71 -6094 -37
rect -6060 -71 -6044 -37
rect -5992 -71 -5976 -37
rect -5942 -71 -5926 -37
rect -5874 -71 -5858 -37
rect -5824 -71 -5808 -37
rect -5756 -71 -5740 -37
rect -5706 -71 -5690 -37
rect -5638 -71 -5622 -37
rect -5588 -71 -5572 -37
rect -5520 -71 -5504 -37
rect -5470 -71 -5454 -37
rect -5402 -71 -5386 -37
rect -5352 -71 -5336 -37
rect -5284 -71 -5268 -37
rect -5234 -71 -5218 -37
rect -5166 -71 -5150 -37
rect -5116 -71 -5100 -37
rect -5048 -71 -5032 -37
rect -4998 -71 -4982 -37
rect -4930 -71 -4914 -37
rect -4880 -71 -4864 -37
rect -4812 -71 -4796 -37
rect -4762 -71 -4746 -37
rect -4694 -71 -4678 -37
rect -4644 -71 -4628 -37
rect -4576 -71 -4560 -37
rect -4526 -71 -4510 -37
rect -4458 -71 -4442 -37
rect -4408 -71 -4392 -37
rect -4340 -71 -4324 -37
rect -4290 -71 -4274 -37
rect -4222 -71 -4206 -37
rect -4172 -71 -4156 -37
rect -4104 -71 -4088 -37
rect -4054 -71 -4038 -37
rect -3986 -71 -3970 -37
rect -3936 -71 -3920 -37
rect -3868 -71 -3852 -37
rect -3818 -71 -3802 -37
rect -3750 -71 -3734 -37
rect -3700 -71 -3684 -37
rect -3632 -71 -3616 -37
rect -3582 -71 -3566 -37
rect -3514 -71 -3498 -37
rect -3464 -71 -3448 -37
rect -3396 -71 -3380 -37
rect -3346 -71 -3330 -37
rect -3278 -71 -3262 -37
rect -3228 -71 -3212 -37
rect -3160 -71 -3144 -37
rect -3110 -71 -3094 -37
rect -3042 -71 -3026 -37
rect -2992 -71 -2976 -37
rect -2924 -71 -2908 -37
rect -2874 -71 -2858 -37
rect -2806 -71 -2790 -37
rect -2756 -71 -2740 -37
rect -2688 -71 -2672 -37
rect -2638 -71 -2622 -37
rect -2570 -71 -2554 -37
rect -2520 -71 -2504 -37
rect -2452 -71 -2436 -37
rect -2402 -71 -2386 -37
rect -2334 -71 -2318 -37
rect -2284 -71 -2268 -37
rect -2216 -71 -2200 -37
rect -2166 -71 -2150 -37
rect -2098 -71 -2082 -37
rect -2048 -71 -2032 -37
rect -1980 -71 -1964 -37
rect -1930 -71 -1914 -37
rect -1862 -71 -1846 -37
rect -1812 -71 -1796 -37
rect -1744 -71 -1728 -37
rect -1694 -71 -1678 -37
rect -1626 -71 -1610 -37
rect -1576 -71 -1560 -37
rect -1508 -71 -1492 -37
rect -1458 -71 -1442 -37
rect -1390 -71 -1374 -37
rect -1340 -71 -1324 -37
rect -1272 -71 -1256 -37
rect -1222 -71 -1206 -37
rect -1154 -71 -1138 -37
rect -1104 -71 -1088 -37
rect -1036 -71 -1020 -37
rect -986 -71 -970 -37
rect -918 -71 -902 -37
rect -868 -71 -852 -37
rect -800 -71 -784 -37
rect -750 -71 -734 -37
rect -682 -71 -666 -37
rect -632 -71 -616 -37
rect -564 -71 -548 -37
rect -514 -71 -498 -37
rect -446 -71 -430 -37
rect -396 -71 -380 -37
rect -328 -71 -312 -37
rect -278 -71 -262 -37
rect -210 -71 -194 -37
rect -160 -71 -144 -37
rect -92 -71 -76 -37
rect -42 -71 -26 -37
rect 26 -71 42 -37
rect 76 -71 92 -37
rect 144 -71 160 -37
rect 194 -71 210 -37
rect 262 -71 278 -37
rect 312 -71 328 -37
rect 380 -71 396 -37
rect 430 -71 446 -37
rect 498 -71 514 -37
rect 548 -71 564 -37
rect 616 -71 632 -37
rect 666 -71 682 -37
rect 734 -71 750 -37
rect 784 -71 800 -37
rect 852 -71 868 -37
rect 902 -71 918 -37
rect 970 -71 986 -37
rect 1020 -71 1036 -37
rect 1088 -71 1104 -37
rect 1138 -71 1154 -37
rect 1206 -71 1222 -37
rect 1256 -71 1272 -37
rect 1324 -71 1340 -37
rect 1374 -71 1390 -37
rect 1442 -71 1458 -37
rect 1492 -71 1508 -37
rect 1560 -71 1576 -37
rect 1610 -71 1626 -37
rect 1678 -71 1694 -37
rect 1728 -71 1744 -37
rect 1796 -71 1812 -37
rect 1846 -71 1862 -37
rect 1914 -71 1930 -37
rect 1964 -71 1980 -37
rect 2032 -71 2048 -37
rect 2082 -71 2098 -37
rect 2150 -71 2166 -37
rect 2200 -71 2216 -37
rect 2268 -71 2284 -37
rect 2318 -71 2334 -37
rect 2386 -71 2402 -37
rect 2436 -71 2452 -37
rect 2504 -71 2520 -37
rect 2554 -71 2570 -37
rect 2622 -71 2638 -37
rect 2672 -71 2688 -37
rect 2740 -71 2756 -37
rect 2790 -71 2806 -37
rect 2858 -71 2874 -37
rect 2908 -71 2924 -37
rect 2976 -71 2992 -37
rect 3026 -71 3042 -37
rect 3094 -71 3110 -37
rect 3144 -71 3160 -37
rect 3212 -71 3228 -37
rect 3262 -71 3278 -37
rect 3330 -71 3346 -37
rect 3380 -71 3396 -37
rect 3448 -71 3464 -37
rect 3498 -71 3514 -37
rect 3566 -71 3582 -37
rect 3616 -71 3632 -37
rect 3684 -71 3700 -37
rect 3734 -71 3750 -37
rect 3802 -71 3818 -37
rect 3852 -71 3868 -37
rect 3920 -71 3936 -37
rect 3970 -71 3986 -37
rect 4038 -71 4054 -37
rect 4088 -71 4104 -37
rect 4156 -71 4172 -37
rect 4206 -71 4222 -37
rect 4274 -71 4290 -37
rect 4324 -71 4340 -37
rect 4392 -71 4408 -37
rect 4442 -71 4458 -37
rect 4510 -71 4526 -37
rect 4560 -71 4576 -37
rect 4628 -71 4644 -37
rect 4678 -71 4694 -37
rect 4746 -71 4762 -37
rect 4796 -71 4812 -37
rect 4864 -71 4880 -37
rect 4914 -71 4930 -37
rect 4982 -71 4998 -37
rect 5032 -71 5048 -37
rect 5100 -71 5116 -37
rect 5150 -71 5166 -37
rect 5218 -71 5234 -37
rect 5268 -71 5284 -37
rect 5336 -71 5352 -37
rect 5386 -71 5402 -37
rect 5454 -71 5470 -37
rect 5504 -71 5520 -37
rect 5572 -71 5588 -37
rect 5622 -71 5638 -37
rect 5690 -71 5706 -37
rect 5740 -71 5756 -37
rect 5808 -71 5824 -37
rect 5858 -71 5874 -37
rect 5926 -71 5942 -37
rect 5976 -71 5992 -37
rect 6044 -71 6060 -37
rect 6094 -71 6110 -37
rect 6162 -71 6178 -37
rect 6212 -71 6228 -37
rect 6280 -71 6296 -37
rect 6330 -71 6346 -37
rect 6398 -71 6414 -37
rect 6448 -71 6464 -37
rect 6516 -71 6532 -37
rect 6566 -71 6582 -37
rect 6634 -71 6650 -37
rect 6684 -71 6700 -37
rect 6752 -71 6768 -37
rect 6802 -71 6818 -37
rect 6870 -71 6886 -37
rect 6920 -71 6936 -37
rect 6988 -71 7004 -37
rect 7038 -71 7054 -37
rect -7097 -130 -7063 -114
rect -7097 -722 -7063 -706
rect -6979 -130 -6945 -114
rect -6979 -722 -6945 -706
rect -6861 -130 -6827 -114
rect -6861 -722 -6827 -706
rect -6743 -130 -6709 -114
rect -6743 -722 -6709 -706
rect -6625 -130 -6591 -114
rect -6625 -722 -6591 -706
rect -6507 -130 -6473 -114
rect -6507 -722 -6473 -706
rect -6389 -130 -6355 -114
rect -6389 -722 -6355 -706
rect -6271 -130 -6237 -114
rect -6271 -722 -6237 -706
rect -6153 -130 -6119 -114
rect -6153 -722 -6119 -706
rect -6035 -130 -6001 -114
rect -6035 -722 -6001 -706
rect -5917 -130 -5883 -114
rect -5917 -722 -5883 -706
rect -5799 -130 -5765 -114
rect -5799 -722 -5765 -706
rect -5681 -130 -5647 -114
rect -5681 -722 -5647 -706
rect -5563 -130 -5529 -114
rect -5563 -722 -5529 -706
rect -5445 -130 -5411 -114
rect -5445 -722 -5411 -706
rect -5327 -130 -5293 -114
rect -5327 -722 -5293 -706
rect -5209 -130 -5175 -114
rect -5209 -722 -5175 -706
rect -5091 -130 -5057 -114
rect -5091 -722 -5057 -706
rect -4973 -130 -4939 -114
rect -4973 -722 -4939 -706
rect -4855 -130 -4821 -114
rect -4855 -722 -4821 -706
rect -4737 -130 -4703 -114
rect -4737 -722 -4703 -706
rect -4619 -130 -4585 -114
rect -4619 -722 -4585 -706
rect -4501 -130 -4467 -114
rect -4501 -722 -4467 -706
rect -4383 -130 -4349 -114
rect -4383 -722 -4349 -706
rect -4265 -130 -4231 -114
rect -4265 -722 -4231 -706
rect -4147 -130 -4113 -114
rect -4147 -722 -4113 -706
rect -4029 -130 -3995 -114
rect -4029 -722 -3995 -706
rect -3911 -130 -3877 -114
rect -3911 -722 -3877 -706
rect -3793 -130 -3759 -114
rect -3793 -722 -3759 -706
rect -3675 -130 -3641 -114
rect -3675 -722 -3641 -706
rect -3557 -130 -3523 -114
rect -3557 -722 -3523 -706
rect -3439 -130 -3405 -114
rect -3439 -722 -3405 -706
rect -3321 -130 -3287 -114
rect -3321 -722 -3287 -706
rect -3203 -130 -3169 -114
rect -3203 -722 -3169 -706
rect -3085 -130 -3051 -114
rect -3085 -722 -3051 -706
rect -2967 -130 -2933 -114
rect -2967 -722 -2933 -706
rect -2849 -130 -2815 -114
rect -2849 -722 -2815 -706
rect -2731 -130 -2697 -114
rect -2731 -722 -2697 -706
rect -2613 -130 -2579 -114
rect -2613 -722 -2579 -706
rect -2495 -130 -2461 -114
rect -2495 -722 -2461 -706
rect -2377 -130 -2343 -114
rect -2377 -722 -2343 -706
rect -2259 -130 -2225 -114
rect -2259 -722 -2225 -706
rect -2141 -130 -2107 -114
rect -2141 -722 -2107 -706
rect -2023 -130 -1989 -114
rect -2023 -722 -1989 -706
rect -1905 -130 -1871 -114
rect -1905 -722 -1871 -706
rect -1787 -130 -1753 -114
rect -1787 -722 -1753 -706
rect -1669 -130 -1635 -114
rect -1669 -722 -1635 -706
rect -1551 -130 -1517 -114
rect -1551 -722 -1517 -706
rect -1433 -130 -1399 -114
rect -1433 -722 -1399 -706
rect -1315 -130 -1281 -114
rect -1315 -722 -1281 -706
rect -1197 -130 -1163 -114
rect -1197 -722 -1163 -706
rect -1079 -130 -1045 -114
rect -1079 -722 -1045 -706
rect -961 -130 -927 -114
rect -961 -722 -927 -706
rect -843 -130 -809 -114
rect -843 -722 -809 -706
rect -725 -130 -691 -114
rect -725 -722 -691 -706
rect -607 -130 -573 -114
rect -607 -722 -573 -706
rect -489 -130 -455 -114
rect -489 -722 -455 -706
rect -371 -130 -337 -114
rect -371 -722 -337 -706
rect -253 -130 -219 -114
rect -253 -722 -219 -706
rect -135 -130 -101 -114
rect -135 -722 -101 -706
rect -17 -130 17 -114
rect -17 -722 17 -706
rect 101 -130 135 -114
rect 101 -722 135 -706
rect 219 -130 253 -114
rect 219 -722 253 -706
rect 337 -130 371 -114
rect 337 -722 371 -706
rect 455 -130 489 -114
rect 455 -722 489 -706
rect 573 -130 607 -114
rect 573 -722 607 -706
rect 691 -130 725 -114
rect 691 -722 725 -706
rect 809 -130 843 -114
rect 809 -722 843 -706
rect 927 -130 961 -114
rect 927 -722 961 -706
rect 1045 -130 1079 -114
rect 1045 -722 1079 -706
rect 1163 -130 1197 -114
rect 1163 -722 1197 -706
rect 1281 -130 1315 -114
rect 1281 -722 1315 -706
rect 1399 -130 1433 -114
rect 1399 -722 1433 -706
rect 1517 -130 1551 -114
rect 1517 -722 1551 -706
rect 1635 -130 1669 -114
rect 1635 -722 1669 -706
rect 1753 -130 1787 -114
rect 1753 -722 1787 -706
rect 1871 -130 1905 -114
rect 1871 -722 1905 -706
rect 1989 -130 2023 -114
rect 1989 -722 2023 -706
rect 2107 -130 2141 -114
rect 2107 -722 2141 -706
rect 2225 -130 2259 -114
rect 2225 -722 2259 -706
rect 2343 -130 2377 -114
rect 2343 -722 2377 -706
rect 2461 -130 2495 -114
rect 2461 -722 2495 -706
rect 2579 -130 2613 -114
rect 2579 -722 2613 -706
rect 2697 -130 2731 -114
rect 2697 -722 2731 -706
rect 2815 -130 2849 -114
rect 2815 -722 2849 -706
rect 2933 -130 2967 -114
rect 2933 -722 2967 -706
rect 3051 -130 3085 -114
rect 3051 -722 3085 -706
rect 3169 -130 3203 -114
rect 3169 -722 3203 -706
rect 3287 -130 3321 -114
rect 3287 -722 3321 -706
rect 3405 -130 3439 -114
rect 3405 -722 3439 -706
rect 3523 -130 3557 -114
rect 3523 -722 3557 -706
rect 3641 -130 3675 -114
rect 3641 -722 3675 -706
rect 3759 -130 3793 -114
rect 3759 -722 3793 -706
rect 3877 -130 3911 -114
rect 3877 -722 3911 -706
rect 3995 -130 4029 -114
rect 3995 -722 4029 -706
rect 4113 -130 4147 -114
rect 4113 -722 4147 -706
rect 4231 -130 4265 -114
rect 4231 -722 4265 -706
rect 4349 -130 4383 -114
rect 4349 -722 4383 -706
rect 4467 -130 4501 -114
rect 4467 -722 4501 -706
rect 4585 -130 4619 -114
rect 4585 -722 4619 -706
rect 4703 -130 4737 -114
rect 4703 -722 4737 -706
rect 4821 -130 4855 -114
rect 4821 -722 4855 -706
rect 4939 -130 4973 -114
rect 4939 -722 4973 -706
rect 5057 -130 5091 -114
rect 5057 -722 5091 -706
rect 5175 -130 5209 -114
rect 5175 -722 5209 -706
rect 5293 -130 5327 -114
rect 5293 -722 5327 -706
rect 5411 -130 5445 -114
rect 5411 -722 5445 -706
rect 5529 -130 5563 -114
rect 5529 -722 5563 -706
rect 5647 -130 5681 -114
rect 5647 -722 5681 -706
rect 5765 -130 5799 -114
rect 5765 -722 5799 -706
rect 5883 -130 5917 -114
rect 5883 -722 5917 -706
rect 6001 -130 6035 -114
rect 6001 -722 6035 -706
rect 6119 -130 6153 -114
rect 6119 -722 6153 -706
rect 6237 -130 6271 -114
rect 6237 -722 6271 -706
rect 6355 -130 6389 -114
rect 6355 -722 6389 -706
rect 6473 -130 6507 -114
rect 6473 -722 6507 -706
rect 6591 -130 6625 -114
rect 6591 -722 6625 -706
rect 6709 -130 6743 -114
rect 6709 -722 6743 -706
rect 6827 -130 6861 -114
rect 6827 -722 6861 -706
rect 6945 -130 6979 -114
rect 6945 -722 6979 -706
rect 7063 -130 7097 -114
rect 7063 -722 7097 -706
rect -7054 -799 -7038 -765
rect -7004 -799 -6988 -765
rect -6936 -799 -6920 -765
rect -6886 -799 -6870 -765
rect -6818 -799 -6802 -765
rect -6768 -799 -6752 -765
rect -6700 -799 -6684 -765
rect -6650 -799 -6634 -765
rect -6582 -799 -6566 -765
rect -6532 -799 -6516 -765
rect -6464 -799 -6448 -765
rect -6414 -799 -6398 -765
rect -6346 -799 -6330 -765
rect -6296 -799 -6280 -765
rect -6228 -799 -6212 -765
rect -6178 -799 -6162 -765
rect -6110 -799 -6094 -765
rect -6060 -799 -6044 -765
rect -5992 -799 -5976 -765
rect -5942 -799 -5926 -765
rect -5874 -799 -5858 -765
rect -5824 -799 -5808 -765
rect -5756 -799 -5740 -765
rect -5706 -799 -5690 -765
rect -5638 -799 -5622 -765
rect -5588 -799 -5572 -765
rect -5520 -799 -5504 -765
rect -5470 -799 -5454 -765
rect -5402 -799 -5386 -765
rect -5352 -799 -5336 -765
rect -5284 -799 -5268 -765
rect -5234 -799 -5218 -765
rect -5166 -799 -5150 -765
rect -5116 -799 -5100 -765
rect -5048 -799 -5032 -765
rect -4998 -799 -4982 -765
rect -4930 -799 -4914 -765
rect -4880 -799 -4864 -765
rect -4812 -799 -4796 -765
rect -4762 -799 -4746 -765
rect -4694 -799 -4678 -765
rect -4644 -799 -4628 -765
rect -4576 -799 -4560 -765
rect -4526 -799 -4510 -765
rect -4458 -799 -4442 -765
rect -4408 -799 -4392 -765
rect -4340 -799 -4324 -765
rect -4290 -799 -4274 -765
rect -4222 -799 -4206 -765
rect -4172 -799 -4156 -765
rect -4104 -799 -4088 -765
rect -4054 -799 -4038 -765
rect -3986 -799 -3970 -765
rect -3936 -799 -3920 -765
rect -3868 -799 -3852 -765
rect -3818 -799 -3802 -765
rect -3750 -799 -3734 -765
rect -3700 -799 -3684 -765
rect -3632 -799 -3616 -765
rect -3582 -799 -3566 -765
rect -3514 -799 -3498 -765
rect -3464 -799 -3448 -765
rect -3396 -799 -3380 -765
rect -3346 -799 -3330 -765
rect -3278 -799 -3262 -765
rect -3228 -799 -3212 -765
rect -3160 -799 -3144 -765
rect -3110 -799 -3094 -765
rect -3042 -799 -3026 -765
rect -2992 -799 -2976 -765
rect -2924 -799 -2908 -765
rect -2874 -799 -2858 -765
rect -2806 -799 -2790 -765
rect -2756 -799 -2740 -765
rect -2688 -799 -2672 -765
rect -2638 -799 -2622 -765
rect -2570 -799 -2554 -765
rect -2520 -799 -2504 -765
rect -2452 -799 -2436 -765
rect -2402 -799 -2386 -765
rect -2334 -799 -2318 -765
rect -2284 -799 -2268 -765
rect -2216 -799 -2200 -765
rect -2166 -799 -2150 -765
rect -2098 -799 -2082 -765
rect -2048 -799 -2032 -765
rect -1980 -799 -1964 -765
rect -1930 -799 -1914 -765
rect -1862 -799 -1846 -765
rect -1812 -799 -1796 -765
rect -1744 -799 -1728 -765
rect -1694 -799 -1678 -765
rect -1626 -799 -1610 -765
rect -1576 -799 -1560 -765
rect -1508 -799 -1492 -765
rect -1458 -799 -1442 -765
rect -1390 -799 -1374 -765
rect -1340 -799 -1324 -765
rect -1272 -799 -1256 -765
rect -1222 -799 -1206 -765
rect -1154 -799 -1138 -765
rect -1104 -799 -1088 -765
rect -1036 -799 -1020 -765
rect -986 -799 -970 -765
rect -918 -799 -902 -765
rect -868 -799 -852 -765
rect -800 -799 -784 -765
rect -750 -799 -734 -765
rect -682 -799 -666 -765
rect -632 -799 -616 -765
rect -564 -799 -548 -765
rect -514 -799 -498 -765
rect -446 -799 -430 -765
rect -396 -799 -380 -765
rect -328 -799 -312 -765
rect -278 -799 -262 -765
rect -210 -799 -194 -765
rect -160 -799 -144 -765
rect -92 -799 -76 -765
rect -42 -799 -26 -765
rect 26 -799 42 -765
rect 76 -799 92 -765
rect 144 -799 160 -765
rect 194 -799 210 -765
rect 262 -799 278 -765
rect 312 -799 328 -765
rect 380 -799 396 -765
rect 430 -799 446 -765
rect 498 -799 514 -765
rect 548 -799 564 -765
rect 616 -799 632 -765
rect 666 -799 682 -765
rect 734 -799 750 -765
rect 784 -799 800 -765
rect 852 -799 868 -765
rect 902 -799 918 -765
rect 970 -799 986 -765
rect 1020 -799 1036 -765
rect 1088 -799 1104 -765
rect 1138 -799 1154 -765
rect 1206 -799 1222 -765
rect 1256 -799 1272 -765
rect 1324 -799 1340 -765
rect 1374 -799 1390 -765
rect 1442 -799 1458 -765
rect 1492 -799 1508 -765
rect 1560 -799 1576 -765
rect 1610 -799 1626 -765
rect 1678 -799 1694 -765
rect 1728 -799 1744 -765
rect 1796 -799 1812 -765
rect 1846 -799 1862 -765
rect 1914 -799 1930 -765
rect 1964 -799 1980 -765
rect 2032 -799 2048 -765
rect 2082 -799 2098 -765
rect 2150 -799 2166 -765
rect 2200 -799 2216 -765
rect 2268 -799 2284 -765
rect 2318 -799 2334 -765
rect 2386 -799 2402 -765
rect 2436 -799 2452 -765
rect 2504 -799 2520 -765
rect 2554 -799 2570 -765
rect 2622 -799 2638 -765
rect 2672 -799 2688 -765
rect 2740 -799 2756 -765
rect 2790 -799 2806 -765
rect 2858 -799 2874 -765
rect 2908 -799 2924 -765
rect 2976 -799 2992 -765
rect 3026 -799 3042 -765
rect 3094 -799 3110 -765
rect 3144 -799 3160 -765
rect 3212 -799 3228 -765
rect 3262 -799 3278 -765
rect 3330 -799 3346 -765
rect 3380 -799 3396 -765
rect 3448 -799 3464 -765
rect 3498 -799 3514 -765
rect 3566 -799 3582 -765
rect 3616 -799 3632 -765
rect 3684 -799 3700 -765
rect 3734 -799 3750 -765
rect 3802 -799 3818 -765
rect 3852 -799 3868 -765
rect 3920 -799 3936 -765
rect 3970 -799 3986 -765
rect 4038 -799 4054 -765
rect 4088 -799 4104 -765
rect 4156 -799 4172 -765
rect 4206 -799 4222 -765
rect 4274 -799 4290 -765
rect 4324 -799 4340 -765
rect 4392 -799 4408 -765
rect 4442 -799 4458 -765
rect 4510 -799 4526 -765
rect 4560 -799 4576 -765
rect 4628 -799 4644 -765
rect 4678 -799 4694 -765
rect 4746 -799 4762 -765
rect 4796 -799 4812 -765
rect 4864 -799 4880 -765
rect 4914 -799 4930 -765
rect 4982 -799 4998 -765
rect 5032 -799 5048 -765
rect 5100 -799 5116 -765
rect 5150 -799 5166 -765
rect 5218 -799 5234 -765
rect 5268 -799 5284 -765
rect 5336 -799 5352 -765
rect 5386 -799 5402 -765
rect 5454 -799 5470 -765
rect 5504 -799 5520 -765
rect 5572 -799 5588 -765
rect 5622 -799 5638 -765
rect 5690 -799 5706 -765
rect 5740 -799 5756 -765
rect 5808 -799 5824 -765
rect 5858 -799 5874 -765
rect 5926 -799 5942 -765
rect 5976 -799 5992 -765
rect 6044 -799 6060 -765
rect 6094 -799 6110 -765
rect 6162 -799 6178 -765
rect 6212 -799 6228 -765
rect 6280 -799 6296 -765
rect 6330 -799 6346 -765
rect 6398 -799 6414 -765
rect 6448 -799 6464 -765
rect 6516 -799 6532 -765
rect 6566 -799 6582 -765
rect 6634 -799 6650 -765
rect 6684 -799 6700 -765
rect 6752 -799 6768 -765
rect 6802 -799 6818 -765
rect 6870 -799 6886 -765
rect 6920 -799 6936 -765
rect 6988 -799 7004 -765
rect 7038 -799 7054 -765
rect -7211 -867 -7177 -805
rect 7177 -867 7211 -805
rect -7211 -901 -7115 -867
rect 7115 -901 7211 -867
<< viali >>
rect -7038 765 -7004 799
rect -6920 765 -6886 799
rect -6802 765 -6768 799
rect -6684 765 -6650 799
rect -6566 765 -6532 799
rect -6448 765 -6414 799
rect -6330 765 -6296 799
rect -6212 765 -6178 799
rect -6094 765 -6060 799
rect -5976 765 -5942 799
rect -5858 765 -5824 799
rect -5740 765 -5706 799
rect -5622 765 -5588 799
rect -5504 765 -5470 799
rect -5386 765 -5352 799
rect -5268 765 -5234 799
rect -5150 765 -5116 799
rect -5032 765 -4998 799
rect -4914 765 -4880 799
rect -4796 765 -4762 799
rect -4678 765 -4644 799
rect -4560 765 -4526 799
rect -4442 765 -4408 799
rect -4324 765 -4290 799
rect -4206 765 -4172 799
rect -4088 765 -4054 799
rect -3970 765 -3936 799
rect -3852 765 -3818 799
rect -3734 765 -3700 799
rect -3616 765 -3582 799
rect -3498 765 -3464 799
rect -3380 765 -3346 799
rect -3262 765 -3228 799
rect -3144 765 -3110 799
rect -3026 765 -2992 799
rect -2908 765 -2874 799
rect -2790 765 -2756 799
rect -2672 765 -2638 799
rect -2554 765 -2520 799
rect -2436 765 -2402 799
rect -2318 765 -2284 799
rect -2200 765 -2166 799
rect -2082 765 -2048 799
rect -1964 765 -1930 799
rect -1846 765 -1812 799
rect -1728 765 -1694 799
rect -1610 765 -1576 799
rect -1492 765 -1458 799
rect -1374 765 -1340 799
rect -1256 765 -1222 799
rect -1138 765 -1104 799
rect -1020 765 -986 799
rect -902 765 -868 799
rect -784 765 -750 799
rect -666 765 -632 799
rect -548 765 -514 799
rect -430 765 -396 799
rect -312 765 -278 799
rect -194 765 -160 799
rect -76 765 -42 799
rect 42 765 76 799
rect 160 765 194 799
rect 278 765 312 799
rect 396 765 430 799
rect 514 765 548 799
rect 632 765 666 799
rect 750 765 784 799
rect 868 765 902 799
rect 986 765 1020 799
rect 1104 765 1138 799
rect 1222 765 1256 799
rect 1340 765 1374 799
rect 1458 765 1492 799
rect 1576 765 1610 799
rect 1694 765 1728 799
rect 1812 765 1846 799
rect 1930 765 1964 799
rect 2048 765 2082 799
rect 2166 765 2200 799
rect 2284 765 2318 799
rect 2402 765 2436 799
rect 2520 765 2554 799
rect 2638 765 2672 799
rect 2756 765 2790 799
rect 2874 765 2908 799
rect 2992 765 3026 799
rect 3110 765 3144 799
rect 3228 765 3262 799
rect 3346 765 3380 799
rect 3464 765 3498 799
rect 3582 765 3616 799
rect 3700 765 3734 799
rect 3818 765 3852 799
rect 3936 765 3970 799
rect 4054 765 4088 799
rect 4172 765 4206 799
rect 4290 765 4324 799
rect 4408 765 4442 799
rect 4526 765 4560 799
rect 4644 765 4678 799
rect 4762 765 4796 799
rect 4880 765 4914 799
rect 4998 765 5032 799
rect 5116 765 5150 799
rect 5234 765 5268 799
rect 5352 765 5386 799
rect 5470 765 5504 799
rect 5588 765 5622 799
rect 5706 765 5740 799
rect 5824 765 5858 799
rect 5942 765 5976 799
rect 6060 765 6094 799
rect 6178 765 6212 799
rect 6296 765 6330 799
rect 6414 765 6448 799
rect 6532 765 6566 799
rect 6650 765 6684 799
rect 6768 765 6802 799
rect 6886 765 6920 799
rect 7004 765 7038 799
rect -7097 130 -7063 706
rect -6979 130 -6945 706
rect -6861 130 -6827 706
rect -6743 130 -6709 706
rect -6625 130 -6591 706
rect -6507 130 -6473 706
rect -6389 130 -6355 706
rect -6271 130 -6237 706
rect -6153 130 -6119 706
rect -6035 130 -6001 706
rect -5917 130 -5883 706
rect -5799 130 -5765 706
rect -5681 130 -5647 706
rect -5563 130 -5529 706
rect -5445 130 -5411 706
rect -5327 130 -5293 706
rect -5209 130 -5175 706
rect -5091 130 -5057 706
rect -4973 130 -4939 706
rect -4855 130 -4821 706
rect -4737 130 -4703 706
rect -4619 130 -4585 706
rect -4501 130 -4467 706
rect -4383 130 -4349 706
rect -4265 130 -4231 706
rect -4147 130 -4113 706
rect -4029 130 -3995 706
rect -3911 130 -3877 706
rect -3793 130 -3759 706
rect -3675 130 -3641 706
rect -3557 130 -3523 706
rect -3439 130 -3405 706
rect -3321 130 -3287 706
rect -3203 130 -3169 706
rect -3085 130 -3051 706
rect -2967 130 -2933 706
rect -2849 130 -2815 706
rect -2731 130 -2697 706
rect -2613 130 -2579 706
rect -2495 130 -2461 706
rect -2377 130 -2343 706
rect -2259 130 -2225 706
rect -2141 130 -2107 706
rect -2023 130 -1989 706
rect -1905 130 -1871 706
rect -1787 130 -1753 706
rect -1669 130 -1635 706
rect -1551 130 -1517 706
rect -1433 130 -1399 706
rect -1315 130 -1281 706
rect -1197 130 -1163 706
rect -1079 130 -1045 706
rect -961 130 -927 706
rect -843 130 -809 706
rect -725 130 -691 706
rect -607 130 -573 706
rect -489 130 -455 706
rect -371 130 -337 706
rect -253 130 -219 706
rect -135 130 -101 706
rect -17 130 17 706
rect 101 130 135 706
rect 219 130 253 706
rect 337 130 371 706
rect 455 130 489 706
rect 573 130 607 706
rect 691 130 725 706
rect 809 130 843 706
rect 927 130 961 706
rect 1045 130 1079 706
rect 1163 130 1197 706
rect 1281 130 1315 706
rect 1399 130 1433 706
rect 1517 130 1551 706
rect 1635 130 1669 706
rect 1753 130 1787 706
rect 1871 130 1905 706
rect 1989 130 2023 706
rect 2107 130 2141 706
rect 2225 130 2259 706
rect 2343 130 2377 706
rect 2461 130 2495 706
rect 2579 130 2613 706
rect 2697 130 2731 706
rect 2815 130 2849 706
rect 2933 130 2967 706
rect 3051 130 3085 706
rect 3169 130 3203 706
rect 3287 130 3321 706
rect 3405 130 3439 706
rect 3523 130 3557 706
rect 3641 130 3675 706
rect 3759 130 3793 706
rect 3877 130 3911 706
rect 3995 130 4029 706
rect 4113 130 4147 706
rect 4231 130 4265 706
rect 4349 130 4383 706
rect 4467 130 4501 706
rect 4585 130 4619 706
rect 4703 130 4737 706
rect 4821 130 4855 706
rect 4939 130 4973 706
rect 5057 130 5091 706
rect 5175 130 5209 706
rect 5293 130 5327 706
rect 5411 130 5445 706
rect 5529 130 5563 706
rect 5647 130 5681 706
rect 5765 130 5799 706
rect 5883 130 5917 706
rect 6001 130 6035 706
rect 6119 130 6153 706
rect 6237 130 6271 706
rect 6355 130 6389 706
rect 6473 130 6507 706
rect 6591 130 6625 706
rect 6709 130 6743 706
rect 6827 130 6861 706
rect 6945 130 6979 706
rect 7063 130 7097 706
rect -7038 37 -7004 71
rect -6920 37 -6886 71
rect -6802 37 -6768 71
rect -6684 37 -6650 71
rect -6566 37 -6532 71
rect -6448 37 -6414 71
rect -6330 37 -6296 71
rect -6212 37 -6178 71
rect -6094 37 -6060 71
rect -5976 37 -5942 71
rect -5858 37 -5824 71
rect -5740 37 -5706 71
rect -5622 37 -5588 71
rect -5504 37 -5470 71
rect -5386 37 -5352 71
rect -5268 37 -5234 71
rect -5150 37 -5116 71
rect -5032 37 -4998 71
rect -4914 37 -4880 71
rect -4796 37 -4762 71
rect -4678 37 -4644 71
rect -4560 37 -4526 71
rect -4442 37 -4408 71
rect -4324 37 -4290 71
rect -4206 37 -4172 71
rect -4088 37 -4054 71
rect -3970 37 -3936 71
rect -3852 37 -3818 71
rect -3734 37 -3700 71
rect -3616 37 -3582 71
rect -3498 37 -3464 71
rect -3380 37 -3346 71
rect -3262 37 -3228 71
rect -3144 37 -3110 71
rect -3026 37 -2992 71
rect -2908 37 -2874 71
rect -2790 37 -2756 71
rect -2672 37 -2638 71
rect -2554 37 -2520 71
rect -2436 37 -2402 71
rect -2318 37 -2284 71
rect -2200 37 -2166 71
rect -2082 37 -2048 71
rect -1964 37 -1930 71
rect -1846 37 -1812 71
rect -1728 37 -1694 71
rect -1610 37 -1576 71
rect -1492 37 -1458 71
rect -1374 37 -1340 71
rect -1256 37 -1222 71
rect -1138 37 -1104 71
rect -1020 37 -986 71
rect -902 37 -868 71
rect -784 37 -750 71
rect -666 37 -632 71
rect -548 37 -514 71
rect -430 37 -396 71
rect -312 37 -278 71
rect -194 37 -160 71
rect -76 37 -42 71
rect 42 37 76 71
rect 160 37 194 71
rect 278 37 312 71
rect 396 37 430 71
rect 514 37 548 71
rect 632 37 666 71
rect 750 37 784 71
rect 868 37 902 71
rect 986 37 1020 71
rect 1104 37 1138 71
rect 1222 37 1256 71
rect 1340 37 1374 71
rect 1458 37 1492 71
rect 1576 37 1610 71
rect 1694 37 1728 71
rect 1812 37 1846 71
rect 1930 37 1964 71
rect 2048 37 2082 71
rect 2166 37 2200 71
rect 2284 37 2318 71
rect 2402 37 2436 71
rect 2520 37 2554 71
rect 2638 37 2672 71
rect 2756 37 2790 71
rect 2874 37 2908 71
rect 2992 37 3026 71
rect 3110 37 3144 71
rect 3228 37 3262 71
rect 3346 37 3380 71
rect 3464 37 3498 71
rect 3582 37 3616 71
rect 3700 37 3734 71
rect 3818 37 3852 71
rect 3936 37 3970 71
rect 4054 37 4088 71
rect 4172 37 4206 71
rect 4290 37 4324 71
rect 4408 37 4442 71
rect 4526 37 4560 71
rect 4644 37 4678 71
rect 4762 37 4796 71
rect 4880 37 4914 71
rect 4998 37 5032 71
rect 5116 37 5150 71
rect 5234 37 5268 71
rect 5352 37 5386 71
rect 5470 37 5504 71
rect 5588 37 5622 71
rect 5706 37 5740 71
rect 5824 37 5858 71
rect 5942 37 5976 71
rect 6060 37 6094 71
rect 6178 37 6212 71
rect 6296 37 6330 71
rect 6414 37 6448 71
rect 6532 37 6566 71
rect 6650 37 6684 71
rect 6768 37 6802 71
rect 6886 37 6920 71
rect 7004 37 7038 71
rect -7038 -71 -7004 -37
rect -6920 -71 -6886 -37
rect -6802 -71 -6768 -37
rect -6684 -71 -6650 -37
rect -6566 -71 -6532 -37
rect -6448 -71 -6414 -37
rect -6330 -71 -6296 -37
rect -6212 -71 -6178 -37
rect -6094 -71 -6060 -37
rect -5976 -71 -5942 -37
rect -5858 -71 -5824 -37
rect -5740 -71 -5706 -37
rect -5622 -71 -5588 -37
rect -5504 -71 -5470 -37
rect -5386 -71 -5352 -37
rect -5268 -71 -5234 -37
rect -5150 -71 -5116 -37
rect -5032 -71 -4998 -37
rect -4914 -71 -4880 -37
rect -4796 -71 -4762 -37
rect -4678 -71 -4644 -37
rect -4560 -71 -4526 -37
rect -4442 -71 -4408 -37
rect -4324 -71 -4290 -37
rect -4206 -71 -4172 -37
rect -4088 -71 -4054 -37
rect -3970 -71 -3936 -37
rect -3852 -71 -3818 -37
rect -3734 -71 -3700 -37
rect -3616 -71 -3582 -37
rect -3498 -71 -3464 -37
rect -3380 -71 -3346 -37
rect -3262 -71 -3228 -37
rect -3144 -71 -3110 -37
rect -3026 -71 -2992 -37
rect -2908 -71 -2874 -37
rect -2790 -71 -2756 -37
rect -2672 -71 -2638 -37
rect -2554 -71 -2520 -37
rect -2436 -71 -2402 -37
rect -2318 -71 -2284 -37
rect -2200 -71 -2166 -37
rect -2082 -71 -2048 -37
rect -1964 -71 -1930 -37
rect -1846 -71 -1812 -37
rect -1728 -71 -1694 -37
rect -1610 -71 -1576 -37
rect -1492 -71 -1458 -37
rect -1374 -71 -1340 -37
rect -1256 -71 -1222 -37
rect -1138 -71 -1104 -37
rect -1020 -71 -986 -37
rect -902 -71 -868 -37
rect -784 -71 -750 -37
rect -666 -71 -632 -37
rect -548 -71 -514 -37
rect -430 -71 -396 -37
rect -312 -71 -278 -37
rect -194 -71 -160 -37
rect -76 -71 -42 -37
rect 42 -71 76 -37
rect 160 -71 194 -37
rect 278 -71 312 -37
rect 396 -71 430 -37
rect 514 -71 548 -37
rect 632 -71 666 -37
rect 750 -71 784 -37
rect 868 -71 902 -37
rect 986 -71 1020 -37
rect 1104 -71 1138 -37
rect 1222 -71 1256 -37
rect 1340 -71 1374 -37
rect 1458 -71 1492 -37
rect 1576 -71 1610 -37
rect 1694 -71 1728 -37
rect 1812 -71 1846 -37
rect 1930 -71 1964 -37
rect 2048 -71 2082 -37
rect 2166 -71 2200 -37
rect 2284 -71 2318 -37
rect 2402 -71 2436 -37
rect 2520 -71 2554 -37
rect 2638 -71 2672 -37
rect 2756 -71 2790 -37
rect 2874 -71 2908 -37
rect 2992 -71 3026 -37
rect 3110 -71 3144 -37
rect 3228 -71 3262 -37
rect 3346 -71 3380 -37
rect 3464 -71 3498 -37
rect 3582 -71 3616 -37
rect 3700 -71 3734 -37
rect 3818 -71 3852 -37
rect 3936 -71 3970 -37
rect 4054 -71 4088 -37
rect 4172 -71 4206 -37
rect 4290 -71 4324 -37
rect 4408 -71 4442 -37
rect 4526 -71 4560 -37
rect 4644 -71 4678 -37
rect 4762 -71 4796 -37
rect 4880 -71 4914 -37
rect 4998 -71 5032 -37
rect 5116 -71 5150 -37
rect 5234 -71 5268 -37
rect 5352 -71 5386 -37
rect 5470 -71 5504 -37
rect 5588 -71 5622 -37
rect 5706 -71 5740 -37
rect 5824 -71 5858 -37
rect 5942 -71 5976 -37
rect 6060 -71 6094 -37
rect 6178 -71 6212 -37
rect 6296 -71 6330 -37
rect 6414 -71 6448 -37
rect 6532 -71 6566 -37
rect 6650 -71 6684 -37
rect 6768 -71 6802 -37
rect 6886 -71 6920 -37
rect 7004 -71 7038 -37
rect -7097 -706 -7063 -130
rect -6979 -706 -6945 -130
rect -6861 -706 -6827 -130
rect -6743 -706 -6709 -130
rect -6625 -706 -6591 -130
rect -6507 -706 -6473 -130
rect -6389 -706 -6355 -130
rect -6271 -706 -6237 -130
rect -6153 -706 -6119 -130
rect -6035 -706 -6001 -130
rect -5917 -706 -5883 -130
rect -5799 -706 -5765 -130
rect -5681 -706 -5647 -130
rect -5563 -706 -5529 -130
rect -5445 -706 -5411 -130
rect -5327 -706 -5293 -130
rect -5209 -706 -5175 -130
rect -5091 -706 -5057 -130
rect -4973 -706 -4939 -130
rect -4855 -706 -4821 -130
rect -4737 -706 -4703 -130
rect -4619 -706 -4585 -130
rect -4501 -706 -4467 -130
rect -4383 -706 -4349 -130
rect -4265 -706 -4231 -130
rect -4147 -706 -4113 -130
rect -4029 -706 -3995 -130
rect -3911 -706 -3877 -130
rect -3793 -706 -3759 -130
rect -3675 -706 -3641 -130
rect -3557 -706 -3523 -130
rect -3439 -706 -3405 -130
rect -3321 -706 -3287 -130
rect -3203 -706 -3169 -130
rect -3085 -706 -3051 -130
rect -2967 -706 -2933 -130
rect -2849 -706 -2815 -130
rect -2731 -706 -2697 -130
rect -2613 -706 -2579 -130
rect -2495 -706 -2461 -130
rect -2377 -706 -2343 -130
rect -2259 -706 -2225 -130
rect -2141 -706 -2107 -130
rect -2023 -706 -1989 -130
rect -1905 -706 -1871 -130
rect -1787 -706 -1753 -130
rect -1669 -706 -1635 -130
rect -1551 -706 -1517 -130
rect -1433 -706 -1399 -130
rect -1315 -706 -1281 -130
rect -1197 -706 -1163 -130
rect -1079 -706 -1045 -130
rect -961 -706 -927 -130
rect -843 -706 -809 -130
rect -725 -706 -691 -130
rect -607 -706 -573 -130
rect -489 -706 -455 -130
rect -371 -706 -337 -130
rect -253 -706 -219 -130
rect -135 -706 -101 -130
rect -17 -706 17 -130
rect 101 -706 135 -130
rect 219 -706 253 -130
rect 337 -706 371 -130
rect 455 -706 489 -130
rect 573 -706 607 -130
rect 691 -706 725 -130
rect 809 -706 843 -130
rect 927 -706 961 -130
rect 1045 -706 1079 -130
rect 1163 -706 1197 -130
rect 1281 -706 1315 -130
rect 1399 -706 1433 -130
rect 1517 -706 1551 -130
rect 1635 -706 1669 -130
rect 1753 -706 1787 -130
rect 1871 -706 1905 -130
rect 1989 -706 2023 -130
rect 2107 -706 2141 -130
rect 2225 -706 2259 -130
rect 2343 -706 2377 -130
rect 2461 -706 2495 -130
rect 2579 -706 2613 -130
rect 2697 -706 2731 -130
rect 2815 -706 2849 -130
rect 2933 -706 2967 -130
rect 3051 -706 3085 -130
rect 3169 -706 3203 -130
rect 3287 -706 3321 -130
rect 3405 -706 3439 -130
rect 3523 -706 3557 -130
rect 3641 -706 3675 -130
rect 3759 -706 3793 -130
rect 3877 -706 3911 -130
rect 3995 -706 4029 -130
rect 4113 -706 4147 -130
rect 4231 -706 4265 -130
rect 4349 -706 4383 -130
rect 4467 -706 4501 -130
rect 4585 -706 4619 -130
rect 4703 -706 4737 -130
rect 4821 -706 4855 -130
rect 4939 -706 4973 -130
rect 5057 -706 5091 -130
rect 5175 -706 5209 -130
rect 5293 -706 5327 -130
rect 5411 -706 5445 -130
rect 5529 -706 5563 -130
rect 5647 -706 5681 -130
rect 5765 -706 5799 -130
rect 5883 -706 5917 -130
rect 6001 -706 6035 -130
rect 6119 -706 6153 -130
rect 6237 -706 6271 -130
rect 6355 -706 6389 -130
rect 6473 -706 6507 -130
rect 6591 -706 6625 -130
rect 6709 -706 6743 -130
rect 6827 -706 6861 -130
rect 6945 -706 6979 -130
rect 7063 -706 7097 -130
rect -7038 -799 -7004 -765
rect -6920 -799 -6886 -765
rect -6802 -799 -6768 -765
rect -6684 -799 -6650 -765
rect -6566 -799 -6532 -765
rect -6448 -799 -6414 -765
rect -6330 -799 -6296 -765
rect -6212 -799 -6178 -765
rect -6094 -799 -6060 -765
rect -5976 -799 -5942 -765
rect -5858 -799 -5824 -765
rect -5740 -799 -5706 -765
rect -5622 -799 -5588 -765
rect -5504 -799 -5470 -765
rect -5386 -799 -5352 -765
rect -5268 -799 -5234 -765
rect -5150 -799 -5116 -765
rect -5032 -799 -4998 -765
rect -4914 -799 -4880 -765
rect -4796 -799 -4762 -765
rect -4678 -799 -4644 -765
rect -4560 -799 -4526 -765
rect -4442 -799 -4408 -765
rect -4324 -799 -4290 -765
rect -4206 -799 -4172 -765
rect -4088 -799 -4054 -765
rect -3970 -799 -3936 -765
rect -3852 -799 -3818 -765
rect -3734 -799 -3700 -765
rect -3616 -799 -3582 -765
rect -3498 -799 -3464 -765
rect -3380 -799 -3346 -765
rect -3262 -799 -3228 -765
rect -3144 -799 -3110 -765
rect -3026 -799 -2992 -765
rect -2908 -799 -2874 -765
rect -2790 -799 -2756 -765
rect -2672 -799 -2638 -765
rect -2554 -799 -2520 -765
rect -2436 -799 -2402 -765
rect -2318 -799 -2284 -765
rect -2200 -799 -2166 -765
rect -2082 -799 -2048 -765
rect -1964 -799 -1930 -765
rect -1846 -799 -1812 -765
rect -1728 -799 -1694 -765
rect -1610 -799 -1576 -765
rect -1492 -799 -1458 -765
rect -1374 -799 -1340 -765
rect -1256 -799 -1222 -765
rect -1138 -799 -1104 -765
rect -1020 -799 -986 -765
rect -902 -799 -868 -765
rect -784 -799 -750 -765
rect -666 -799 -632 -765
rect -548 -799 -514 -765
rect -430 -799 -396 -765
rect -312 -799 -278 -765
rect -194 -799 -160 -765
rect -76 -799 -42 -765
rect 42 -799 76 -765
rect 160 -799 194 -765
rect 278 -799 312 -765
rect 396 -799 430 -765
rect 514 -799 548 -765
rect 632 -799 666 -765
rect 750 -799 784 -765
rect 868 -799 902 -765
rect 986 -799 1020 -765
rect 1104 -799 1138 -765
rect 1222 -799 1256 -765
rect 1340 -799 1374 -765
rect 1458 -799 1492 -765
rect 1576 -799 1610 -765
rect 1694 -799 1728 -765
rect 1812 -799 1846 -765
rect 1930 -799 1964 -765
rect 2048 -799 2082 -765
rect 2166 -799 2200 -765
rect 2284 -799 2318 -765
rect 2402 -799 2436 -765
rect 2520 -799 2554 -765
rect 2638 -799 2672 -765
rect 2756 -799 2790 -765
rect 2874 -799 2908 -765
rect 2992 -799 3026 -765
rect 3110 -799 3144 -765
rect 3228 -799 3262 -765
rect 3346 -799 3380 -765
rect 3464 -799 3498 -765
rect 3582 -799 3616 -765
rect 3700 -799 3734 -765
rect 3818 -799 3852 -765
rect 3936 -799 3970 -765
rect 4054 -799 4088 -765
rect 4172 -799 4206 -765
rect 4290 -799 4324 -765
rect 4408 -799 4442 -765
rect 4526 -799 4560 -765
rect 4644 -799 4678 -765
rect 4762 -799 4796 -765
rect 4880 -799 4914 -765
rect 4998 -799 5032 -765
rect 5116 -799 5150 -765
rect 5234 -799 5268 -765
rect 5352 -799 5386 -765
rect 5470 -799 5504 -765
rect 5588 -799 5622 -765
rect 5706 -799 5740 -765
rect 5824 -799 5858 -765
rect 5942 -799 5976 -765
rect 6060 -799 6094 -765
rect 6178 -799 6212 -765
rect 6296 -799 6330 -765
rect 6414 -799 6448 -765
rect 6532 -799 6566 -765
rect 6650 -799 6684 -765
rect 6768 -799 6802 -765
rect 6886 -799 6920 -765
rect 7004 -799 7038 -765
<< metal1 >>
rect -7050 799 -6992 805
rect -7050 765 -7038 799
rect -7004 765 -6992 799
rect -7050 759 -6992 765
rect -6932 799 -6874 805
rect -6932 765 -6920 799
rect -6886 765 -6874 799
rect -6932 759 -6874 765
rect -6814 799 -6756 805
rect -6814 765 -6802 799
rect -6768 765 -6756 799
rect -6814 759 -6756 765
rect -6696 799 -6638 805
rect -6696 765 -6684 799
rect -6650 765 -6638 799
rect -6696 759 -6638 765
rect -6578 799 -6520 805
rect -6578 765 -6566 799
rect -6532 765 -6520 799
rect -6578 759 -6520 765
rect -6460 799 -6402 805
rect -6460 765 -6448 799
rect -6414 765 -6402 799
rect -6460 759 -6402 765
rect -6342 799 -6284 805
rect -6342 765 -6330 799
rect -6296 765 -6284 799
rect -6342 759 -6284 765
rect -6224 799 -6166 805
rect -6224 765 -6212 799
rect -6178 765 -6166 799
rect -6224 759 -6166 765
rect -6106 799 -6048 805
rect -6106 765 -6094 799
rect -6060 765 -6048 799
rect -6106 759 -6048 765
rect -5988 799 -5930 805
rect -5988 765 -5976 799
rect -5942 765 -5930 799
rect -5988 759 -5930 765
rect -5870 799 -5812 805
rect -5870 765 -5858 799
rect -5824 765 -5812 799
rect -5870 759 -5812 765
rect -5752 799 -5694 805
rect -5752 765 -5740 799
rect -5706 765 -5694 799
rect -5752 759 -5694 765
rect -5634 799 -5576 805
rect -5634 765 -5622 799
rect -5588 765 -5576 799
rect -5634 759 -5576 765
rect -5516 799 -5458 805
rect -5516 765 -5504 799
rect -5470 765 -5458 799
rect -5516 759 -5458 765
rect -5398 799 -5340 805
rect -5398 765 -5386 799
rect -5352 765 -5340 799
rect -5398 759 -5340 765
rect -5280 799 -5222 805
rect -5280 765 -5268 799
rect -5234 765 -5222 799
rect -5280 759 -5222 765
rect -5162 799 -5104 805
rect -5162 765 -5150 799
rect -5116 765 -5104 799
rect -5162 759 -5104 765
rect -5044 799 -4986 805
rect -5044 765 -5032 799
rect -4998 765 -4986 799
rect -5044 759 -4986 765
rect -4926 799 -4868 805
rect -4926 765 -4914 799
rect -4880 765 -4868 799
rect -4926 759 -4868 765
rect -4808 799 -4750 805
rect -4808 765 -4796 799
rect -4762 765 -4750 799
rect -4808 759 -4750 765
rect -4690 799 -4632 805
rect -4690 765 -4678 799
rect -4644 765 -4632 799
rect -4690 759 -4632 765
rect -4572 799 -4514 805
rect -4572 765 -4560 799
rect -4526 765 -4514 799
rect -4572 759 -4514 765
rect -4454 799 -4396 805
rect -4454 765 -4442 799
rect -4408 765 -4396 799
rect -4454 759 -4396 765
rect -4336 799 -4278 805
rect -4336 765 -4324 799
rect -4290 765 -4278 799
rect -4336 759 -4278 765
rect -4218 799 -4160 805
rect -4218 765 -4206 799
rect -4172 765 -4160 799
rect -4218 759 -4160 765
rect -4100 799 -4042 805
rect -4100 765 -4088 799
rect -4054 765 -4042 799
rect -4100 759 -4042 765
rect -3982 799 -3924 805
rect -3982 765 -3970 799
rect -3936 765 -3924 799
rect -3982 759 -3924 765
rect -3864 799 -3806 805
rect -3864 765 -3852 799
rect -3818 765 -3806 799
rect -3864 759 -3806 765
rect -3746 799 -3688 805
rect -3746 765 -3734 799
rect -3700 765 -3688 799
rect -3746 759 -3688 765
rect -3628 799 -3570 805
rect -3628 765 -3616 799
rect -3582 765 -3570 799
rect -3628 759 -3570 765
rect -3510 799 -3452 805
rect -3510 765 -3498 799
rect -3464 765 -3452 799
rect -3510 759 -3452 765
rect -3392 799 -3334 805
rect -3392 765 -3380 799
rect -3346 765 -3334 799
rect -3392 759 -3334 765
rect -3274 799 -3216 805
rect -3274 765 -3262 799
rect -3228 765 -3216 799
rect -3274 759 -3216 765
rect -3156 799 -3098 805
rect -3156 765 -3144 799
rect -3110 765 -3098 799
rect -3156 759 -3098 765
rect -3038 799 -2980 805
rect -3038 765 -3026 799
rect -2992 765 -2980 799
rect -3038 759 -2980 765
rect -2920 799 -2862 805
rect -2920 765 -2908 799
rect -2874 765 -2862 799
rect -2920 759 -2862 765
rect -2802 799 -2744 805
rect -2802 765 -2790 799
rect -2756 765 -2744 799
rect -2802 759 -2744 765
rect -2684 799 -2626 805
rect -2684 765 -2672 799
rect -2638 765 -2626 799
rect -2684 759 -2626 765
rect -2566 799 -2508 805
rect -2566 765 -2554 799
rect -2520 765 -2508 799
rect -2566 759 -2508 765
rect -2448 799 -2390 805
rect -2448 765 -2436 799
rect -2402 765 -2390 799
rect -2448 759 -2390 765
rect -2330 799 -2272 805
rect -2330 765 -2318 799
rect -2284 765 -2272 799
rect -2330 759 -2272 765
rect -2212 799 -2154 805
rect -2212 765 -2200 799
rect -2166 765 -2154 799
rect -2212 759 -2154 765
rect -2094 799 -2036 805
rect -2094 765 -2082 799
rect -2048 765 -2036 799
rect -2094 759 -2036 765
rect -1976 799 -1918 805
rect -1976 765 -1964 799
rect -1930 765 -1918 799
rect -1976 759 -1918 765
rect -1858 799 -1800 805
rect -1858 765 -1846 799
rect -1812 765 -1800 799
rect -1858 759 -1800 765
rect -1740 799 -1682 805
rect -1740 765 -1728 799
rect -1694 765 -1682 799
rect -1740 759 -1682 765
rect -1622 799 -1564 805
rect -1622 765 -1610 799
rect -1576 765 -1564 799
rect -1622 759 -1564 765
rect -1504 799 -1446 805
rect -1504 765 -1492 799
rect -1458 765 -1446 799
rect -1504 759 -1446 765
rect -1386 799 -1328 805
rect -1386 765 -1374 799
rect -1340 765 -1328 799
rect -1386 759 -1328 765
rect -1268 799 -1210 805
rect -1268 765 -1256 799
rect -1222 765 -1210 799
rect -1268 759 -1210 765
rect -1150 799 -1092 805
rect -1150 765 -1138 799
rect -1104 765 -1092 799
rect -1150 759 -1092 765
rect -1032 799 -974 805
rect -1032 765 -1020 799
rect -986 765 -974 799
rect -1032 759 -974 765
rect -914 799 -856 805
rect -914 765 -902 799
rect -868 765 -856 799
rect -914 759 -856 765
rect -796 799 -738 805
rect -796 765 -784 799
rect -750 765 -738 799
rect -796 759 -738 765
rect -678 799 -620 805
rect -678 765 -666 799
rect -632 765 -620 799
rect -678 759 -620 765
rect -560 799 -502 805
rect -560 765 -548 799
rect -514 765 -502 799
rect -560 759 -502 765
rect -442 799 -384 805
rect -442 765 -430 799
rect -396 765 -384 799
rect -442 759 -384 765
rect -324 799 -266 805
rect -324 765 -312 799
rect -278 765 -266 799
rect -324 759 -266 765
rect -206 799 -148 805
rect -206 765 -194 799
rect -160 765 -148 799
rect -206 759 -148 765
rect -88 799 -30 805
rect -88 765 -76 799
rect -42 765 -30 799
rect -88 759 -30 765
rect 30 799 88 805
rect 30 765 42 799
rect 76 765 88 799
rect 30 759 88 765
rect 148 799 206 805
rect 148 765 160 799
rect 194 765 206 799
rect 148 759 206 765
rect 266 799 324 805
rect 266 765 278 799
rect 312 765 324 799
rect 266 759 324 765
rect 384 799 442 805
rect 384 765 396 799
rect 430 765 442 799
rect 384 759 442 765
rect 502 799 560 805
rect 502 765 514 799
rect 548 765 560 799
rect 502 759 560 765
rect 620 799 678 805
rect 620 765 632 799
rect 666 765 678 799
rect 620 759 678 765
rect 738 799 796 805
rect 738 765 750 799
rect 784 765 796 799
rect 738 759 796 765
rect 856 799 914 805
rect 856 765 868 799
rect 902 765 914 799
rect 856 759 914 765
rect 974 799 1032 805
rect 974 765 986 799
rect 1020 765 1032 799
rect 974 759 1032 765
rect 1092 799 1150 805
rect 1092 765 1104 799
rect 1138 765 1150 799
rect 1092 759 1150 765
rect 1210 799 1268 805
rect 1210 765 1222 799
rect 1256 765 1268 799
rect 1210 759 1268 765
rect 1328 799 1386 805
rect 1328 765 1340 799
rect 1374 765 1386 799
rect 1328 759 1386 765
rect 1446 799 1504 805
rect 1446 765 1458 799
rect 1492 765 1504 799
rect 1446 759 1504 765
rect 1564 799 1622 805
rect 1564 765 1576 799
rect 1610 765 1622 799
rect 1564 759 1622 765
rect 1682 799 1740 805
rect 1682 765 1694 799
rect 1728 765 1740 799
rect 1682 759 1740 765
rect 1800 799 1858 805
rect 1800 765 1812 799
rect 1846 765 1858 799
rect 1800 759 1858 765
rect 1918 799 1976 805
rect 1918 765 1930 799
rect 1964 765 1976 799
rect 1918 759 1976 765
rect 2036 799 2094 805
rect 2036 765 2048 799
rect 2082 765 2094 799
rect 2036 759 2094 765
rect 2154 799 2212 805
rect 2154 765 2166 799
rect 2200 765 2212 799
rect 2154 759 2212 765
rect 2272 799 2330 805
rect 2272 765 2284 799
rect 2318 765 2330 799
rect 2272 759 2330 765
rect 2390 799 2448 805
rect 2390 765 2402 799
rect 2436 765 2448 799
rect 2390 759 2448 765
rect 2508 799 2566 805
rect 2508 765 2520 799
rect 2554 765 2566 799
rect 2508 759 2566 765
rect 2626 799 2684 805
rect 2626 765 2638 799
rect 2672 765 2684 799
rect 2626 759 2684 765
rect 2744 799 2802 805
rect 2744 765 2756 799
rect 2790 765 2802 799
rect 2744 759 2802 765
rect 2862 799 2920 805
rect 2862 765 2874 799
rect 2908 765 2920 799
rect 2862 759 2920 765
rect 2980 799 3038 805
rect 2980 765 2992 799
rect 3026 765 3038 799
rect 2980 759 3038 765
rect 3098 799 3156 805
rect 3098 765 3110 799
rect 3144 765 3156 799
rect 3098 759 3156 765
rect 3216 799 3274 805
rect 3216 765 3228 799
rect 3262 765 3274 799
rect 3216 759 3274 765
rect 3334 799 3392 805
rect 3334 765 3346 799
rect 3380 765 3392 799
rect 3334 759 3392 765
rect 3452 799 3510 805
rect 3452 765 3464 799
rect 3498 765 3510 799
rect 3452 759 3510 765
rect 3570 799 3628 805
rect 3570 765 3582 799
rect 3616 765 3628 799
rect 3570 759 3628 765
rect 3688 799 3746 805
rect 3688 765 3700 799
rect 3734 765 3746 799
rect 3688 759 3746 765
rect 3806 799 3864 805
rect 3806 765 3818 799
rect 3852 765 3864 799
rect 3806 759 3864 765
rect 3924 799 3982 805
rect 3924 765 3936 799
rect 3970 765 3982 799
rect 3924 759 3982 765
rect 4042 799 4100 805
rect 4042 765 4054 799
rect 4088 765 4100 799
rect 4042 759 4100 765
rect 4160 799 4218 805
rect 4160 765 4172 799
rect 4206 765 4218 799
rect 4160 759 4218 765
rect 4278 799 4336 805
rect 4278 765 4290 799
rect 4324 765 4336 799
rect 4278 759 4336 765
rect 4396 799 4454 805
rect 4396 765 4408 799
rect 4442 765 4454 799
rect 4396 759 4454 765
rect 4514 799 4572 805
rect 4514 765 4526 799
rect 4560 765 4572 799
rect 4514 759 4572 765
rect 4632 799 4690 805
rect 4632 765 4644 799
rect 4678 765 4690 799
rect 4632 759 4690 765
rect 4750 799 4808 805
rect 4750 765 4762 799
rect 4796 765 4808 799
rect 4750 759 4808 765
rect 4868 799 4926 805
rect 4868 765 4880 799
rect 4914 765 4926 799
rect 4868 759 4926 765
rect 4986 799 5044 805
rect 4986 765 4998 799
rect 5032 765 5044 799
rect 4986 759 5044 765
rect 5104 799 5162 805
rect 5104 765 5116 799
rect 5150 765 5162 799
rect 5104 759 5162 765
rect 5222 799 5280 805
rect 5222 765 5234 799
rect 5268 765 5280 799
rect 5222 759 5280 765
rect 5340 799 5398 805
rect 5340 765 5352 799
rect 5386 765 5398 799
rect 5340 759 5398 765
rect 5458 799 5516 805
rect 5458 765 5470 799
rect 5504 765 5516 799
rect 5458 759 5516 765
rect 5576 799 5634 805
rect 5576 765 5588 799
rect 5622 765 5634 799
rect 5576 759 5634 765
rect 5694 799 5752 805
rect 5694 765 5706 799
rect 5740 765 5752 799
rect 5694 759 5752 765
rect 5812 799 5870 805
rect 5812 765 5824 799
rect 5858 765 5870 799
rect 5812 759 5870 765
rect 5930 799 5988 805
rect 5930 765 5942 799
rect 5976 765 5988 799
rect 5930 759 5988 765
rect 6048 799 6106 805
rect 6048 765 6060 799
rect 6094 765 6106 799
rect 6048 759 6106 765
rect 6166 799 6224 805
rect 6166 765 6178 799
rect 6212 765 6224 799
rect 6166 759 6224 765
rect 6284 799 6342 805
rect 6284 765 6296 799
rect 6330 765 6342 799
rect 6284 759 6342 765
rect 6402 799 6460 805
rect 6402 765 6414 799
rect 6448 765 6460 799
rect 6402 759 6460 765
rect 6520 799 6578 805
rect 6520 765 6532 799
rect 6566 765 6578 799
rect 6520 759 6578 765
rect 6638 799 6696 805
rect 6638 765 6650 799
rect 6684 765 6696 799
rect 6638 759 6696 765
rect 6756 799 6814 805
rect 6756 765 6768 799
rect 6802 765 6814 799
rect 6756 759 6814 765
rect 6874 799 6932 805
rect 6874 765 6886 799
rect 6920 765 6932 799
rect 6874 759 6932 765
rect 6992 799 7050 805
rect 6992 765 7004 799
rect 7038 765 7050 799
rect 6992 759 7050 765
rect -7103 706 -7057 718
rect -7103 130 -7097 706
rect -7063 130 -7057 706
rect -7103 118 -7057 130
rect -6985 706 -6939 718
rect -6985 130 -6979 706
rect -6945 130 -6939 706
rect -6985 118 -6939 130
rect -6867 706 -6821 718
rect -6867 130 -6861 706
rect -6827 130 -6821 706
rect -6867 118 -6821 130
rect -6749 706 -6703 718
rect -6749 130 -6743 706
rect -6709 130 -6703 706
rect -6749 118 -6703 130
rect -6631 706 -6585 718
rect -6631 130 -6625 706
rect -6591 130 -6585 706
rect -6631 118 -6585 130
rect -6513 706 -6467 718
rect -6513 130 -6507 706
rect -6473 130 -6467 706
rect -6513 118 -6467 130
rect -6395 706 -6349 718
rect -6395 130 -6389 706
rect -6355 130 -6349 706
rect -6395 118 -6349 130
rect -6277 706 -6231 718
rect -6277 130 -6271 706
rect -6237 130 -6231 706
rect -6277 118 -6231 130
rect -6159 706 -6113 718
rect -6159 130 -6153 706
rect -6119 130 -6113 706
rect -6159 118 -6113 130
rect -6041 706 -5995 718
rect -6041 130 -6035 706
rect -6001 130 -5995 706
rect -6041 118 -5995 130
rect -5923 706 -5877 718
rect -5923 130 -5917 706
rect -5883 130 -5877 706
rect -5923 118 -5877 130
rect -5805 706 -5759 718
rect -5805 130 -5799 706
rect -5765 130 -5759 706
rect -5805 118 -5759 130
rect -5687 706 -5641 718
rect -5687 130 -5681 706
rect -5647 130 -5641 706
rect -5687 118 -5641 130
rect -5569 706 -5523 718
rect -5569 130 -5563 706
rect -5529 130 -5523 706
rect -5569 118 -5523 130
rect -5451 706 -5405 718
rect -5451 130 -5445 706
rect -5411 130 -5405 706
rect -5451 118 -5405 130
rect -5333 706 -5287 718
rect -5333 130 -5327 706
rect -5293 130 -5287 706
rect -5333 118 -5287 130
rect -5215 706 -5169 718
rect -5215 130 -5209 706
rect -5175 130 -5169 706
rect -5215 118 -5169 130
rect -5097 706 -5051 718
rect -5097 130 -5091 706
rect -5057 130 -5051 706
rect -5097 118 -5051 130
rect -4979 706 -4933 718
rect -4979 130 -4973 706
rect -4939 130 -4933 706
rect -4979 118 -4933 130
rect -4861 706 -4815 718
rect -4861 130 -4855 706
rect -4821 130 -4815 706
rect -4861 118 -4815 130
rect -4743 706 -4697 718
rect -4743 130 -4737 706
rect -4703 130 -4697 706
rect -4743 118 -4697 130
rect -4625 706 -4579 718
rect -4625 130 -4619 706
rect -4585 130 -4579 706
rect -4625 118 -4579 130
rect -4507 706 -4461 718
rect -4507 130 -4501 706
rect -4467 130 -4461 706
rect -4507 118 -4461 130
rect -4389 706 -4343 718
rect -4389 130 -4383 706
rect -4349 130 -4343 706
rect -4389 118 -4343 130
rect -4271 706 -4225 718
rect -4271 130 -4265 706
rect -4231 130 -4225 706
rect -4271 118 -4225 130
rect -4153 706 -4107 718
rect -4153 130 -4147 706
rect -4113 130 -4107 706
rect -4153 118 -4107 130
rect -4035 706 -3989 718
rect -4035 130 -4029 706
rect -3995 130 -3989 706
rect -4035 118 -3989 130
rect -3917 706 -3871 718
rect -3917 130 -3911 706
rect -3877 130 -3871 706
rect -3917 118 -3871 130
rect -3799 706 -3753 718
rect -3799 130 -3793 706
rect -3759 130 -3753 706
rect -3799 118 -3753 130
rect -3681 706 -3635 718
rect -3681 130 -3675 706
rect -3641 130 -3635 706
rect -3681 118 -3635 130
rect -3563 706 -3517 718
rect -3563 130 -3557 706
rect -3523 130 -3517 706
rect -3563 118 -3517 130
rect -3445 706 -3399 718
rect -3445 130 -3439 706
rect -3405 130 -3399 706
rect -3445 118 -3399 130
rect -3327 706 -3281 718
rect -3327 130 -3321 706
rect -3287 130 -3281 706
rect -3327 118 -3281 130
rect -3209 706 -3163 718
rect -3209 130 -3203 706
rect -3169 130 -3163 706
rect -3209 118 -3163 130
rect -3091 706 -3045 718
rect -3091 130 -3085 706
rect -3051 130 -3045 706
rect -3091 118 -3045 130
rect -2973 706 -2927 718
rect -2973 130 -2967 706
rect -2933 130 -2927 706
rect -2973 118 -2927 130
rect -2855 706 -2809 718
rect -2855 130 -2849 706
rect -2815 130 -2809 706
rect -2855 118 -2809 130
rect -2737 706 -2691 718
rect -2737 130 -2731 706
rect -2697 130 -2691 706
rect -2737 118 -2691 130
rect -2619 706 -2573 718
rect -2619 130 -2613 706
rect -2579 130 -2573 706
rect -2619 118 -2573 130
rect -2501 706 -2455 718
rect -2501 130 -2495 706
rect -2461 130 -2455 706
rect -2501 118 -2455 130
rect -2383 706 -2337 718
rect -2383 130 -2377 706
rect -2343 130 -2337 706
rect -2383 118 -2337 130
rect -2265 706 -2219 718
rect -2265 130 -2259 706
rect -2225 130 -2219 706
rect -2265 118 -2219 130
rect -2147 706 -2101 718
rect -2147 130 -2141 706
rect -2107 130 -2101 706
rect -2147 118 -2101 130
rect -2029 706 -1983 718
rect -2029 130 -2023 706
rect -1989 130 -1983 706
rect -2029 118 -1983 130
rect -1911 706 -1865 718
rect -1911 130 -1905 706
rect -1871 130 -1865 706
rect -1911 118 -1865 130
rect -1793 706 -1747 718
rect -1793 130 -1787 706
rect -1753 130 -1747 706
rect -1793 118 -1747 130
rect -1675 706 -1629 718
rect -1675 130 -1669 706
rect -1635 130 -1629 706
rect -1675 118 -1629 130
rect -1557 706 -1511 718
rect -1557 130 -1551 706
rect -1517 130 -1511 706
rect -1557 118 -1511 130
rect -1439 706 -1393 718
rect -1439 130 -1433 706
rect -1399 130 -1393 706
rect -1439 118 -1393 130
rect -1321 706 -1275 718
rect -1321 130 -1315 706
rect -1281 130 -1275 706
rect -1321 118 -1275 130
rect -1203 706 -1157 718
rect -1203 130 -1197 706
rect -1163 130 -1157 706
rect -1203 118 -1157 130
rect -1085 706 -1039 718
rect -1085 130 -1079 706
rect -1045 130 -1039 706
rect -1085 118 -1039 130
rect -967 706 -921 718
rect -967 130 -961 706
rect -927 130 -921 706
rect -967 118 -921 130
rect -849 706 -803 718
rect -849 130 -843 706
rect -809 130 -803 706
rect -849 118 -803 130
rect -731 706 -685 718
rect -731 130 -725 706
rect -691 130 -685 706
rect -731 118 -685 130
rect -613 706 -567 718
rect -613 130 -607 706
rect -573 130 -567 706
rect -613 118 -567 130
rect -495 706 -449 718
rect -495 130 -489 706
rect -455 130 -449 706
rect -495 118 -449 130
rect -377 706 -331 718
rect -377 130 -371 706
rect -337 130 -331 706
rect -377 118 -331 130
rect -259 706 -213 718
rect -259 130 -253 706
rect -219 130 -213 706
rect -259 118 -213 130
rect -141 706 -95 718
rect -141 130 -135 706
rect -101 130 -95 706
rect -141 118 -95 130
rect -23 706 23 718
rect -23 130 -17 706
rect 17 130 23 706
rect -23 118 23 130
rect 95 706 141 718
rect 95 130 101 706
rect 135 130 141 706
rect 95 118 141 130
rect 213 706 259 718
rect 213 130 219 706
rect 253 130 259 706
rect 213 118 259 130
rect 331 706 377 718
rect 331 130 337 706
rect 371 130 377 706
rect 331 118 377 130
rect 449 706 495 718
rect 449 130 455 706
rect 489 130 495 706
rect 449 118 495 130
rect 567 706 613 718
rect 567 130 573 706
rect 607 130 613 706
rect 567 118 613 130
rect 685 706 731 718
rect 685 130 691 706
rect 725 130 731 706
rect 685 118 731 130
rect 803 706 849 718
rect 803 130 809 706
rect 843 130 849 706
rect 803 118 849 130
rect 921 706 967 718
rect 921 130 927 706
rect 961 130 967 706
rect 921 118 967 130
rect 1039 706 1085 718
rect 1039 130 1045 706
rect 1079 130 1085 706
rect 1039 118 1085 130
rect 1157 706 1203 718
rect 1157 130 1163 706
rect 1197 130 1203 706
rect 1157 118 1203 130
rect 1275 706 1321 718
rect 1275 130 1281 706
rect 1315 130 1321 706
rect 1275 118 1321 130
rect 1393 706 1439 718
rect 1393 130 1399 706
rect 1433 130 1439 706
rect 1393 118 1439 130
rect 1511 706 1557 718
rect 1511 130 1517 706
rect 1551 130 1557 706
rect 1511 118 1557 130
rect 1629 706 1675 718
rect 1629 130 1635 706
rect 1669 130 1675 706
rect 1629 118 1675 130
rect 1747 706 1793 718
rect 1747 130 1753 706
rect 1787 130 1793 706
rect 1747 118 1793 130
rect 1865 706 1911 718
rect 1865 130 1871 706
rect 1905 130 1911 706
rect 1865 118 1911 130
rect 1983 706 2029 718
rect 1983 130 1989 706
rect 2023 130 2029 706
rect 1983 118 2029 130
rect 2101 706 2147 718
rect 2101 130 2107 706
rect 2141 130 2147 706
rect 2101 118 2147 130
rect 2219 706 2265 718
rect 2219 130 2225 706
rect 2259 130 2265 706
rect 2219 118 2265 130
rect 2337 706 2383 718
rect 2337 130 2343 706
rect 2377 130 2383 706
rect 2337 118 2383 130
rect 2455 706 2501 718
rect 2455 130 2461 706
rect 2495 130 2501 706
rect 2455 118 2501 130
rect 2573 706 2619 718
rect 2573 130 2579 706
rect 2613 130 2619 706
rect 2573 118 2619 130
rect 2691 706 2737 718
rect 2691 130 2697 706
rect 2731 130 2737 706
rect 2691 118 2737 130
rect 2809 706 2855 718
rect 2809 130 2815 706
rect 2849 130 2855 706
rect 2809 118 2855 130
rect 2927 706 2973 718
rect 2927 130 2933 706
rect 2967 130 2973 706
rect 2927 118 2973 130
rect 3045 706 3091 718
rect 3045 130 3051 706
rect 3085 130 3091 706
rect 3045 118 3091 130
rect 3163 706 3209 718
rect 3163 130 3169 706
rect 3203 130 3209 706
rect 3163 118 3209 130
rect 3281 706 3327 718
rect 3281 130 3287 706
rect 3321 130 3327 706
rect 3281 118 3327 130
rect 3399 706 3445 718
rect 3399 130 3405 706
rect 3439 130 3445 706
rect 3399 118 3445 130
rect 3517 706 3563 718
rect 3517 130 3523 706
rect 3557 130 3563 706
rect 3517 118 3563 130
rect 3635 706 3681 718
rect 3635 130 3641 706
rect 3675 130 3681 706
rect 3635 118 3681 130
rect 3753 706 3799 718
rect 3753 130 3759 706
rect 3793 130 3799 706
rect 3753 118 3799 130
rect 3871 706 3917 718
rect 3871 130 3877 706
rect 3911 130 3917 706
rect 3871 118 3917 130
rect 3989 706 4035 718
rect 3989 130 3995 706
rect 4029 130 4035 706
rect 3989 118 4035 130
rect 4107 706 4153 718
rect 4107 130 4113 706
rect 4147 130 4153 706
rect 4107 118 4153 130
rect 4225 706 4271 718
rect 4225 130 4231 706
rect 4265 130 4271 706
rect 4225 118 4271 130
rect 4343 706 4389 718
rect 4343 130 4349 706
rect 4383 130 4389 706
rect 4343 118 4389 130
rect 4461 706 4507 718
rect 4461 130 4467 706
rect 4501 130 4507 706
rect 4461 118 4507 130
rect 4579 706 4625 718
rect 4579 130 4585 706
rect 4619 130 4625 706
rect 4579 118 4625 130
rect 4697 706 4743 718
rect 4697 130 4703 706
rect 4737 130 4743 706
rect 4697 118 4743 130
rect 4815 706 4861 718
rect 4815 130 4821 706
rect 4855 130 4861 706
rect 4815 118 4861 130
rect 4933 706 4979 718
rect 4933 130 4939 706
rect 4973 130 4979 706
rect 4933 118 4979 130
rect 5051 706 5097 718
rect 5051 130 5057 706
rect 5091 130 5097 706
rect 5051 118 5097 130
rect 5169 706 5215 718
rect 5169 130 5175 706
rect 5209 130 5215 706
rect 5169 118 5215 130
rect 5287 706 5333 718
rect 5287 130 5293 706
rect 5327 130 5333 706
rect 5287 118 5333 130
rect 5405 706 5451 718
rect 5405 130 5411 706
rect 5445 130 5451 706
rect 5405 118 5451 130
rect 5523 706 5569 718
rect 5523 130 5529 706
rect 5563 130 5569 706
rect 5523 118 5569 130
rect 5641 706 5687 718
rect 5641 130 5647 706
rect 5681 130 5687 706
rect 5641 118 5687 130
rect 5759 706 5805 718
rect 5759 130 5765 706
rect 5799 130 5805 706
rect 5759 118 5805 130
rect 5877 706 5923 718
rect 5877 130 5883 706
rect 5917 130 5923 706
rect 5877 118 5923 130
rect 5995 706 6041 718
rect 5995 130 6001 706
rect 6035 130 6041 706
rect 5995 118 6041 130
rect 6113 706 6159 718
rect 6113 130 6119 706
rect 6153 130 6159 706
rect 6113 118 6159 130
rect 6231 706 6277 718
rect 6231 130 6237 706
rect 6271 130 6277 706
rect 6231 118 6277 130
rect 6349 706 6395 718
rect 6349 130 6355 706
rect 6389 130 6395 706
rect 6349 118 6395 130
rect 6467 706 6513 718
rect 6467 130 6473 706
rect 6507 130 6513 706
rect 6467 118 6513 130
rect 6585 706 6631 718
rect 6585 130 6591 706
rect 6625 130 6631 706
rect 6585 118 6631 130
rect 6703 706 6749 718
rect 6703 130 6709 706
rect 6743 130 6749 706
rect 6703 118 6749 130
rect 6821 706 6867 718
rect 6821 130 6827 706
rect 6861 130 6867 706
rect 6821 118 6867 130
rect 6939 706 6985 718
rect 6939 130 6945 706
rect 6979 130 6985 706
rect 6939 118 6985 130
rect 7057 706 7103 718
rect 7057 130 7063 706
rect 7097 130 7103 706
rect 7057 118 7103 130
rect -7050 71 -6992 77
rect -7050 37 -7038 71
rect -7004 37 -6992 71
rect -7050 31 -6992 37
rect -6932 71 -6874 77
rect -6932 37 -6920 71
rect -6886 37 -6874 71
rect -6932 31 -6874 37
rect -6814 71 -6756 77
rect -6814 37 -6802 71
rect -6768 37 -6756 71
rect -6814 31 -6756 37
rect -6696 71 -6638 77
rect -6696 37 -6684 71
rect -6650 37 -6638 71
rect -6696 31 -6638 37
rect -6578 71 -6520 77
rect -6578 37 -6566 71
rect -6532 37 -6520 71
rect -6578 31 -6520 37
rect -6460 71 -6402 77
rect -6460 37 -6448 71
rect -6414 37 -6402 71
rect -6460 31 -6402 37
rect -6342 71 -6284 77
rect -6342 37 -6330 71
rect -6296 37 -6284 71
rect -6342 31 -6284 37
rect -6224 71 -6166 77
rect -6224 37 -6212 71
rect -6178 37 -6166 71
rect -6224 31 -6166 37
rect -6106 71 -6048 77
rect -6106 37 -6094 71
rect -6060 37 -6048 71
rect -6106 31 -6048 37
rect -5988 71 -5930 77
rect -5988 37 -5976 71
rect -5942 37 -5930 71
rect -5988 31 -5930 37
rect -5870 71 -5812 77
rect -5870 37 -5858 71
rect -5824 37 -5812 71
rect -5870 31 -5812 37
rect -5752 71 -5694 77
rect -5752 37 -5740 71
rect -5706 37 -5694 71
rect -5752 31 -5694 37
rect -5634 71 -5576 77
rect -5634 37 -5622 71
rect -5588 37 -5576 71
rect -5634 31 -5576 37
rect -5516 71 -5458 77
rect -5516 37 -5504 71
rect -5470 37 -5458 71
rect -5516 31 -5458 37
rect -5398 71 -5340 77
rect -5398 37 -5386 71
rect -5352 37 -5340 71
rect -5398 31 -5340 37
rect -5280 71 -5222 77
rect -5280 37 -5268 71
rect -5234 37 -5222 71
rect -5280 31 -5222 37
rect -5162 71 -5104 77
rect -5162 37 -5150 71
rect -5116 37 -5104 71
rect -5162 31 -5104 37
rect -5044 71 -4986 77
rect -5044 37 -5032 71
rect -4998 37 -4986 71
rect -5044 31 -4986 37
rect -4926 71 -4868 77
rect -4926 37 -4914 71
rect -4880 37 -4868 71
rect -4926 31 -4868 37
rect -4808 71 -4750 77
rect -4808 37 -4796 71
rect -4762 37 -4750 71
rect -4808 31 -4750 37
rect -4690 71 -4632 77
rect -4690 37 -4678 71
rect -4644 37 -4632 71
rect -4690 31 -4632 37
rect -4572 71 -4514 77
rect -4572 37 -4560 71
rect -4526 37 -4514 71
rect -4572 31 -4514 37
rect -4454 71 -4396 77
rect -4454 37 -4442 71
rect -4408 37 -4396 71
rect -4454 31 -4396 37
rect -4336 71 -4278 77
rect -4336 37 -4324 71
rect -4290 37 -4278 71
rect -4336 31 -4278 37
rect -4218 71 -4160 77
rect -4218 37 -4206 71
rect -4172 37 -4160 71
rect -4218 31 -4160 37
rect -4100 71 -4042 77
rect -4100 37 -4088 71
rect -4054 37 -4042 71
rect -4100 31 -4042 37
rect -3982 71 -3924 77
rect -3982 37 -3970 71
rect -3936 37 -3924 71
rect -3982 31 -3924 37
rect -3864 71 -3806 77
rect -3864 37 -3852 71
rect -3818 37 -3806 71
rect -3864 31 -3806 37
rect -3746 71 -3688 77
rect -3746 37 -3734 71
rect -3700 37 -3688 71
rect -3746 31 -3688 37
rect -3628 71 -3570 77
rect -3628 37 -3616 71
rect -3582 37 -3570 71
rect -3628 31 -3570 37
rect -3510 71 -3452 77
rect -3510 37 -3498 71
rect -3464 37 -3452 71
rect -3510 31 -3452 37
rect -3392 71 -3334 77
rect -3392 37 -3380 71
rect -3346 37 -3334 71
rect -3392 31 -3334 37
rect -3274 71 -3216 77
rect -3274 37 -3262 71
rect -3228 37 -3216 71
rect -3274 31 -3216 37
rect -3156 71 -3098 77
rect -3156 37 -3144 71
rect -3110 37 -3098 71
rect -3156 31 -3098 37
rect -3038 71 -2980 77
rect -3038 37 -3026 71
rect -2992 37 -2980 71
rect -3038 31 -2980 37
rect -2920 71 -2862 77
rect -2920 37 -2908 71
rect -2874 37 -2862 71
rect -2920 31 -2862 37
rect -2802 71 -2744 77
rect -2802 37 -2790 71
rect -2756 37 -2744 71
rect -2802 31 -2744 37
rect -2684 71 -2626 77
rect -2684 37 -2672 71
rect -2638 37 -2626 71
rect -2684 31 -2626 37
rect -2566 71 -2508 77
rect -2566 37 -2554 71
rect -2520 37 -2508 71
rect -2566 31 -2508 37
rect -2448 71 -2390 77
rect -2448 37 -2436 71
rect -2402 37 -2390 71
rect -2448 31 -2390 37
rect -2330 71 -2272 77
rect -2330 37 -2318 71
rect -2284 37 -2272 71
rect -2330 31 -2272 37
rect -2212 71 -2154 77
rect -2212 37 -2200 71
rect -2166 37 -2154 71
rect -2212 31 -2154 37
rect -2094 71 -2036 77
rect -2094 37 -2082 71
rect -2048 37 -2036 71
rect -2094 31 -2036 37
rect -1976 71 -1918 77
rect -1976 37 -1964 71
rect -1930 37 -1918 71
rect -1976 31 -1918 37
rect -1858 71 -1800 77
rect -1858 37 -1846 71
rect -1812 37 -1800 71
rect -1858 31 -1800 37
rect -1740 71 -1682 77
rect -1740 37 -1728 71
rect -1694 37 -1682 71
rect -1740 31 -1682 37
rect -1622 71 -1564 77
rect -1622 37 -1610 71
rect -1576 37 -1564 71
rect -1622 31 -1564 37
rect -1504 71 -1446 77
rect -1504 37 -1492 71
rect -1458 37 -1446 71
rect -1504 31 -1446 37
rect -1386 71 -1328 77
rect -1386 37 -1374 71
rect -1340 37 -1328 71
rect -1386 31 -1328 37
rect -1268 71 -1210 77
rect -1268 37 -1256 71
rect -1222 37 -1210 71
rect -1268 31 -1210 37
rect -1150 71 -1092 77
rect -1150 37 -1138 71
rect -1104 37 -1092 71
rect -1150 31 -1092 37
rect -1032 71 -974 77
rect -1032 37 -1020 71
rect -986 37 -974 71
rect -1032 31 -974 37
rect -914 71 -856 77
rect -914 37 -902 71
rect -868 37 -856 71
rect -914 31 -856 37
rect -796 71 -738 77
rect -796 37 -784 71
rect -750 37 -738 71
rect -796 31 -738 37
rect -678 71 -620 77
rect -678 37 -666 71
rect -632 37 -620 71
rect -678 31 -620 37
rect -560 71 -502 77
rect -560 37 -548 71
rect -514 37 -502 71
rect -560 31 -502 37
rect -442 71 -384 77
rect -442 37 -430 71
rect -396 37 -384 71
rect -442 31 -384 37
rect -324 71 -266 77
rect -324 37 -312 71
rect -278 37 -266 71
rect -324 31 -266 37
rect -206 71 -148 77
rect -206 37 -194 71
rect -160 37 -148 71
rect -206 31 -148 37
rect -88 71 -30 77
rect -88 37 -76 71
rect -42 37 -30 71
rect -88 31 -30 37
rect 30 71 88 77
rect 30 37 42 71
rect 76 37 88 71
rect 30 31 88 37
rect 148 71 206 77
rect 148 37 160 71
rect 194 37 206 71
rect 148 31 206 37
rect 266 71 324 77
rect 266 37 278 71
rect 312 37 324 71
rect 266 31 324 37
rect 384 71 442 77
rect 384 37 396 71
rect 430 37 442 71
rect 384 31 442 37
rect 502 71 560 77
rect 502 37 514 71
rect 548 37 560 71
rect 502 31 560 37
rect 620 71 678 77
rect 620 37 632 71
rect 666 37 678 71
rect 620 31 678 37
rect 738 71 796 77
rect 738 37 750 71
rect 784 37 796 71
rect 738 31 796 37
rect 856 71 914 77
rect 856 37 868 71
rect 902 37 914 71
rect 856 31 914 37
rect 974 71 1032 77
rect 974 37 986 71
rect 1020 37 1032 71
rect 974 31 1032 37
rect 1092 71 1150 77
rect 1092 37 1104 71
rect 1138 37 1150 71
rect 1092 31 1150 37
rect 1210 71 1268 77
rect 1210 37 1222 71
rect 1256 37 1268 71
rect 1210 31 1268 37
rect 1328 71 1386 77
rect 1328 37 1340 71
rect 1374 37 1386 71
rect 1328 31 1386 37
rect 1446 71 1504 77
rect 1446 37 1458 71
rect 1492 37 1504 71
rect 1446 31 1504 37
rect 1564 71 1622 77
rect 1564 37 1576 71
rect 1610 37 1622 71
rect 1564 31 1622 37
rect 1682 71 1740 77
rect 1682 37 1694 71
rect 1728 37 1740 71
rect 1682 31 1740 37
rect 1800 71 1858 77
rect 1800 37 1812 71
rect 1846 37 1858 71
rect 1800 31 1858 37
rect 1918 71 1976 77
rect 1918 37 1930 71
rect 1964 37 1976 71
rect 1918 31 1976 37
rect 2036 71 2094 77
rect 2036 37 2048 71
rect 2082 37 2094 71
rect 2036 31 2094 37
rect 2154 71 2212 77
rect 2154 37 2166 71
rect 2200 37 2212 71
rect 2154 31 2212 37
rect 2272 71 2330 77
rect 2272 37 2284 71
rect 2318 37 2330 71
rect 2272 31 2330 37
rect 2390 71 2448 77
rect 2390 37 2402 71
rect 2436 37 2448 71
rect 2390 31 2448 37
rect 2508 71 2566 77
rect 2508 37 2520 71
rect 2554 37 2566 71
rect 2508 31 2566 37
rect 2626 71 2684 77
rect 2626 37 2638 71
rect 2672 37 2684 71
rect 2626 31 2684 37
rect 2744 71 2802 77
rect 2744 37 2756 71
rect 2790 37 2802 71
rect 2744 31 2802 37
rect 2862 71 2920 77
rect 2862 37 2874 71
rect 2908 37 2920 71
rect 2862 31 2920 37
rect 2980 71 3038 77
rect 2980 37 2992 71
rect 3026 37 3038 71
rect 2980 31 3038 37
rect 3098 71 3156 77
rect 3098 37 3110 71
rect 3144 37 3156 71
rect 3098 31 3156 37
rect 3216 71 3274 77
rect 3216 37 3228 71
rect 3262 37 3274 71
rect 3216 31 3274 37
rect 3334 71 3392 77
rect 3334 37 3346 71
rect 3380 37 3392 71
rect 3334 31 3392 37
rect 3452 71 3510 77
rect 3452 37 3464 71
rect 3498 37 3510 71
rect 3452 31 3510 37
rect 3570 71 3628 77
rect 3570 37 3582 71
rect 3616 37 3628 71
rect 3570 31 3628 37
rect 3688 71 3746 77
rect 3688 37 3700 71
rect 3734 37 3746 71
rect 3688 31 3746 37
rect 3806 71 3864 77
rect 3806 37 3818 71
rect 3852 37 3864 71
rect 3806 31 3864 37
rect 3924 71 3982 77
rect 3924 37 3936 71
rect 3970 37 3982 71
rect 3924 31 3982 37
rect 4042 71 4100 77
rect 4042 37 4054 71
rect 4088 37 4100 71
rect 4042 31 4100 37
rect 4160 71 4218 77
rect 4160 37 4172 71
rect 4206 37 4218 71
rect 4160 31 4218 37
rect 4278 71 4336 77
rect 4278 37 4290 71
rect 4324 37 4336 71
rect 4278 31 4336 37
rect 4396 71 4454 77
rect 4396 37 4408 71
rect 4442 37 4454 71
rect 4396 31 4454 37
rect 4514 71 4572 77
rect 4514 37 4526 71
rect 4560 37 4572 71
rect 4514 31 4572 37
rect 4632 71 4690 77
rect 4632 37 4644 71
rect 4678 37 4690 71
rect 4632 31 4690 37
rect 4750 71 4808 77
rect 4750 37 4762 71
rect 4796 37 4808 71
rect 4750 31 4808 37
rect 4868 71 4926 77
rect 4868 37 4880 71
rect 4914 37 4926 71
rect 4868 31 4926 37
rect 4986 71 5044 77
rect 4986 37 4998 71
rect 5032 37 5044 71
rect 4986 31 5044 37
rect 5104 71 5162 77
rect 5104 37 5116 71
rect 5150 37 5162 71
rect 5104 31 5162 37
rect 5222 71 5280 77
rect 5222 37 5234 71
rect 5268 37 5280 71
rect 5222 31 5280 37
rect 5340 71 5398 77
rect 5340 37 5352 71
rect 5386 37 5398 71
rect 5340 31 5398 37
rect 5458 71 5516 77
rect 5458 37 5470 71
rect 5504 37 5516 71
rect 5458 31 5516 37
rect 5576 71 5634 77
rect 5576 37 5588 71
rect 5622 37 5634 71
rect 5576 31 5634 37
rect 5694 71 5752 77
rect 5694 37 5706 71
rect 5740 37 5752 71
rect 5694 31 5752 37
rect 5812 71 5870 77
rect 5812 37 5824 71
rect 5858 37 5870 71
rect 5812 31 5870 37
rect 5930 71 5988 77
rect 5930 37 5942 71
rect 5976 37 5988 71
rect 5930 31 5988 37
rect 6048 71 6106 77
rect 6048 37 6060 71
rect 6094 37 6106 71
rect 6048 31 6106 37
rect 6166 71 6224 77
rect 6166 37 6178 71
rect 6212 37 6224 71
rect 6166 31 6224 37
rect 6284 71 6342 77
rect 6284 37 6296 71
rect 6330 37 6342 71
rect 6284 31 6342 37
rect 6402 71 6460 77
rect 6402 37 6414 71
rect 6448 37 6460 71
rect 6402 31 6460 37
rect 6520 71 6578 77
rect 6520 37 6532 71
rect 6566 37 6578 71
rect 6520 31 6578 37
rect 6638 71 6696 77
rect 6638 37 6650 71
rect 6684 37 6696 71
rect 6638 31 6696 37
rect 6756 71 6814 77
rect 6756 37 6768 71
rect 6802 37 6814 71
rect 6756 31 6814 37
rect 6874 71 6932 77
rect 6874 37 6886 71
rect 6920 37 6932 71
rect 6874 31 6932 37
rect 6992 71 7050 77
rect 6992 37 7004 71
rect 7038 37 7050 71
rect 6992 31 7050 37
rect -7050 -37 -6992 -31
rect -7050 -71 -7038 -37
rect -7004 -71 -6992 -37
rect -7050 -77 -6992 -71
rect -6932 -37 -6874 -31
rect -6932 -71 -6920 -37
rect -6886 -71 -6874 -37
rect -6932 -77 -6874 -71
rect -6814 -37 -6756 -31
rect -6814 -71 -6802 -37
rect -6768 -71 -6756 -37
rect -6814 -77 -6756 -71
rect -6696 -37 -6638 -31
rect -6696 -71 -6684 -37
rect -6650 -71 -6638 -37
rect -6696 -77 -6638 -71
rect -6578 -37 -6520 -31
rect -6578 -71 -6566 -37
rect -6532 -71 -6520 -37
rect -6578 -77 -6520 -71
rect -6460 -37 -6402 -31
rect -6460 -71 -6448 -37
rect -6414 -71 -6402 -37
rect -6460 -77 -6402 -71
rect -6342 -37 -6284 -31
rect -6342 -71 -6330 -37
rect -6296 -71 -6284 -37
rect -6342 -77 -6284 -71
rect -6224 -37 -6166 -31
rect -6224 -71 -6212 -37
rect -6178 -71 -6166 -37
rect -6224 -77 -6166 -71
rect -6106 -37 -6048 -31
rect -6106 -71 -6094 -37
rect -6060 -71 -6048 -37
rect -6106 -77 -6048 -71
rect -5988 -37 -5930 -31
rect -5988 -71 -5976 -37
rect -5942 -71 -5930 -37
rect -5988 -77 -5930 -71
rect -5870 -37 -5812 -31
rect -5870 -71 -5858 -37
rect -5824 -71 -5812 -37
rect -5870 -77 -5812 -71
rect -5752 -37 -5694 -31
rect -5752 -71 -5740 -37
rect -5706 -71 -5694 -37
rect -5752 -77 -5694 -71
rect -5634 -37 -5576 -31
rect -5634 -71 -5622 -37
rect -5588 -71 -5576 -37
rect -5634 -77 -5576 -71
rect -5516 -37 -5458 -31
rect -5516 -71 -5504 -37
rect -5470 -71 -5458 -37
rect -5516 -77 -5458 -71
rect -5398 -37 -5340 -31
rect -5398 -71 -5386 -37
rect -5352 -71 -5340 -37
rect -5398 -77 -5340 -71
rect -5280 -37 -5222 -31
rect -5280 -71 -5268 -37
rect -5234 -71 -5222 -37
rect -5280 -77 -5222 -71
rect -5162 -37 -5104 -31
rect -5162 -71 -5150 -37
rect -5116 -71 -5104 -37
rect -5162 -77 -5104 -71
rect -5044 -37 -4986 -31
rect -5044 -71 -5032 -37
rect -4998 -71 -4986 -37
rect -5044 -77 -4986 -71
rect -4926 -37 -4868 -31
rect -4926 -71 -4914 -37
rect -4880 -71 -4868 -37
rect -4926 -77 -4868 -71
rect -4808 -37 -4750 -31
rect -4808 -71 -4796 -37
rect -4762 -71 -4750 -37
rect -4808 -77 -4750 -71
rect -4690 -37 -4632 -31
rect -4690 -71 -4678 -37
rect -4644 -71 -4632 -37
rect -4690 -77 -4632 -71
rect -4572 -37 -4514 -31
rect -4572 -71 -4560 -37
rect -4526 -71 -4514 -37
rect -4572 -77 -4514 -71
rect -4454 -37 -4396 -31
rect -4454 -71 -4442 -37
rect -4408 -71 -4396 -37
rect -4454 -77 -4396 -71
rect -4336 -37 -4278 -31
rect -4336 -71 -4324 -37
rect -4290 -71 -4278 -37
rect -4336 -77 -4278 -71
rect -4218 -37 -4160 -31
rect -4218 -71 -4206 -37
rect -4172 -71 -4160 -37
rect -4218 -77 -4160 -71
rect -4100 -37 -4042 -31
rect -4100 -71 -4088 -37
rect -4054 -71 -4042 -37
rect -4100 -77 -4042 -71
rect -3982 -37 -3924 -31
rect -3982 -71 -3970 -37
rect -3936 -71 -3924 -37
rect -3982 -77 -3924 -71
rect -3864 -37 -3806 -31
rect -3864 -71 -3852 -37
rect -3818 -71 -3806 -37
rect -3864 -77 -3806 -71
rect -3746 -37 -3688 -31
rect -3746 -71 -3734 -37
rect -3700 -71 -3688 -37
rect -3746 -77 -3688 -71
rect -3628 -37 -3570 -31
rect -3628 -71 -3616 -37
rect -3582 -71 -3570 -37
rect -3628 -77 -3570 -71
rect -3510 -37 -3452 -31
rect -3510 -71 -3498 -37
rect -3464 -71 -3452 -37
rect -3510 -77 -3452 -71
rect -3392 -37 -3334 -31
rect -3392 -71 -3380 -37
rect -3346 -71 -3334 -37
rect -3392 -77 -3334 -71
rect -3274 -37 -3216 -31
rect -3274 -71 -3262 -37
rect -3228 -71 -3216 -37
rect -3274 -77 -3216 -71
rect -3156 -37 -3098 -31
rect -3156 -71 -3144 -37
rect -3110 -71 -3098 -37
rect -3156 -77 -3098 -71
rect -3038 -37 -2980 -31
rect -3038 -71 -3026 -37
rect -2992 -71 -2980 -37
rect -3038 -77 -2980 -71
rect -2920 -37 -2862 -31
rect -2920 -71 -2908 -37
rect -2874 -71 -2862 -37
rect -2920 -77 -2862 -71
rect -2802 -37 -2744 -31
rect -2802 -71 -2790 -37
rect -2756 -71 -2744 -37
rect -2802 -77 -2744 -71
rect -2684 -37 -2626 -31
rect -2684 -71 -2672 -37
rect -2638 -71 -2626 -37
rect -2684 -77 -2626 -71
rect -2566 -37 -2508 -31
rect -2566 -71 -2554 -37
rect -2520 -71 -2508 -37
rect -2566 -77 -2508 -71
rect -2448 -37 -2390 -31
rect -2448 -71 -2436 -37
rect -2402 -71 -2390 -37
rect -2448 -77 -2390 -71
rect -2330 -37 -2272 -31
rect -2330 -71 -2318 -37
rect -2284 -71 -2272 -37
rect -2330 -77 -2272 -71
rect -2212 -37 -2154 -31
rect -2212 -71 -2200 -37
rect -2166 -71 -2154 -37
rect -2212 -77 -2154 -71
rect -2094 -37 -2036 -31
rect -2094 -71 -2082 -37
rect -2048 -71 -2036 -37
rect -2094 -77 -2036 -71
rect -1976 -37 -1918 -31
rect -1976 -71 -1964 -37
rect -1930 -71 -1918 -37
rect -1976 -77 -1918 -71
rect -1858 -37 -1800 -31
rect -1858 -71 -1846 -37
rect -1812 -71 -1800 -37
rect -1858 -77 -1800 -71
rect -1740 -37 -1682 -31
rect -1740 -71 -1728 -37
rect -1694 -71 -1682 -37
rect -1740 -77 -1682 -71
rect -1622 -37 -1564 -31
rect -1622 -71 -1610 -37
rect -1576 -71 -1564 -37
rect -1622 -77 -1564 -71
rect -1504 -37 -1446 -31
rect -1504 -71 -1492 -37
rect -1458 -71 -1446 -37
rect -1504 -77 -1446 -71
rect -1386 -37 -1328 -31
rect -1386 -71 -1374 -37
rect -1340 -71 -1328 -37
rect -1386 -77 -1328 -71
rect -1268 -37 -1210 -31
rect -1268 -71 -1256 -37
rect -1222 -71 -1210 -37
rect -1268 -77 -1210 -71
rect -1150 -37 -1092 -31
rect -1150 -71 -1138 -37
rect -1104 -71 -1092 -37
rect -1150 -77 -1092 -71
rect -1032 -37 -974 -31
rect -1032 -71 -1020 -37
rect -986 -71 -974 -37
rect -1032 -77 -974 -71
rect -914 -37 -856 -31
rect -914 -71 -902 -37
rect -868 -71 -856 -37
rect -914 -77 -856 -71
rect -796 -37 -738 -31
rect -796 -71 -784 -37
rect -750 -71 -738 -37
rect -796 -77 -738 -71
rect -678 -37 -620 -31
rect -678 -71 -666 -37
rect -632 -71 -620 -37
rect -678 -77 -620 -71
rect -560 -37 -502 -31
rect -560 -71 -548 -37
rect -514 -71 -502 -37
rect -560 -77 -502 -71
rect -442 -37 -384 -31
rect -442 -71 -430 -37
rect -396 -71 -384 -37
rect -442 -77 -384 -71
rect -324 -37 -266 -31
rect -324 -71 -312 -37
rect -278 -71 -266 -37
rect -324 -77 -266 -71
rect -206 -37 -148 -31
rect -206 -71 -194 -37
rect -160 -71 -148 -37
rect -206 -77 -148 -71
rect -88 -37 -30 -31
rect -88 -71 -76 -37
rect -42 -71 -30 -37
rect -88 -77 -30 -71
rect 30 -37 88 -31
rect 30 -71 42 -37
rect 76 -71 88 -37
rect 30 -77 88 -71
rect 148 -37 206 -31
rect 148 -71 160 -37
rect 194 -71 206 -37
rect 148 -77 206 -71
rect 266 -37 324 -31
rect 266 -71 278 -37
rect 312 -71 324 -37
rect 266 -77 324 -71
rect 384 -37 442 -31
rect 384 -71 396 -37
rect 430 -71 442 -37
rect 384 -77 442 -71
rect 502 -37 560 -31
rect 502 -71 514 -37
rect 548 -71 560 -37
rect 502 -77 560 -71
rect 620 -37 678 -31
rect 620 -71 632 -37
rect 666 -71 678 -37
rect 620 -77 678 -71
rect 738 -37 796 -31
rect 738 -71 750 -37
rect 784 -71 796 -37
rect 738 -77 796 -71
rect 856 -37 914 -31
rect 856 -71 868 -37
rect 902 -71 914 -37
rect 856 -77 914 -71
rect 974 -37 1032 -31
rect 974 -71 986 -37
rect 1020 -71 1032 -37
rect 974 -77 1032 -71
rect 1092 -37 1150 -31
rect 1092 -71 1104 -37
rect 1138 -71 1150 -37
rect 1092 -77 1150 -71
rect 1210 -37 1268 -31
rect 1210 -71 1222 -37
rect 1256 -71 1268 -37
rect 1210 -77 1268 -71
rect 1328 -37 1386 -31
rect 1328 -71 1340 -37
rect 1374 -71 1386 -37
rect 1328 -77 1386 -71
rect 1446 -37 1504 -31
rect 1446 -71 1458 -37
rect 1492 -71 1504 -37
rect 1446 -77 1504 -71
rect 1564 -37 1622 -31
rect 1564 -71 1576 -37
rect 1610 -71 1622 -37
rect 1564 -77 1622 -71
rect 1682 -37 1740 -31
rect 1682 -71 1694 -37
rect 1728 -71 1740 -37
rect 1682 -77 1740 -71
rect 1800 -37 1858 -31
rect 1800 -71 1812 -37
rect 1846 -71 1858 -37
rect 1800 -77 1858 -71
rect 1918 -37 1976 -31
rect 1918 -71 1930 -37
rect 1964 -71 1976 -37
rect 1918 -77 1976 -71
rect 2036 -37 2094 -31
rect 2036 -71 2048 -37
rect 2082 -71 2094 -37
rect 2036 -77 2094 -71
rect 2154 -37 2212 -31
rect 2154 -71 2166 -37
rect 2200 -71 2212 -37
rect 2154 -77 2212 -71
rect 2272 -37 2330 -31
rect 2272 -71 2284 -37
rect 2318 -71 2330 -37
rect 2272 -77 2330 -71
rect 2390 -37 2448 -31
rect 2390 -71 2402 -37
rect 2436 -71 2448 -37
rect 2390 -77 2448 -71
rect 2508 -37 2566 -31
rect 2508 -71 2520 -37
rect 2554 -71 2566 -37
rect 2508 -77 2566 -71
rect 2626 -37 2684 -31
rect 2626 -71 2638 -37
rect 2672 -71 2684 -37
rect 2626 -77 2684 -71
rect 2744 -37 2802 -31
rect 2744 -71 2756 -37
rect 2790 -71 2802 -37
rect 2744 -77 2802 -71
rect 2862 -37 2920 -31
rect 2862 -71 2874 -37
rect 2908 -71 2920 -37
rect 2862 -77 2920 -71
rect 2980 -37 3038 -31
rect 2980 -71 2992 -37
rect 3026 -71 3038 -37
rect 2980 -77 3038 -71
rect 3098 -37 3156 -31
rect 3098 -71 3110 -37
rect 3144 -71 3156 -37
rect 3098 -77 3156 -71
rect 3216 -37 3274 -31
rect 3216 -71 3228 -37
rect 3262 -71 3274 -37
rect 3216 -77 3274 -71
rect 3334 -37 3392 -31
rect 3334 -71 3346 -37
rect 3380 -71 3392 -37
rect 3334 -77 3392 -71
rect 3452 -37 3510 -31
rect 3452 -71 3464 -37
rect 3498 -71 3510 -37
rect 3452 -77 3510 -71
rect 3570 -37 3628 -31
rect 3570 -71 3582 -37
rect 3616 -71 3628 -37
rect 3570 -77 3628 -71
rect 3688 -37 3746 -31
rect 3688 -71 3700 -37
rect 3734 -71 3746 -37
rect 3688 -77 3746 -71
rect 3806 -37 3864 -31
rect 3806 -71 3818 -37
rect 3852 -71 3864 -37
rect 3806 -77 3864 -71
rect 3924 -37 3982 -31
rect 3924 -71 3936 -37
rect 3970 -71 3982 -37
rect 3924 -77 3982 -71
rect 4042 -37 4100 -31
rect 4042 -71 4054 -37
rect 4088 -71 4100 -37
rect 4042 -77 4100 -71
rect 4160 -37 4218 -31
rect 4160 -71 4172 -37
rect 4206 -71 4218 -37
rect 4160 -77 4218 -71
rect 4278 -37 4336 -31
rect 4278 -71 4290 -37
rect 4324 -71 4336 -37
rect 4278 -77 4336 -71
rect 4396 -37 4454 -31
rect 4396 -71 4408 -37
rect 4442 -71 4454 -37
rect 4396 -77 4454 -71
rect 4514 -37 4572 -31
rect 4514 -71 4526 -37
rect 4560 -71 4572 -37
rect 4514 -77 4572 -71
rect 4632 -37 4690 -31
rect 4632 -71 4644 -37
rect 4678 -71 4690 -37
rect 4632 -77 4690 -71
rect 4750 -37 4808 -31
rect 4750 -71 4762 -37
rect 4796 -71 4808 -37
rect 4750 -77 4808 -71
rect 4868 -37 4926 -31
rect 4868 -71 4880 -37
rect 4914 -71 4926 -37
rect 4868 -77 4926 -71
rect 4986 -37 5044 -31
rect 4986 -71 4998 -37
rect 5032 -71 5044 -37
rect 4986 -77 5044 -71
rect 5104 -37 5162 -31
rect 5104 -71 5116 -37
rect 5150 -71 5162 -37
rect 5104 -77 5162 -71
rect 5222 -37 5280 -31
rect 5222 -71 5234 -37
rect 5268 -71 5280 -37
rect 5222 -77 5280 -71
rect 5340 -37 5398 -31
rect 5340 -71 5352 -37
rect 5386 -71 5398 -37
rect 5340 -77 5398 -71
rect 5458 -37 5516 -31
rect 5458 -71 5470 -37
rect 5504 -71 5516 -37
rect 5458 -77 5516 -71
rect 5576 -37 5634 -31
rect 5576 -71 5588 -37
rect 5622 -71 5634 -37
rect 5576 -77 5634 -71
rect 5694 -37 5752 -31
rect 5694 -71 5706 -37
rect 5740 -71 5752 -37
rect 5694 -77 5752 -71
rect 5812 -37 5870 -31
rect 5812 -71 5824 -37
rect 5858 -71 5870 -37
rect 5812 -77 5870 -71
rect 5930 -37 5988 -31
rect 5930 -71 5942 -37
rect 5976 -71 5988 -37
rect 5930 -77 5988 -71
rect 6048 -37 6106 -31
rect 6048 -71 6060 -37
rect 6094 -71 6106 -37
rect 6048 -77 6106 -71
rect 6166 -37 6224 -31
rect 6166 -71 6178 -37
rect 6212 -71 6224 -37
rect 6166 -77 6224 -71
rect 6284 -37 6342 -31
rect 6284 -71 6296 -37
rect 6330 -71 6342 -37
rect 6284 -77 6342 -71
rect 6402 -37 6460 -31
rect 6402 -71 6414 -37
rect 6448 -71 6460 -37
rect 6402 -77 6460 -71
rect 6520 -37 6578 -31
rect 6520 -71 6532 -37
rect 6566 -71 6578 -37
rect 6520 -77 6578 -71
rect 6638 -37 6696 -31
rect 6638 -71 6650 -37
rect 6684 -71 6696 -37
rect 6638 -77 6696 -71
rect 6756 -37 6814 -31
rect 6756 -71 6768 -37
rect 6802 -71 6814 -37
rect 6756 -77 6814 -71
rect 6874 -37 6932 -31
rect 6874 -71 6886 -37
rect 6920 -71 6932 -37
rect 6874 -77 6932 -71
rect 6992 -37 7050 -31
rect 6992 -71 7004 -37
rect 7038 -71 7050 -37
rect 6992 -77 7050 -71
rect -7103 -130 -7057 -118
rect -7103 -706 -7097 -130
rect -7063 -706 -7057 -130
rect -7103 -718 -7057 -706
rect -6985 -130 -6939 -118
rect -6985 -706 -6979 -130
rect -6945 -706 -6939 -130
rect -6985 -718 -6939 -706
rect -6867 -130 -6821 -118
rect -6867 -706 -6861 -130
rect -6827 -706 -6821 -130
rect -6867 -718 -6821 -706
rect -6749 -130 -6703 -118
rect -6749 -706 -6743 -130
rect -6709 -706 -6703 -130
rect -6749 -718 -6703 -706
rect -6631 -130 -6585 -118
rect -6631 -706 -6625 -130
rect -6591 -706 -6585 -130
rect -6631 -718 -6585 -706
rect -6513 -130 -6467 -118
rect -6513 -706 -6507 -130
rect -6473 -706 -6467 -130
rect -6513 -718 -6467 -706
rect -6395 -130 -6349 -118
rect -6395 -706 -6389 -130
rect -6355 -706 -6349 -130
rect -6395 -718 -6349 -706
rect -6277 -130 -6231 -118
rect -6277 -706 -6271 -130
rect -6237 -706 -6231 -130
rect -6277 -718 -6231 -706
rect -6159 -130 -6113 -118
rect -6159 -706 -6153 -130
rect -6119 -706 -6113 -130
rect -6159 -718 -6113 -706
rect -6041 -130 -5995 -118
rect -6041 -706 -6035 -130
rect -6001 -706 -5995 -130
rect -6041 -718 -5995 -706
rect -5923 -130 -5877 -118
rect -5923 -706 -5917 -130
rect -5883 -706 -5877 -130
rect -5923 -718 -5877 -706
rect -5805 -130 -5759 -118
rect -5805 -706 -5799 -130
rect -5765 -706 -5759 -130
rect -5805 -718 -5759 -706
rect -5687 -130 -5641 -118
rect -5687 -706 -5681 -130
rect -5647 -706 -5641 -130
rect -5687 -718 -5641 -706
rect -5569 -130 -5523 -118
rect -5569 -706 -5563 -130
rect -5529 -706 -5523 -130
rect -5569 -718 -5523 -706
rect -5451 -130 -5405 -118
rect -5451 -706 -5445 -130
rect -5411 -706 -5405 -130
rect -5451 -718 -5405 -706
rect -5333 -130 -5287 -118
rect -5333 -706 -5327 -130
rect -5293 -706 -5287 -130
rect -5333 -718 -5287 -706
rect -5215 -130 -5169 -118
rect -5215 -706 -5209 -130
rect -5175 -706 -5169 -130
rect -5215 -718 -5169 -706
rect -5097 -130 -5051 -118
rect -5097 -706 -5091 -130
rect -5057 -706 -5051 -130
rect -5097 -718 -5051 -706
rect -4979 -130 -4933 -118
rect -4979 -706 -4973 -130
rect -4939 -706 -4933 -130
rect -4979 -718 -4933 -706
rect -4861 -130 -4815 -118
rect -4861 -706 -4855 -130
rect -4821 -706 -4815 -130
rect -4861 -718 -4815 -706
rect -4743 -130 -4697 -118
rect -4743 -706 -4737 -130
rect -4703 -706 -4697 -130
rect -4743 -718 -4697 -706
rect -4625 -130 -4579 -118
rect -4625 -706 -4619 -130
rect -4585 -706 -4579 -130
rect -4625 -718 -4579 -706
rect -4507 -130 -4461 -118
rect -4507 -706 -4501 -130
rect -4467 -706 -4461 -130
rect -4507 -718 -4461 -706
rect -4389 -130 -4343 -118
rect -4389 -706 -4383 -130
rect -4349 -706 -4343 -130
rect -4389 -718 -4343 -706
rect -4271 -130 -4225 -118
rect -4271 -706 -4265 -130
rect -4231 -706 -4225 -130
rect -4271 -718 -4225 -706
rect -4153 -130 -4107 -118
rect -4153 -706 -4147 -130
rect -4113 -706 -4107 -130
rect -4153 -718 -4107 -706
rect -4035 -130 -3989 -118
rect -4035 -706 -4029 -130
rect -3995 -706 -3989 -130
rect -4035 -718 -3989 -706
rect -3917 -130 -3871 -118
rect -3917 -706 -3911 -130
rect -3877 -706 -3871 -130
rect -3917 -718 -3871 -706
rect -3799 -130 -3753 -118
rect -3799 -706 -3793 -130
rect -3759 -706 -3753 -130
rect -3799 -718 -3753 -706
rect -3681 -130 -3635 -118
rect -3681 -706 -3675 -130
rect -3641 -706 -3635 -130
rect -3681 -718 -3635 -706
rect -3563 -130 -3517 -118
rect -3563 -706 -3557 -130
rect -3523 -706 -3517 -130
rect -3563 -718 -3517 -706
rect -3445 -130 -3399 -118
rect -3445 -706 -3439 -130
rect -3405 -706 -3399 -130
rect -3445 -718 -3399 -706
rect -3327 -130 -3281 -118
rect -3327 -706 -3321 -130
rect -3287 -706 -3281 -130
rect -3327 -718 -3281 -706
rect -3209 -130 -3163 -118
rect -3209 -706 -3203 -130
rect -3169 -706 -3163 -130
rect -3209 -718 -3163 -706
rect -3091 -130 -3045 -118
rect -3091 -706 -3085 -130
rect -3051 -706 -3045 -130
rect -3091 -718 -3045 -706
rect -2973 -130 -2927 -118
rect -2973 -706 -2967 -130
rect -2933 -706 -2927 -130
rect -2973 -718 -2927 -706
rect -2855 -130 -2809 -118
rect -2855 -706 -2849 -130
rect -2815 -706 -2809 -130
rect -2855 -718 -2809 -706
rect -2737 -130 -2691 -118
rect -2737 -706 -2731 -130
rect -2697 -706 -2691 -130
rect -2737 -718 -2691 -706
rect -2619 -130 -2573 -118
rect -2619 -706 -2613 -130
rect -2579 -706 -2573 -130
rect -2619 -718 -2573 -706
rect -2501 -130 -2455 -118
rect -2501 -706 -2495 -130
rect -2461 -706 -2455 -130
rect -2501 -718 -2455 -706
rect -2383 -130 -2337 -118
rect -2383 -706 -2377 -130
rect -2343 -706 -2337 -130
rect -2383 -718 -2337 -706
rect -2265 -130 -2219 -118
rect -2265 -706 -2259 -130
rect -2225 -706 -2219 -130
rect -2265 -718 -2219 -706
rect -2147 -130 -2101 -118
rect -2147 -706 -2141 -130
rect -2107 -706 -2101 -130
rect -2147 -718 -2101 -706
rect -2029 -130 -1983 -118
rect -2029 -706 -2023 -130
rect -1989 -706 -1983 -130
rect -2029 -718 -1983 -706
rect -1911 -130 -1865 -118
rect -1911 -706 -1905 -130
rect -1871 -706 -1865 -130
rect -1911 -718 -1865 -706
rect -1793 -130 -1747 -118
rect -1793 -706 -1787 -130
rect -1753 -706 -1747 -130
rect -1793 -718 -1747 -706
rect -1675 -130 -1629 -118
rect -1675 -706 -1669 -130
rect -1635 -706 -1629 -130
rect -1675 -718 -1629 -706
rect -1557 -130 -1511 -118
rect -1557 -706 -1551 -130
rect -1517 -706 -1511 -130
rect -1557 -718 -1511 -706
rect -1439 -130 -1393 -118
rect -1439 -706 -1433 -130
rect -1399 -706 -1393 -130
rect -1439 -718 -1393 -706
rect -1321 -130 -1275 -118
rect -1321 -706 -1315 -130
rect -1281 -706 -1275 -130
rect -1321 -718 -1275 -706
rect -1203 -130 -1157 -118
rect -1203 -706 -1197 -130
rect -1163 -706 -1157 -130
rect -1203 -718 -1157 -706
rect -1085 -130 -1039 -118
rect -1085 -706 -1079 -130
rect -1045 -706 -1039 -130
rect -1085 -718 -1039 -706
rect -967 -130 -921 -118
rect -967 -706 -961 -130
rect -927 -706 -921 -130
rect -967 -718 -921 -706
rect -849 -130 -803 -118
rect -849 -706 -843 -130
rect -809 -706 -803 -130
rect -849 -718 -803 -706
rect -731 -130 -685 -118
rect -731 -706 -725 -130
rect -691 -706 -685 -130
rect -731 -718 -685 -706
rect -613 -130 -567 -118
rect -613 -706 -607 -130
rect -573 -706 -567 -130
rect -613 -718 -567 -706
rect -495 -130 -449 -118
rect -495 -706 -489 -130
rect -455 -706 -449 -130
rect -495 -718 -449 -706
rect -377 -130 -331 -118
rect -377 -706 -371 -130
rect -337 -706 -331 -130
rect -377 -718 -331 -706
rect -259 -130 -213 -118
rect -259 -706 -253 -130
rect -219 -706 -213 -130
rect -259 -718 -213 -706
rect -141 -130 -95 -118
rect -141 -706 -135 -130
rect -101 -706 -95 -130
rect -141 -718 -95 -706
rect -23 -130 23 -118
rect -23 -706 -17 -130
rect 17 -706 23 -130
rect -23 -718 23 -706
rect 95 -130 141 -118
rect 95 -706 101 -130
rect 135 -706 141 -130
rect 95 -718 141 -706
rect 213 -130 259 -118
rect 213 -706 219 -130
rect 253 -706 259 -130
rect 213 -718 259 -706
rect 331 -130 377 -118
rect 331 -706 337 -130
rect 371 -706 377 -130
rect 331 -718 377 -706
rect 449 -130 495 -118
rect 449 -706 455 -130
rect 489 -706 495 -130
rect 449 -718 495 -706
rect 567 -130 613 -118
rect 567 -706 573 -130
rect 607 -706 613 -130
rect 567 -718 613 -706
rect 685 -130 731 -118
rect 685 -706 691 -130
rect 725 -706 731 -130
rect 685 -718 731 -706
rect 803 -130 849 -118
rect 803 -706 809 -130
rect 843 -706 849 -130
rect 803 -718 849 -706
rect 921 -130 967 -118
rect 921 -706 927 -130
rect 961 -706 967 -130
rect 921 -718 967 -706
rect 1039 -130 1085 -118
rect 1039 -706 1045 -130
rect 1079 -706 1085 -130
rect 1039 -718 1085 -706
rect 1157 -130 1203 -118
rect 1157 -706 1163 -130
rect 1197 -706 1203 -130
rect 1157 -718 1203 -706
rect 1275 -130 1321 -118
rect 1275 -706 1281 -130
rect 1315 -706 1321 -130
rect 1275 -718 1321 -706
rect 1393 -130 1439 -118
rect 1393 -706 1399 -130
rect 1433 -706 1439 -130
rect 1393 -718 1439 -706
rect 1511 -130 1557 -118
rect 1511 -706 1517 -130
rect 1551 -706 1557 -130
rect 1511 -718 1557 -706
rect 1629 -130 1675 -118
rect 1629 -706 1635 -130
rect 1669 -706 1675 -130
rect 1629 -718 1675 -706
rect 1747 -130 1793 -118
rect 1747 -706 1753 -130
rect 1787 -706 1793 -130
rect 1747 -718 1793 -706
rect 1865 -130 1911 -118
rect 1865 -706 1871 -130
rect 1905 -706 1911 -130
rect 1865 -718 1911 -706
rect 1983 -130 2029 -118
rect 1983 -706 1989 -130
rect 2023 -706 2029 -130
rect 1983 -718 2029 -706
rect 2101 -130 2147 -118
rect 2101 -706 2107 -130
rect 2141 -706 2147 -130
rect 2101 -718 2147 -706
rect 2219 -130 2265 -118
rect 2219 -706 2225 -130
rect 2259 -706 2265 -130
rect 2219 -718 2265 -706
rect 2337 -130 2383 -118
rect 2337 -706 2343 -130
rect 2377 -706 2383 -130
rect 2337 -718 2383 -706
rect 2455 -130 2501 -118
rect 2455 -706 2461 -130
rect 2495 -706 2501 -130
rect 2455 -718 2501 -706
rect 2573 -130 2619 -118
rect 2573 -706 2579 -130
rect 2613 -706 2619 -130
rect 2573 -718 2619 -706
rect 2691 -130 2737 -118
rect 2691 -706 2697 -130
rect 2731 -706 2737 -130
rect 2691 -718 2737 -706
rect 2809 -130 2855 -118
rect 2809 -706 2815 -130
rect 2849 -706 2855 -130
rect 2809 -718 2855 -706
rect 2927 -130 2973 -118
rect 2927 -706 2933 -130
rect 2967 -706 2973 -130
rect 2927 -718 2973 -706
rect 3045 -130 3091 -118
rect 3045 -706 3051 -130
rect 3085 -706 3091 -130
rect 3045 -718 3091 -706
rect 3163 -130 3209 -118
rect 3163 -706 3169 -130
rect 3203 -706 3209 -130
rect 3163 -718 3209 -706
rect 3281 -130 3327 -118
rect 3281 -706 3287 -130
rect 3321 -706 3327 -130
rect 3281 -718 3327 -706
rect 3399 -130 3445 -118
rect 3399 -706 3405 -130
rect 3439 -706 3445 -130
rect 3399 -718 3445 -706
rect 3517 -130 3563 -118
rect 3517 -706 3523 -130
rect 3557 -706 3563 -130
rect 3517 -718 3563 -706
rect 3635 -130 3681 -118
rect 3635 -706 3641 -130
rect 3675 -706 3681 -130
rect 3635 -718 3681 -706
rect 3753 -130 3799 -118
rect 3753 -706 3759 -130
rect 3793 -706 3799 -130
rect 3753 -718 3799 -706
rect 3871 -130 3917 -118
rect 3871 -706 3877 -130
rect 3911 -706 3917 -130
rect 3871 -718 3917 -706
rect 3989 -130 4035 -118
rect 3989 -706 3995 -130
rect 4029 -706 4035 -130
rect 3989 -718 4035 -706
rect 4107 -130 4153 -118
rect 4107 -706 4113 -130
rect 4147 -706 4153 -130
rect 4107 -718 4153 -706
rect 4225 -130 4271 -118
rect 4225 -706 4231 -130
rect 4265 -706 4271 -130
rect 4225 -718 4271 -706
rect 4343 -130 4389 -118
rect 4343 -706 4349 -130
rect 4383 -706 4389 -130
rect 4343 -718 4389 -706
rect 4461 -130 4507 -118
rect 4461 -706 4467 -130
rect 4501 -706 4507 -130
rect 4461 -718 4507 -706
rect 4579 -130 4625 -118
rect 4579 -706 4585 -130
rect 4619 -706 4625 -130
rect 4579 -718 4625 -706
rect 4697 -130 4743 -118
rect 4697 -706 4703 -130
rect 4737 -706 4743 -130
rect 4697 -718 4743 -706
rect 4815 -130 4861 -118
rect 4815 -706 4821 -130
rect 4855 -706 4861 -130
rect 4815 -718 4861 -706
rect 4933 -130 4979 -118
rect 4933 -706 4939 -130
rect 4973 -706 4979 -130
rect 4933 -718 4979 -706
rect 5051 -130 5097 -118
rect 5051 -706 5057 -130
rect 5091 -706 5097 -130
rect 5051 -718 5097 -706
rect 5169 -130 5215 -118
rect 5169 -706 5175 -130
rect 5209 -706 5215 -130
rect 5169 -718 5215 -706
rect 5287 -130 5333 -118
rect 5287 -706 5293 -130
rect 5327 -706 5333 -130
rect 5287 -718 5333 -706
rect 5405 -130 5451 -118
rect 5405 -706 5411 -130
rect 5445 -706 5451 -130
rect 5405 -718 5451 -706
rect 5523 -130 5569 -118
rect 5523 -706 5529 -130
rect 5563 -706 5569 -130
rect 5523 -718 5569 -706
rect 5641 -130 5687 -118
rect 5641 -706 5647 -130
rect 5681 -706 5687 -130
rect 5641 -718 5687 -706
rect 5759 -130 5805 -118
rect 5759 -706 5765 -130
rect 5799 -706 5805 -130
rect 5759 -718 5805 -706
rect 5877 -130 5923 -118
rect 5877 -706 5883 -130
rect 5917 -706 5923 -130
rect 5877 -718 5923 -706
rect 5995 -130 6041 -118
rect 5995 -706 6001 -130
rect 6035 -706 6041 -130
rect 5995 -718 6041 -706
rect 6113 -130 6159 -118
rect 6113 -706 6119 -130
rect 6153 -706 6159 -130
rect 6113 -718 6159 -706
rect 6231 -130 6277 -118
rect 6231 -706 6237 -130
rect 6271 -706 6277 -130
rect 6231 -718 6277 -706
rect 6349 -130 6395 -118
rect 6349 -706 6355 -130
rect 6389 -706 6395 -130
rect 6349 -718 6395 -706
rect 6467 -130 6513 -118
rect 6467 -706 6473 -130
rect 6507 -706 6513 -130
rect 6467 -718 6513 -706
rect 6585 -130 6631 -118
rect 6585 -706 6591 -130
rect 6625 -706 6631 -130
rect 6585 -718 6631 -706
rect 6703 -130 6749 -118
rect 6703 -706 6709 -130
rect 6743 -706 6749 -130
rect 6703 -718 6749 -706
rect 6821 -130 6867 -118
rect 6821 -706 6827 -130
rect 6861 -706 6867 -130
rect 6821 -718 6867 -706
rect 6939 -130 6985 -118
rect 6939 -706 6945 -130
rect 6979 -706 6985 -130
rect 6939 -718 6985 -706
rect 7057 -130 7103 -118
rect 7057 -706 7063 -130
rect 7097 -706 7103 -130
rect 7057 -718 7103 -706
rect -7050 -765 -6992 -759
rect -7050 -799 -7038 -765
rect -7004 -799 -6992 -765
rect -7050 -805 -6992 -799
rect -6932 -765 -6874 -759
rect -6932 -799 -6920 -765
rect -6886 -799 -6874 -765
rect -6932 -805 -6874 -799
rect -6814 -765 -6756 -759
rect -6814 -799 -6802 -765
rect -6768 -799 -6756 -765
rect -6814 -805 -6756 -799
rect -6696 -765 -6638 -759
rect -6696 -799 -6684 -765
rect -6650 -799 -6638 -765
rect -6696 -805 -6638 -799
rect -6578 -765 -6520 -759
rect -6578 -799 -6566 -765
rect -6532 -799 -6520 -765
rect -6578 -805 -6520 -799
rect -6460 -765 -6402 -759
rect -6460 -799 -6448 -765
rect -6414 -799 -6402 -765
rect -6460 -805 -6402 -799
rect -6342 -765 -6284 -759
rect -6342 -799 -6330 -765
rect -6296 -799 -6284 -765
rect -6342 -805 -6284 -799
rect -6224 -765 -6166 -759
rect -6224 -799 -6212 -765
rect -6178 -799 -6166 -765
rect -6224 -805 -6166 -799
rect -6106 -765 -6048 -759
rect -6106 -799 -6094 -765
rect -6060 -799 -6048 -765
rect -6106 -805 -6048 -799
rect -5988 -765 -5930 -759
rect -5988 -799 -5976 -765
rect -5942 -799 -5930 -765
rect -5988 -805 -5930 -799
rect -5870 -765 -5812 -759
rect -5870 -799 -5858 -765
rect -5824 -799 -5812 -765
rect -5870 -805 -5812 -799
rect -5752 -765 -5694 -759
rect -5752 -799 -5740 -765
rect -5706 -799 -5694 -765
rect -5752 -805 -5694 -799
rect -5634 -765 -5576 -759
rect -5634 -799 -5622 -765
rect -5588 -799 -5576 -765
rect -5634 -805 -5576 -799
rect -5516 -765 -5458 -759
rect -5516 -799 -5504 -765
rect -5470 -799 -5458 -765
rect -5516 -805 -5458 -799
rect -5398 -765 -5340 -759
rect -5398 -799 -5386 -765
rect -5352 -799 -5340 -765
rect -5398 -805 -5340 -799
rect -5280 -765 -5222 -759
rect -5280 -799 -5268 -765
rect -5234 -799 -5222 -765
rect -5280 -805 -5222 -799
rect -5162 -765 -5104 -759
rect -5162 -799 -5150 -765
rect -5116 -799 -5104 -765
rect -5162 -805 -5104 -799
rect -5044 -765 -4986 -759
rect -5044 -799 -5032 -765
rect -4998 -799 -4986 -765
rect -5044 -805 -4986 -799
rect -4926 -765 -4868 -759
rect -4926 -799 -4914 -765
rect -4880 -799 -4868 -765
rect -4926 -805 -4868 -799
rect -4808 -765 -4750 -759
rect -4808 -799 -4796 -765
rect -4762 -799 -4750 -765
rect -4808 -805 -4750 -799
rect -4690 -765 -4632 -759
rect -4690 -799 -4678 -765
rect -4644 -799 -4632 -765
rect -4690 -805 -4632 -799
rect -4572 -765 -4514 -759
rect -4572 -799 -4560 -765
rect -4526 -799 -4514 -765
rect -4572 -805 -4514 -799
rect -4454 -765 -4396 -759
rect -4454 -799 -4442 -765
rect -4408 -799 -4396 -765
rect -4454 -805 -4396 -799
rect -4336 -765 -4278 -759
rect -4336 -799 -4324 -765
rect -4290 -799 -4278 -765
rect -4336 -805 -4278 -799
rect -4218 -765 -4160 -759
rect -4218 -799 -4206 -765
rect -4172 -799 -4160 -765
rect -4218 -805 -4160 -799
rect -4100 -765 -4042 -759
rect -4100 -799 -4088 -765
rect -4054 -799 -4042 -765
rect -4100 -805 -4042 -799
rect -3982 -765 -3924 -759
rect -3982 -799 -3970 -765
rect -3936 -799 -3924 -765
rect -3982 -805 -3924 -799
rect -3864 -765 -3806 -759
rect -3864 -799 -3852 -765
rect -3818 -799 -3806 -765
rect -3864 -805 -3806 -799
rect -3746 -765 -3688 -759
rect -3746 -799 -3734 -765
rect -3700 -799 -3688 -765
rect -3746 -805 -3688 -799
rect -3628 -765 -3570 -759
rect -3628 -799 -3616 -765
rect -3582 -799 -3570 -765
rect -3628 -805 -3570 -799
rect -3510 -765 -3452 -759
rect -3510 -799 -3498 -765
rect -3464 -799 -3452 -765
rect -3510 -805 -3452 -799
rect -3392 -765 -3334 -759
rect -3392 -799 -3380 -765
rect -3346 -799 -3334 -765
rect -3392 -805 -3334 -799
rect -3274 -765 -3216 -759
rect -3274 -799 -3262 -765
rect -3228 -799 -3216 -765
rect -3274 -805 -3216 -799
rect -3156 -765 -3098 -759
rect -3156 -799 -3144 -765
rect -3110 -799 -3098 -765
rect -3156 -805 -3098 -799
rect -3038 -765 -2980 -759
rect -3038 -799 -3026 -765
rect -2992 -799 -2980 -765
rect -3038 -805 -2980 -799
rect -2920 -765 -2862 -759
rect -2920 -799 -2908 -765
rect -2874 -799 -2862 -765
rect -2920 -805 -2862 -799
rect -2802 -765 -2744 -759
rect -2802 -799 -2790 -765
rect -2756 -799 -2744 -765
rect -2802 -805 -2744 -799
rect -2684 -765 -2626 -759
rect -2684 -799 -2672 -765
rect -2638 -799 -2626 -765
rect -2684 -805 -2626 -799
rect -2566 -765 -2508 -759
rect -2566 -799 -2554 -765
rect -2520 -799 -2508 -765
rect -2566 -805 -2508 -799
rect -2448 -765 -2390 -759
rect -2448 -799 -2436 -765
rect -2402 -799 -2390 -765
rect -2448 -805 -2390 -799
rect -2330 -765 -2272 -759
rect -2330 -799 -2318 -765
rect -2284 -799 -2272 -765
rect -2330 -805 -2272 -799
rect -2212 -765 -2154 -759
rect -2212 -799 -2200 -765
rect -2166 -799 -2154 -765
rect -2212 -805 -2154 -799
rect -2094 -765 -2036 -759
rect -2094 -799 -2082 -765
rect -2048 -799 -2036 -765
rect -2094 -805 -2036 -799
rect -1976 -765 -1918 -759
rect -1976 -799 -1964 -765
rect -1930 -799 -1918 -765
rect -1976 -805 -1918 -799
rect -1858 -765 -1800 -759
rect -1858 -799 -1846 -765
rect -1812 -799 -1800 -765
rect -1858 -805 -1800 -799
rect -1740 -765 -1682 -759
rect -1740 -799 -1728 -765
rect -1694 -799 -1682 -765
rect -1740 -805 -1682 -799
rect -1622 -765 -1564 -759
rect -1622 -799 -1610 -765
rect -1576 -799 -1564 -765
rect -1622 -805 -1564 -799
rect -1504 -765 -1446 -759
rect -1504 -799 -1492 -765
rect -1458 -799 -1446 -765
rect -1504 -805 -1446 -799
rect -1386 -765 -1328 -759
rect -1386 -799 -1374 -765
rect -1340 -799 -1328 -765
rect -1386 -805 -1328 -799
rect -1268 -765 -1210 -759
rect -1268 -799 -1256 -765
rect -1222 -799 -1210 -765
rect -1268 -805 -1210 -799
rect -1150 -765 -1092 -759
rect -1150 -799 -1138 -765
rect -1104 -799 -1092 -765
rect -1150 -805 -1092 -799
rect -1032 -765 -974 -759
rect -1032 -799 -1020 -765
rect -986 -799 -974 -765
rect -1032 -805 -974 -799
rect -914 -765 -856 -759
rect -914 -799 -902 -765
rect -868 -799 -856 -765
rect -914 -805 -856 -799
rect -796 -765 -738 -759
rect -796 -799 -784 -765
rect -750 -799 -738 -765
rect -796 -805 -738 -799
rect -678 -765 -620 -759
rect -678 -799 -666 -765
rect -632 -799 -620 -765
rect -678 -805 -620 -799
rect -560 -765 -502 -759
rect -560 -799 -548 -765
rect -514 -799 -502 -765
rect -560 -805 -502 -799
rect -442 -765 -384 -759
rect -442 -799 -430 -765
rect -396 -799 -384 -765
rect -442 -805 -384 -799
rect -324 -765 -266 -759
rect -324 -799 -312 -765
rect -278 -799 -266 -765
rect -324 -805 -266 -799
rect -206 -765 -148 -759
rect -206 -799 -194 -765
rect -160 -799 -148 -765
rect -206 -805 -148 -799
rect -88 -765 -30 -759
rect -88 -799 -76 -765
rect -42 -799 -30 -765
rect -88 -805 -30 -799
rect 30 -765 88 -759
rect 30 -799 42 -765
rect 76 -799 88 -765
rect 30 -805 88 -799
rect 148 -765 206 -759
rect 148 -799 160 -765
rect 194 -799 206 -765
rect 148 -805 206 -799
rect 266 -765 324 -759
rect 266 -799 278 -765
rect 312 -799 324 -765
rect 266 -805 324 -799
rect 384 -765 442 -759
rect 384 -799 396 -765
rect 430 -799 442 -765
rect 384 -805 442 -799
rect 502 -765 560 -759
rect 502 -799 514 -765
rect 548 -799 560 -765
rect 502 -805 560 -799
rect 620 -765 678 -759
rect 620 -799 632 -765
rect 666 -799 678 -765
rect 620 -805 678 -799
rect 738 -765 796 -759
rect 738 -799 750 -765
rect 784 -799 796 -765
rect 738 -805 796 -799
rect 856 -765 914 -759
rect 856 -799 868 -765
rect 902 -799 914 -765
rect 856 -805 914 -799
rect 974 -765 1032 -759
rect 974 -799 986 -765
rect 1020 -799 1032 -765
rect 974 -805 1032 -799
rect 1092 -765 1150 -759
rect 1092 -799 1104 -765
rect 1138 -799 1150 -765
rect 1092 -805 1150 -799
rect 1210 -765 1268 -759
rect 1210 -799 1222 -765
rect 1256 -799 1268 -765
rect 1210 -805 1268 -799
rect 1328 -765 1386 -759
rect 1328 -799 1340 -765
rect 1374 -799 1386 -765
rect 1328 -805 1386 -799
rect 1446 -765 1504 -759
rect 1446 -799 1458 -765
rect 1492 -799 1504 -765
rect 1446 -805 1504 -799
rect 1564 -765 1622 -759
rect 1564 -799 1576 -765
rect 1610 -799 1622 -765
rect 1564 -805 1622 -799
rect 1682 -765 1740 -759
rect 1682 -799 1694 -765
rect 1728 -799 1740 -765
rect 1682 -805 1740 -799
rect 1800 -765 1858 -759
rect 1800 -799 1812 -765
rect 1846 -799 1858 -765
rect 1800 -805 1858 -799
rect 1918 -765 1976 -759
rect 1918 -799 1930 -765
rect 1964 -799 1976 -765
rect 1918 -805 1976 -799
rect 2036 -765 2094 -759
rect 2036 -799 2048 -765
rect 2082 -799 2094 -765
rect 2036 -805 2094 -799
rect 2154 -765 2212 -759
rect 2154 -799 2166 -765
rect 2200 -799 2212 -765
rect 2154 -805 2212 -799
rect 2272 -765 2330 -759
rect 2272 -799 2284 -765
rect 2318 -799 2330 -765
rect 2272 -805 2330 -799
rect 2390 -765 2448 -759
rect 2390 -799 2402 -765
rect 2436 -799 2448 -765
rect 2390 -805 2448 -799
rect 2508 -765 2566 -759
rect 2508 -799 2520 -765
rect 2554 -799 2566 -765
rect 2508 -805 2566 -799
rect 2626 -765 2684 -759
rect 2626 -799 2638 -765
rect 2672 -799 2684 -765
rect 2626 -805 2684 -799
rect 2744 -765 2802 -759
rect 2744 -799 2756 -765
rect 2790 -799 2802 -765
rect 2744 -805 2802 -799
rect 2862 -765 2920 -759
rect 2862 -799 2874 -765
rect 2908 -799 2920 -765
rect 2862 -805 2920 -799
rect 2980 -765 3038 -759
rect 2980 -799 2992 -765
rect 3026 -799 3038 -765
rect 2980 -805 3038 -799
rect 3098 -765 3156 -759
rect 3098 -799 3110 -765
rect 3144 -799 3156 -765
rect 3098 -805 3156 -799
rect 3216 -765 3274 -759
rect 3216 -799 3228 -765
rect 3262 -799 3274 -765
rect 3216 -805 3274 -799
rect 3334 -765 3392 -759
rect 3334 -799 3346 -765
rect 3380 -799 3392 -765
rect 3334 -805 3392 -799
rect 3452 -765 3510 -759
rect 3452 -799 3464 -765
rect 3498 -799 3510 -765
rect 3452 -805 3510 -799
rect 3570 -765 3628 -759
rect 3570 -799 3582 -765
rect 3616 -799 3628 -765
rect 3570 -805 3628 -799
rect 3688 -765 3746 -759
rect 3688 -799 3700 -765
rect 3734 -799 3746 -765
rect 3688 -805 3746 -799
rect 3806 -765 3864 -759
rect 3806 -799 3818 -765
rect 3852 -799 3864 -765
rect 3806 -805 3864 -799
rect 3924 -765 3982 -759
rect 3924 -799 3936 -765
rect 3970 -799 3982 -765
rect 3924 -805 3982 -799
rect 4042 -765 4100 -759
rect 4042 -799 4054 -765
rect 4088 -799 4100 -765
rect 4042 -805 4100 -799
rect 4160 -765 4218 -759
rect 4160 -799 4172 -765
rect 4206 -799 4218 -765
rect 4160 -805 4218 -799
rect 4278 -765 4336 -759
rect 4278 -799 4290 -765
rect 4324 -799 4336 -765
rect 4278 -805 4336 -799
rect 4396 -765 4454 -759
rect 4396 -799 4408 -765
rect 4442 -799 4454 -765
rect 4396 -805 4454 -799
rect 4514 -765 4572 -759
rect 4514 -799 4526 -765
rect 4560 -799 4572 -765
rect 4514 -805 4572 -799
rect 4632 -765 4690 -759
rect 4632 -799 4644 -765
rect 4678 -799 4690 -765
rect 4632 -805 4690 -799
rect 4750 -765 4808 -759
rect 4750 -799 4762 -765
rect 4796 -799 4808 -765
rect 4750 -805 4808 -799
rect 4868 -765 4926 -759
rect 4868 -799 4880 -765
rect 4914 -799 4926 -765
rect 4868 -805 4926 -799
rect 4986 -765 5044 -759
rect 4986 -799 4998 -765
rect 5032 -799 5044 -765
rect 4986 -805 5044 -799
rect 5104 -765 5162 -759
rect 5104 -799 5116 -765
rect 5150 -799 5162 -765
rect 5104 -805 5162 -799
rect 5222 -765 5280 -759
rect 5222 -799 5234 -765
rect 5268 -799 5280 -765
rect 5222 -805 5280 -799
rect 5340 -765 5398 -759
rect 5340 -799 5352 -765
rect 5386 -799 5398 -765
rect 5340 -805 5398 -799
rect 5458 -765 5516 -759
rect 5458 -799 5470 -765
rect 5504 -799 5516 -765
rect 5458 -805 5516 -799
rect 5576 -765 5634 -759
rect 5576 -799 5588 -765
rect 5622 -799 5634 -765
rect 5576 -805 5634 -799
rect 5694 -765 5752 -759
rect 5694 -799 5706 -765
rect 5740 -799 5752 -765
rect 5694 -805 5752 -799
rect 5812 -765 5870 -759
rect 5812 -799 5824 -765
rect 5858 -799 5870 -765
rect 5812 -805 5870 -799
rect 5930 -765 5988 -759
rect 5930 -799 5942 -765
rect 5976 -799 5988 -765
rect 5930 -805 5988 -799
rect 6048 -765 6106 -759
rect 6048 -799 6060 -765
rect 6094 -799 6106 -765
rect 6048 -805 6106 -799
rect 6166 -765 6224 -759
rect 6166 -799 6178 -765
rect 6212 -799 6224 -765
rect 6166 -805 6224 -799
rect 6284 -765 6342 -759
rect 6284 -799 6296 -765
rect 6330 -799 6342 -765
rect 6284 -805 6342 -799
rect 6402 -765 6460 -759
rect 6402 -799 6414 -765
rect 6448 -799 6460 -765
rect 6402 -805 6460 -799
rect 6520 -765 6578 -759
rect 6520 -799 6532 -765
rect 6566 -799 6578 -765
rect 6520 -805 6578 -799
rect 6638 -765 6696 -759
rect 6638 -799 6650 -765
rect 6684 -799 6696 -765
rect 6638 -805 6696 -799
rect 6756 -765 6814 -759
rect 6756 -799 6768 -765
rect 6802 -799 6814 -765
rect 6756 -805 6814 -799
rect 6874 -765 6932 -759
rect 6874 -799 6886 -765
rect 6920 -799 6932 -765
rect 6874 -805 6932 -799
rect 6992 -765 7050 -759
rect 6992 -799 7004 -765
rect 7038 -799 7050 -765
rect 6992 -805 7050 -799
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -7194 -884 7194 884
string parameters w 3 l 0.3 m 2 nf 120 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
