magic
tech sky130A
magscale 12 1
timestamp 1598766404
<< metal5 >>
rect 0 15 15 105
rect 0 0 45 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
