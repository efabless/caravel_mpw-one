magic
tech sky130A
magscale 1 2
timestamp 1622226225
<< obsli1 >>
rect 48 197 14951 39549
<< obsm1 >>
rect 24 0 15000 39561
rect 15049 6891 17239 7665
rect 3331 -7 11313 0
rect 4099 -163 11313 -7
rect 15240 -163 17187 6891
rect 4099 -203 17187 -163
tri 3331 -603 3731 -203 se
rect 3731 -603 17187 -203
rect 3331 -1307 17187 -603
rect 3331 -1707 16387 -1307
tri 3331 -2107 3731 -1707 ne
rect 3731 -2107 16387 -1707
tri 16387 -2107 17187 -1307 nw
<< obsm2 >>
rect 98 8840 15000 38879
rect 98 7910 17228 8840
rect 98 0 15000 7910
rect 15049 6891 17239 7665
rect 100 -7 4099 0
rect 4185 -7 10707 0
rect 10819 -7 14940 0
<< metal3 >>
rect 100 -7 4900 1373
rect 10151 -7 14940 1373
<< obsm3 >>
rect 98 1453 15000 38714
rect 15121 7910 17228 8840
rect 15088 6939 17228 7632
rect 4980 0 10071 1453
rect 5200 -7 7376 0
rect 7676 -7 9851 0
<< metal4 >>
rect 0 34750 254 39593
rect 14746 34750 15000 39593
rect 0 13600 254 18593
rect 14746 13600 15000 18593
rect 0 12410 254 13300
rect 14746 12410 15000 13300
rect 0 11240 254 12130
rect 14746 11240 15000 12130
rect 0 10874 15000 10940
rect 0 10218 15000 10814
rect 0 9922 254 10158
rect 14746 9922 15000 10158
rect 0 9266 15000 9862
rect 0 9140 15000 9206
rect 0 7910 254 8840
rect 14746 7910 15000 8840
rect 0 6940 254 7630
rect 14746 6940 15000 7630
rect 0 5970 254 6660
rect 14746 5970 15000 6660
rect 0 4760 254 5690
rect 14746 4760 15000 5690
rect 0 3550 254 4480
rect 14746 3550 15000 4480
rect 0 2580 193 3270
rect 14807 2580 15000 3270
rect 0 1370 254 2300
rect 14746 1370 15000 2300
rect 0 0 254 1090
rect 14746 0 15000 1090
<< obsm4 >>
rect 334 34670 14666 39593
rect 193 18673 15000 34670
rect 334 13520 14666 18673
rect 193 13380 15000 13520
rect 334 12330 14666 13380
rect 193 12210 15000 12330
rect 334 11160 14666 12210
rect 193 11020 15000 11160
rect 334 9942 14666 10138
rect 193 8920 15000 9060
rect 334 7830 14666 8920
rect 15000 7910 17228 8840
rect 193 7710 15000 7830
rect 334 6860 14666 7710
rect 15000 6940 17233 7630
rect 193 6740 15000 6860
rect 334 5890 14666 6740
rect 193 5770 15000 5890
rect 334 4680 14666 5770
rect 193 4560 15000 4680
rect 334 3470 14666 4560
rect 193 3350 15000 3470
rect 273 2500 14727 3350
rect 193 2380 15000 2500
rect 334 1290 14666 2380
rect 193 1170 15000 1290
rect 334 0 14666 1170
<< metal5 >>
rect 2054 19973 12934 33426
rect 0 13600 254 18590
rect 0 12430 254 13280
rect 0 11260 254 12110
rect 0 9140 254 10940
rect 0 7930 254 8820
rect 0 6961 254 7610
rect 14746 13600 15000 18590
rect 14746 12430 15000 13280
rect 14746 11260 15000 12110
rect 14746 9140 15000 10940
rect 14746 7930 15000 8820
rect 14746 6961 15000 7610
rect 0 5990 254 6640
rect 0 4780 254 5670
rect 0 3570 254 4460
rect 14746 5990 15000 6640
rect 14746 4780 15000 5670
rect 14746 3570 15000 4460
rect 0 2600 193 3250
rect 14807 2600 15000 3250
rect 0 1390 254 2280
rect 0 20 254 1070
rect 14746 1390 15000 2280
rect 14746 20 15000 1070
<< obsm5 >>
rect 0 33746 15000 39593
rect 0 19653 1734 33746
rect 13254 19653 15000 33746
rect 0 18910 15000 19653
rect 574 6961 14426 18910
rect 0 6960 15000 6961
rect 574 3250 14426 6960
rect 513 2600 14487 3250
rect 574 20 14426 2600
<< labels >>
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VCCD
port 9 nsew power bidirectional
rlabel metal3 s 10151 -7 14940 1373 6 VCCD
port 9 nsew power bidirectional
rlabel metal3 s 100 -7 4900 1373 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 14845 34750 15000 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 34750 141 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 11 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 11 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 11 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 11 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 12 nsew ground bidirectional
<< properties >>
string LEFclass PAD POWER
string FIXED_BBOX 0 0 15000 39593
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 1552532
string GDS_END 1565676
string LEFview TRUE
<< end >>
