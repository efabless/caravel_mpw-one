magic
tech sky130A
magscale 1 2
timestamp 1606431493
<< metal3 >>
rect -5943 3222 -2061 3250
rect -5943 78 -2145 3222
rect -2081 78 -2061 3222
rect -5943 50 -2061 78
rect -1941 3222 1941 3250
rect -1941 78 1857 3222
rect 1921 78 1941 3222
rect -1941 50 1941 78
rect 2061 3222 5943 3250
rect 2061 78 5859 3222
rect 5923 78 5943 3222
rect 2061 50 5943 78
rect -5943 -78 -2061 -50
rect -5943 -3222 -2145 -78
rect -2081 -3222 -2061 -78
rect -5943 -3250 -2061 -3222
rect -1941 -78 1941 -50
rect -1941 -3222 1857 -78
rect 1921 -3222 1941 -78
rect -1941 -3250 1941 -3222
rect 2061 -78 5943 -50
rect 2061 -3222 5859 -78
rect 5923 -3222 5943 -78
rect 2061 -3250 5943 -3222
<< via3 >>
rect -2145 78 -2081 3222
rect 1857 78 1921 3222
rect 5859 78 5923 3222
rect -2145 -3222 -2081 -78
rect 1857 -3222 1921 -78
rect 5859 -3222 5923 -78
<< mimcap >>
rect -5843 3110 -2333 3150
rect -5843 190 -5803 3110
rect -2373 190 -2333 3110
rect -5843 150 -2333 190
rect -1841 3110 1669 3150
rect -1841 190 -1801 3110
rect 1629 190 1669 3110
rect -1841 150 1669 190
rect 2161 3110 5671 3150
rect 2161 190 2201 3110
rect 5631 190 5671 3110
rect 2161 150 5671 190
rect -5843 -190 -2333 -150
rect -5843 -3110 -5803 -190
rect -2373 -3110 -2333 -190
rect -5843 -3150 -2333 -3110
rect -1841 -190 1669 -150
rect -1841 -3110 -1801 -190
rect 1629 -3110 1669 -190
rect -1841 -3150 1669 -3110
rect 2161 -190 5671 -150
rect 2161 -3110 2201 -190
rect 5631 -3110 5671 -190
rect 2161 -3150 5671 -3110
<< mimcapcontact >>
rect -5803 190 -2373 3110
rect -1801 190 1629 3110
rect 2201 190 5631 3110
rect -5803 -3110 -2373 -190
rect -1801 -3110 1629 -190
rect 2201 -3110 5631 -190
<< metal4 >>
rect -4140 3111 -4036 3300
rect -2165 3222 -2061 3300
rect -5804 3110 -2372 3111
rect -5804 190 -5803 3110
rect -2373 190 -2372 3110
rect -5804 189 -2372 190
rect -4140 -189 -4036 189
rect -2165 78 -2145 3222
rect -2081 78 -2061 3222
rect -138 3111 -34 3300
rect 1837 3222 1941 3300
rect -1802 3110 1630 3111
rect -1802 190 -1801 3110
rect 1629 190 1630 3110
rect -1802 189 1630 190
rect -2165 -78 -2061 78
rect -5804 -190 -2372 -189
rect -5804 -3110 -5803 -190
rect -2373 -3110 -2372 -190
rect -5804 -3111 -2372 -3110
rect -4140 -3300 -4036 -3111
rect -2165 -3222 -2145 -78
rect -2081 -3222 -2061 -78
rect -138 -189 -34 189
rect 1837 78 1857 3222
rect 1921 78 1941 3222
rect 3864 3111 3968 3300
rect 5839 3222 5943 3300
rect 2200 3110 5632 3111
rect 2200 190 2201 3110
rect 5631 190 5632 3110
rect 2200 189 5632 190
rect 1837 -78 1941 78
rect -1802 -190 1630 -189
rect -1802 -3110 -1801 -190
rect 1629 -3110 1630 -190
rect -1802 -3111 1630 -3110
rect -2165 -3300 -2061 -3222
rect -138 -3300 -34 -3111
rect 1837 -3222 1857 -78
rect 1921 -3222 1941 -78
rect 3864 -189 3968 189
rect 5839 78 5859 3222
rect 5923 78 5943 3222
rect 5839 -78 5943 78
rect 2200 -190 5632 -189
rect 2200 -3110 2201 -190
rect 5631 -3110 5632 -190
rect 2200 -3111 5632 -3110
rect 1837 -3300 1941 -3222
rect 3864 -3300 3968 -3111
rect 5839 -3222 5859 -78
rect 5923 -3222 5943 -78
rect 5839 -3300 5943 -3222
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 2061 50 5771 3250
string parameters w 17.55 l 15.0 val 274.317 carea 1.00 cperi 0.17 nx 3 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string library sky130
<< end >>
