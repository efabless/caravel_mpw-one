magic
tech sky130A
magscale 1 2
timestamp 1607953902
<< obsli1 >>
rect 65257 17969 65659 18003
rect 65625 17940 65659 17969
rect 90649 17969 94639 18003
rect 90649 17940 90683 17969
rect 94605 17940 94639 17969
rect 1104 1071 198812 17940
<< obsm1 >>
rect 59262 18000 59326 18012
rect 65245 18000 65303 18009
rect 59262 17972 65303 18000
rect 59262 17960 59326 17972
rect 65245 17963 65303 17972
rect 65334 18000 65398 18012
rect 120166 18000 120230 18012
rect 65334 17972 120230 18000
rect 65334 17960 65398 17972
rect 120166 17960 120230 17972
rect 26510 17940 26574 17944
rect 94501 17940 94559 17941
rect 94593 17940 94651 17941
rect 95145 17940 95203 17941
rect 95234 17940 95298 17944
rect 150802 17940 150866 17944
rect 198 620 199810 17940
<< metal2 >>
rect 202 17940 258 18400
rect 570 17940 626 18400
rect 1030 17940 1086 18400
rect 1490 17940 1546 18400
rect 1858 17940 1914 18400
rect 2318 17940 2374 18400
rect 2778 17940 2834 18400
rect 3238 17940 3294 18400
rect 3606 17940 3662 18400
rect 4066 17940 4122 18400
rect 4526 17940 4582 18400
rect 4986 17940 5042 18400
rect 5354 17940 5410 18400
rect 5814 17940 5870 18400
rect 6274 17940 6330 18400
rect 6734 17940 6790 18400
rect 7102 17940 7158 18400
rect 7562 17940 7618 18400
rect 8022 17940 8078 18400
rect 8390 17940 8446 18400
rect 8850 17940 8906 18400
rect 9310 17940 9366 18400
rect 9770 17940 9826 18400
rect 10138 17940 10194 18400
rect 10598 17940 10654 18400
rect 11058 17940 11114 18400
rect 11518 17940 11574 18400
rect 11886 17940 11942 18400
rect 12346 17940 12402 18400
rect 12806 17940 12862 18400
rect 13266 17940 13322 18400
rect 13634 17940 13690 18400
rect 14094 17940 14150 18400
rect 14554 17940 14610 18400
rect 15014 17940 15070 18400
rect 15382 17940 15438 18400
rect 15842 17940 15898 18400
rect 16302 17940 16358 18400
rect 16670 17940 16726 18400
rect 17130 17940 17186 18400
rect 17590 17940 17646 18400
rect 18050 17940 18106 18400
rect 18418 17940 18474 18400
rect 18878 17940 18934 18400
rect 19338 17940 19394 18400
rect 19798 17940 19854 18400
rect 20166 17940 20222 18400
rect 20626 17940 20682 18400
rect 21086 17940 21142 18400
rect 21546 17940 21602 18400
rect 21914 17940 21970 18400
rect 22374 17940 22430 18400
rect 22834 17940 22890 18400
rect 23294 17940 23350 18400
rect 23662 17940 23718 18400
rect 24122 17940 24178 18400
rect 24582 17940 24638 18400
rect 24950 17940 25006 18400
rect 25410 17940 25466 18400
rect 25870 17940 25926 18400
rect 26330 17940 26386 18400
rect 26698 17940 26754 18400
rect 27158 17940 27214 18400
rect 27618 17940 27674 18400
rect 28078 17940 28134 18400
rect 28446 17940 28502 18400
rect 28906 17940 28962 18400
rect 29366 17940 29422 18400
rect 29826 17940 29882 18400
rect 30194 17940 30250 18400
rect 30654 17940 30710 18400
rect 31114 17940 31170 18400
rect 31574 17940 31630 18400
rect 31942 17940 31998 18400
rect 32402 17940 32458 18400
rect 32862 17940 32918 18400
rect 33230 17940 33286 18400
rect 33690 17940 33746 18400
rect 34150 17940 34206 18400
rect 34610 17940 34666 18400
rect 34978 17940 35034 18400
rect 35438 17940 35494 18400
rect 35898 17940 35954 18400
rect 36358 17940 36414 18400
rect 36726 17940 36782 18400
rect 37186 17940 37242 18400
rect 37646 17940 37702 18400
rect 38106 17940 38162 18400
rect 38474 17940 38530 18400
rect 38934 17940 38990 18400
rect 39394 17940 39450 18400
rect 39854 17940 39910 18400
rect 40222 17940 40278 18400
rect 40682 17940 40738 18400
rect 41142 17940 41198 18400
rect 41510 17940 41566 18400
rect 41970 17940 42026 18400
rect 42430 17940 42486 18400
rect 42890 17940 42946 18400
rect 43258 17940 43314 18400
rect 43718 17940 43774 18400
rect 44178 17940 44234 18400
rect 44638 17940 44694 18400
rect 45006 17940 45062 18400
rect 45466 17940 45522 18400
rect 45926 17940 45982 18400
rect 46386 17940 46442 18400
rect 46754 17940 46810 18400
rect 47214 17940 47270 18400
rect 47674 17940 47730 18400
rect 48134 17940 48190 18400
rect 48502 17940 48558 18400
rect 48962 17940 49018 18400
rect 49422 17940 49478 18400
rect 49790 17940 49846 18400
rect 50250 17940 50306 18400
rect 50710 17940 50766 18400
rect 51170 17940 51226 18400
rect 51538 17940 51594 18400
rect 51998 17940 52054 18400
rect 52458 17940 52514 18400
rect 52918 17940 52974 18400
rect 53286 17940 53342 18400
rect 53746 17940 53802 18400
rect 54206 17940 54262 18400
rect 54666 17940 54722 18400
rect 55034 17940 55090 18400
rect 55494 17940 55550 18400
rect 55954 17940 56010 18400
rect 56322 17940 56378 18400
rect 56782 17940 56838 18400
rect 57242 17940 57298 18400
rect 57702 17940 57758 18400
rect 58070 17940 58126 18400
rect 58530 17940 58586 18400
rect 58990 17940 59046 18400
rect 59450 17940 59506 18400
rect 59818 17940 59874 18400
rect 60278 17940 60334 18400
rect 60738 17940 60794 18400
rect 61198 17940 61254 18400
rect 61566 17940 61622 18400
rect 62026 17940 62082 18400
rect 62486 17940 62542 18400
rect 62946 17940 63002 18400
rect 63314 17940 63370 18400
rect 63774 17940 63830 18400
rect 64234 17940 64290 18400
rect 64602 17940 64658 18400
rect 65062 17940 65118 18400
rect 65522 17940 65578 18400
rect 65982 17940 66038 18400
rect 66350 17940 66406 18400
rect 66810 17940 66866 18400
rect 67270 17940 67326 18400
rect 67730 17940 67786 18400
rect 68098 17940 68154 18400
rect 68558 17940 68614 18400
rect 69018 17940 69074 18400
rect 69478 17940 69534 18400
rect 69846 17940 69902 18400
rect 70306 17940 70362 18400
rect 70766 17940 70822 18400
rect 71226 17940 71282 18400
rect 71594 17940 71650 18400
rect 72054 17940 72110 18400
rect 72514 17940 72570 18400
rect 72882 17940 72938 18400
rect 73342 17940 73398 18400
rect 73802 17940 73858 18400
rect 74262 17940 74318 18400
rect 74630 17940 74686 18400
rect 75090 17940 75146 18400
rect 75550 17940 75606 18400
rect 76010 17940 76066 18400
rect 76378 17940 76434 18400
rect 76838 17940 76894 18400
rect 77298 17940 77354 18400
rect 77758 17940 77814 18400
rect 78126 17940 78182 18400
rect 78586 17940 78642 18400
rect 79046 17940 79102 18400
rect 79506 17940 79562 18400
rect 79874 17940 79930 18400
rect 80334 17940 80390 18400
rect 80794 17940 80850 18400
rect 81162 17940 81218 18400
rect 81622 17940 81678 18400
rect 82082 17940 82138 18400
rect 82542 17940 82598 18400
rect 82910 17940 82966 18400
rect 83370 17940 83426 18400
rect 83830 17940 83886 18400
rect 84290 17940 84346 18400
rect 84658 17940 84714 18400
rect 85118 17940 85174 18400
rect 85578 17940 85634 18400
rect 86038 17940 86094 18400
rect 86406 17940 86462 18400
rect 86866 17940 86922 18400
rect 87326 17940 87382 18400
rect 87786 17940 87842 18400
rect 88154 17940 88210 18400
rect 88614 17940 88670 18400
rect 89074 17940 89130 18400
rect 89442 17940 89498 18400
rect 89902 17940 89958 18400
rect 90362 17940 90418 18400
rect 90822 17940 90878 18400
rect 91190 17940 91246 18400
rect 91650 17940 91706 18400
rect 92110 17940 92166 18400
rect 92570 17940 92626 18400
rect 92938 17940 92994 18400
rect 93398 17940 93454 18400
rect 93858 17940 93914 18400
rect 94318 17940 94374 18400
rect 94686 17940 94742 18400
rect 95146 17940 95202 18400
rect 95606 17940 95662 18400
rect 96066 17940 96122 18400
rect 96434 17940 96490 18400
rect 96894 17940 96950 18400
rect 97354 17940 97410 18400
rect 97722 17940 97778 18400
rect 98182 17940 98238 18400
rect 98642 17940 98698 18400
rect 99102 17940 99158 18400
rect 99470 17940 99526 18400
rect 99930 17940 99986 18400
rect 100390 17940 100446 18400
rect 100850 17940 100906 18400
rect 101218 17940 101274 18400
rect 101678 17940 101734 18400
rect 102138 17940 102194 18400
rect 102598 17940 102654 18400
rect 102966 17940 103022 18400
rect 103426 17940 103482 18400
rect 103886 17940 103942 18400
rect 104254 17940 104310 18400
rect 104714 17940 104770 18400
rect 105174 17940 105230 18400
rect 105634 17940 105690 18400
rect 106002 17940 106058 18400
rect 106462 17940 106518 18400
rect 106922 17940 106978 18400
rect 107382 17940 107438 18400
rect 107750 17940 107806 18400
rect 108210 17940 108266 18400
rect 108670 17940 108726 18400
rect 109130 17940 109186 18400
rect 109498 17940 109554 18400
rect 109958 17940 110014 18400
rect 110418 17940 110474 18400
rect 110878 17940 110934 18400
rect 111246 17940 111302 18400
rect 111706 17940 111762 18400
rect 112166 17940 112222 18400
rect 112534 17940 112590 18400
rect 112994 17940 113050 18400
rect 113454 17940 113510 18400
rect 113914 17940 113970 18400
rect 114282 17940 114338 18400
rect 114742 17940 114798 18400
rect 115202 17940 115258 18400
rect 115662 17940 115718 18400
rect 116030 17940 116086 18400
rect 116490 17940 116546 18400
rect 116950 17940 117006 18400
rect 117410 17940 117466 18400
rect 117778 17940 117834 18400
rect 118238 17940 118294 18400
rect 118698 17940 118754 18400
rect 119158 17940 119214 18400
rect 119526 17940 119582 18400
rect 119986 17940 120042 18400
rect 120446 17940 120502 18400
rect 120814 17940 120870 18400
rect 121274 17940 121330 18400
rect 121734 17940 121790 18400
rect 122194 17940 122250 18400
rect 122562 17940 122618 18400
rect 123022 17940 123078 18400
rect 123482 17940 123538 18400
rect 123942 17940 123998 18400
rect 124310 17940 124366 18400
rect 124770 17940 124826 18400
rect 125230 17940 125286 18400
rect 125690 17940 125746 18400
rect 126058 17940 126114 18400
rect 126518 17940 126574 18400
rect 126978 17940 127034 18400
rect 127438 17940 127494 18400
rect 127806 17940 127862 18400
rect 128266 17940 128322 18400
rect 128726 17940 128782 18400
rect 129094 17940 129150 18400
rect 129554 17940 129610 18400
rect 130014 17940 130070 18400
rect 130474 17940 130530 18400
rect 130842 17940 130898 18400
rect 131302 17940 131358 18400
rect 131762 17940 131818 18400
rect 132222 17940 132278 18400
rect 132590 17940 132646 18400
rect 133050 17940 133106 18400
rect 133510 17940 133566 18400
rect 133970 17940 134026 18400
rect 134338 17940 134394 18400
rect 134798 17940 134854 18400
rect 135258 17940 135314 18400
rect 135718 17940 135774 18400
rect 136086 17940 136142 18400
rect 136546 17940 136602 18400
rect 137006 17940 137062 18400
rect 137374 17940 137430 18400
rect 137834 17940 137890 18400
rect 138294 17940 138350 18400
rect 138754 17940 138810 18400
rect 139122 17940 139178 18400
rect 139582 17940 139638 18400
rect 140042 17940 140098 18400
rect 140502 17940 140558 18400
rect 140870 17940 140926 18400
rect 141330 17940 141386 18400
rect 141790 17940 141846 18400
rect 142250 17940 142306 18400
rect 142618 17940 142674 18400
rect 143078 17940 143134 18400
rect 143538 17940 143594 18400
rect 143998 17940 144054 18400
rect 144366 17940 144422 18400
rect 144826 17940 144882 18400
rect 145286 17940 145342 18400
rect 145654 17940 145710 18400
rect 146114 17940 146170 18400
rect 146574 17940 146630 18400
rect 147034 17940 147090 18400
rect 147402 17940 147458 18400
rect 147862 17940 147918 18400
rect 148322 17940 148378 18400
rect 148782 17940 148838 18400
rect 149150 17940 149206 18400
rect 149610 17940 149666 18400
rect 150070 17940 150126 18400
rect 150530 17940 150586 18400
rect 150898 17940 150954 18400
rect 151358 17940 151414 18400
rect 151818 17940 151874 18400
rect 152186 17940 152242 18400
rect 152646 17940 152702 18400
rect 153106 17940 153162 18400
rect 153566 17940 153622 18400
rect 153934 17940 153990 18400
rect 154394 17940 154450 18400
rect 154854 17940 154910 18400
rect 155314 17940 155370 18400
rect 155682 17940 155738 18400
rect 156142 17940 156198 18400
rect 156602 17940 156658 18400
rect 157062 17940 157118 18400
rect 157430 17940 157486 18400
rect 157890 17940 157946 18400
rect 158350 17940 158406 18400
rect 158810 17940 158866 18400
rect 159178 17940 159234 18400
rect 159638 17940 159694 18400
rect 160098 17940 160154 18400
rect 160466 17940 160522 18400
rect 160926 17940 160982 18400
rect 161386 17940 161442 18400
rect 161846 17940 161902 18400
rect 162214 17940 162270 18400
rect 162674 17940 162730 18400
rect 163134 17940 163190 18400
rect 163594 17940 163650 18400
rect 163962 17940 164018 18400
rect 164422 17940 164478 18400
rect 164882 17940 164938 18400
rect 165342 17940 165398 18400
rect 165710 17940 165766 18400
rect 166170 17940 166226 18400
rect 166630 17940 166686 18400
rect 167090 17940 167146 18400
rect 167458 17940 167514 18400
rect 167918 17940 167974 18400
rect 168378 17940 168434 18400
rect 168746 17940 168802 18400
rect 169206 17940 169262 18400
rect 169666 17940 169722 18400
rect 170126 17940 170182 18400
rect 170494 17940 170550 18400
rect 170954 17940 171010 18400
rect 171414 17940 171470 18400
rect 171874 17940 171930 18400
rect 172242 17940 172298 18400
rect 172702 17940 172758 18400
rect 173162 17940 173218 18400
rect 173622 17940 173678 18400
rect 173990 17940 174046 18400
rect 174450 17940 174506 18400
rect 174910 17940 174966 18400
rect 175370 17940 175426 18400
rect 175738 17940 175794 18400
rect 176198 17940 176254 18400
rect 176658 17940 176714 18400
rect 177026 17940 177082 18400
rect 177486 17940 177542 18400
rect 177946 17940 178002 18400
rect 178406 17940 178462 18400
rect 178774 17940 178830 18400
rect 179234 17940 179290 18400
rect 179694 17940 179750 18400
rect 180154 17940 180210 18400
rect 180522 17940 180578 18400
rect 180982 17940 181038 18400
rect 181442 17940 181498 18400
rect 181902 17940 181958 18400
rect 182270 17940 182326 18400
rect 182730 17940 182786 18400
rect 183190 17940 183246 18400
rect 183650 17940 183706 18400
rect 184018 17940 184074 18400
rect 184478 17940 184534 18400
rect 184938 17940 184994 18400
rect 185306 17940 185362 18400
rect 185766 17940 185822 18400
rect 186226 17940 186282 18400
rect 186686 17940 186742 18400
rect 187054 17940 187110 18400
rect 187514 17940 187570 18400
rect 187974 17940 188030 18400
rect 188434 17940 188490 18400
rect 188802 17940 188858 18400
rect 189262 17940 189318 18400
rect 189722 17940 189778 18400
rect 190182 17940 190238 18400
rect 190550 17940 190606 18400
rect 191010 17940 191066 18400
rect 191470 17940 191526 18400
rect 191930 17940 191986 18400
rect 192298 17940 192354 18400
rect 192758 17940 192814 18400
rect 193218 17940 193274 18400
rect 193586 17940 193642 18400
rect 194046 17940 194102 18400
rect 194506 17940 194562 18400
rect 194966 17940 195022 18400
rect 195334 17940 195390 18400
rect 195794 17940 195850 18400
rect 196254 17940 196310 18400
rect 196714 17940 196770 18400
rect 197082 17940 197138 18400
rect 197542 17940 197598 18400
rect 198002 17940 198058 18400
rect 198462 17940 198518 18400
rect 198830 17940 198886 18400
rect 199290 17940 199346 18400
rect 199750 17940 199806 18400
rect 202 -400 258 60
rect 570 -400 626 60
rect 1030 -400 1086 60
rect 1490 -400 1546 60
rect 1858 -400 1914 60
rect 2318 -400 2374 60
rect 2778 -400 2834 60
rect 3238 -400 3294 60
rect 3606 -400 3662 60
rect 4066 -400 4122 60
rect 4526 -400 4582 60
rect 4986 -400 5042 60
rect 5354 -400 5410 60
rect 5814 -400 5870 60
rect 6274 -400 6330 60
rect 6734 -400 6790 60
rect 7102 -400 7158 60
rect 7562 -400 7618 60
rect 8022 -400 8078 60
rect 8390 -400 8446 60
rect 8850 -400 8906 60
rect 9310 -400 9366 60
rect 9770 -400 9826 60
rect 10138 -400 10194 60
rect 10598 -400 10654 60
rect 11058 -400 11114 60
rect 11518 -400 11574 60
rect 11886 -400 11942 60
rect 12346 -400 12402 60
rect 12806 -400 12862 60
rect 13266 -400 13322 60
rect 13634 -400 13690 60
rect 14094 -400 14150 60
rect 14554 -400 14610 60
rect 15014 -400 15070 60
rect 15382 -400 15438 60
rect 15842 -400 15898 60
rect 16302 -400 16358 60
rect 16670 -400 16726 60
rect 17130 -400 17186 60
rect 17590 -400 17646 60
rect 18050 -400 18106 60
rect 18418 -400 18474 60
rect 18878 -400 18934 60
rect 19338 -400 19394 60
rect 19798 -400 19854 60
rect 20166 -400 20222 60
rect 20626 -400 20682 60
rect 21086 -400 21142 60
rect 21546 -400 21602 60
rect 21914 -400 21970 60
rect 22374 -400 22430 60
rect 22834 -400 22890 60
rect 23294 -400 23350 60
rect 23662 -400 23718 60
rect 24122 -400 24178 60
rect 24582 -400 24638 60
rect 24950 -400 25006 60
rect 25410 -400 25466 60
rect 25870 -400 25926 60
rect 26330 -400 26386 60
rect 26698 -400 26754 60
rect 27158 -400 27214 60
rect 27618 -400 27674 60
rect 28078 -400 28134 60
rect 28446 -400 28502 60
rect 28906 -400 28962 60
rect 29366 -400 29422 60
rect 29826 -400 29882 60
rect 30194 -400 30250 60
rect 30654 -400 30710 60
rect 31114 -400 31170 60
rect 31574 -400 31630 60
rect 31942 -400 31998 60
rect 32402 -400 32458 60
rect 32862 -400 32918 60
rect 33230 -400 33286 60
rect 33690 -400 33746 60
rect 34150 -400 34206 60
rect 34610 -400 34666 60
rect 34978 -400 35034 60
rect 35438 -400 35494 60
rect 35898 -400 35954 60
rect 36358 -400 36414 60
rect 36726 -400 36782 60
rect 37186 -400 37242 60
rect 37646 -400 37702 60
rect 38106 -400 38162 60
rect 38474 -400 38530 60
rect 38934 -400 38990 60
rect 39394 -400 39450 60
rect 39854 -400 39910 60
rect 40222 -400 40278 60
rect 40682 -400 40738 60
rect 41142 -400 41198 60
rect 41510 -400 41566 60
rect 41970 -400 42026 60
rect 42430 -400 42486 60
rect 42890 -400 42946 60
rect 43258 -400 43314 60
rect 43718 -400 43774 60
rect 44178 -400 44234 60
rect 44638 -400 44694 60
rect 45006 -400 45062 60
rect 45466 -400 45522 60
rect 45926 -400 45982 60
rect 46386 -400 46442 60
rect 46754 -400 46810 60
rect 47214 -400 47270 60
rect 47674 -400 47730 60
rect 48134 -400 48190 60
rect 48502 -400 48558 60
rect 48962 -400 49018 60
rect 49422 -400 49478 60
rect 49790 -400 49846 60
rect 50250 -400 50306 60
rect 50710 -400 50766 60
rect 51170 -400 51226 60
rect 51538 -400 51594 60
rect 51998 -400 52054 60
rect 52458 -400 52514 60
rect 52918 -400 52974 60
rect 53286 -400 53342 60
rect 53746 -400 53802 60
rect 54206 -400 54262 60
rect 54666 -400 54722 60
rect 55034 -400 55090 60
rect 55494 -400 55550 60
rect 55954 -400 56010 60
rect 56322 -400 56378 60
rect 56782 -400 56838 60
rect 57242 -400 57298 60
rect 57702 -400 57758 60
rect 58070 -400 58126 60
rect 58530 -400 58586 60
rect 58990 -400 59046 60
rect 59450 -400 59506 60
rect 59818 -400 59874 60
rect 60278 -400 60334 60
rect 60738 -400 60794 60
rect 61198 -400 61254 60
rect 61566 -400 61622 60
rect 62026 -400 62082 60
rect 62486 -400 62542 60
rect 62946 -400 63002 60
rect 63314 -400 63370 60
rect 63774 -400 63830 60
rect 64234 -400 64290 60
rect 64602 -400 64658 60
rect 65062 -400 65118 60
rect 65522 -400 65578 60
rect 65982 -400 66038 60
rect 66350 -400 66406 60
rect 66810 -400 66866 60
rect 67270 -400 67326 60
rect 67730 -400 67786 60
rect 68098 -400 68154 60
rect 68558 -400 68614 60
rect 69018 -400 69074 60
rect 69478 -400 69534 60
rect 69846 -400 69902 60
rect 70306 -400 70362 60
rect 70766 -400 70822 60
rect 71226 -400 71282 60
rect 71594 -400 71650 60
rect 72054 -400 72110 60
rect 72514 -400 72570 60
rect 72882 -400 72938 60
rect 73342 -400 73398 60
rect 73802 -400 73858 60
rect 74262 -400 74318 60
rect 74630 -400 74686 60
rect 75090 -400 75146 60
rect 75550 -400 75606 60
rect 76010 -400 76066 60
rect 76378 -400 76434 60
rect 76838 -400 76894 60
rect 77298 -400 77354 60
rect 77758 -400 77814 60
rect 78126 -400 78182 60
rect 78586 -400 78642 60
rect 79046 -400 79102 60
rect 79506 -400 79562 60
rect 79874 -400 79930 60
rect 80334 -400 80390 60
rect 80794 -400 80850 60
rect 81162 -400 81218 60
rect 81622 -400 81678 60
rect 82082 -400 82138 60
rect 82542 -400 82598 60
rect 82910 -400 82966 60
rect 83370 -400 83426 60
rect 83830 -400 83886 60
rect 84290 -400 84346 60
rect 84658 -400 84714 60
rect 85118 -400 85174 60
rect 85578 -400 85634 60
rect 86038 -400 86094 60
rect 86406 -400 86462 60
rect 86866 -400 86922 60
rect 87326 -400 87382 60
rect 87786 -400 87842 60
rect 88154 -400 88210 60
rect 88614 -400 88670 60
rect 89074 -400 89130 60
rect 89442 -400 89498 60
rect 89902 -400 89958 60
rect 90362 -400 90418 60
rect 90822 -400 90878 60
rect 91190 -400 91246 60
rect 91650 -400 91706 60
rect 92110 -400 92166 60
rect 92570 -400 92626 60
rect 92938 -400 92994 60
rect 93398 -400 93454 60
rect 93858 -400 93914 60
rect 94318 -400 94374 60
rect 94686 -400 94742 60
rect 95146 -400 95202 60
rect 95606 -400 95662 60
rect 96066 -400 96122 60
rect 96434 -400 96490 60
rect 96894 -400 96950 60
rect 97354 -400 97410 60
rect 97722 -400 97778 60
rect 98182 -400 98238 60
rect 98642 -400 98698 60
rect 99102 -400 99158 60
rect 99470 -400 99526 60
rect 99930 -400 99986 60
rect 100390 -400 100446 60
rect 100850 -400 100906 60
rect 101218 -400 101274 60
rect 101678 -400 101734 60
rect 102138 -400 102194 60
rect 102598 -400 102654 60
rect 102966 -400 103022 60
rect 103426 -400 103482 60
rect 103886 -400 103942 60
rect 104254 -400 104310 60
rect 104714 -400 104770 60
rect 105174 -400 105230 60
rect 105634 -400 105690 60
rect 106002 -400 106058 60
rect 106462 -400 106518 60
rect 106922 -400 106978 60
rect 107382 -400 107438 60
rect 107750 -400 107806 60
rect 108210 -400 108266 60
rect 108670 -400 108726 60
rect 109130 -400 109186 60
rect 109498 -400 109554 60
rect 109958 -400 110014 60
rect 110418 -400 110474 60
rect 110878 -400 110934 60
rect 111246 -400 111302 60
rect 111706 -400 111762 60
rect 112166 -400 112222 60
rect 112534 -400 112590 60
rect 112994 -400 113050 60
rect 113454 -400 113510 60
rect 113914 -400 113970 60
rect 114282 -400 114338 60
rect 114742 -400 114798 60
rect 115202 -400 115258 60
rect 115662 -400 115718 60
rect 116030 -400 116086 60
rect 116490 -400 116546 60
rect 116950 -400 117006 60
rect 117410 -400 117466 60
rect 117778 -400 117834 60
rect 118238 -400 118294 60
rect 118698 -400 118754 60
rect 119158 -400 119214 60
rect 119526 -400 119582 60
rect 119986 -400 120042 60
rect 120446 -400 120502 60
rect 120814 -400 120870 60
rect 121274 -400 121330 60
rect 121734 -400 121790 60
rect 122194 -400 122250 60
rect 122562 -400 122618 60
rect 123022 -400 123078 60
rect 123482 -400 123538 60
rect 123942 -400 123998 60
rect 124310 -400 124366 60
rect 124770 -400 124826 60
rect 125230 -400 125286 60
rect 125690 -400 125746 60
rect 126058 -400 126114 60
rect 126518 -400 126574 60
rect 126978 -400 127034 60
rect 127438 -400 127494 60
rect 127806 -400 127862 60
rect 128266 -400 128322 60
rect 128726 -400 128782 60
rect 129094 -400 129150 60
rect 129554 -400 129610 60
rect 130014 -400 130070 60
rect 130474 -400 130530 60
rect 130842 -400 130898 60
rect 131302 -400 131358 60
rect 131762 -400 131818 60
rect 132222 -400 132278 60
rect 132590 -400 132646 60
rect 133050 -400 133106 60
rect 133510 -400 133566 60
rect 133970 -400 134026 60
rect 134338 -400 134394 60
rect 134798 -400 134854 60
rect 135258 -400 135314 60
rect 135718 -400 135774 60
rect 136086 -400 136142 60
rect 136546 -400 136602 60
rect 137006 -400 137062 60
rect 137374 -400 137430 60
rect 137834 -400 137890 60
rect 138294 -400 138350 60
rect 138754 -400 138810 60
rect 139122 -400 139178 60
rect 139582 -400 139638 60
rect 140042 -400 140098 60
rect 140502 -400 140558 60
rect 140870 -400 140926 60
rect 141330 -400 141386 60
rect 141790 -400 141846 60
rect 142250 -400 142306 60
rect 142618 -400 142674 60
rect 143078 -400 143134 60
rect 143538 -400 143594 60
rect 143998 -400 144054 60
rect 144366 -400 144422 60
rect 144826 -400 144882 60
rect 145286 -400 145342 60
rect 145654 -400 145710 60
rect 146114 -400 146170 60
rect 146574 -400 146630 60
rect 147034 -400 147090 60
rect 147402 -400 147458 60
rect 147862 -400 147918 60
rect 148322 -400 148378 60
rect 148782 -400 148838 60
rect 149150 -400 149206 60
rect 149610 -400 149666 60
rect 150070 -400 150126 60
rect 150530 -400 150586 60
rect 150898 -400 150954 60
rect 151358 -400 151414 60
rect 151818 -400 151874 60
rect 152186 -400 152242 60
rect 152646 -400 152702 60
rect 153106 -400 153162 60
rect 153566 -400 153622 60
rect 153934 -400 153990 60
rect 154394 -400 154450 60
rect 154854 -400 154910 60
rect 155314 -400 155370 60
rect 155682 -400 155738 60
rect 156142 -400 156198 60
rect 156602 -400 156658 60
rect 157062 -400 157118 60
rect 157430 -400 157486 60
rect 157890 -400 157946 60
rect 158350 -400 158406 60
rect 158810 -400 158866 60
rect 159178 -400 159234 60
rect 159638 -400 159694 60
rect 160098 -400 160154 60
rect 160466 -400 160522 60
rect 160926 -400 160982 60
rect 161386 -400 161442 60
rect 161846 -400 161902 60
rect 162214 -400 162270 60
rect 162674 -400 162730 60
rect 163134 -400 163190 60
rect 163594 -400 163650 60
rect 163962 -400 164018 60
rect 164422 -400 164478 60
rect 164882 -400 164938 60
rect 165342 -400 165398 60
rect 165710 -400 165766 60
rect 166170 -400 166226 60
rect 166630 -400 166686 60
rect 167090 -400 167146 60
rect 167458 -400 167514 60
rect 167918 -400 167974 60
rect 168378 -400 168434 60
rect 168746 -400 168802 60
rect 169206 -400 169262 60
rect 169666 -400 169722 60
rect 170126 -400 170182 60
rect 170494 -400 170550 60
rect 170954 -400 171010 60
rect 171414 -400 171470 60
rect 171874 -400 171930 60
rect 172242 -400 172298 60
rect 172702 -400 172758 60
rect 173162 -400 173218 60
rect 173622 -400 173678 60
rect 173990 -400 174046 60
rect 174450 -400 174506 60
rect 174910 -400 174966 60
rect 175370 -400 175426 60
rect 175738 -400 175794 60
rect 176198 -400 176254 60
rect 176658 -400 176714 60
rect 177026 -400 177082 60
rect 177486 -400 177542 60
rect 177946 -400 178002 60
rect 178406 -400 178462 60
rect 178774 -400 178830 60
rect 179234 -400 179290 60
rect 179694 -400 179750 60
rect 180154 -400 180210 60
rect 180522 -400 180578 60
rect 180982 -400 181038 60
rect 181442 -400 181498 60
rect 181902 -400 181958 60
rect 182270 -400 182326 60
rect 182730 -400 182786 60
rect 183190 -400 183246 60
rect 183650 -400 183706 60
rect 184018 -400 184074 60
rect 184478 -400 184534 60
rect 184938 -400 184994 60
rect 185306 -400 185362 60
rect 185766 -400 185822 60
rect 186226 -400 186282 60
rect 186686 -400 186742 60
rect 187054 -400 187110 60
rect 187514 -400 187570 60
rect 187974 -400 188030 60
rect 188434 -400 188490 60
rect 188802 -400 188858 60
rect 189262 -400 189318 60
rect 189722 -400 189778 60
rect 190182 -400 190238 60
rect 190550 -400 190606 60
rect 191010 -400 191066 60
rect 191470 -400 191526 60
rect 191930 -400 191986 60
rect 192298 -400 192354 60
rect 192758 -400 192814 60
rect 193218 -400 193274 60
rect 193586 -400 193642 60
rect 194046 -400 194102 60
rect 194506 -400 194562 60
rect 194966 -400 195022 60
rect 195334 -400 195390 60
rect 195794 -400 195850 60
rect 196254 -400 196310 60
rect 196714 -400 196770 60
rect 197082 -400 197138 60
rect 197542 -400 197598 60
rect 198002 -400 198058 60
rect 198462 -400 198518 60
rect 198830 -400 198886 60
rect 199290 -400 199346 60
rect 199750 -400 199806 60
<< obsm2 >>
rect 26516 17940 26568 17950
rect 59268 17954 59320 18018
rect 59280 17940 59308 17954
rect 65340 17954 65392 18018
rect 65352 17940 65380 17954
rect 95240 17940 95292 17950
rect 120172 17954 120224 18018
rect 120184 17940 120212 17954
rect 150808 17940 150860 17950
rect 202 60 199806 17940
<< metal3 >>
rect 22504 19554 22512 19556
rect -1586 19494 22512 19554
rect 22504 19492 22512 19494
rect 22576 19492 22592 19556
rect 22656 19492 22672 19556
rect 22736 19554 22744 19556
rect 52504 19554 52512 19556
rect 22736 19494 52512 19554
rect 22736 19492 22744 19494
rect 52504 19492 52512 19494
rect 52576 19492 52592 19556
rect 52656 19492 52672 19556
rect 52736 19554 52744 19556
rect 82504 19554 82512 19556
rect 52736 19494 82512 19554
rect 52736 19492 52744 19494
rect 82504 19492 82512 19494
rect 82576 19492 82592 19556
rect 82656 19492 82672 19556
rect 82736 19554 82744 19556
rect 112504 19554 112512 19556
rect 82736 19494 112512 19554
rect 82736 19492 82744 19494
rect 112504 19492 112512 19494
rect 112576 19492 112592 19556
rect 112656 19492 112672 19556
rect 112736 19554 112744 19556
rect 142504 19554 142512 19556
rect 112736 19494 142512 19554
rect 112736 19492 112744 19494
rect 142504 19492 142512 19494
rect 142576 19492 142592 19556
rect 142656 19492 142672 19556
rect 142736 19554 142744 19556
rect 172504 19554 172512 19556
rect 142736 19494 172512 19554
rect 142736 19492 142744 19494
rect 172504 19492 172512 19494
rect 172576 19492 172592 19556
rect 172656 19492 172672 19556
rect 172736 19554 172744 19556
rect 172736 19494 201502 19554
rect 172736 19492 172744 19494
rect 7504 19414 7512 19416
rect -1446 19354 7512 19414
rect 7504 19352 7512 19354
rect 7576 19352 7592 19416
rect 7656 19352 7672 19416
rect 7736 19414 7744 19416
rect 37504 19414 37512 19416
rect 7736 19354 37512 19414
rect 7736 19352 7744 19354
rect 37504 19352 37512 19354
rect 37576 19352 37592 19416
rect 37656 19352 37672 19416
rect 37736 19414 37744 19416
rect 67504 19414 67512 19416
rect 37736 19354 67512 19414
rect 37736 19352 37744 19354
rect 67504 19352 67512 19354
rect 67576 19352 67592 19416
rect 67656 19352 67672 19416
rect 67736 19414 67744 19416
rect 97504 19414 97512 19416
rect 67736 19354 97512 19414
rect 67736 19352 67744 19354
rect 97504 19352 97512 19354
rect 97576 19352 97592 19416
rect 97656 19352 97672 19416
rect 97736 19414 97744 19416
rect 127504 19414 127512 19416
rect 97736 19354 127512 19414
rect 97736 19352 97744 19354
rect 127504 19352 127512 19354
rect 127576 19352 127592 19416
rect 127656 19352 127672 19416
rect 127736 19414 127744 19416
rect 157504 19414 157512 19416
rect 127736 19354 157512 19414
rect 127736 19352 127744 19354
rect 157504 19352 157512 19354
rect 157576 19352 157592 19416
rect 157656 19352 157672 19416
rect 157736 19414 157744 19416
rect 187504 19414 187512 19416
rect 157736 19354 187512 19414
rect 157736 19352 157744 19354
rect 187504 19352 187512 19354
rect 187576 19352 187592 19416
rect 187656 19352 187672 19416
rect 187736 19414 187744 19416
rect 187736 19354 201362 19414
rect 187736 19352 187744 19354
rect 21624 19274 21632 19276
rect -1306 19214 21632 19274
rect 21624 19212 21632 19214
rect 21696 19212 21712 19276
rect 21776 19212 21792 19276
rect 21856 19274 21864 19276
rect 51624 19274 51632 19276
rect 21856 19214 51632 19274
rect 21856 19212 21864 19214
rect 51624 19212 51632 19214
rect 51696 19212 51712 19276
rect 51776 19212 51792 19276
rect 51856 19274 51864 19276
rect 81624 19274 81632 19276
rect 51856 19214 81632 19274
rect 51856 19212 51864 19214
rect 81624 19212 81632 19214
rect 81696 19212 81712 19276
rect 81776 19212 81792 19276
rect 81856 19274 81864 19276
rect 111624 19274 111632 19276
rect 81856 19214 111632 19274
rect 81856 19212 81864 19214
rect 111624 19212 111632 19214
rect 111696 19212 111712 19276
rect 111776 19212 111792 19276
rect 111856 19274 111864 19276
rect 141624 19274 141632 19276
rect 111856 19214 141632 19274
rect 111856 19212 111864 19214
rect 141624 19212 141632 19214
rect 141696 19212 141712 19276
rect 141776 19212 141792 19276
rect 141856 19274 141864 19276
rect 171624 19274 171632 19276
rect 141856 19214 171632 19274
rect 141856 19212 141864 19214
rect 171624 19212 171632 19214
rect 171696 19212 171712 19276
rect 171776 19212 171792 19276
rect 171856 19274 171864 19276
rect 171856 19214 201222 19274
rect 171856 19212 171864 19214
rect 6624 19134 6632 19136
rect -1166 19074 6632 19134
rect 6624 19072 6632 19074
rect 6696 19072 6712 19136
rect 6776 19072 6792 19136
rect 6856 19134 6864 19136
rect 36624 19134 36632 19136
rect 6856 19074 36632 19134
rect 6856 19072 6864 19074
rect 36624 19072 36632 19074
rect 36696 19072 36712 19136
rect 36776 19072 36792 19136
rect 36856 19134 36864 19136
rect 66624 19134 66632 19136
rect 36856 19074 66632 19134
rect 36856 19072 36864 19074
rect 66624 19072 66632 19074
rect 66696 19072 66712 19136
rect 66776 19072 66792 19136
rect 66856 19134 66864 19136
rect 96624 19134 96632 19136
rect 66856 19074 96632 19134
rect 66856 19072 66864 19074
rect 96624 19072 96632 19074
rect 96696 19072 96712 19136
rect 96776 19072 96792 19136
rect 96856 19134 96864 19136
rect 126624 19134 126632 19136
rect 96856 19074 126632 19134
rect 96856 19072 96864 19074
rect 126624 19072 126632 19074
rect 126696 19072 126712 19136
rect 126776 19072 126792 19136
rect 126856 19134 126864 19136
rect 156624 19134 156632 19136
rect 126856 19074 156632 19134
rect 126856 19072 126864 19074
rect 156624 19072 156632 19074
rect 156696 19072 156712 19136
rect 156776 19072 156792 19136
rect 156856 19134 156864 19136
rect 186624 19134 186632 19136
rect 156856 19074 186632 19134
rect 156856 19072 156864 19074
rect 186624 19072 186632 19074
rect 186696 19072 186712 19136
rect 186776 19072 186792 19136
rect 186856 19134 186864 19136
rect 186856 19074 201082 19134
rect 186856 19072 186864 19074
rect 20744 18994 20752 18996
rect -1026 18934 20752 18994
rect 20744 18932 20752 18934
rect 20816 18932 20832 18996
rect 20896 18932 20912 18996
rect 20976 18994 20984 18996
rect 50744 18994 50752 18996
rect 20976 18934 50752 18994
rect 20976 18932 20984 18934
rect 50744 18932 50752 18934
rect 50816 18932 50832 18996
rect 50896 18932 50912 18996
rect 50976 18994 50984 18996
rect 80744 18994 80752 18996
rect 50976 18934 80752 18994
rect 50976 18932 50984 18934
rect 80744 18932 80752 18934
rect 80816 18932 80832 18996
rect 80896 18932 80912 18996
rect 80976 18994 80984 18996
rect 110744 18994 110752 18996
rect 80976 18934 110752 18994
rect 80976 18932 80984 18934
rect 110744 18932 110752 18934
rect 110816 18932 110832 18996
rect 110896 18932 110912 18996
rect 110976 18994 110984 18996
rect 140744 18994 140752 18996
rect 110976 18934 140752 18994
rect 110976 18932 110984 18934
rect 140744 18932 140752 18934
rect 140816 18932 140832 18996
rect 140896 18932 140912 18996
rect 140976 18994 140984 18996
rect 170744 18994 170752 18996
rect 140976 18934 170752 18994
rect 140976 18932 140984 18934
rect 170744 18932 170752 18934
rect 170816 18932 170832 18996
rect 170896 18932 170912 18996
rect 170976 18994 170984 18996
rect 170976 18934 200942 18994
rect 170976 18932 170984 18934
rect 5744 18854 5752 18856
rect -886 18794 5752 18854
rect 5744 18792 5752 18794
rect 5816 18792 5832 18856
rect 5896 18792 5912 18856
rect 5976 18854 5984 18856
rect 35744 18854 35752 18856
rect 5976 18794 35752 18854
rect 5976 18792 5984 18794
rect 35744 18792 35752 18794
rect 35816 18792 35832 18856
rect 35896 18792 35912 18856
rect 35976 18854 35984 18856
rect 65744 18854 65752 18856
rect 35976 18794 65752 18854
rect 35976 18792 35984 18794
rect 65744 18792 65752 18794
rect 65816 18792 65832 18856
rect 65896 18792 65912 18856
rect 65976 18854 65984 18856
rect 95744 18854 95752 18856
rect 65976 18794 95752 18854
rect 65976 18792 65984 18794
rect 95744 18792 95752 18794
rect 95816 18792 95832 18856
rect 95896 18792 95912 18856
rect 95976 18854 95984 18856
rect 125744 18854 125752 18856
rect 95976 18794 125752 18854
rect 95976 18792 95984 18794
rect 125744 18792 125752 18794
rect 125816 18792 125832 18856
rect 125896 18792 125912 18856
rect 125976 18854 125984 18856
rect 155744 18854 155752 18856
rect 125976 18794 155752 18854
rect 125976 18792 125984 18794
rect 155744 18792 155752 18794
rect 155816 18792 155832 18856
rect 155896 18792 155912 18856
rect 155976 18854 155984 18856
rect 185744 18854 185752 18856
rect 155976 18794 185752 18854
rect 155976 18792 155984 18794
rect 185744 18792 185752 18794
rect 185816 18792 185832 18856
rect 185896 18792 185912 18856
rect 185976 18854 185984 18856
rect 185976 18794 200802 18854
rect 185976 18792 185984 18794
rect 19864 18714 19872 18716
rect -746 18654 19872 18714
rect 19864 18652 19872 18654
rect 19936 18652 19952 18716
rect 20016 18652 20032 18716
rect 20096 18714 20104 18716
rect 49864 18714 49872 18716
rect 20096 18654 49872 18714
rect 20096 18652 20104 18654
rect 49864 18652 49872 18654
rect 49936 18652 49952 18716
rect 50016 18652 50032 18716
rect 50096 18714 50104 18716
rect 79864 18714 79872 18716
rect 50096 18654 79872 18714
rect 50096 18652 50104 18654
rect 79864 18652 79872 18654
rect 79936 18652 79952 18716
rect 80016 18652 80032 18716
rect 80096 18714 80104 18716
rect 109864 18714 109872 18716
rect 80096 18654 109872 18714
rect 80096 18652 80104 18654
rect 109864 18652 109872 18654
rect 109936 18652 109952 18716
rect 110016 18652 110032 18716
rect 110096 18714 110104 18716
rect 139864 18714 139872 18716
rect 110096 18654 139872 18714
rect 110096 18652 110104 18654
rect 139864 18652 139872 18654
rect 139936 18652 139952 18716
rect 140016 18652 140032 18716
rect 140096 18714 140104 18716
rect 169864 18714 169872 18716
rect 140096 18654 169872 18714
rect 140096 18652 140104 18654
rect 169864 18652 169872 18654
rect 169936 18652 169952 18716
rect 170016 18652 170032 18716
rect 170096 18714 170104 18716
rect 170096 18654 200662 18714
rect 170096 18652 170104 18654
rect 4864 18574 4872 18576
rect -606 18514 4872 18574
rect 4864 18512 4872 18514
rect 4936 18512 4952 18576
rect 5016 18512 5032 18576
rect 5096 18574 5104 18576
rect 34864 18574 34872 18576
rect 5096 18514 34872 18574
rect 5096 18512 5104 18514
rect 34864 18512 34872 18514
rect 34936 18512 34952 18576
rect 35016 18512 35032 18576
rect 35096 18574 35104 18576
rect 64864 18574 64872 18576
rect 35096 18514 64872 18574
rect 35096 18512 35104 18514
rect 64864 18512 64872 18514
rect 64936 18512 64952 18576
rect 65016 18512 65032 18576
rect 65096 18574 65104 18576
rect 94864 18574 94872 18576
rect 65096 18514 94872 18574
rect 65096 18512 65104 18514
rect 94864 18512 94872 18514
rect 94936 18512 94952 18576
rect 95016 18512 95032 18576
rect 95096 18574 95104 18576
rect 124864 18574 124872 18576
rect 95096 18514 124872 18574
rect 95096 18512 95104 18514
rect 124864 18512 124872 18514
rect 124936 18512 124952 18576
rect 125016 18512 125032 18576
rect 125096 18574 125104 18576
rect 154864 18574 154872 18576
rect 125096 18514 154872 18574
rect 125096 18512 125104 18514
rect 154864 18512 154872 18514
rect 154936 18512 154952 18576
rect 155016 18512 155032 18576
rect 155096 18574 155104 18576
rect 184864 18574 184872 18576
rect 155096 18514 184872 18574
rect 155096 18512 155104 18514
rect 184864 18512 184872 18514
rect 184936 18512 184952 18576
rect 185016 18512 185032 18576
rect 185096 18574 185104 18576
rect 185096 18514 200522 18574
rect 185096 18512 185104 18514
rect 18984 18434 18992 18436
rect -466 18374 18992 18434
rect 18984 18372 18992 18374
rect 19056 18372 19072 18436
rect 19136 18372 19152 18436
rect 19216 18434 19224 18436
rect 48984 18434 48992 18436
rect 19216 18374 48992 18434
rect 19216 18372 19224 18374
rect 48984 18372 48992 18374
rect 49056 18372 49072 18436
rect 49136 18372 49152 18436
rect 49216 18434 49224 18436
rect 78984 18434 78992 18436
rect 49216 18374 78992 18434
rect 49216 18372 49224 18374
rect 78984 18372 78992 18374
rect 79056 18372 79072 18436
rect 79136 18372 79152 18436
rect 79216 18434 79224 18436
rect 108984 18434 108992 18436
rect 79216 18374 108992 18434
rect 79216 18372 79224 18374
rect 108984 18372 108992 18374
rect 109056 18372 109072 18436
rect 109136 18372 109152 18436
rect 109216 18434 109224 18436
rect 138984 18434 138992 18436
rect 109216 18374 138992 18434
rect 109216 18372 109224 18374
rect 138984 18372 138992 18374
rect 139056 18372 139072 18436
rect 139136 18372 139152 18436
rect 139216 18434 139224 18436
rect 168984 18434 168992 18436
rect 139216 18374 168992 18434
rect 139216 18372 139224 18374
rect 168984 18372 168992 18374
rect 169056 18372 169072 18436
rect 169136 18372 169152 18436
rect 169216 18434 169224 18436
rect 169216 18374 200382 18434
rect 169216 18372 169224 18374
rect 3984 18294 3992 18296
rect -326 18234 3992 18294
rect 3984 18232 3992 18234
rect 4056 18232 4072 18296
rect 4136 18232 4152 18296
rect 4216 18294 4224 18296
rect 33984 18294 33992 18296
rect 4216 18234 33992 18294
rect 4216 18232 4224 18234
rect 33984 18232 33992 18234
rect 34056 18232 34072 18296
rect 34136 18232 34152 18296
rect 34216 18294 34224 18296
rect 63984 18294 63992 18296
rect 34216 18234 63992 18294
rect 34216 18232 34224 18234
rect 63984 18232 63992 18234
rect 64056 18232 64072 18296
rect 64136 18232 64152 18296
rect 64216 18294 64224 18296
rect 93984 18294 93992 18296
rect 64216 18234 93992 18294
rect 64216 18232 64224 18234
rect 93984 18232 93992 18234
rect 94056 18232 94072 18296
rect 94136 18232 94152 18296
rect 94216 18294 94224 18296
rect 123984 18294 123992 18296
rect 94216 18234 123992 18294
rect 94216 18232 94224 18234
rect 123984 18232 123992 18234
rect 124056 18232 124072 18296
rect 124136 18232 124152 18296
rect 124216 18294 124224 18296
rect 153984 18294 153992 18296
rect 124216 18234 153992 18294
rect 124216 18232 124224 18234
rect 153984 18232 153992 18234
rect 154056 18232 154072 18296
rect 154136 18232 154152 18296
rect 154216 18294 154224 18296
rect 183984 18294 183992 18296
rect 154216 18234 183992 18294
rect 154216 18232 154224 18234
rect 183984 18232 183992 18234
rect 184056 18232 184072 18296
rect 184136 18232 184152 18296
rect 184216 18294 184224 18296
rect 184216 18234 200242 18294
rect 184216 18232 184224 18234
rect -400 14968 60 15088
rect -400 8984 60 9104
rect -400 3000 60 3120
rect 3984 -282 3992 -280
rect -326 -342 3992 -282
rect 3984 -344 3992 -342
rect 4056 -344 4072 -280
rect 4136 -344 4152 -280
rect 4216 -282 4224 -280
rect 33984 -282 33992 -280
rect 4216 -342 33992 -282
rect 4216 -344 4224 -342
rect 33984 -344 33992 -342
rect 34056 -344 34072 -280
rect 34136 -344 34152 -280
rect 34216 -282 34224 -280
rect 63984 -282 63992 -280
rect 34216 -342 63992 -282
rect 34216 -344 34224 -342
rect 63984 -344 63992 -342
rect 64056 -344 64072 -280
rect 64136 -344 64152 -280
rect 64216 -282 64224 -280
rect 93984 -282 93992 -280
rect 64216 -342 93992 -282
rect 64216 -344 64224 -342
rect 93984 -344 93992 -342
rect 94056 -344 94072 -280
rect 94136 -344 94152 -280
rect 94216 -282 94224 -280
rect 123984 -282 123992 -280
rect 94216 -342 123992 -282
rect 94216 -344 94224 -342
rect 123984 -344 123992 -342
rect 124056 -344 124072 -280
rect 124136 -344 124152 -280
rect 124216 -282 124224 -280
rect 153984 -282 153992 -280
rect 124216 -342 153992 -282
rect 124216 -344 124224 -342
rect 153984 -344 153992 -342
rect 154056 -344 154072 -280
rect 154136 -344 154152 -280
rect 154216 -282 154224 -280
rect 183984 -282 183992 -280
rect 154216 -342 183992 -282
rect 154216 -344 154224 -342
rect 183984 -344 183992 -342
rect 184056 -344 184072 -280
rect 184136 -344 184152 -280
rect 184216 -282 184224 -280
rect 184216 -342 200242 -282
rect 184216 -344 184224 -342
rect 18984 -422 18992 -420
rect -466 -482 18992 -422
rect 18984 -484 18992 -482
rect 19056 -484 19072 -420
rect 19136 -484 19152 -420
rect 19216 -422 19224 -420
rect 48984 -422 48992 -420
rect 19216 -482 48992 -422
rect 19216 -484 19224 -482
rect 48984 -484 48992 -482
rect 49056 -484 49072 -420
rect 49136 -484 49152 -420
rect 49216 -422 49224 -420
rect 78984 -422 78992 -420
rect 49216 -482 78992 -422
rect 49216 -484 49224 -482
rect 78984 -484 78992 -482
rect 79056 -484 79072 -420
rect 79136 -484 79152 -420
rect 79216 -422 79224 -420
rect 108984 -422 108992 -420
rect 79216 -482 108992 -422
rect 79216 -484 79224 -482
rect 108984 -484 108992 -482
rect 109056 -484 109072 -420
rect 109136 -484 109152 -420
rect 109216 -422 109224 -420
rect 138984 -422 138992 -420
rect 109216 -482 138992 -422
rect 109216 -484 109224 -482
rect 138984 -484 138992 -482
rect 139056 -484 139072 -420
rect 139136 -484 139152 -420
rect 139216 -422 139224 -420
rect 168984 -422 168992 -420
rect 139216 -482 168992 -422
rect 139216 -484 139224 -482
rect 168984 -484 168992 -482
rect 169056 -484 169072 -420
rect 169136 -484 169152 -420
rect 169216 -422 169224 -420
rect 169216 -482 200382 -422
rect 169216 -484 169224 -482
rect 4864 -562 4872 -560
rect -606 -622 4872 -562
rect 4864 -624 4872 -622
rect 4936 -624 4952 -560
rect 5016 -624 5032 -560
rect 5096 -562 5104 -560
rect 34864 -562 34872 -560
rect 5096 -622 34872 -562
rect 5096 -624 5104 -622
rect 34864 -624 34872 -622
rect 34936 -624 34952 -560
rect 35016 -624 35032 -560
rect 35096 -562 35104 -560
rect 64864 -562 64872 -560
rect 35096 -622 64872 -562
rect 35096 -624 35104 -622
rect 64864 -624 64872 -622
rect 64936 -624 64952 -560
rect 65016 -624 65032 -560
rect 65096 -562 65104 -560
rect 94864 -562 94872 -560
rect 65096 -622 94872 -562
rect 65096 -624 65104 -622
rect 94864 -624 94872 -622
rect 94936 -624 94952 -560
rect 95016 -624 95032 -560
rect 95096 -562 95104 -560
rect 124864 -562 124872 -560
rect 95096 -622 124872 -562
rect 95096 -624 95104 -622
rect 124864 -624 124872 -622
rect 124936 -624 124952 -560
rect 125016 -624 125032 -560
rect 125096 -562 125104 -560
rect 154864 -562 154872 -560
rect 125096 -622 154872 -562
rect 125096 -624 125104 -622
rect 154864 -624 154872 -622
rect 154936 -624 154952 -560
rect 155016 -624 155032 -560
rect 155096 -562 155104 -560
rect 184864 -562 184872 -560
rect 155096 -622 184872 -562
rect 155096 -624 155104 -622
rect 184864 -624 184872 -622
rect 184936 -624 184952 -560
rect 185016 -624 185032 -560
rect 185096 -562 185104 -560
rect 185096 -622 200522 -562
rect 185096 -624 185104 -622
rect 19864 -702 19872 -700
rect -746 -762 19872 -702
rect 19864 -764 19872 -762
rect 19936 -764 19952 -700
rect 20016 -764 20032 -700
rect 20096 -702 20104 -700
rect 49864 -702 49872 -700
rect 20096 -762 49872 -702
rect 20096 -764 20104 -762
rect 49864 -764 49872 -762
rect 49936 -764 49952 -700
rect 50016 -764 50032 -700
rect 50096 -702 50104 -700
rect 79864 -702 79872 -700
rect 50096 -762 79872 -702
rect 50096 -764 50104 -762
rect 79864 -764 79872 -762
rect 79936 -764 79952 -700
rect 80016 -764 80032 -700
rect 80096 -702 80104 -700
rect 109864 -702 109872 -700
rect 80096 -762 109872 -702
rect 80096 -764 80104 -762
rect 109864 -764 109872 -762
rect 109936 -764 109952 -700
rect 110016 -764 110032 -700
rect 110096 -702 110104 -700
rect 139864 -702 139872 -700
rect 110096 -762 139872 -702
rect 110096 -764 110104 -762
rect 139864 -764 139872 -762
rect 139936 -764 139952 -700
rect 140016 -764 140032 -700
rect 140096 -702 140104 -700
rect 169864 -702 169872 -700
rect 140096 -762 169872 -702
rect 140096 -764 140104 -762
rect 169864 -764 169872 -762
rect 169936 -764 169952 -700
rect 170016 -764 170032 -700
rect 170096 -702 170104 -700
rect 170096 -762 200662 -702
rect 170096 -764 170104 -762
rect 5744 -842 5752 -840
rect -886 -902 5752 -842
rect 5744 -904 5752 -902
rect 5816 -904 5832 -840
rect 5896 -904 5912 -840
rect 5976 -842 5984 -840
rect 35744 -842 35752 -840
rect 5976 -902 35752 -842
rect 5976 -904 5984 -902
rect 35744 -904 35752 -902
rect 35816 -904 35832 -840
rect 35896 -904 35912 -840
rect 35976 -842 35984 -840
rect 65744 -842 65752 -840
rect 35976 -902 65752 -842
rect 35976 -904 35984 -902
rect 65744 -904 65752 -902
rect 65816 -904 65832 -840
rect 65896 -904 65912 -840
rect 65976 -842 65984 -840
rect 95744 -842 95752 -840
rect 65976 -902 95752 -842
rect 65976 -904 65984 -902
rect 95744 -904 95752 -902
rect 95816 -904 95832 -840
rect 95896 -904 95912 -840
rect 95976 -842 95984 -840
rect 125744 -842 125752 -840
rect 95976 -902 125752 -842
rect 95976 -904 95984 -902
rect 125744 -904 125752 -902
rect 125816 -904 125832 -840
rect 125896 -904 125912 -840
rect 125976 -842 125984 -840
rect 155744 -842 155752 -840
rect 125976 -902 155752 -842
rect 125976 -904 125984 -902
rect 155744 -904 155752 -902
rect 155816 -904 155832 -840
rect 155896 -904 155912 -840
rect 155976 -842 155984 -840
rect 185744 -842 185752 -840
rect 155976 -902 185752 -842
rect 155976 -904 155984 -902
rect 185744 -904 185752 -902
rect 185816 -904 185832 -840
rect 185896 -904 185912 -840
rect 185976 -842 185984 -840
rect 185976 -902 200802 -842
rect 185976 -904 185984 -902
rect 20744 -982 20752 -980
rect -1026 -1042 20752 -982
rect 20744 -1044 20752 -1042
rect 20816 -1044 20832 -980
rect 20896 -1044 20912 -980
rect 20976 -982 20984 -980
rect 50744 -982 50752 -980
rect 20976 -1042 50752 -982
rect 20976 -1044 20984 -1042
rect 50744 -1044 50752 -1042
rect 50816 -1044 50832 -980
rect 50896 -1044 50912 -980
rect 50976 -982 50984 -980
rect 80744 -982 80752 -980
rect 50976 -1042 80752 -982
rect 50976 -1044 50984 -1042
rect 80744 -1044 80752 -1042
rect 80816 -1044 80832 -980
rect 80896 -1044 80912 -980
rect 80976 -982 80984 -980
rect 110744 -982 110752 -980
rect 80976 -1042 110752 -982
rect 80976 -1044 80984 -1042
rect 110744 -1044 110752 -1042
rect 110816 -1044 110832 -980
rect 110896 -1044 110912 -980
rect 110976 -982 110984 -980
rect 140744 -982 140752 -980
rect 110976 -1042 140752 -982
rect 110976 -1044 110984 -1042
rect 140744 -1044 140752 -1042
rect 140816 -1044 140832 -980
rect 140896 -1044 140912 -980
rect 140976 -982 140984 -980
rect 170744 -982 170752 -980
rect 140976 -1042 170752 -982
rect 140976 -1044 140984 -1042
rect 170744 -1044 170752 -1042
rect 170816 -1044 170832 -980
rect 170896 -1044 170912 -980
rect 170976 -982 170984 -980
rect 170976 -1042 200942 -982
rect 170976 -1044 170984 -1042
rect 6624 -1122 6632 -1120
rect -1166 -1182 6632 -1122
rect 6624 -1184 6632 -1182
rect 6696 -1184 6712 -1120
rect 6776 -1184 6792 -1120
rect 6856 -1122 6864 -1120
rect 36624 -1122 36632 -1120
rect 6856 -1182 36632 -1122
rect 6856 -1184 6864 -1182
rect 36624 -1184 36632 -1182
rect 36696 -1184 36712 -1120
rect 36776 -1184 36792 -1120
rect 36856 -1122 36864 -1120
rect 66624 -1122 66632 -1120
rect 36856 -1182 66632 -1122
rect 36856 -1184 36864 -1182
rect 66624 -1184 66632 -1182
rect 66696 -1184 66712 -1120
rect 66776 -1184 66792 -1120
rect 66856 -1122 66864 -1120
rect 96624 -1122 96632 -1120
rect 66856 -1182 96632 -1122
rect 66856 -1184 66864 -1182
rect 96624 -1184 96632 -1182
rect 96696 -1184 96712 -1120
rect 96776 -1184 96792 -1120
rect 96856 -1122 96864 -1120
rect 126624 -1122 126632 -1120
rect 96856 -1182 126632 -1122
rect 96856 -1184 96864 -1182
rect 126624 -1184 126632 -1182
rect 126696 -1184 126712 -1120
rect 126776 -1184 126792 -1120
rect 126856 -1122 126864 -1120
rect 156624 -1122 156632 -1120
rect 126856 -1182 156632 -1122
rect 126856 -1184 126864 -1182
rect 156624 -1184 156632 -1182
rect 156696 -1184 156712 -1120
rect 156776 -1184 156792 -1120
rect 156856 -1122 156864 -1120
rect 186624 -1122 186632 -1120
rect 156856 -1182 186632 -1122
rect 156856 -1184 156864 -1182
rect 186624 -1184 186632 -1182
rect 186696 -1184 186712 -1120
rect 186776 -1184 186792 -1120
rect 186856 -1122 186864 -1120
rect 186856 -1182 201082 -1122
rect 186856 -1184 186864 -1182
rect 21624 -1262 21632 -1260
rect -1306 -1322 21632 -1262
rect 21624 -1324 21632 -1322
rect 21696 -1324 21712 -1260
rect 21776 -1324 21792 -1260
rect 21856 -1262 21864 -1260
rect 51624 -1262 51632 -1260
rect 21856 -1322 51632 -1262
rect 21856 -1324 21864 -1322
rect 51624 -1324 51632 -1322
rect 51696 -1324 51712 -1260
rect 51776 -1324 51792 -1260
rect 51856 -1262 51864 -1260
rect 81624 -1262 81632 -1260
rect 51856 -1322 81632 -1262
rect 51856 -1324 51864 -1322
rect 81624 -1324 81632 -1322
rect 81696 -1324 81712 -1260
rect 81776 -1324 81792 -1260
rect 81856 -1262 81864 -1260
rect 111624 -1262 111632 -1260
rect 81856 -1322 111632 -1262
rect 81856 -1324 81864 -1322
rect 111624 -1324 111632 -1322
rect 111696 -1324 111712 -1260
rect 111776 -1324 111792 -1260
rect 111856 -1262 111864 -1260
rect 141624 -1262 141632 -1260
rect 111856 -1322 141632 -1262
rect 111856 -1324 111864 -1322
rect 141624 -1324 141632 -1322
rect 141696 -1324 141712 -1260
rect 141776 -1324 141792 -1260
rect 141856 -1262 141864 -1260
rect 171624 -1262 171632 -1260
rect 141856 -1322 171632 -1262
rect 141856 -1324 141864 -1322
rect 171624 -1324 171632 -1322
rect 171696 -1324 171712 -1260
rect 171776 -1324 171792 -1260
rect 171856 -1262 171864 -1260
rect 171856 -1322 201222 -1262
rect 171856 -1324 171864 -1322
rect 7504 -1402 7512 -1400
rect -1446 -1462 7512 -1402
rect 7504 -1464 7512 -1462
rect 7576 -1464 7592 -1400
rect 7656 -1464 7672 -1400
rect 7736 -1402 7744 -1400
rect 37504 -1402 37512 -1400
rect 7736 -1462 37512 -1402
rect 7736 -1464 7744 -1462
rect 37504 -1464 37512 -1462
rect 37576 -1464 37592 -1400
rect 37656 -1464 37672 -1400
rect 37736 -1402 37744 -1400
rect 67504 -1402 67512 -1400
rect 37736 -1462 67512 -1402
rect 37736 -1464 37744 -1462
rect 67504 -1464 67512 -1462
rect 67576 -1464 67592 -1400
rect 67656 -1464 67672 -1400
rect 67736 -1402 67744 -1400
rect 97504 -1402 97512 -1400
rect 67736 -1462 97512 -1402
rect 67736 -1464 67744 -1462
rect 97504 -1464 97512 -1462
rect 97576 -1464 97592 -1400
rect 97656 -1464 97672 -1400
rect 97736 -1402 97744 -1400
rect 127504 -1402 127512 -1400
rect 97736 -1462 127512 -1402
rect 97736 -1464 97744 -1462
rect 127504 -1464 127512 -1462
rect 127576 -1464 127592 -1400
rect 127656 -1464 127672 -1400
rect 127736 -1402 127744 -1400
rect 157504 -1402 157512 -1400
rect 127736 -1462 157512 -1402
rect 127736 -1464 127744 -1462
rect 157504 -1464 157512 -1462
rect 157576 -1464 157592 -1400
rect 157656 -1464 157672 -1400
rect 157736 -1402 157744 -1400
rect 187504 -1402 187512 -1400
rect 157736 -1462 187512 -1402
rect 157736 -1464 157744 -1462
rect 187504 -1464 187512 -1462
rect 187576 -1464 187592 -1400
rect 187656 -1464 187672 -1400
rect 187736 -1402 187744 -1400
rect 187736 -1462 201362 -1402
rect 187736 -1464 187744 -1462
rect 22504 -1542 22512 -1540
rect -1586 -1602 22512 -1542
rect 22504 -1604 22512 -1602
rect 22576 -1604 22592 -1540
rect 22656 -1604 22672 -1540
rect 22736 -1542 22744 -1540
rect 52504 -1542 52512 -1540
rect 22736 -1602 52512 -1542
rect 22736 -1604 22744 -1602
rect 52504 -1604 52512 -1602
rect 52576 -1604 52592 -1540
rect 52656 -1604 52672 -1540
rect 52736 -1542 52744 -1540
rect 82504 -1542 82512 -1540
rect 52736 -1602 82512 -1542
rect 52736 -1604 52744 -1602
rect 82504 -1604 82512 -1602
rect 82576 -1604 82592 -1540
rect 82656 -1604 82672 -1540
rect 82736 -1542 82744 -1540
rect 112504 -1542 112512 -1540
rect 82736 -1602 112512 -1542
rect 82736 -1604 82744 -1602
rect 112504 -1604 112512 -1602
rect 112576 -1604 112592 -1540
rect 112656 -1604 112672 -1540
rect 112736 -1542 112744 -1540
rect 142504 -1542 142512 -1540
rect 112736 -1602 142512 -1542
rect 112736 -1604 112744 -1602
rect 142504 -1604 142512 -1602
rect 142576 -1604 142592 -1540
rect 142656 -1604 142672 -1540
rect 142736 -1542 142744 -1540
rect 172504 -1542 172512 -1540
rect 142736 -1602 172512 -1542
rect 142736 -1604 142744 -1602
rect 172504 -1604 172512 -1602
rect 172576 -1604 172592 -1540
rect 172656 -1604 172672 -1540
rect 172736 -1542 172744 -1540
rect 172736 -1602 201502 -1542
rect 172736 -1604 172744 -1602
<< obsm3 >>
rect 60 851 194659 17917
<< via3 >>
rect 22512 19492 22576 19556
rect 22592 19492 22656 19556
rect 22672 19492 22736 19556
rect 52512 19492 52576 19556
rect 52592 19492 52656 19556
rect 52672 19492 52736 19556
rect 82512 19492 82576 19556
rect 82592 19492 82656 19556
rect 82672 19492 82736 19556
rect 112512 19492 112576 19556
rect 112592 19492 112656 19556
rect 112672 19492 112736 19556
rect 142512 19492 142576 19556
rect 142592 19492 142656 19556
rect 142672 19492 142736 19556
rect 172512 19492 172576 19556
rect 172592 19492 172656 19556
rect 172672 19492 172736 19556
rect 7512 19352 7576 19416
rect 7592 19352 7656 19416
rect 7672 19352 7736 19416
rect 37512 19352 37576 19416
rect 37592 19352 37656 19416
rect 37672 19352 37736 19416
rect 67512 19352 67576 19416
rect 67592 19352 67656 19416
rect 67672 19352 67736 19416
rect 97512 19352 97576 19416
rect 97592 19352 97656 19416
rect 97672 19352 97736 19416
rect 127512 19352 127576 19416
rect 127592 19352 127656 19416
rect 127672 19352 127736 19416
rect 157512 19352 157576 19416
rect 157592 19352 157656 19416
rect 157672 19352 157736 19416
rect 187512 19352 187576 19416
rect 187592 19352 187656 19416
rect 187672 19352 187736 19416
rect 21632 19212 21696 19276
rect 21712 19212 21776 19276
rect 21792 19212 21856 19276
rect 51632 19212 51696 19276
rect 51712 19212 51776 19276
rect 51792 19212 51856 19276
rect 81632 19212 81696 19276
rect 81712 19212 81776 19276
rect 81792 19212 81856 19276
rect 111632 19212 111696 19276
rect 111712 19212 111776 19276
rect 111792 19212 111856 19276
rect 141632 19212 141696 19276
rect 141712 19212 141776 19276
rect 141792 19212 141856 19276
rect 171632 19212 171696 19276
rect 171712 19212 171776 19276
rect 171792 19212 171856 19276
rect 6632 19072 6696 19136
rect 6712 19072 6776 19136
rect 6792 19072 6856 19136
rect 36632 19072 36696 19136
rect 36712 19072 36776 19136
rect 36792 19072 36856 19136
rect 66632 19072 66696 19136
rect 66712 19072 66776 19136
rect 66792 19072 66856 19136
rect 96632 19072 96696 19136
rect 96712 19072 96776 19136
rect 96792 19072 96856 19136
rect 126632 19072 126696 19136
rect 126712 19072 126776 19136
rect 126792 19072 126856 19136
rect 156632 19072 156696 19136
rect 156712 19072 156776 19136
rect 156792 19072 156856 19136
rect 186632 19072 186696 19136
rect 186712 19072 186776 19136
rect 186792 19072 186856 19136
rect 20752 18932 20816 18996
rect 20832 18932 20896 18996
rect 20912 18932 20976 18996
rect 50752 18932 50816 18996
rect 50832 18932 50896 18996
rect 50912 18932 50976 18996
rect 80752 18932 80816 18996
rect 80832 18932 80896 18996
rect 80912 18932 80976 18996
rect 110752 18932 110816 18996
rect 110832 18932 110896 18996
rect 110912 18932 110976 18996
rect 140752 18932 140816 18996
rect 140832 18932 140896 18996
rect 140912 18932 140976 18996
rect 170752 18932 170816 18996
rect 170832 18932 170896 18996
rect 170912 18932 170976 18996
rect 5752 18792 5816 18856
rect 5832 18792 5896 18856
rect 5912 18792 5976 18856
rect 35752 18792 35816 18856
rect 35832 18792 35896 18856
rect 35912 18792 35976 18856
rect 65752 18792 65816 18856
rect 65832 18792 65896 18856
rect 65912 18792 65976 18856
rect 95752 18792 95816 18856
rect 95832 18792 95896 18856
rect 95912 18792 95976 18856
rect 125752 18792 125816 18856
rect 125832 18792 125896 18856
rect 125912 18792 125976 18856
rect 155752 18792 155816 18856
rect 155832 18792 155896 18856
rect 155912 18792 155976 18856
rect 185752 18792 185816 18856
rect 185832 18792 185896 18856
rect 185912 18792 185976 18856
rect 19872 18652 19936 18716
rect 19952 18652 20016 18716
rect 20032 18652 20096 18716
rect 49872 18652 49936 18716
rect 49952 18652 50016 18716
rect 50032 18652 50096 18716
rect 79872 18652 79936 18716
rect 79952 18652 80016 18716
rect 80032 18652 80096 18716
rect 109872 18652 109936 18716
rect 109952 18652 110016 18716
rect 110032 18652 110096 18716
rect 139872 18652 139936 18716
rect 139952 18652 140016 18716
rect 140032 18652 140096 18716
rect 169872 18652 169936 18716
rect 169952 18652 170016 18716
rect 170032 18652 170096 18716
rect 4872 18512 4936 18576
rect 4952 18512 5016 18576
rect 5032 18512 5096 18576
rect 34872 18512 34936 18576
rect 34952 18512 35016 18576
rect 35032 18512 35096 18576
rect 64872 18512 64936 18576
rect 64952 18512 65016 18576
rect 65032 18512 65096 18576
rect 94872 18512 94936 18576
rect 94952 18512 95016 18576
rect 95032 18512 95096 18576
rect 124872 18512 124936 18576
rect 124952 18512 125016 18576
rect 125032 18512 125096 18576
rect 154872 18512 154936 18576
rect 154952 18512 155016 18576
rect 155032 18512 155096 18576
rect 184872 18512 184936 18576
rect 184952 18512 185016 18576
rect 185032 18512 185096 18576
rect 18992 18372 19056 18436
rect 19072 18372 19136 18436
rect 19152 18372 19216 18436
rect 48992 18372 49056 18436
rect 49072 18372 49136 18436
rect 49152 18372 49216 18436
rect 78992 18372 79056 18436
rect 79072 18372 79136 18436
rect 79152 18372 79216 18436
rect 108992 18372 109056 18436
rect 109072 18372 109136 18436
rect 109152 18372 109216 18436
rect 138992 18372 139056 18436
rect 139072 18372 139136 18436
rect 139152 18372 139216 18436
rect 168992 18372 169056 18436
rect 169072 18372 169136 18436
rect 169152 18372 169216 18436
rect 3992 18232 4056 18296
rect 4072 18232 4136 18296
rect 4152 18232 4216 18296
rect 33992 18232 34056 18296
rect 34072 18232 34136 18296
rect 34152 18232 34216 18296
rect 63992 18232 64056 18296
rect 64072 18232 64136 18296
rect 64152 18232 64216 18296
rect 93992 18232 94056 18296
rect 94072 18232 94136 18296
rect 94152 18232 94216 18296
rect 123992 18232 124056 18296
rect 124072 18232 124136 18296
rect 124152 18232 124216 18296
rect 153992 18232 154056 18296
rect 154072 18232 154136 18296
rect 154152 18232 154216 18296
rect 183992 18232 184056 18296
rect 184072 18232 184136 18296
rect 184152 18232 184216 18296
rect 3992 -344 4056 -280
rect 4072 -344 4136 -280
rect 4152 -344 4216 -280
rect 33992 -344 34056 -280
rect 34072 -344 34136 -280
rect 34152 -344 34216 -280
rect 63992 -344 64056 -280
rect 64072 -344 64136 -280
rect 64152 -344 64216 -280
rect 93992 -344 94056 -280
rect 94072 -344 94136 -280
rect 94152 -344 94216 -280
rect 123992 -344 124056 -280
rect 124072 -344 124136 -280
rect 124152 -344 124216 -280
rect 153992 -344 154056 -280
rect 154072 -344 154136 -280
rect 154152 -344 154216 -280
rect 183992 -344 184056 -280
rect 184072 -344 184136 -280
rect 184152 -344 184216 -280
rect 18992 -484 19056 -420
rect 19072 -484 19136 -420
rect 19152 -484 19216 -420
rect 48992 -484 49056 -420
rect 49072 -484 49136 -420
rect 49152 -484 49216 -420
rect 78992 -484 79056 -420
rect 79072 -484 79136 -420
rect 79152 -484 79216 -420
rect 108992 -484 109056 -420
rect 109072 -484 109136 -420
rect 109152 -484 109216 -420
rect 138992 -484 139056 -420
rect 139072 -484 139136 -420
rect 139152 -484 139216 -420
rect 168992 -484 169056 -420
rect 169072 -484 169136 -420
rect 169152 -484 169216 -420
rect 4872 -624 4936 -560
rect 4952 -624 5016 -560
rect 5032 -624 5096 -560
rect 34872 -624 34936 -560
rect 34952 -624 35016 -560
rect 35032 -624 35096 -560
rect 64872 -624 64936 -560
rect 64952 -624 65016 -560
rect 65032 -624 65096 -560
rect 94872 -624 94936 -560
rect 94952 -624 95016 -560
rect 95032 -624 95096 -560
rect 124872 -624 124936 -560
rect 124952 -624 125016 -560
rect 125032 -624 125096 -560
rect 154872 -624 154936 -560
rect 154952 -624 155016 -560
rect 155032 -624 155096 -560
rect 184872 -624 184936 -560
rect 184952 -624 185016 -560
rect 185032 -624 185096 -560
rect 19872 -764 19936 -700
rect 19952 -764 20016 -700
rect 20032 -764 20096 -700
rect 49872 -764 49936 -700
rect 49952 -764 50016 -700
rect 50032 -764 50096 -700
rect 79872 -764 79936 -700
rect 79952 -764 80016 -700
rect 80032 -764 80096 -700
rect 109872 -764 109936 -700
rect 109952 -764 110016 -700
rect 110032 -764 110096 -700
rect 139872 -764 139936 -700
rect 139952 -764 140016 -700
rect 140032 -764 140096 -700
rect 169872 -764 169936 -700
rect 169952 -764 170016 -700
rect 170032 -764 170096 -700
rect 5752 -904 5816 -840
rect 5832 -904 5896 -840
rect 5912 -904 5976 -840
rect 35752 -904 35816 -840
rect 35832 -904 35896 -840
rect 35912 -904 35976 -840
rect 65752 -904 65816 -840
rect 65832 -904 65896 -840
rect 65912 -904 65976 -840
rect 95752 -904 95816 -840
rect 95832 -904 95896 -840
rect 95912 -904 95976 -840
rect 125752 -904 125816 -840
rect 125832 -904 125896 -840
rect 125912 -904 125976 -840
rect 155752 -904 155816 -840
rect 155832 -904 155896 -840
rect 155912 -904 155976 -840
rect 185752 -904 185816 -840
rect 185832 -904 185896 -840
rect 185912 -904 185976 -840
rect 20752 -1044 20816 -980
rect 20832 -1044 20896 -980
rect 20912 -1044 20976 -980
rect 50752 -1044 50816 -980
rect 50832 -1044 50896 -980
rect 50912 -1044 50976 -980
rect 80752 -1044 80816 -980
rect 80832 -1044 80896 -980
rect 80912 -1044 80976 -980
rect 110752 -1044 110816 -980
rect 110832 -1044 110896 -980
rect 110912 -1044 110976 -980
rect 140752 -1044 140816 -980
rect 140832 -1044 140896 -980
rect 140912 -1044 140976 -980
rect 170752 -1044 170816 -980
rect 170832 -1044 170896 -980
rect 170912 -1044 170976 -980
rect 6632 -1184 6696 -1120
rect 6712 -1184 6776 -1120
rect 6792 -1184 6856 -1120
rect 36632 -1184 36696 -1120
rect 36712 -1184 36776 -1120
rect 36792 -1184 36856 -1120
rect 66632 -1184 66696 -1120
rect 66712 -1184 66776 -1120
rect 66792 -1184 66856 -1120
rect 96632 -1184 96696 -1120
rect 96712 -1184 96776 -1120
rect 96792 -1184 96856 -1120
rect 126632 -1184 126696 -1120
rect 126712 -1184 126776 -1120
rect 126792 -1184 126856 -1120
rect 156632 -1184 156696 -1120
rect 156712 -1184 156776 -1120
rect 156792 -1184 156856 -1120
rect 186632 -1184 186696 -1120
rect 186712 -1184 186776 -1120
rect 186792 -1184 186856 -1120
rect 21632 -1324 21696 -1260
rect 21712 -1324 21776 -1260
rect 21792 -1324 21856 -1260
rect 51632 -1324 51696 -1260
rect 51712 -1324 51776 -1260
rect 51792 -1324 51856 -1260
rect 81632 -1324 81696 -1260
rect 81712 -1324 81776 -1260
rect 81792 -1324 81856 -1260
rect 111632 -1324 111696 -1260
rect 111712 -1324 111776 -1260
rect 111792 -1324 111856 -1260
rect 141632 -1324 141696 -1260
rect 141712 -1324 141776 -1260
rect 141792 -1324 141856 -1260
rect 171632 -1324 171696 -1260
rect 171712 -1324 171776 -1260
rect 171792 -1324 171856 -1260
rect 7512 -1464 7576 -1400
rect 7592 -1464 7656 -1400
rect 7672 -1464 7736 -1400
rect 37512 -1464 37576 -1400
rect 37592 -1464 37656 -1400
rect 37672 -1464 37736 -1400
rect 67512 -1464 67576 -1400
rect 67592 -1464 67656 -1400
rect 67672 -1464 67736 -1400
rect 97512 -1464 97576 -1400
rect 97592 -1464 97656 -1400
rect 97672 -1464 97736 -1400
rect 127512 -1464 127576 -1400
rect 127592 -1464 127656 -1400
rect 127672 -1464 127736 -1400
rect 157512 -1464 157576 -1400
rect 157592 -1464 157656 -1400
rect 157672 -1464 157736 -1400
rect 187512 -1464 187576 -1400
rect 187592 -1464 187656 -1400
rect 187672 -1464 187736 -1400
rect 22512 -1604 22576 -1540
rect 22592 -1604 22656 -1540
rect 22672 -1604 22736 -1540
rect 52512 -1604 52576 -1540
rect 52592 -1604 52656 -1540
rect 52672 -1604 52736 -1540
rect 82512 -1604 82576 -1540
rect 82592 -1604 82656 -1540
rect 82672 -1604 82736 -1540
rect 112512 -1604 112576 -1540
rect 112592 -1604 112656 -1540
rect 112672 -1604 112736 -1540
rect 142512 -1604 142576 -1540
rect 142592 -1604 142656 -1540
rect 142672 -1604 142736 -1540
rect 172512 -1604 172576 -1540
rect 172592 -1604 172656 -1540
rect 172672 -1604 172736 -1540
<< metal4 >>
rect 22504 19556 22744 19557
rect -1586 -1602 -1526 19554
rect 7504 19416 7744 19554
rect -1446 -1462 -1386 19414
rect 7504 19352 7512 19416
rect 7576 19352 7592 19416
rect 7656 19352 7672 19416
rect 7736 19352 7744 19416
rect -1306 -1322 -1246 19274
rect 6624 19136 6864 19274
rect -1166 -1182 -1106 19134
rect 6624 19072 6632 19136
rect 6696 19072 6712 19136
rect 6776 19072 6792 19136
rect 6856 19072 6864 19136
rect -1026 -1042 -966 18994
rect 5744 18856 5984 18994
rect -886 -902 -826 18854
rect 5744 18792 5752 18856
rect 5816 18792 5832 18856
rect 5896 18792 5912 18856
rect 5976 18792 5984 18856
rect -746 -762 -686 18714
rect 4864 18576 5104 18714
rect -606 -622 -546 18574
rect 4864 18512 4872 18576
rect 4936 18512 4952 18576
rect 5016 18512 5032 18576
rect 5096 18512 5104 18576
rect -466 -482 -406 18434
rect 3984 18296 4224 18434
rect -326 -342 -266 18294
rect 3984 18232 3992 18296
rect 4056 18232 4072 18296
rect 4136 18232 4152 18296
rect 4216 18232 4224 18296
rect 3984 17940 4224 18232
rect 4864 17940 5104 18512
rect 5744 17940 5984 18792
rect 6624 17940 6864 19072
rect 7504 17940 7744 19352
rect 22504 19492 22512 19556
rect 22576 19492 22592 19556
rect 22656 19492 22672 19556
rect 22736 19492 22744 19556
rect 52504 19556 52744 19557
rect 21624 19276 21864 19277
rect 21624 19212 21632 19276
rect 21696 19212 21712 19276
rect 21776 19212 21792 19276
rect 21856 19212 21864 19276
rect 20744 18996 20984 18997
rect 20744 18932 20752 18996
rect 20816 18932 20832 18996
rect 20896 18932 20912 18996
rect 20976 18932 20984 18996
rect 19864 18716 20104 18717
rect 19864 18652 19872 18716
rect 19936 18652 19952 18716
rect 20016 18652 20032 18716
rect 20096 18652 20104 18716
rect 18984 18436 19224 18437
rect 18984 18372 18992 18436
rect 19056 18372 19072 18436
rect 19136 18372 19152 18436
rect 19216 18372 19224 18436
rect 18984 17940 19224 18372
rect 19864 17940 20104 18652
rect 20744 17940 20984 18932
rect 21624 17940 21864 19212
rect 22504 17940 22744 19492
rect 37504 19416 37744 19554
rect 37504 19352 37512 19416
rect 37576 19352 37592 19416
rect 37656 19352 37672 19416
rect 37736 19352 37744 19416
rect 36624 19136 36864 19274
rect 36624 19072 36632 19136
rect 36696 19072 36712 19136
rect 36776 19072 36792 19136
rect 36856 19072 36864 19136
rect 35744 18856 35984 18994
rect 35744 18792 35752 18856
rect 35816 18792 35832 18856
rect 35896 18792 35912 18856
rect 35976 18792 35984 18856
rect 34864 18576 35104 18714
rect 34864 18512 34872 18576
rect 34936 18512 34952 18576
rect 35016 18512 35032 18576
rect 35096 18512 35104 18576
rect 33984 18296 34224 18434
rect 33984 18232 33992 18296
rect 34056 18232 34072 18296
rect 34136 18232 34152 18296
rect 34216 18232 34224 18296
rect 33984 17940 34224 18232
rect 34864 17940 35104 18512
rect 35744 17940 35984 18792
rect 36624 17940 36864 19072
rect 37504 17940 37744 19352
rect 52504 19492 52512 19556
rect 52576 19492 52592 19556
rect 52656 19492 52672 19556
rect 52736 19492 52744 19556
rect 82504 19556 82744 19557
rect 51624 19276 51864 19277
rect 51624 19212 51632 19276
rect 51696 19212 51712 19276
rect 51776 19212 51792 19276
rect 51856 19212 51864 19276
rect 50744 18996 50984 18997
rect 50744 18932 50752 18996
rect 50816 18932 50832 18996
rect 50896 18932 50912 18996
rect 50976 18932 50984 18996
rect 49864 18716 50104 18717
rect 49864 18652 49872 18716
rect 49936 18652 49952 18716
rect 50016 18652 50032 18716
rect 50096 18652 50104 18716
rect 48984 18436 49224 18437
rect 48984 18372 48992 18436
rect 49056 18372 49072 18436
rect 49136 18372 49152 18436
rect 49216 18372 49224 18436
rect 48984 17940 49224 18372
rect 49864 17940 50104 18652
rect 50744 17940 50984 18932
rect 51624 17940 51864 19212
rect 52504 17940 52744 19492
rect 67504 19416 67744 19554
rect 67504 19352 67512 19416
rect 67576 19352 67592 19416
rect 67656 19352 67672 19416
rect 67736 19352 67744 19416
rect 66624 19136 66864 19274
rect 66624 19072 66632 19136
rect 66696 19072 66712 19136
rect 66776 19072 66792 19136
rect 66856 19072 66864 19136
rect 65744 18856 65984 18994
rect 65744 18792 65752 18856
rect 65816 18792 65832 18856
rect 65896 18792 65912 18856
rect 65976 18792 65984 18856
rect 64864 18576 65104 18714
rect 64864 18512 64872 18576
rect 64936 18512 64952 18576
rect 65016 18512 65032 18576
rect 65096 18512 65104 18576
rect 63984 18296 64224 18434
rect 63984 18232 63992 18296
rect 64056 18232 64072 18296
rect 64136 18232 64152 18296
rect 64216 18232 64224 18296
rect 63984 17940 64224 18232
rect 64864 17940 65104 18512
rect 65744 17940 65984 18792
rect 66624 17940 66864 19072
rect 67504 17940 67744 19352
rect 82504 19492 82512 19556
rect 82576 19492 82592 19556
rect 82656 19492 82672 19556
rect 82736 19492 82744 19556
rect 112504 19556 112744 19557
rect 81624 19276 81864 19277
rect 81624 19212 81632 19276
rect 81696 19212 81712 19276
rect 81776 19212 81792 19276
rect 81856 19212 81864 19276
rect 80744 18996 80984 18997
rect 80744 18932 80752 18996
rect 80816 18932 80832 18996
rect 80896 18932 80912 18996
rect 80976 18932 80984 18996
rect 79864 18716 80104 18717
rect 79864 18652 79872 18716
rect 79936 18652 79952 18716
rect 80016 18652 80032 18716
rect 80096 18652 80104 18716
rect 78984 18436 79224 18437
rect 78984 18372 78992 18436
rect 79056 18372 79072 18436
rect 79136 18372 79152 18436
rect 79216 18372 79224 18436
rect 78984 17940 79224 18372
rect 79864 17940 80104 18652
rect 80744 17940 80984 18932
rect 81624 17940 81864 19212
rect 82504 17940 82744 19492
rect 97504 19416 97744 19554
rect 97504 19352 97512 19416
rect 97576 19352 97592 19416
rect 97656 19352 97672 19416
rect 97736 19352 97744 19416
rect 96624 19136 96864 19274
rect 96624 19072 96632 19136
rect 96696 19072 96712 19136
rect 96776 19072 96792 19136
rect 96856 19072 96864 19136
rect 95744 18856 95984 18994
rect 95744 18792 95752 18856
rect 95816 18792 95832 18856
rect 95896 18792 95912 18856
rect 95976 18792 95984 18856
rect 94864 18576 95104 18714
rect 94864 18512 94872 18576
rect 94936 18512 94952 18576
rect 95016 18512 95032 18576
rect 95096 18512 95104 18576
rect 93984 18296 94224 18434
rect 93984 18232 93992 18296
rect 94056 18232 94072 18296
rect 94136 18232 94152 18296
rect 94216 18232 94224 18296
rect 93984 17940 94224 18232
rect 94864 17940 95104 18512
rect 95744 17940 95984 18792
rect 96624 17940 96864 19072
rect 97504 17940 97744 19352
rect 112504 19492 112512 19556
rect 112576 19492 112592 19556
rect 112656 19492 112672 19556
rect 112736 19492 112744 19556
rect 142504 19556 142744 19557
rect 111624 19276 111864 19277
rect 111624 19212 111632 19276
rect 111696 19212 111712 19276
rect 111776 19212 111792 19276
rect 111856 19212 111864 19276
rect 110744 18996 110984 18997
rect 110744 18932 110752 18996
rect 110816 18932 110832 18996
rect 110896 18932 110912 18996
rect 110976 18932 110984 18996
rect 109864 18716 110104 18717
rect 109864 18652 109872 18716
rect 109936 18652 109952 18716
rect 110016 18652 110032 18716
rect 110096 18652 110104 18716
rect 108984 18436 109224 18437
rect 108984 18372 108992 18436
rect 109056 18372 109072 18436
rect 109136 18372 109152 18436
rect 109216 18372 109224 18436
rect 108984 17940 109224 18372
rect 109864 17940 110104 18652
rect 110744 17940 110984 18932
rect 111624 17940 111864 19212
rect 112504 17940 112744 19492
rect 127504 19416 127744 19554
rect 127504 19352 127512 19416
rect 127576 19352 127592 19416
rect 127656 19352 127672 19416
rect 127736 19352 127744 19416
rect 126624 19136 126864 19274
rect 126624 19072 126632 19136
rect 126696 19072 126712 19136
rect 126776 19072 126792 19136
rect 126856 19072 126864 19136
rect 125744 18856 125984 18994
rect 125744 18792 125752 18856
rect 125816 18792 125832 18856
rect 125896 18792 125912 18856
rect 125976 18792 125984 18856
rect 124864 18576 125104 18714
rect 124864 18512 124872 18576
rect 124936 18512 124952 18576
rect 125016 18512 125032 18576
rect 125096 18512 125104 18576
rect 123984 18296 124224 18434
rect 123984 18232 123992 18296
rect 124056 18232 124072 18296
rect 124136 18232 124152 18296
rect 124216 18232 124224 18296
rect 123984 17940 124224 18232
rect 124864 17940 125104 18512
rect 125744 17940 125984 18792
rect 126624 17940 126864 19072
rect 127504 17940 127744 19352
rect 142504 19492 142512 19556
rect 142576 19492 142592 19556
rect 142656 19492 142672 19556
rect 142736 19492 142744 19556
rect 172504 19556 172744 19557
rect 141624 19276 141864 19277
rect 141624 19212 141632 19276
rect 141696 19212 141712 19276
rect 141776 19212 141792 19276
rect 141856 19212 141864 19276
rect 140744 18996 140984 18997
rect 140744 18932 140752 18996
rect 140816 18932 140832 18996
rect 140896 18932 140912 18996
rect 140976 18932 140984 18996
rect 139864 18716 140104 18717
rect 139864 18652 139872 18716
rect 139936 18652 139952 18716
rect 140016 18652 140032 18716
rect 140096 18652 140104 18716
rect 138984 18436 139224 18437
rect 138984 18372 138992 18436
rect 139056 18372 139072 18436
rect 139136 18372 139152 18436
rect 139216 18372 139224 18436
rect 138984 17940 139224 18372
rect 139864 17940 140104 18652
rect 140744 17940 140984 18932
rect 141624 17940 141864 19212
rect 142504 17940 142744 19492
rect 157504 19416 157744 19554
rect 157504 19352 157512 19416
rect 157576 19352 157592 19416
rect 157656 19352 157672 19416
rect 157736 19352 157744 19416
rect 156624 19136 156864 19274
rect 156624 19072 156632 19136
rect 156696 19072 156712 19136
rect 156776 19072 156792 19136
rect 156856 19072 156864 19136
rect 155744 18856 155984 18994
rect 155744 18792 155752 18856
rect 155816 18792 155832 18856
rect 155896 18792 155912 18856
rect 155976 18792 155984 18856
rect 154864 18576 155104 18714
rect 154864 18512 154872 18576
rect 154936 18512 154952 18576
rect 155016 18512 155032 18576
rect 155096 18512 155104 18576
rect 153984 18296 154224 18434
rect 153984 18232 153992 18296
rect 154056 18232 154072 18296
rect 154136 18232 154152 18296
rect 154216 18232 154224 18296
rect 153984 17940 154224 18232
rect 154864 17940 155104 18512
rect 155744 17940 155984 18792
rect 156624 17940 156864 19072
rect 157504 17940 157744 19352
rect 172504 19492 172512 19556
rect 172576 19492 172592 19556
rect 172656 19492 172672 19556
rect 172736 19492 172744 19556
rect 171624 19276 171864 19277
rect 171624 19212 171632 19276
rect 171696 19212 171712 19276
rect 171776 19212 171792 19276
rect 171856 19212 171864 19276
rect 170744 18996 170984 18997
rect 170744 18932 170752 18996
rect 170816 18932 170832 18996
rect 170896 18932 170912 18996
rect 170976 18932 170984 18996
rect 169864 18716 170104 18717
rect 169864 18652 169872 18716
rect 169936 18652 169952 18716
rect 170016 18652 170032 18716
rect 170096 18652 170104 18716
rect 168984 18436 169224 18437
rect 168984 18372 168992 18436
rect 169056 18372 169072 18436
rect 169136 18372 169152 18436
rect 169216 18372 169224 18436
rect 168984 17940 169224 18372
rect 169864 17940 170104 18652
rect 170744 17940 170984 18932
rect 171624 17940 171864 19212
rect 172504 17940 172744 19492
rect 187504 19416 187744 19554
rect 187504 19352 187512 19416
rect 187576 19352 187592 19416
rect 187656 19352 187672 19416
rect 187736 19352 187744 19416
rect 186624 19136 186864 19274
rect 186624 19072 186632 19136
rect 186696 19072 186712 19136
rect 186776 19072 186792 19136
rect 186856 19072 186864 19136
rect 185744 18856 185984 18994
rect 185744 18792 185752 18856
rect 185816 18792 185832 18856
rect 185896 18792 185912 18856
rect 185976 18792 185984 18856
rect 184864 18576 185104 18714
rect 184864 18512 184872 18576
rect 184936 18512 184952 18576
rect 185016 18512 185032 18576
rect 185096 18512 185104 18576
rect 183984 18296 184224 18434
rect 183984 18232 183992 18296
rect 184056 18232 184072 18296
rect 184136 18232 184152 18296
rect 184216 18232 184224 18296
rect 183984 17940 184224 18232
rect 184864 17940 185104 18512
rect 185744 17940 185984 18792
rect 186624 17940 186864 19072
rect 187504 17940 187744 19352
rect 3984 -280 4224 60
rect 3984 -344 3992 -280
rect 4056 -344 4072 -280
rect 4136 -344 4152 -280
rect 4216 -344 4224 -280
rect 3984 -482 4224 -344
rect 4864 -560 5104 60
rect 4864 -624 4872 -560
rect 4936 -624 4952 -560
rect 5016 -624 5032 -560
rect 5096 -624 5104 -560
rect 4864 -762 5104 -624
rect 5744 -840 5984 60
rect 5744 -904 5752 -840
rect 5816 -904 5832 -840
rect 5896 -904 5912 -840
rect 5976 -904 5984 -840
rect 5744 -1042 5984 -904
rect 6624 -1120 6864 60
rect 6624 -1184 6632 -1120
rect 6696 -1184 6712 -1120
rect 6776 -1184 6792 -1120
rect 6856 -1184 6864 -1120
rect 6624 -1322 6864 -1184
rect 7504 -1400 7744 60
rect 18984 -420 19224 60
rect 18984 -484 18992 -420
rect 19056 -484 19072 -420
rect 19136 -484 19152 -420
rect 19216 -484 19224 -420
rect 18984 -485 19224 -484
rect 19864 -700 20104 60
rect 19864 -764 19872 -700
rect 19936 -764 19952 -700
rect 20016 -764 20032 -700
rect 20096 -764 20104 -700
rect 19864 -765 20104 -764
rect 20744 -980 20984 60
rect 20744 -1044 20752 -980
rect 20816 -1044 20832 -980
rect 20896 -1044 20912 -980
rect 20976 -1044 20984 -980
rect 20744 -1045 20984 -1044
rect 21624 -1260 21864 60
rect 21624 -1324 21632 -1260
rect 21696 -1324 21712 -1260
rect 21776 -1324 21792 -1260
rect 21856 -1324 21864 -1260
rect 21624 -1325 21864 -1324
rect 7504 -1464 7512 -1400
rect 7576 -1464 7592 -1400
rect 7656 -1464 7672 -1400
rect 7736 -1464 7744 -1400
rect 7504 -1602 7744 -1464
rect 22504 -1540 22744 60
rect 33984 -280 34224 60
rect 33984 -344 33992 -280
rect 34056 -344 34072 -280
rect 34136 -344 34152 -280
rect 34216 -344 34224 -280
rect 33984 -482 34224 -344
rect 34864 -560 35104 60
rect 34864 -624 34872 -560
rect 34936 -624 34952 -560
rect 35016 -624 35032 -560
rect 35096 -624 35104 -560
rect 34864 -762 35104 -624
rect 35744 -840 35984 60
rect 35744 -904 35752 -840
rect 35816 -904 35832 -840
rect 35896 -904 35912 -840
rect 35976 -904 35984 -840
rect 35744 -1042 35984 -904
rect 36624 -1120 36864 60
rect 36624 -1184 36632 -1120
rect 36696 -1184 36712 -1120
rect 36776 -1184 36792 -1120
rect 36856 -1184 36864 -1120
rect 36624 -1322 36864 -1184
rect 22504 -1604 22512 -1540
rect 22576 -1604 22592 -1540
rect 22656 -1604 22672 -1540
rect 22736 -1604 22744 -1540
rect 37504 -1400 37744 60
rect 48984 -420 49224 60
rect 48984 -484 48992 -420
rect 49056 -484 49072 -420
rect 49136 -484 49152 -420
rect 49216 -484 49224 -420
rect 48984 -485 49224 -484
rect 49864 -700 50104 60
rect 49864 -764 49872 -700
rect 49936 -764 49952 -700
rect 50016 -764 50032 -700
rect 50096 -764 50104 -700
rect 49864 -765 50104 -764
rect 50744 -980 50984 60
rect 50744 -1044 50752 -980
rect 50816 -1044 50832 -980
rect 50896 -1044 50912 -980
rect 50976 -1044 50984 -980
rect 50744 -1045 50984 -1044
rect 51624 -1260 51864 60
rect 51624 -1324 51632 -1260
rect 51696 -1324 51712 -1260
rect 51776 -1324 51792 -1260
rect 51856 -1324 51864 -1260
rect 51624 -1325 51864 -1324
rect 37504 -1464 37512 -1400
rect 37576 -1464 37592 -1400
rect 37656 -1464 37672 -1400
rect 37736 -1464 37744 -1400
rect 37504 -1602 37744 -1464
rect 52504 -1540 52744 60
rect 63984 -280 64224 60
rect 63984 -344 63992 -280
rect 64056 -344 64072 -280
rect 64136 -344 64152 -280
rect 64216 -344 64224 -280
rect 63984 -482 64224 -344
rect 64864 -560 65104 60
rect 64864 -624 64872 -560
rect 64936 -624 64952 -560
rect 65016 -624 65032 -560
rect 65096 -624 65104 -560
rect 64864 -762 65104 -624
rect 65744 -840 65984 60
rect 65744 -904 65752 -840
rect 65816 -904 65832 -840
rect 65896 -904 65912 -840
rect 65976 -904 65984 -840
rect 65744 -1042 65984 -904
rect 66624 -1120 66864 60
rect 66624 -1184 66632 -1120
rect 66696 -1184 66712 -1120
rect 66776 -1184 66792 -1120
rect 66856 -1184 66864 -1120
rect 66624 -1322 66864 -1184
rect 22504 -1605 22744 -1604
rect 52504 -1604 52512 -1540
rect 52576 -1604 52592 -1540
rect 52656 -1604 52672 -1540
rect 52736 -1604 52744 -1540
rect 67504 -1400 67744 60
rect 78984 -420 79224 60
rect 78984 -484 78992 -420
rect 79056 -484 79072 -420
rect 79136 -484 79152 -420
rect 79216 -484 79224 -420
rect 78984 -485 79224 -484
rect 79864 -700 80104 60
rect 79864 -764 79872 -700
rect 79936 -764 79952 -700
rect 80016 -764 80032 -700
rect 80096 -764 80104 -700
rect 79864 -765 80104 -764
rect 80744 -980 80984 60
rect 80744 -1044 80752 -980
rect 80816 -1044 80832 -980
rect 80896 -1044 80912 -980
rect 80976 -1044 80984 -980
rect 80744 -1045 80984 -1044
rect 81624 -1260 81864 60
rect 81624 -1324 81632 -1260
rect 81696 -1324 81712 -1260
rect 81776 -1324 81792 -1260
rect 81856 -1324 81864 -1260
rect 81624 -1325 81864 -1324
rect 67504 -1464 67512 -1400
rect 67576 -1464 67592 -1400
rect 67656 -1464 67672 -1400
rect 67736 -1464 67744 -1400
rect 67504 -1602 67744 -1464
rect 82504 -1540 82744 60
rect 93984 -280 94224 60
rect 93984 -344 93992 -280
rect 94056 -344 94072 -280
rect 94136 -344 94152 -280
rect 94216 -344 94224 -280
rect 93984 -482 94224 -344
rect 94864 -560 95104 60
rect 94864 -624 94872 -560
rect 94936 -624 94952 -560
rect 95016 -624 95032 -560
rect 95096 -624 95104 -560
rect 94864 -762 95104 -624
rect 95744 -840 95984 60
rect 95744 -904 95752 -840
rect 95816 -904 95832 -840
rect 95896 -904 95912 -840
rect 95976 -904 95984 -840
rect 95744 -1042 95984 -904
rect 96624 -1120 96864 60
rect 96624 -1184 96632 -1120
rect 96696 -1184 96712 -1120
rect 96776 -1184 96792 -1120
rect 96856 -1184 96864 -1120
rect 96624 -1322 96864 -1184
rect 52504 -1605 52744 -1604
rect 82504 -1604 82512 -1540
rect 82576 -1604 82592 -1540
rect 82656 -1604 82672 -1540
rect 82736 -1604 82744 -1540
rect 97504 -1400 97744 60
rect 108984 -420 109224 60
rect 108984 -484 108992 -420
rect 109056 -484 109072 -420
rect 109136 -484 109152 -420
rect 109216 -484 109224 -420
rect 108984 -485 109224 -484
rect 109864 -700 110104 60
rect 109864 -764 109872 -700
rect 109936 -764 109952 -700
rect 110016 -764 110032 -700
rect 110096 -764 110104 -700
rect 109864 -765 110104 -764
rect 110744 -980 110984 60
rect 110744 -1044 110752 -980
rect 110816 -1044 110832 -980
rect 110896 -1044 110912 -980
rect 110976 -1044 110984 -980
rect 110744 -1045 110984 -1044
rect 111624 -1260 111864 60
rect 111624 -1324 111632 -1260
rect 111696 -1324 111712 -1260
rect 111776 -1324 111792 -1260
rect 111856 -1324 111864 -1260
rect 111624 -1325 111864 -1324
rect 97504 -1464 97512 -1400
rect 97576 -1464 97592 -1400
rect 97656 -1464 97672 -1400
rect 97736 -1464 97744 -1400
rect 97504 -1602 97744 -1464
rect 112504 -1540 112744 60
rect 123984 -280 124224 60
rect 123984 -344 123992 -280
rect 124056 -344 124072 -280
rect 124136 -344 124152 -280
rect 124216 -344 124224 -280
rect 123984 -482 124224 -344
rect 124864 -560 125104 60
rect 124864 -624 124872 -560
rect 124936 -624 124952 -560
rect 125016 -624 125032 -560
rect 125096 -624 125104 -560
rect 124864 -762 125104 -624
rect 125744 -840 125984 60
rect 125744 -904 125752 -840
rect 125816 -904 125832 -840
rect 125896 -904 125912 -840
rect 125976 -904 125984 -840
rect 125744 -1042 125984 -904
rect 126624 -1120 126864 60
rect 126624 -1184 126632 -1120
rect 126696 -1184 126712 -1120
rect 126776 -1184 126792 -1120
rect 126856 -1184 126864 -1120
rect 126624 -1322 126864 -1184
rect 82504 -1605 82744 -1604
rect 112504 -1604 112512 -1540
rect 112576 -1604 112592 -1540
rect 112656 -1604 112672 -1540
rect 112736 -1604 112744 -1540
rect 127504 -1400 127744 60
rect 138984 -420 139224 60
rect 138984 -484 138992 -420
rect 139056 -484 139072 -420
rect 139136 -484 139152 -420
rect 139216 -484 139224 -420
rect 138984 -485 139224 -484
rect 139864 -700 140104 60
rect 139864 -764 139872 -700
rect 139936 -764 139952 -700
rect 140016 -764 140032 -700
rect 140096 -764 140104 -700
rect 139864 -765 140104 -764
rect 140744 -980 140984 60
rect 140744 -1044 140752 -980
rect 140816 -1044 140832 -980
rect 140896 -1044 140912 -980
rect 140976 -1044 140984 -980
rect 140744 -1045 140984 -1044
rect 141624 -1260 141864 60
rect 141624 -1324 141632 -1260
rect 141696 -1324 141712 -1260
rect 141776 -1324 141792 -1260
rect 141856 -1324 141864 -1260
rect 141624 -1325 141864 -1324
rect 127504 -1464 127512 -1400
rect 127576 -1464 127592 -1400
rect 127656 -1464 127672 -1400
rect 127736 -1464 127744 -1400
rect 127504 -1602 127744 -1464
rect 142504 -1540 142744 60
rect 153984 -280 154224 60
rect 153984 -344 153992 -280
rect 154056 -344 154072 -280
rect 154136 -344 154152 -280
rect 154216 -344 154224 -280
rect 153984 -482 154224 -344
rect 154864 -560 155104 60
rect 154864 -624 154872 -560
rect 154936 -624 154952 -560
rect 155016 -624 155032 -560
rect 155096 -624 155104 -560
rect 154864 -762 155104 -624
rect 155744 -840 155984 60
rect 155744 -904 155752 -840
rect 155816 -904 155832 -840
rect 155896 -904 155912 -840
rect 155976 -904 155984 -840
rect 155744 -1042 155984 -904
rect 156624 -1120 156864 60
rect 156624 -1184 156632 -1120
rect 156696 -1184 156712 -1120
rect 156776 -1184 156792 -1120
rect 156856 -1184 156864 -1120
rect 156624 -1322 156864 -1184
rect 112504 -1605 112744 -1604
rect 142504 -1604 142512 -1540
rect 142576 -1604 142592 -1540
rect 142656 -1604 142672 -1540
rect 142736 -1604 142744 -1540
rect 157504 -1400 157744 60
rect 168984 -420 169224 60
rect 168984 -484 168992 -420
rect 169056 -484 169072 -420
rect 169136 -484 169152 -420
rect 169216 -484 169224 -420
rect 168984 -485 169224 -484
rect 169864 -700 170104 60
rect 169864 -764 169872 -700
rect 169936 -764 169952 -700
rect 170016 -764 170032 -700
rect 170096 -764 170104 -700
rect 169864 -765 170104 -764
rect 170744 -980 170984 60
rect 170744 -1044 170752 -980
rect 170816 -1044 170832 -980
rect 170896 -1044 170912 -980
rect 170976 -1044 170984 -980
rect 170744 -1045 170984 -1044
rect 171624 -1260 171864 60
rect 171624 -1324 171632 -1260
rect 171696 -1324 171712 -1260
rect 171776 -1324 171792 -1260
rect 171856 -1324 171864 -1260
rect 171624 -1325 171864 -1324
rect 157504 -1464 157512 -1400
rect 157576 -1464 157592 -1400
rect 157656 -1464 157672 -1400
rect 157736 -1464 157744 -1400
rect 157504 -1602 157744 -1464
rect 172504 -1540 172744 60
rect 183984 -280 184224 60
rect 183984 -344 183992 -280
rect 184056 -344 184072 -280
rect 184136 -344 184152 -280
rect 184216 -344 184224 -280
rect 183984 -482 184224 -344
rect 184864 -560 185104 60
rect 184864 -624 184872 -560
rect 184936 -624 184952 -560
rect 185016 -624 185032 -560
rect 185096 -624 185104 -560
rect 184864 -762 185104 -624
rect 185744 -840 185984 60
rect 185744 -904 185752 -840
rect 185816 -904 185832 -840
rect 185896 -904 185912 -840
rect 185976 -904 185984 -840
rect 185744 -1042 185984 -904
rect 186624 -1120 186864 60
rect 186624 -1184 186632 -1120
rect 186696 -1184 186712 -1120
rect 186776 -1184 186792 -1120
rect 186856 -1184 186864 -1120
rect 186624 -1322 186864 -1184
rect 142504 -1605 142744 -1604
rect 172504 -1604 172512 -1540
rect 172576 -1604 172592 -1540
rect 172656 -1604 172672 -1540
rect 172736 -1604 172744 -1540
rect 187504 -1400 187744 60
rect 200182 -342 200242 18294
rect 200322 -482 200382 18434
rect 200462 -622 200522 18574
rect 200602 -762 200662 18714
rect 200742 -902 200802 18854
rect 200882 -1042 200942 18994
rect 201022 -1182 201082 19134
rect 201162 -1322 201222 19274
rect 187504 -1464 187512 -1400
rect 187576 -1464 187592 -1400
rect 187656 -1464 187672 -1400
rect 187736 -1464 187744 -1400
rect 201302 -1462 201362 19414
rect 187504 -1602 187744 -1464
rect 201442 -1602 201502 19554
rect 172504 -1605 172744 -1604
<< obsm4 >>
rect 3984 60 187744 17940
<< labels >>
rlabel metal3 s -400 3000 60 3120 4 caravel_clk
port 1 nsew signal input
rlabel metal3 s -400 8984 60 9104 4 caravel_clk2
port 2 nsew signal input
rlabel metal3 s -400 14968 60 15088 4 caravel_rstn
port 3 nsew signal input
rlabel metal2 s 1858 17940 1914 18400 6 la_data_in_core[0]
port 4 nsew signal output
rlabel metal2 s 45466 17940 45522 18400 6 la_data_in_core[100]
port 5 nsew signal output
rlabel metal2 s 45926 17940 45982 18400 6 la_data_in_core[101]
port 6 nsew signal output
rlabel metal2 s 46386 17940 46442 18400 6 la_data_in_core[102]
port 7 nsew signal output
rlabel metal2 s 46754 17940 46810 18400 6 la_data_in_core[103]
port 8 nsew signal output
rlabel metal2 s 47214 17940 47270 18400 6 la_data_in_core[104]
port 9 nsew signal output
rlabel metal2 s 47674 17940 47730 18400 6 la_data_in_core[105]
port 10 nsew signal output
rlabel metal2 s 48134 17940 48190 18400 6 la_data_in_core[106]
port 11 nsew signal output
rlabel metal2 s 48502 17940 48558 18400 6 la_data_in_core[107]
port 12 nsew signal output
rlabel metal2 s 48962 17940 49018 18400 6 la_data_in_core[108]
port 13 nsew signal output
rlabel metal2 s 49422 17940 49478 18400 6 la_data_in_core[109]
port 14 nsew signal output
rlabel metal2 s 6274 17940 6330 18400 6 la_data_in_core[10]
port 15 nsew signal output
rlabel metal2 s 49790 17940 49846 18400 6 la_data_in_core[110]
port 16 nsew signal output
rlabel metal2 s 50250 17940 50306 18400 6 la_data_in_core[111]
port 17 nsew signal output
rlabel metal2 s 50710 17940 50766 18400 6 la_data_in_core[112]
port 18 nsew signal output
rlabel metal2 s 51170 17940 51226 18400 6 la_data_in_core[113]
port 19 nsew signal output
rlabel metal2 s 51538 17940 51594 18400 6 la_data_in_core[114]
port 20 nsew signal output
rlabel metal2 s 51998 17940 52054 18400 6 la_data_in_core[115]
port 21 nsew signal output
rlabel metal2 s 52458 17940 52514 18400 6 la_data_in_core[116]
port 22 nsew signal output
rlabel metal2 s 52918 17940 52974 18400 6 la_data_in_core[117]
port 23 nsew signal output
rlabel metal2 s 53286 17940 53342 18400 6 la_data_in_core[118]
port 24 nsew signal output
rlabel metal2 s 53746 17940 53802 18400 6 la_data_in_core[119]
port 25 nsew signal output
rlabel metal2 s 6734 17940 6790 18400 6 la_data_in_core[11]
port 26 nsew signal output
rlabel metal2 s 54206 17940 54262 18400 6 la_data_in_core[120]
port 27 nsew signal output
rlabel metal2 s 54666 17940 54722 18400 6 la_data_in_core[121]
port 28 nsew signal output
rlabel metal2 s 55034 17940 55090 18400 6 la_data_in_core[122]
port 29 nsew signal output
rlabel metal2 s 55494 17940 55550 18400 6 la_data_in_core[123]
port 30 nsew signal output
rlabel metal2 s 55954 17940 56010 18400 6 la_data_in_core[124]
port 31 nsew signal output
rlabel metal2 s 56322 17940 56378 18400 6 la_data_in_core[125]
port 32 nsew signal output
rlabel metal2 s 56782 17940 56838 18400 6 la_data_in_core[126]
port 33 nsew signal output
rlabel metal2 s 57242 17940 57298 18400 6 la_data_in_core[127]
port 34 nsew signal output
rlabel metal2 s 7102 17940 7158 18400 6 la_data_in_core[12]
port 35 nsew signal output
rlabel metal2 s 7562 17940 7618 18400 6 la_data_in_core[13]
port 36 nsew signal output
rlabel metal2 s 8022 17940 8078 18400 6 la_data_in_core[14]
port 37 nsew signal output
rlabel metal2 s 8390 17940 8446 18400 6 la_data_in_core[15]
port 38 nsew signal output
rlabel metal2 s 8850 17940 8906 18400 6 la_data_in_core[16]
port 39 nsew signal output
rlabel metal2 s 9310 17940 9366 18400 6 la_data_in_core[17]
port 40 nsew signal output
rlabel metal2 s 9770 17940 9826 18400 6 la_data_in_core[18]
port 41 nsew signal output
rlabel metal2 s 10138 17940 10194 18400 6 la_data_in_core[19]
port 42 nsew signal output
rlabel metal2 s 2318 17940 2374 18400 6 la_data_in_core[1]
port 43 nsew signal output
rlabel metal2 s 10598 17940 10654 18400 6 la_data_in_core[20]
port 44 nsew signal output
rlabel metal2 s 11058 17940 11114 18400 6 la_data_in_core[21]
port 45 nsew signal output
rlabel metal2 s 11518 17940 11574 18400 6 la_data_in_core[22]
port 46 nsew signal output
rlabel metal2 s 11886 17940 11942 18400 6 la_data_in_core[23]
port 47 nsew signal output
rlabel metal2 s 12346 17940 12402 18400 6 la_data_in_core[24]
port 48 nsew signal output
rlabel metal2 s 12806 17940 12862 18400 6 la_data_in_core[25]
port 49 nsew signal output
rlabel metal2 s 13266 17940 13322 18400 6 la_data_in_core[26]
port 50 nsew signal output
rlabel metal2 s 13634 17940 13690 18400 6 la_data_in_core[27]
port 51 nsew signal output
rlabel metal2 s 14094 17940 14150 18400 6 la_data_in_core[28]
port 52 nsew signal output
rlabel metal2 s 14554 17940 14610 18400 6 la_data_in_core[29]
port 53 nsew signal output
rlabel metal2 s 2778 17940 2834 18400 6 la_data_in_core[2]
port 54 nsew signal output
rlabel metal2 s 15014 17940 15070 18400 6 la_data_in_core[30]
port 55 nsew signal output
rlabel metal2 s 15382 17940 15438 18400 6 la_data_in_core[31]
port 56 nsew signal output
rlabel metal2 s 15842 17940 15898 18400 6 la_data_in_core[32]
port 57 nsew signal output
rlabel metal2 s 16302 17940 16358 18400 6 la_data_in_core[33]
port 58 nsew signal output
rlabel metal2 s 16670 17940 16726 18400 6 la_data_in_core[34]
port 59 nsew signal output
rlabel metal2 s 17130 17940 17186 18400 6 la_data_in_core[35]
port 60 nsew signal output
rlabel metal2 s 17590 17940 17646 18400 6 la_data_in_core[36]
port 61 nsew signal output
rlabel metal2 s 18050 17940 18106 18400 6 la_data_in_core[37]
port 62 nsew signal output
rlabel metal2 s 18418 17940 18474 18400 6 la_data_in_core[38]
port 63 nsew signal output
rlabel metal2 s 18878 17940 18934 18400 6 la_data_in_core[39]
port 64 nsew signal output
rlabel metal2 s 3238 17940 3294 18400 6 la_data_in_core[3]
port 65 nsew signal output
rlabel metal2 s 19338 17940 19394 18400 6 la_data_in_core[40]
port 66 nsew signal output
rlabel metal2 s 19798 17940 19854 18400 6 la_data_in_core[41]
port 67 nsew signal output
rlabel metal2 s 20166 17940 20222 18400 6 la_data_in_core[42]
port 68 nsew signal output
rlabel metal2 s 20626 17940 20682 18400 6 la_data_in_core[43]
port 69 nsew signal output
rlabel metal2 s 21086 17940 21142 18400 6 la_data_in_core[44]
port 70 nsew signal output
rlabel metal2 s 21546 17940 21602 18400 6 la_data_in_core[45]
port 71 nsew signal output
rlabel metal2 s 21914 17940 21970 18400 6 la_data_in_core[46]
port 72 nsew signal output
rlabel metal2 s 22374 17940 22430 18400 6 la_data_in_core[47]
port 73 nsew signal output
rlabel metal2 s 22834 17940 22890 18400 6 la_data_in_core[48]
port 74 nsew signal output
rlabel metal2 s 23294 17940 23350 18400 6 la_data_in_core[49]
port 75 nsew signal output
rlabel metal2 s 3606 17940 3662 18400 6 la_data_in_core[4]
port 76 nsew signal output
rlabel metal2 s 23662 17940 23718 18400 6 la_data_in_core[50]
port 77 nsew signal output
rlabel metal2 s 24122 17940 24178 18400 6 la_data_in_core[51]
port 78 nsew signal output
rlabel metal2 s 24582 17940 24638 18400 6 la_data_in_core[52]
port 79 nsew signal output
rlabel metal2 s 24950 17940 25006 18400 6 la_data_in_core[53]
port 80 nsew signal output
rlabel metal2 s 25410 17940 25466 18400 6 la_data_in_core[54]
port 81 nsew signal output
rlabel metal2 s 25870 17940 25926 18400 6 la_data_in_core[55]
port 82 nsew signal output
rlabel metal2 s 26330 17940 26386 18400 6 la_data_in_core[56]
port 83 nsew signal output
rlabel metal2 s 26698 17940 26754 18400 6 la_data_in_core[57]
port 84 nsew signal output
rlabel metal2 s 27158 17940 27214 18400 6 la_data_in_core[58]
port 85 nsew signal output
rlabel metal2 s 27618 17940 27674 18400 6 la_data_in_core[59]
port 86 nsew signal output
rlabel metal2 s 4066 17940 4122 18400 6 la_data_in_core[5]
port 87 nsew signal output
rlabel metal2 s 28078 17940 28134 18400 6 la_data_in_core[60]
port 88 nsew signal output
rlabel metal2 s 28446 17940 28502 18400 6 la_data_in_core[61]
port 89 nsew signal output
rlabel metal2 s 28906 17940 28962 18400 6 la_data_in_core[62]
port 90 nsew signal output
rlabel metal2 s 29366 17940 29422 18400 6 la_data_in_core[63]
port 91 nsew signal output
rlabel metal2 s 29826 17940 29882 18400 6 la_data_in_core[64]
port 92 nsew signal output
rlabel metal2 s 30194 17940 30250 18400 6 la_data_in_core[65]
port 93 nsew signal output
rlabel metal2 s 30654 17940 30710 18400 6 la_data_in_core[66]
port 94 nsew signal output
rlabel metal2 s 31114 17940 31170 18400 6 la_data_in_core[67]
port 95 nsew signal output
rlabel metal2 s 31574 17940 31630 18400 6 la_data_in_core[68]
port 96 nsew signal output
rlabel metal2 s 31942 17940 31998 18400 6 la_data_in_core[69]
port 97 nsew signal output
rlabel metal2 s 4526 17940 4582 18400 6 la_data_in_core[6]
port 98 nsew signal output
rlabel metal2 s 32402 17940 32458 18400 6 la_data_in_core[70]
port 99 nsew signal output
rlabel metal2 s 32862 17940 32918 18400 6 la_data_in_core[71]
port 100 nsew signal output
rlabel metal2 s 33230 17940 33286 18400 6 la_data_in_core[72]
port 101 nsew signal output
rlabel metal2 s 33690 17940 33746 18400 6 la_data_in_core[73]
port 102 nsew signal output
rlabel metal2 s 34150 17940 34206 18400 6 la_data_in_core[74]
port 103 nsew signal output
rlabel metal2 s 34610 17940 34666 18400 6 la_data_in_core[75]
port 104 nsew signal output
rlabel metal2 s 34978 17940 35034 18400 6 la_data_in_core[76]
port 105 nsew signal output
rlabel metal2 s 35438 17940 35494 18400 6 la_data_in_core[77]
port 106 nsew signal output
rlabel metal2 s 35898 17940 35954 18400 6 la_data_in_core[78]
port 107 nsew signal output
rlabel metal2 s 36358 17940 36414 18400 6 la_data_in_core[79]
port 108 nsew signal output
rlabel metal2 s 4986 17940 5042 18400 6 la_data_in_core[7]
port 109 nsew signal output
rlabel metal2 s 36726 17940 36782 18400 6 la_data_in_core[80]
port 110 nsew signal output
rlabel metal2 s 37186 17940 37242 18400 6 la_data_in_core[81]
port 111 nsew signal output
rlabel metal2 s 37646 17940 37702 18400 6 la_data_in_core[82]
port 112 nsew signal output
rlabel metal2 s 38106 17940 38162 18400 6 la_data_in_core[83]
port 113 nsew signal output
rlabel metal2 s 38474 17940 38530 18400 6 la_data_in_core[84]
port 114 nsew signal output
rlabel metal2 s 38934 17940 38990 18400 6 la_data_in_core[85]
port 115 nsew signal output
rlabel metal2 s 39394 17940 39450 18400 6 la_data_in_core[86]
port 116 nsew signal output
rlabel metal2 s 39854 17940 39910 18400 6 la_data_in_core[87]
port 117 nsew signal output
rlabel metal2 s 40222 17940 40278 18400 6 la_data_in_core[88]
port 118 nsew signal output
rlabel metal2 s 40682 17940 40738 18400 6 la_data_in_core[89]
port 119 nsew signal output
rlabel metal2 s 5354 17940 5410 18400 6 la_data_in_core[8]
port 120 nsew signal output
rlabel metal2 s 41142 17940 41198 18400 6 la_data_in_core[90]
port 121 nsew signal output
rlabel metal2 s 41510 17940 41566 18400 6 la_data_in_core[91]
port 122 nsew signal output
rlabel metal2 s 41970 17940 42026 18400 6 la_data_in_core[92]
port 123 nsew signal output
rlabel metal2 s 42430 17940 42486 18400 6 la_data_in_core[93]
port 124 nsew signal output
rlabel metal2 s 42890 17940 42946 18400 6 la_data_in_core[94]
port 125 nsew signal output
rlabel metal2 s 43258 17940 43314 18400 6 la_data_in_core[95]
port 126 nsew signal output
rlabel metal2 s 43718 17940 43774 18400 6 la_data_in_core[96]
port 127 nsew signal output
rlabel metal2 s 44178 17940 44234 18400 6 la_data_in_core[97]
port 128 nsew signal output
rlabel metal2 s 44638 17940 44694 18400 6 la_data_in_core[98]
port 129 nsew signal output
rlabel metal2 s 45006 17940 45062 18400 6 la_data_in_core[99]
port 130 nsew signal output
rlabel metal2 s 5814 17940 5870 18400 6 la_data_in_core[9]
port 131 nsew signal output
rlabel metal2 s 55954 -400 56010 60 8 la_data_in_mprj[0]
port 132 nsew signal output
rlabel metal2 s 99470 -400 99526 60 8 la_data_in_mprj[100]
port 133 nsew signal output
rlabel metal2 s 99930 -400 99986 60 8 la_data_in_mprj[101]
port 134 nsew signal output
rlabel metal2 s 100390 -400 100446 60 8 la_data_in_mprj[102]
port 135 nsew signal output
rlabel metal2 s 100850 -400 100906 60 8 la_data_in_mprj[103]
port 136 nsew signal output
rlabel metal2 s 101218 -400 101274 60 8 la_data_in_mprj[104]
port 137 nsew signal output
rlabel metal2 s 101678 -400 101734 60 8 la_data_in_mprj[105]
port 138 nsew signal output
rlabel metal2 s 102138 -400 102194 60 8 la_data_in_mprj[106]
port 139 nsew signal output
rlabel metal2 s 102598 -400 102654 60 8 la_data_in_mprj[107]
port 140 nsew signal output
rlabel metal2 s 102966 -400 103022 60 8 la_data_in_mprj[108]
port 141 nsew signal output
rlabel metal2 s 103426 -400 103482 60 8 la_data_in_mprj[109]
port 142 nsew signal output
rlabel metal2 s 60278 -400 60334 60 8 la_data_in_mprj[10]
port 143 nsew signal output
rlabel metal2 s 103886 -400 103942 60 8 la_data_in_mprj[110]
port 144 nsew signal output
rlabel metal2 s 104254 -400 104310 60 8 la_data_in_mprj[111]
port 145 nsew signal output
rlabel metal2 s 104714 -400 104770 60 8 la_data_in_mprj[112]
port 146 nsew signal output
rlabel metal2 s 105174 -400 105230 60 8 la_data_in_mprj[113]
port 147 nsew signal output
rlabel metal2 s 105634 -400 105690 60 8 la_data_in_mprj[114]
port 148 nsew signal output
rlabel metal2 s 106002 -400 106058 60 8 la_data_in_mprj[115]
port 149 nsew signal output
rlabel metal2 s 106462 -400 106518 60 8 la_data_in_mprj[116]
port 150 nsew signal output
rlabel metal2 s 106922 -400 106978 60 8 la_data_in_mprj[117]
port 151 nsew signal output
rlabel metal2 s 107382 -400 107438 60 8 la_data_in_mprj[118]
port 152 nsew signal output
rlabel metal2 s 107750 -400 107806 60 8 la_data_in_mprj[119]
port 153 nsew signal output
rlabel metal2 s 60738 -400 60794 60 8 la_data_in_mprj[11]
port 154 nsew signal output
rlabel metal2 s 108210 -400 108266 60 8 la_data_in_mprj[120]
port 155 nsew signal output
rlabel metal2 s 108670 -400 108726 60 8 la_data_in_mprj[121]
port 156 nsew signal output
rlabel metal2 s 109130 -400 109186 60 8 la_data_in_mprj[122]
port 157 nsew signal output
rlabel metal2 s 109498 -400 109554 60 8 la_data_in_mprj[123]
port 158 nsew signal output
rlabel metal2 s 109958 -400 110014 60 8 la_data_in_mprj[124]
port 159 nsew signal output
rlabel metal2 s 110418 -400 110474 60 8 la_data_in_mprj[125]
port 160 nsew signal output
rlabel metal2 s 110878 -400 110934 60 8 la_data_in_mprj[126]
port 161 nsew signal output
rlabel metal2 s 111246 -400 111302 60 8 la_data_in_mprj[127]
port 162 nsew signal output
rlabel metal2 s 61198 -400 61254 60 8 la_data_in_mprj[12]
port 163 nsew signal output
rlabel metal2 s 61566 -400 61622 60 8 la_data_in_mprj[13]
port 164 nsew signal output
rlabel metal2 s 62026 -400 62082 60 8 la_data_in_mprj[14]
port 165 nsew signal output
rlabel metal2 s 62486 -400 62542 60 8 la_data_in_mprj[15]
port 166 nsew signal output
rlabel metal2 s 62946 -400 63002 60 8 la_data_in_mprj[16]
port 167 nsew signal output
rlabel metal2 s 63314 -400 63370 60 8 la_data_in_mprj[17]
port 168 nsew signal output
rlabel metal2 s 63774 -400 63830 60 8 la_data_in_mprj[18]
port 169 nsew signal output
rlabel metal2 s 64234 -400 64290 60 8 la_data_in_mprj[19]
port 170 nsew signal output
rlabel metal2 s 56322 -400 56378 60 8 la_data_in_mprj[1]
port 171 nsew signal output
rlabel metal2 s 64602 -400 64658 60 8 la_data_in_mprj[20]
port 172 nsew signal output
rlabel metal2 s 65062 -400 65118 60 8 la_data_in_mprj[21]
port 173 nsew signal output
rlabel metal2 s 65522 -400 65578 60 8 la_data_in_mprj[22]
port 174 nsew signal output
rlabel metal2 s 65982 -400 66038 60 8 la_data_in_mprj[23]
port 175 nsew signal output
rlabel metal2 s 66350 -400 66406 60 8 la_data_in_mprj[24]
port 176 nsew signal output
rlabel metal2 s 66810 -400 66866 60 8 la_data_in_mprj[25]
port 177 nsew signal output
rlabel metal2 s 67270 -400 67326 60 8 la_data_in_mprj[26]
port 178 nsew signal output
rlabel metal2 s 67730 -400 67786 60 8 la_data_in_mprj[27]
port 179 nsew signal output
rlabel metal2 s 68098 -400 68154 60 8 la_data_in_mprj[28]
port 180 nsew signal output
rlabel metal2 s 68558 -400 68614 60 8 la_data_in_mprj[29]
port 181 nsew signal output
rlabel metal2 s 56782 -400 56838 60 8 la_data_in_mprj[2]
port 182 nsew signal output
rlabel metal2 s 69018 -400 69074 60 8 la_data_in_mprj[30]
port 183 nsew signal output
rlabel metal2 s 69478 -400 69534 60 8 la_data_in_mprj[31]
port 184 nsew signal output
rlabel metal2 s 69846 -400 69902 60 8 la_data_in_mprj[32]
port 185 nsew signal output
rlabel metal2 s 70306 -400 70362 60 8 la_data_in_mprj[33]
port 186 nsew signal output
rlabel metal2 s 70766 -400 70822 60 8 la_data_in_mprj[34]
port 187 nsew signal output
rlabel metal2 s 71226 -400 71282 60 8 la_data_in_mprj[35]
port 188 nsew signal output
rlabel metal2 s 71594 -400 71650 60 8 la_data_in_mprj[36]
port 189 nsew signal output
rlabel metal2 s 72054 -400 72110 60 8 la_data_in_mprj[37]
port 190 nsew signal output
rlabel metal2 s 72514 -400 72570 60 8 la_data_in_mprj[38]
port 191 nsew signal output
rlabel metal2 s 72882 -400 72938 60 8 la_data_in_mprj[39]
port 192 nsew signal output
rlabel metal2 s 57242 -400 57298 60 8 la_data_in_mprj[3]
port 193 nsew signal output
rlabel metal2 s 73342 -400 73398 60 8 la_data_in_mprj[40]
port 194 nsew signal output
rlabel metal2 s 73802 -400 73858 60 8 la_data_in_mprj[41]
port 195 nsew signal output
rlabel metal2 s 74262 -400 74318 60 8 la_data_in_mprj[42]
port 196 nsew signal output
rlabel metal2 s 74630 -400 74686 60 8 la_data_in_mprj[43]
port 197 nsew signal output
rlabel metal2 s 75090 -400 75146 60 8 la_data_in_mprj[44]
port 198 nsew signal output
rlabel metal2 s 75550 -400 75606 60 8 la_data_in_mprj[45]
port 199 nsew signal output
rlabel metal2 s 76010 -400 76066 60 8 la_data_in_mprj[46]
port 200 nsew signal output
rlabel metal2 s 76378 -400 76434 60 8 la_data_in_mprj[47]
port 201 nsew signal output
rlabel metal2 s 76838 -400 76894 60 8 la_data_in_mprj[48]
port 202 nsew signal output
rlabel metal2 s 77298 -400 77354 60 8 la_data_in_mprj[49]
port 203 nsew signal output
rlabel metal2 s 57702 -400 57758 60 8 la_data_in_mprj[4]
port 204 nsew signal output
rlabel metal2 s 77758 -400 77814 60 8 la_data_in_mprj[50]
port 205 nsew signal output
rlabel metal2 s 78126 -400 78182 60 8 la_data_in_mprj[51]
port 206 nsew signal output
rlabel metal2 s 78586 -400 78642 60 8 la_data_in_mprj[52]
port 207 nsew signal output
rlabel metal2 s 79046 -400 79102 60 8 la_data_in_mprj[53]
port 208 nsew signal output
rlabel metal2 s 79506 -400 79562 60 8 la_data_in_mprj[54]
port 209 nsew signal output
rlabel metal2 s 79874 -400 79930 60 8 la_data_in_mprj[55]
port 210 nsew signal output
rlabel metal2 s 80334 -400 80390 60 8 la_data_in_mprj[56]
port 211 nsew signal output
rlabel metal2 s 80794 -400 80850 60 8 la_data_in_mprj[57]
port 212 nsew signal output
rlabel metal2 s 81162 -400 81218 60 8 la_data_in_mprj[58]
port 213 nsew signal output
rlabel metal2 s 81622 -400 81678 60 8 la_data_in_mprj[59]
port 214 nsew signal output
rlabel metal2 s 58070 -400 58126 60 8 la_data_in_mprj[5]
port 215 nsew signal output
rlabel metal2 s 82082 -400 82138 60 8 la_data_in_mprj[60]
port 216 nsew signal output
rlabel metal2 s 82542 -400 82598 60 8 la_data_in_mprj[61]
port 217 nsew signal output
rlabel metal2 s 82910 -400 82966 60 8 la_data_in_mprj[62]
port 218 nsew signal output
rlabel metal2 s 83370 -400 83426 60 8 la_data_in_mprj[63]
port 219 nsew signal output
rlabel metal2 s 83830 -400 83886 60 8 la_data_in_mprj[64]
port 220 nsew signal output
rlabel metal2 s 84290 -400 84346 60 8 la_data_in_mprj[65]
port 221 nsew signal output
rlabel metal2 s 84658 -400 84714 60 8 la_data_in_mprj[66]
port 222 nsew signal output
rlabel metal2 s 85118 -400 85174 60 8 la_data_in_mprj[67]
port 223 nsew signal output
rlabel metal2 s 85578 -400 85634 60 8 la_data_in_mprj[68]
port 224 nsew signal output
rlabel metal2 s 86038 -400 86094 60 8 la_data_in_mprj[69]
port 225 nsew signal output
rlabel metal2 s 58530 -400 58586 60 8 la_data_in_mprj[6]
port 226 nsew signal output
rlabel metal2 s 86406 -400 86462 60 8 la_data_in_mprj[70]
port 227 nsew signal output
rlabel metal2 s 86866 -400 86922 60 8 la_data_in_mprj[71]
port 228 nsew signal output
rlabel metal2 s 87326 -400 87382 60 8 la_data_in_mprj[72]
port 229 nsew signal output
rlabel metal2 s 87786 -400 87842 60 8 la_data_in_mprj[73]
port 230 nsew signal output
rlabel metal2 s 88154 -400 88210 60 8 la_data_in_mprj[74]
port 231 nsew signal output
rlabel metal2 s 88614 -400 88670 60 8 la_data_in_mprj[75]
port 232 nsew signal output
rlabel metal2 s 89074 -400 89130 60 8 la_data_in_mprj[76]
port 233 nsew signal output
rlabel metal2 s 89442 -400 89498 60 8 la_data_in_mprj[77]
port 234 nsew signal output
rlabel metal2 s 89902 -400 89958 60 8 la_data_in_mprj[78]
port 235 nsew signal output
rlabel metal2 s 90362 -400 90418 60 8 la_data_in_mprj[79]
port 236 nsew signal output
rlabel metal2 s 58990 -400 59046 60 8 la_data_in_mprj[7]
port 237 nsew signal output
rlabel metal2 s 90822 -400 90878 60 8 la_data_in_mprj[80]
port 238 nsew signal output
rlabel metal2 s 91190 -400 91246 60 8 la_data_in_mprj[81]
port 239 nsew signal output
rlabel metal2 s 91650 -400 91706 60 8 la_data_in_mprj[82]
port 240 nsew signal output
rlabel metal2 s 92110 -400 92166 60 8 la_data_in_mprj[83]
port 241 nsew signal output
rlabel metal2 s 92570 -400 92626 60 8 la_data_in_mprj[84]
port 242 nsew signal output
rlabel metal2 s 92938 -400 92994 60 8 la_data_in_mprj[85]
port 243 nsew signal output
rlabel metal2 s 93398 -400 93454 60 8 la_data_in_mprj[86]
port 244 nsew signal output
rlabel metal2 s 93858 -400 93914 60 8 la_data_in_mprj[87]
port 245 nsew signal output
rlabel metal2 s 94318 -400 94374 60 8 la_data_in_mprj[88]
port 246 nsew signal output
rlabel metal2 s 94686 -400 94742 60 8 la_data_in_mprj[89]
port 247 nsew signal output
rlabel metal2 s 59450 -400 59506 60 8 la_data_in_mprj[8]
port 248 nsew signal output
rlabel metal2 s 95146 -400 95202 60 8 la_data_in_mprj[90]
port 249 nsew signal output
rlabel metal2 s 95606 -400 95662 60 8 la_data_in_mprj[91]
port 250 nsew signal output
rlabel metal2 s 96066 -400 96122 60 8 la_data_in_mprj[92]
port 251 nsew signal output
rlabel metal2 s 96434 -400 96490 60 8 la_data_in_mprj[93]
port 252 nsew signal output
rlabel metal2 s 96894 -400 96950 60 8 la_data_in_mprj[94]
port 253 nsew signal output
rlabel metal2 s 97354 -400 97410 60 8 la_data_in_mprj[95]
port 254 nsew signal output
rlabel metal2 s 97722 -400 97778 60 8 la_data_in_mprj[96]
port 255 nsew signal output
rlabel metal2 s 98182 -400 98238 60 8 la_data_in_mprj[97]
port 256 nsew signal output
rlabel metal2 s 98642 -400 98698 60 8 la_data_in_mprj[98]
port 257 nsew signal output
rlabel metal2 s 99102 -400 99158 60 8 la_data_in_mprj[99]
port 258 nsew signal output
rlabel metal2 s 59818 -400 59874 60 8 la_data_in_mprj[9]
port 259 nsew signal output
rlabel metal2 s 57702 17940 57758 18400 6 la_data_out_core[0]
port 260 nsew signal input
rlabel metal2 s 101218 17940 101274 18400 6 la_data_out_core[100]
port 261 nsew signal input
rlabel metal2 s 101678 17940 101734 18400 6 la_data_out_core[101]
port 262 nsew signal input
rlabel metal2 s 102138 17940 102194 18400 6 la_data_out_core[102]
port 263 nsew signal input
rlabel metal2 s 102598 17940 102654 18400 6 la_data_out_core[103]
port 264 nsew signal input
rlabel metal2 s 102966 17940 103022 18400 6 la_data_out_core[104]
port 265 nsew signal input
rlabel metal2 s 103426 17940 103482 18400 6 la_data_out_core[105]
port 266 nsew signal input
rlabel metal2 s 103886 17940 103942 18400 6 la_data_out_core[106]
port 267 nsew signal input
rlabel metal2 s 104254 17940 104310 18400 6 la_data_out_core[107]
port 268 nsew signal input
rlabel metal2 s 104714 17940 104770 18400 6 la_data_out_core[108]
port 269 nsew signal input
rlabel metal2 s 105174 17940 105230 18400 6 la_data_out_core[109]
port 270 nsew signal input
rlabel metal2 s 62026 17940 62082 18400 6 la_data_out_core[10]
port 271 nsew signal input
rlabel metal2 s 105634 17940 105690 18400 6 la_data_out_core[110]
port 272 nsew signal input
rlabel metal2 s 106002 17940 106058 18400 6 la_data_out_core[111]
port 273 nsew signal input
rlabel metal2 s 106462 17940 106518 18400 6 la_data_out_core[112]
port 274 nsew signal input
rlabel metal2 s 106922 17940 106978 18400 6 la_data_out_core[113]
port 275 nsew signal input
rlabel metal2 s 107382 17940 107438 18400 6 la_data_out_core[114]
port 276 nsew signal input
rlabel metal2 s 107750 17940 107806 18400 6 la_data_out_core[115]
port 277 nsew signal input
rlabel metal2 s 108210 17940 108266 18400 6 la_data_out_core[116]
port 278 nsew signal input
rlabel metal2 s 108670 17940 108726 18400 6 la_data_out_core[117]
port 279 nsew signal input
rlabel metal2 s 109130 17940 109186 18400 6 la_data_out_core[118]
port 280 nsew signal input
rlabel metal2 s 109498 17940 109554 18400 6 la_data_out_core[119]
port 281 nsew signal input
rlabel metal2 s 62486 17940 62542 18400 6 la_data_out_core[11]
port 282 nsew signal input
rlabel metal2 s 109958 17940 110014 18400 6 la_data_out_core[120]
port 283 nsew signal input
rlabel metal2 s 110418 17940 110474 18400 6 la_data_out_core[121]
port 284 nsew signal input
rlabel metal2 s 110878 17940 110934 18400 6 la_data_out_core[122]
port 285 nsew signal input
rlabel metal2 s 111246 17940 111302 18400 6 la_data_out_core[123]
port 286 nsew signal input
rlabel metal2 s 111706 17940 111762 18400 6 la_data_out_core[124]
port 287 nsew signal input
rlabel metal2 s 112166 17940 112222 18400 6 la_data_out_core[125]
port 288 nsew signal input
rlabel metal2 s 112534 17940 112590 18400 6 la_data_out_core[126]
port 289 nsew signal input
rlabel metal2 s 112994 17940 113050 18400 6 la_data_out_core[127]
port 290 nsew signal input
rlabel metal2 s 62946 17940 63002 18400 6 la_data_out_core[12]
port 291 nsew signal input
rlabel metal2 s 63314 17940 63370 18400 6 la_data_out_core[13]
port 292 nsew signal input
rlabel metal2 s 63774 17940 63830 18400 6 la_data_out_core[14]
port 293 nsew signal input
rlabel metal2 s 64234 17940 64290 18400 6 la_data_out_core[15]
port 294 nsew signal input
rlabel metal2 s 64602 17940 64658 18400 6 la_data_out_core[16]
port 295 nsew signal input
rlabel metal2 s 65062 17940 65118 18400 6 la_data_out_core[17]
port 296 nsew signal input
rlabel metal2 s 65522 17940 65578 18400 6 la_data_out_core[18]
port 297 nsew signal input
rlabel metal2 s 65982 17940 66038 18400 6 la_data_out_core[19]
port 298 nsew signal input
rlabel metal2 s 58070 17940 58126 18400 6 la_data_out_core[1]
port 299 nsew signal input
rlabel metal2 s 66350 17940 66406 18400 6 la_data_out_core[20]
port 300 nsew signal input
rlabel metal2 s 66810 17940 66866 18400 6 la_data_out_core[21]
port 301 nsew signal input
rlabel metal2 s 67270 17940 67326 18400 6 la_data_out_core[22]
port 302 nsew signal input
rlabel metal2 s 67730 17940 67786 18400 6 la_data_out_core[23]
port 303 nsew signal input
rlabel metal2 s 68098 17940 68154 18400 6 la_data_out_core[24]
port 304 nsew signal input
rlabel metal2 s 68558 17940 68614 18400 6 la_data_out_core[25]
port 305 nsew signal input
rlabel metal2 s 69018 17940 69074 18400 6 la_data_out_core[26]
port 306 nsew signal input
rlabel metal2 s 69478 17940 69534 18400 6 la_data_out_core[27]
port 307 nsew signal input
rlabel metal2 s 69846 17940 69902 18400 6 la_data_out_core[28]
port 308 nsew signal input
rlabel metal2 s 70306 17940 70362 18400 6 la_data_out_core[29]
port 309 nsew signal input
rlabel metal2 s 58530 17940 58586 18400 6 la_data_out_core[2]
port 310 nsew signal input
rlabel metal2 s 70766 17940 70822 18400 6 la_data_out_core[30]
port 311 nsew signal input
rlabel metal2 s 71226 17940 71282 18400 6 la_data_out_core[31]
port 312 nsew signal input
rlabel metal2 s 71594 17940 71650 18400 6 la_data_out_core[32]
port 313 nsew signal input
rlabel metal2 s 72054 17940 72110 18400 6 la_data_out_core[33]
port 314 nsew signal input
rlabel metal2 s 72514 17940 72570 18400 6 la_data_out_core[34]
port 315 nsew signal input
rlabel metal2 s 72882 17940 72938 18400 6 la_data_out_core[35]
port 316 nsew signal input
rlabel metal2 s 73342 17940 73398 18400 6 la_data_out_core[36]
port 317 nsew signal input
rlabel metal2 s 73802 17940 73858 18400 6 la_data_out_core[37]
port 318 nsew signal input
rlabel metal2 s 74262 17940 74318 18400 6 la_data_out_core[38]
port 319 nsew signal input
rlabel metal2 s 74630 17940 74686 18400 6 la_data_out_core[39]
port 320 nsew signal input
rlabel metal2 s 58990 17940 59046 18400 6 la_data_out_core[3]
port 321 nsew signal input
rlabel metal2 s 75090 17940 75146 18400 6 la_data_out_core[40]
port 322 nsew signal input
rlabel metal2 s 75550 17940 75606 18400 6 la_data_out_core[41]
port 323 nsew signal input
rlabel metal2 s 76010 17940 76066 18400 6 la_data_out_core[42]
port 324 nsew signal input
rlabel metal2 s 76378 17940 76434 18400 6 la_data_out_core[43]
port 325 nsew signal input
rlabel metal2 s 76838 17940 76894 18400 6 la_data_out_core[44]
port 326 nsew signal input
rlabel metal2 s 77298 17940 77354 18400 6 la_data_out_core[45]
port 327 nsew signal input
rlabel metal2 s 77758 17940 77814 18400 6 la_data_out_core[46]
port 328 nsew signal input
rlabel metal2 s 78126 17940 78182 18400 6 la_data_out_core[47]
port 329 nsew signal input
rlabel metal2 s 78586 17940 78642 18400 6 la_data_out_core[48]
port 330 nsew signal input
rlabel metal2 s 79046 17940 79102 18400 6 la_data_out_core[49]
port 331 nsew signal input
rlabel metal2 s 59450 17940 59506 18400 6 la_data_out_core[4]
port 332 nsew signal input
rlabel metal2 s 79506 17940 79562 18400 6 la_data_out_core[50]
port 333 nsew signal input
rlabel metal2 s 79874 17940 79930 18400 6 la_data_out_core[51]
port 334 nsew signal input
rlabel metal2 s 80334 17940 80390 18400 6 la_data_out_core[52]
port 335 nsew signal input
rlabel metal2 s 80794 17940 80850 18400 6 la_data_out_core[53]
port 336 nsew signal input
rlabel metal2 s 81162 17940 81218 18400 6 la_data_out_core[54]
port 337 nsew signal input
rlabel metal2 s 81622 17940 81678 18400 6 la_data_out_core[55]
port 338 nsew signal input
rlabel metal2 s 82082 17940 82138 18400 6 la_data_out_core[56]
port 339 nsew signal input
rlabel metal2 s 82542 17940 82598 18400 6 la_data_out_core[57]
port 340 nsew signal input
rlabel metal2 s 82910 17940 82966 18400 6 la_data_out_core[58]
port 341 nsew signal input
rlabel metal2 s 83370 17940 83426 18400 6 la_data_out_core[59]
port 342 nsew signal input
rlabel metal2 s 59818 17940 59874 18400 6 la_data_out_core[5]
port 343 nsew signal input
rlabel metal2 s 83830 17940 83886 18400 6 la_data_out_core[60]
port 344 nsew signal input
rlabel metal2 s 84290 17940 84346 18400 6 la_data_out_core[61]
port 345 nsew signal input
rlabel metal2 s 84658 17940 84714 18400 6 la_data_out_core[62]
port 346 nsew signal input
rlabel metal2 s 85118 17940 85174 18400 6 la_data_out_core[63]
port 347 nsew signal input
rlabel metal2 s 85578 17940 85634 18400 6 la_data_out_core[64]
port 348 nsew signal input
rlabel metal2 s 86038 17940 86094 18400 6 la_data_out_core[65]
port 349 nsew signal input
rlabel metal2 s 86406 17940 86462 18400 6 la_data_out_core[66]
port 350 nsew signal input
rlabel metal2 s 86866 17940 86922 18400 6 la_data_out_core[67]
port 351 nsew signal input
rlabel metal2 s 87326 17940 87382 18400 6 la_data_out_core[68]
port 352 nsew signal input
rlabel metal2 s 87786 17940 87842 18400 6 la_data_out_core[69]
port 353 nsew signal input
rlabel metal2 s 60278 17940 60334 18400 6 la_data_out_core[6]
port 354 nsew signal input
rlabel metal2 s 88154 17940 88210 18400 6 la_data_out_core[70]
port 355 nsew signal input
rlabel metal2 s 88614 17940 88670 18400 6 la_data_out_core[71]
port 356 nsew signal input
rlabel metal2 s 89074 17940 89130 18400 6 la_data_out_core[72]
port 357 nsew signal input
rlabel metal2 s 89442 17940 89498 18400 6 la_data_out_core[73]
port 358 nsew signal input
rlabel metal2 s 89902 17940 89958 18400 6 la_data_out_core[74]
port 359 nsew signal input
rlabel metal2 s 90362 17940 90418 18400 6 la_data_out_core[75]
port 360 nsew signal input
rlabel metal2 s 90822 17940 90878 18400 6 la_data_out_core[76]
port 361 nsew signal input
rlabel metal2 s 91190 17940 91246 18400 6 la_data_out_core[77]
port 362 nsew signal input
rlabel metal2 s 91650 17940 91706 18400 6 la_data_out_core[78]
port 363 nsew signal input
rlabel metal2 s 92110 17940 92166 18400 6 la_data_out_core[79]
port 364 nsew signal input
rlabel metal2 s 60738 17940 60794 18400 6 la_data_out_core[7]
port 365 nsew signal input
rlabel metal2 s 92570 17940 92626 18400 6 la_data_out_core[80]
port 366 nsew signal input
rlabel metal2 s 92938 17940 92994 18400 6 la_data_out_core[81]
port 367 nsew signal input
rlabel metal2 s 93398 17940 93454 18400 6 la_data_out_core[82]
port 368 nsew signal input
rlabel metal2 s 93858 17940 93914 18400 6 la_data_out_core[83]
port 369 nsew signal input
rlabel metal2 s 94318 17940 94374 18400 6 la_data_out_core[84]
port 370 nsew signal input
rlabel metal2 s 94686 17940 94742 18400 6 la_data_out_core[85]
port 371 nsew signal input
rlabel metal2 s 95146 17940 95202 18400 6 la_data_out_core[86]
port 372 nsew signal input
rlabel metal2 s 95606 17940 95662 18400 6 la_data_out_core[87]
port 373 nsew signal input
rlabel metal2 s 96066 17940 96122 18400 6 la_data_out_core[88]
port 374 nsew signal input
rlabel metal2 s 96434 17940 96490 18400 6 la_data_out_core[89]
port 375 nsew signal input
rlabel metal2 s 61198 17940 61254 18400 6 la_data_out_core[8]
port 376 nsew signal input
rlabel metal2 s 96894 17940 96950 18400 6 la_data_out_core[90]
port 377 nsew signal input
rlabel metal2 s 97354 17940 97410 18400 6 la_data_out_core[91]
port 378 nsew signal input
rlabel metal2 s 97722 17940 97778 18400 6 la_data_out_core[92]
port 379 nsew signal input
rlabel metal2 s 98182 17940 98238 18400 6 la_data_out_core[93]
port 380 nsew signal input
rlabel metal2 s 98642 17940 98698 18400 6 la_data_out_core[94]
port 381 nsew signal input
rlabel metal2 s 99102 17940 99158 18400 6 la_data_out_core[95]
port 382 nsew signal input
rlabel metal2 s 99470 17940 99526 18400 6 la_data_out_core[96]
port 383 nsew signal input
rlabel metal2 s 99930 17940 99986 18400 6 la_data_out_core[97]
port 384 nsew signal input
rlabel metal2 s 100390 17940 100446 18400 6 la_data_out_core[98]
port 385 nsew signal input
rlabel metal2 s 100850 17940 100906 18400 6 la_data_out_core[99]
port 386 nsew signal input
rlabel metal2 s 61566 17940 61622 18400 6 la_data_out_core[9]
port 387 nsew signal input
rlabel metal2 s 202 -400 258 60 8 la_data_out_mprj[0]
port 388 nsew signal input
rlabel metal2 s 43718 -400 43774 60 8 la_data_out_mprj[100]
port 389 nsew signal input
rlabel metal2 s 44178 -400 44234 60 8 la_data_out_mprj[101]
port 390 nsew signal input
rlabel metal2 s 44638 -400 44694 60 8 la_data_out_mprj[102]
port 391 nsew signal input
rlabel metal2 s 45006 -400 45062 60 8 la_data_out_mprj[103]
port 392 nsew signal input
rlabel metal2 s 45466 -400 45522 60 8 la_data_out_mprj[104]
port 393 nsew signal input
rlabel metal2 s 45926 -400 45982 60 8 la_data_out_mprj[105]
port 394 nsew signal input
rlabel metal2 s 46386 -400 46442 60 8 la_data_out_mprj[106]
port 395 nsew signal input
rlabel metal2 s 46754 -400 46810 60 8 la_data_out_mprj[107]
port 396 nsew signal input
rlabel metal2 s 47214 -400 47270 60 8 la_data_out_mprj[108]
port 397 nsew signal input
rlabel metal2 s 47674 -400 47730 60 8 la_data_out_mprj[109]
port 398 nsew signal input
rlabel metal2 s 4526 -400 4582 60 8 la_data_out_mprj[10]
port 399 nsew signal input
rlabel metal2 s 48134 -400 48190 60 8 la_data_out_mprj[110]
port 400 nsew signal input
rlabel metal2 s 48502 -400 48558 60 8 la_data_out_mprj[111]
port 401 nsew signal input
rlabel metal2 s 48962 -400 49018 60 8 la_data_out_mprj[112]
port 402 nsew signal input
rlabel metal2 s 49422 -400 49478 60 8 la_data_out_mprj[113]
port 403 nsew signal input
rlabel metal2 s 49790 -400 49846 60 8 la_data_out_mprj[114]
port 404 nsew signal input
rlabel metal2 s 50250 -400 50306 60 8 la_data_out_mprj[115]
port 405 nsew signal input
rlabel metal2 s 50710 -400 50766 60 8 la_data_out_mprj[116]
port 406 nsew signal input
rlabel metal2 s 51170 -400 51226 60 8 la_data_out_mprj[117]
port 407 nsew signal input
rlabel metal2 s 51538 -400 51594 60 8 la_data_out_mprj[118]
port 408 nsew signal input
rlabel metal2 s 51998 -400 52054 60 8 la_data_out_mprj[119]
port 409 nsew signal input
rlabel metal2 s 4986 -400 5042 60 8 la_data_out_mprj[11]
port 410 nsew signal input
rlabel metal2 s 52458 -400 52514 60 8 la_data_out_mprj[120]
port 411 nsew signal input
rlabel metal2 s 52918 -400 52974 60 8 la_data_out_mprj[121]
port 412 nsew signal input
rlabel metal2 s 53286 -400 53342 60 8 la_data_out_mprj[122]
port 413 nsew signal input
rlabel metal2 s 53746 -400 53802 60 8 la_data_out_mprj[123]
port 414 nsew signal input
rlabel metal2 s 54206 -400 54262 60 8 la_data_out_mprj[124]
port 415 nsew signal input
rlabel metal2 s 54666 -400 54722 60 8 la_data_out_mprj[125]
port 416 nsew signal input
rlabel metal2 s 55034 -400 55090 60 8 la_data_out_mprj[126]
port 417 nsew signal input
rlabel metal2 s 55494 -400 55550 60 8 la_data_out_mprj[127]
port 418 nsew signal input
rlabel metal2 s 5354 -400 5410 60 8 la_data_out_mprj[12]
port 419 nsew signal input
rlabel metal2 s 5814 -400 5870 60 8 la_data_out_mprj[13]
port 420 nsew signal input
rlabel metal2 s 6274 -400 6330 60 8 la_data_out_mprj[14]
port 421 nsew signal input
rlabel metal2 s 6734 -400 6790 60 8 la_data_out_mprj[15]
port 422 nsew signal input
rlabel metal2 s 7102 -400 7158 60 8 la_data_out_mprj[16]
port 423 nsew signal input
rlabel metal2 s 7562 -400 7618 60 8 la_data_out_mprj[17]
port 424 nsew signal input
rlabel metal2 s 8022 -400 8078 60 8 la_data_out_mprj[18]
port 425 nsew signal input
rlabel metal2 s 8390 -400 8446 60 8 la_data_out_mprj[19]
port 426 nsew signal input
rlabel metal2 s 570 -400 626 60 8 la_data_out_mprj[1]
port 427 nsew signal input
rlabel metal2 s 8850 -400 8906 60 8 la_data_out_mprj[20]
port 428 nsew signal input
rlabel metal2 s 9310 -400 9366 60 8 la_data_out_mprj[21]
port 429 nsew signal input
rlabel metal2 s 9770 -400 9826 60 8 la_data_out_mprj[22]
port 430 nsew signal input
rlabel metal2 s 10138 -400 10194 60 8 la_data_out_mprj[23]
port 431 nsew signal input
rlabel metal2 s 10598 -400 10654 60 8 la_data_out_mprj[24]
port 432 nsew signal input
rlabel metal2 s 11058 -400 11114 60 8 la_data_out_mprj[25]
port 433 nsew signal input
rlabel metal2 s 11518 -400 11574 60 8 la_data_out_mprj[26]
port 434 nsew signal input
rlabel metal2 s 11886 -400 11942 60 8 la_data_out_mprj[27]
port 435 nsew signal input
rlabel metal2 s 12346 -400 12402 60 8 la_data_out_mprj[28]
port 436 nsew signal input
rlabel metal2 s 12806 -400 12862 60 8 la_data_out_mprj[29]
port 437 nsew signal input
rlabel metal2 s 1030 -400 1086 60 8 la_data_out_mprj[2]
port 438 nsew signal input
rlabel metal2 s 13266 -400 13322 60 8 la_data_out_mprj[30]
port 439 nsew signal input
rlabel metal2 s 13634 -400 13690 60 8 la_data_out_mprj[31]
port 440 nsew signal input
rlabel metal2 s 14094 -400 14150 60 8 la_data_out_mprj[32]
port 441 nsew signal input
rlabel metal2 s 14554 -400 14610 60 8 la_data_out_mprj[33]
port 442 nsew signal input
rlabel metal2 s 15014 -400 15070 60 8 la_data_out_mprj[34]
port 443 nsew signal input
rlabel metal2 s 15382 -400 15438 60 8 la_data_out_mprj[35]
port 444 nsew signal input
rlabel metal2 s 15842 -400 15898 60 8 la_data_out_mprj[36]
port 445 nsew signal input
rlabel metal2 s 16302 -400 16358 60 8 la_data_out_mprj[37]
port 446 nsew signal input
rlabel metal2 s 16670 -400 16726 60 8 la_data_out_mprj[38]
port 447 nsew signal input
rlabel metal2 s 17130 -400 17186 60 8 la_data_out_mprj[39]
port 448 nsew signal input
rlabel metal2 s 1490 -400 1546 60 8 la_data_out_mprj[3]
port 449 nsew signal input
rlabel metal2 s 17590 -400 17646 60 8 la_data_out_mprj[40]
port 450 nsew signal input
rlabel metal2 s 18050 -400 18106 60 8 la_data_out_mprj[41]
port 451 nsew signal input
rlabel metal2 s 18418 -400 18474 60 8 la_data_out_mprj[42]
port 452 nsew signal input
rlabel metal2 s 18878 -400 18934 60 8 la_data_out_mprj[43]
port 453 nsew signal input
rlabel metal2 s 19338 -400 19394 60 8 la_data_out_mprj[44]
port 454 nsew signal input
rlabel metal2 s 19798 -400 19854 60 8 la_data_out_mprj[45]
port 455 nsew signal input
rlabel metal2 s 20166 -400 20222 60 8 la_data_out_mprj[46]
port 456 nsew signal input
rlabel metal2 s 20626 -400 20682 60 8 la_data_out_mprj[47]
port 457 nsew signal input
rlabel metal2 s 21086 -400 21142 60 8 la_data_out_mprj[48]
port 458 nsew signal input
rlabel metal2 s 21546 -400 21602 60 8 la_data_out_mprj[49]
port 459 nsew signal input
rlabel metal2 s 1858 -400 1914 60 8 la_data_out_mprj[4]
port 460 nsew signal input
rlabel metal2 s 21914 -400 21970 60 8 la_data_out_mprj[50]
port 461 nsew signal input
rlabel metal2 s 22374 -400 22430 60 8 la_data_out_mprj[51]
port 462 nsew signal input
rlabel metal2 s 22834 -400 22890 60 8 la_data_out_mprj[52]
port 463 nsew signal input
rlabel metal2 s 23294 -400 23350 60 8 la_data_out_mprj[53]
port 464 nsew signal input
rlabel metal2 s 23662 -400 23718 60 8 la_data_out_mprj[54]
port 465 nsew signal input
rlabel metal2 s 24122 -400 24178 60 8 la_data_out_mprj[55]
port 466 nsew signal input
rlabel metal2 s 24582 -400 24638 60 8 la_data_out_mprj[56]
port 467 nsew signal input
rlabel metal2 s 24950 -400 25006 60 8 la_data_out_mprj[57]
port 468 nsew signal input
rlabel metal2 s 25410 -400 25466 60 8 la_data_out_mprj[58]
port 469 nsew signal input
rlabel metal2 s 25870 -400 25926 60 8 la_data_out_mprj[59]
port 470 nsew signal input
rlabel metal2 s 2318 -400 2374 60 8 la_data_out_mprj[5]
port 471 nsew signal input
rlabel metal2 s 26330 -400 26386 60 8 la_data_out_mprj[60]
port 472 nsew signal input
rlabel metal2 s 26698 -400 26754 60 8 la_data_out_mprj[61]
port 473 nsew signal input
rlabel metal2 s 27158 -400 27214 60 8 la_data_out_mprj[62]
port 474 nsew signal input
rlabel metal2 s 27618 -400 27674 60 8 la_data_out_mprj[63]
port 475 nsew signal input
rlabel metal2 s 28078 -400 28134 60 8 la_data_out_mprj[64]
port 476 nsew signal input
rlabel metal2 s 28446 -400 28502 60 8 la_data_out_mprj[65]
port 477 nsew signal input
rlabel metal2 s 28906 -400 28962 60 8 la_data_out_mprj[66]
port 478 nsew signal input
rlabel metal2 s 29366 -400 29422 60 8 la_data_out_mprj[67]
port 479 nsew signal input
rlabel metal2 s 29826 -400 29882 60 8 la_data_out_mprj[68]
port 480 nsew signal input
rlabel metal2 s 30194 -400 30250 60 8 la_data_out_mprj[69]
port 481 nsew signal input
rlabel metal2 s 2778 -400 2834 60 8 la_data_out_mprj[6]
port 482 nsew signal input
rlabel metal2 s 30654 -400 30710 60 8 la_data_out_mprj[70]
port 483 nsew signal input
rlabel metal2 s 31114 -400 31170 60 8 la_data_out_mprj[71]
port 484 nsew signal input
rlabel metal2 s 31574 -400 31630 60 8 la_data_out_mprj[72]
port 485 nsew signal input
rlabel metal2 s 31942 -400 31998 60 8 la_data_out_mprj[73]
port 486 nsew signal input
rlabel metal2 s 32402 -400 32458 60 8 la_data_out_mprj[74]
port 487 nsew signal input
rlabel metal2 s 32862 -400 32918 60 8 la_data_out_mprj[75]
port 488 nsew signal input
rlabel metal2 s 33230 -400 33286 60 8 la_data_out_mprj[76]
port 489 nsew signal input
rlabel metal2 s 33690 -400 33746 60 8 la_data_out_mprj[77]
port 490 nsew signal input
rlabel metal2 s 34150 -400 34206 60 8 la_data_out_mprj[78]
port 491 nsew signal input
rlabel metal2 s 34610 -400 34666 60 8 la_data_out_mprj[79]
port 492 nsew signal input
rlabel metal2 s 3238 -400 3294 60 8 la_data_out_mprj[7]
port 493 nsew signal input
rlabel metal2 s 34978 -400 35034 60 8 la_data_out_mprj[80]
port 494 nsew signal input
rlabel metal2 s 35438 -400 35494 60 8 la_data_out_mprj[81]
port 495 nsew signal input
rlabel metal2 s 35898 -400 35954 60 8 la_data_out_mprj[82]
port 496 nsew signal input
rlabel metal2 s 36358 -400 36414 60 8 la_data_out_mprj[83]
port 497 nsew signal input
rlabel metal2 s 36726 -400 36782 60 8 la_data_out_mprj[84]
port 498 nsew signal input
rlabel metal2 s 37186 -400 37242 60 8 la_data_out_mprj[85]
port 499 nsew signal input
rlabel metal2 s 37646 -400 37702 60 8 la_data_out_mprj[86]
port 500 nsew signal input
rlabel metal2 s 38106 -400 38162 60 8 la_data_out_mprj[87]
port 501 nsew signal input
rlabel metal2 s 38474 -400 38530 60 8 la_data_out_mprj[88]
port 502 nsew signal input
rlabel metal2 s 38934 -400 38990 60 8 la_data_out_mprj[89]
port 503 nsew signal input
rlabel metal2 s 3606 -400 3662 60 8 la_data_out_mprj[8]
port 504 nsew signal input
rlabel metal2 s 39394 -400 39450 60 8 la_data_out_mprj[90]
port 505 nsew signal input
rlabel metal2 s 39854 -400 39910 60 8 la_data_out_mprj[91]
port 506 nsew signal input
rlabel metal2 s 40222 -400 40278 60 8 la_data_out_mprj[92]
port 507 nsew signal input
rlabel metal2 s 40682 -400 40738 60 8 la_data_out_mprj[93]
port 508 nsew signal input
rlabel metal2 s 41142 -400 41198 60 8 la_data_out_mprj[94]
port 509 nsew signal input
rlabel metal2 s 41510 -400 41566 60 8 la_data_out_mprj[95]
port 510 nsew signal input
rlabel metal2 s 41970 -400 42026 60 8 la_data_out_mprj[96]
port 511 nsew signal input
rlabel metal2 s 42430 -400 42486 60 8 la_data_out_mprj[97]
port 512 nsew signal input
rlabel metal2 s 42890 -400 42946 60 8 la_data_out_mprj[98]
port 513 nsew signal input
rlabel metal2 s 43258 -400 43314 60 8 la_data_out_mprj[99]
port 514 nsew signal input
rlabel metal2 s 4066 -400 4122 60 8 la_data_out_mprj[9]
port 515 nsew signal input
rlabel metal2 s 113454 17940 113510 18400 6 la_oen_core[0]
port 516 nsew signal output
rlabel metal2 s 157062 17940 157118 18400 6 la_oen_core[100]
port 517 nsew signal output
rlabel metal2 s 157430 17940 157486 18400 6 la_oen_core[101]
port 518 nsew signal output
rlabel metal2 s 157890 17940 157946 18400 6 la_oen_core[102]
port 519 nsew signal output
rlabel metal2 s 158350 17940 158406 18400 6 la_oen_core[103]
port 520 nsew signal output
rlabel metal2 s 158810 17940 158866 18400 6 la_oen_core[104]
port 521 nsew signal output
rlabel metal2 s 159178 17940 159234 18400 6 la_oen_core[105]
port 522 nsew signal output
rlabel metal2 s 159638 17940 159694 18400 6 la_oen_core[106]
port 523 nsew signal output
rlabel metal2 s 160098 17940 160154 18400 6 la_oen_core[107]
port 524 nsew signal output
rlabel metal2 s 160466 17940 160522 18400 6 la_oen_core[108]
port 525 nsew signal output
rlabel metal2 s 160926 17940 160982 18400 6 la_oen_core[109]
port 526 nsew signal output
rlabel metal2 s 117778 17940 117834 18400 6 la_oen_core[10]
port 527 nsew signal output
rlabel metal2 s 161386 17940 161442 18400 6 la_oen_core[110]
port 528 nsew signal output
rlabel metal2 s 161846 17940 161902 18400 6 la_oen_core[111]
port 529 nsew signal output
rlabel metal2 s 162214 17940 162270 18400 6 la_oen_core[112]
port 530 nsew signal output
rlabel metal2 s 162674 17940 162730 18400 6 la_oen_core[113]
port 531 nsew signal output
rlabel metal2 s 163134 17940 163190 18400 6 la_oen_core[114]
port 532 nsew signal output
rlabel metal2 s 163594 17940 163650 18400 6 la_oen_core[115]
port 533 nsew signal output
rlabel metal2 s 163962 17940 164018 18400 6 la_oen_core[116]
port 534 nsew signal output
rlabel metal2 s 164422 17940 164478 18400 6 la_oen_core[117]
port 535 nsew signal output
rlabel metal2 s 164882 17940 164938 18400 6 la_oen_core[118]
port 536 nsew signal output
rlabel metal2 s 165342 17940 165398 18400 6 la_oen_core[119]
port 537 nsew signal output
rlabel metal2 s 118238 17940 118294 18400 6 la_oen_core[11]
port 538 nsew signal output
rlabel metal2 s 165710 17940 165766 18400 6 la_oen_core[120]
port 539 nsew signal output
rlabel metal2 s 166170 17940 166226 18400 6 la_oen_core[121]
port 540 nsew signal output
rlabel metal2 s 166630 17940 166686 18400 6 la_oen_core[122]
port 541 nsew signal output
rlabel metal2 s 167090 17940 167146 18400 6 la_oen_core[123]
port 542 nsew signal output
rlabel metal2 s 167458 17940 167514 18400 6 la_oen_core[124]
port 543 nsew signal output
rlabel metal2 s 167918 17940 167974 18400 6 la_oen_core[125]
port 544 nsew signal output
rlabel metal2 s 168378 17940 168434 18400 6 la_oen_core[126]
port 545 nsew signal output
rlabel metal2 s 168746 17940 168802 18400 6 la_oen_core[127]
port 546 nsew signal output
rlabel metal2 s 118698 17940 118754 18400 6 la_oen_core[12]
port 547 nsew signal output
rlabel metal2 s 119158 17940 119214 18400 6 la_oen_core[13]
port 548 nsew signal output
rlabel metal2 s 119526 17940 119582 18400 6 la_oen_core[14]
port 549 nsew signal output
rlabel metal2 s 119986 17940 120042 18400 6 la_oen_core[15]
port 550 nsew signal output
rlabel metal2 s 120446 17940 120502 18400 6 la_oen_core[16]
port 551 nsew signal output
rlabel metal2 s 120814 17940 120870 18400 6 la_oen_core[17]
port 552 nsew signal output
rlabel metal2 s 121274 17940 121330 18400 6 la_oen_core[18]
port 553 nsew signal output
rlabel metal2 s 121734 17940 121790 18400 6 la_oen_core[19]
port 554 nsew signal output
rlabel metal2 s 113914 17940 113970 18400 6 la_oen_core[1]
port 555 nsew signal output
rlabel metal2 s 122194 17940 122250 18400 6 la_oen_core[20]
port 556 nsew signal output
rlabel metal2 s 122562 17940 122618 18400 6 la_oen_core[21]
port 557 nsew signal output
rlabel metal2 s 123022 17940 123078 18400 6 la_oen_core[22]
port 558 nsew signal output
rlabel metal2 s 123482 17940 123538 18400 6 la_oen_core[23]
port 559 nsew signal output
rlabel metal2 s 123942 17940 123998 18400 6 la_oen_core[24]
port 560 nsew signal output
rlabel metal2 s 124310 17940 124366 18400 6 la_oen_core[25]
port 561 nsew signal output
rlabel metal2 s 124770 17940 124826 18400 6 la_oen_core[26]
port 562 nsew signal output
rlabel metal2 s 125230 17940 125286 18400 6 la_oen_core[27]
port 563 nsew signal output
rlabel metal2 s 125690 17940 125746 18400 6 la_oen_core[28]
port 564 nsew signal output
rlabel metal2 s 126058 17940 126114 18400 6 la_oen_core[29]
port 565 nsew signal output
rlabel metal2 s 114282 17940 114338 18400 6 la_oen_core[2]
port 566 nsew signal output
rlabel metal2 s 126518 17940 126574 18400 6 la_oen_core[30]
port 567 nsew signal output
rlabel metal2 s 126978 17940 127034 18400 6 la_oen_core[31]
port 568 nsew signal output
rlabel metal2 s 127438 17940 127494 18400 6 la_oen_core[32]
port 569 nsew signal output
rlabel metal2 s 127806 17940 127862 18400 6 la_oen_core[33]
port 570 nsew signal output
rlabel metal2 s 128266 17940 128322 18400 6 la_oen_core[34]
port 571 nsew signal output
rlabel metal2 s 128726 17940 128782 18400 6 la_oen_core[35]
port 572 nsew signal output
rlabel metal2 s 129094 17940 129150 18400 6 la_oen_core[36]
port 573 nsew signal output
rlabel metal2 s 129554 17940 129610 18400 6 la_oen_core[37]
port 574 nsew signal output
rlabel metal2 s 130014 17940 130070 18400 6 la_oen_core[38]
port 575 nsew signal output
rlabel metal2 s 130474 17940 130530 18400 6 la_oen_core[39]
port 576 nsew signal output
rlabel metal2 s 114742 17940 114798 18400 6 la_oen_core[3]
port 577 nsew signal output
rlabel metal2 s 130842 17940 130898 18400 6 la_oen_core[40]
port 578 nsew signal output
rlabel metal2 s 131302 17940 131358 18400 6 la_oen_core[41]
port 579 nsew signal output
rlabel metal2 s 131762 17940 131818 18400 6 la_oen_core[42]
port 580 nsew signal output
rlabel metal2 s 132222 17940 132278 18400 6 la_oen_core[43]
port 581 nsew signal output
rlabel metal2 s 132590 17940 132646 18400 6 la_oen_core[44]
port 582 nsew signal output
rlabel metal2 s 133050 17940 133106 18400 6 la_oen_core[45]
port 583 nsew signal output
rlabel metal2 s 133510 17940 133566 18400 6 la_oen_core[46]
port 584 nsew signal output
rlabel metal2 s 133970 17940 134026 18400 6 la_oen_core[47]
port 585 nsew signal output
rlabel metal2 s 134338 17940 134394 18400 6 la_oen_core[48]
port 586 nsew signal output
rlabel metal2 s 134798 17940 134854 18400 6 la_oen_core[49]
port 587 nsew signal output
rlabel metal2 s 115202 17940 115258 18400 6 la_oen_core[4]
port 588 nsew signal output
rlabel metal2 s 135258 17940 135314 18400 6 la_oen_core[50]
port 589 nsew signal output
rlabel metal2 s 135718 17940 135774 18400 6 la_oen_core[51]
port 590 nsew signal output
rlabel metal2 s 136086 17940 136142 18400 6 la_oen_core[52]
port 591 nsew signal output
rlabel metal2 s 136546 17940 136602 18400 6 la_oen_core[53]
port 592 nsew signal output
rlabel metal2 s 137006 17940 137062 18400 6 la_oen_core[54]
port 593 nsew signal output
rlabel metal2 s 137374 17940 137430 18400 6 la_oen_core[55]
port 594 nsew signal output
rlabel metal2 s 137834 17940 137890 18400 6 la_oen_core[56]
port 595 nsew signal output
rlabel metal2 s 138294 17940 138350 18400 6 la_oen_core[57]
port 596 nsew signal output
rlabel metal2 s 138754 17940 138810 18400 6 la_oen_core[58]
port 597 nsew signal output
rlabel metal2 s 139122 17940 139178 18400 6 la_oen_core[59]
port 598 nsew signal output
rlabel metal2 s 115662 17940 115718 18400 6 la_oen_core[5]
port 599 nsew signal output
rlabel metal2 s 139582 17940 139638 18400 6 la_oen_core[60]
port 600 nsew signal output
rlabel metal2 s 140042 17940 140098 18400 6 la_oen_core[61]
port 601 nsew signal output
rlabel metal2 s 140502 17940 140558 18400 6 la_oen_core[62]
port 602 nsew signal output
rlabel metal2 s 140870 17940 140926 18400 6 la_oen_core[63]
port 603 nsew signal output
rlabel metal2 s 141330 17940 141386 18400 6 la_oen_core[64]
port 604 nsew signal output
rlabel metal2 s 141790 17940 141846 18400 6 la_oen_core[65]
port 605 nsew signal output
rlabel metal2 s 142250 17940 142306 18400 6 la_oen_core[66]
port 606 nsew signal output
rlabel metal2 s 142618 17940 142674 18400 6 la_oen_core[67]
port 607 nsew signal output
rlabel metal2 s 143078 17940 143134 18400 6 la_oen_core[68]
port 608 nsew signal output
rlabel metal2 s 143538 17940 143594 18400 6 la_oen_core[69]
port 609 nsew signal output
rlabel metal2 s 116030 17940 116086 18400 6 la_oen_core[6]
port 610 nsew signal output
rlabel metal2 s 143998 17940 144054 18400 6 la_oen_core[70]
port 611 nsew signal output
rlabel metal2 s 144366 17940 144422 18400 6 la_oen_core[71]
port 612 nsew signal output
rlabel metal2 s 144826 17940 144882 18400 6 la_oen_core[72]
port 613 nsew signal output
rlabel metal2 s 145286 17940 145342 18400 6 la_oen_core[73]
port 614 nsew signal output
rlabel metal2 s 145654 17940 145710 18400 6 la_oen_core[74]
port 615 nsew signal output
rlabel metal2 s 146114 17940 146170 18400 6 la_oen_core[75]
port 616 nsew signal output
rlabel metal2 s 146574 17940 146630 18400 6 la_oen_core[76]
port 617 nsew signal output
rlabel metal2 s 147034 17940 147090 18400 6 la_oen_core[77]
port 618 nsew signal output
rlabel metal2 s 147402 17940 147458 18400 6 la_oen_core[78]
port 619 nsew signal output
rlabel metal2 s 147862 17940 147918 18400 6 la_oen_core[79]
port 620 nsew signal output
rlabel metal2 s 116490 17940 116546 18400 6 la_oen_core[7]
port 621 nsew signal output
rlabel metal2 s 148322 17940 148378 18400 6 la_oen_core[80]
port 622 nsew signal output
rlabel metal2 s 148782 17940 148838 18400 6 la_oen_core[81]
port 623 nsew signal output
rlabel metal2 s 149150 17940 149206 18400 6 la_oen_core[82]
port 624 nsew signal output
rlabel metal2 s 149610 17940 149666 18400 6 la_oen_core[83]
port 625 nsew signal output
rlabel metal2 s 150070 17940 150126 18400 6 la_oen_core[84]
port 626 nsew signal output
rlabel metal2 s 150530 17940 150586 18400 6 la_oen_core[85]
port 627 nsew signal output
rlabel metal2 s 150898 17940 150954 18400 6 la_oen_core[86]
port 628 nsew signal output
rlabel metal2 s 151358 17940 151414 18400 6 la_oen_core[87]
port 629 nsew signal output
rlabel metal2 s 151818 17940 151874 18400 6 la_oen_core[88]
port 630 nsew signal output
rlabel metal2 s 152186 17940 152242 18400 6 la_oen_core[89]
port 631 nsew signal output
rlabel metal2 s 116950 17940 117006 18400 6 la_oen_core[8]
port 632 nsew signal output
rlabel metal2 s 152646 17940 152702 18400 6 la_oen_core[90]
port 633 nsew signal output
rlabel metal2 s 153106 17940 153162 18400 6 la_oen_core[91]
port 634 nsew signal output
rlabel metal2 s 153566 17940 153622 18400 6 la_oen_core[92]
port 635 nsew signal output
rlabel metal2 s 153934 17940 153990 18400 6 la_oen_core[93]
port 636 nsew signal output
rlabel metal2 s 154394 17940 154450 18400 6 la_oen_core[94]
port 637 nsew signal output
rlabel metal2 s 154854 17940 154910 18400 6 la_oen_core[95]
port 638 nsew signal output
rlabel metal2 s 155314 17940 155370 18400 6 la_oen_core[96]
port 639 nsew signal output
rlabel metal2 s 155682 17940 155738 18400 6 la_oen_core[97]
port 640 nsew signal output
rlabel metal2 s 156142 17940 156198 18400 6 la_oen_core[98]
port 641 nsew signal output
rlabel metal2 s 156602 17940 156658 18400 6 la_oen_core[99]
port 642 nsew signal output
rlabel metal2 s 117410 17940 117466 18400 6 la_oen_core[9]
port 643 nsew signal output
rlabel metal2 s 111706 -400 111762 60 8 la_oen_mprj[0]
port 644 nsew signal input
rlabel metal2 s 155314 -400 155370 60 8 la_oen_mprj[100]
port 645 nsew signal input
rlabel metal2 s 155682 -400 155738 60 8 la_oen_mprj[101]
port 646 nsew signal input
rlabel metal2 s 156142 -400 156198 60 8 la_oen_mprj[102]
port 647 nsew signal input
rlabel metal2 s 156602 -400 156658 60 8 la_oen_mprj[103]
port 648 nsew signal input
rlabel metal2 s 157062 -400 157118 60 8 la_oen_mprj[104]
port 649 nsew signal input
rlabel metal2 s 157430 -400 157486 60 8 la_oen_mprj[105]
port 650 nsew signal input
rlabel metal2 s 157890 -400 157946 60 8 la_oen_mprj[106]
port 651 nsew signal input
rlabel metal2 s 158350 -400 158406 60 8 la_oen_mprj[107]
port 652 nsew signal input
rlabel metal2 s 158810 -400 158866 60 8 la_oen_mprj[108]
port 653 nsew signal input
rlabel metal2 s 159178 -400 159234 60 8 la_oen_mprj[109]
port 654 nsew signal input
rlabel metal2 s 116030 -400 116086 60 8 la_oen_mprj[10]
port 655 nsew signal input
rlabel metal2 s 159638 -400 159694 60 8 la_oen_mprj[110]
port 656 nsew signal input
rlabel metal2 s 160098 -400 160154 60 8 la_oen_mprj[111]
port 657 nsew signal input
rlabel metal2 s 160466 -400 160522 60 8 la_oen_mprj[112]
port 658 nsew signal input
rlabel metal2 s 160926 -400 160982 60 8 la_oen_mprj[113]
port 659 nsew signal input
rlabel metal2 s 161386 -400 161442 60 8 la_oen_mprj[114]
port 660 nsew signal input
rlabel metal2 s 161846 -400 161902 60 8 la_oen_mprj[115]
port 661 nsew signal input
rlabel metal2 s 162214 -400 162270 60 8 la_oen_mprj[116]
port 662 nsew signal input
rlabel metal2 s 162674 -400 162730 60 8 la_oen_mprj[117]
port 663 nsew signal input
rlabel metal2 s 163134 -400 163190 60 8 la_oen_mprj[118]
port 664 nsew signal input
rlabel metal2 s 163594 -400 163650 60 8 la_oen_mprj[119]
port 665 nsew signal input
rlabel metal2 s 116490 -400 116546 60 8 la_oen_mprj[11]
port 666 nsew signal input
rlabel metal2 s 163962 -400 164018 60 8 la_oen_mprj[120]
port 667 nsew signal input
rlabel metal2 s 164422 -400 164478 60 8 la_oen_mprj[121]
port 668 nsew signal input
rlabel metal2 s 164882 -400 164938 60 8 la_oen_mprj[122]
port 669 nsew signal input
rlabel metal2 s 165342 -400 165398 60 8 la_oen_mprj[123]
port 670 nsew signal input
rlabel metal2 s 165710 -400 165766 60 8 la_oen_mprj[124]
port 671 nsew signal input
rlabel metal2 s 166170 -400 166226 60 8 la_oen_mprj[125]
port 672 nsew signal input
rlabel metal2 s 166630 -400 166686 60 8 la_oen_mprj[126]
port 673 nsew signal input
rlabel metal2 s 167090 -400 167146 60 8 la_oen_mprj[127]
port 674 nsew signal input
rlabel metal2 s 116950 -400 117006 60 8 la_oen_mprj[12]
port 675 nsew signal input
rlabel metal2 s 117410 -400 117466 60 8 la_oen_mprj[13]
port 676 nsew signal input
rlabel metal2 s 117778 -400 117834 60 8 la_oen_mprj[14]
port 677 nsew signal input
rlabel metal2 s 118238 -400 118294 60 8 la_oen_mprj[15]
port 678 nsew signal input
rlabel metal2 s 118698 -400 118754 60 8 la_oen_mprj[16]
port 679 nsew signal input
rlabel metal2 s 119158 -400 119214 60 8 la_oen_mprj[17]
port 680 nsew signal input
rlabel metal2 s 119526 -400 119582 60 8 la_oen_mprj[18]
port 681 nsew signal input
rlabel metal2 s 119986 -400 120042 60 8 la_oen_mprj[19]
port 682 nsew signal input
rlabel metal2 s 112166 -400 112222 60 8 la_oen_mprj[1]
port 683 nsew signal input
rlabel metal2 s 120446 -400 120502 60 8 la_oen_mprj[20]
port 684 nsew signal input
rlabel metal2 s 120814 -400 120870 60 8 la_oen_mprj[21]
port 685 nsew signal input
rlabel metal2 s 121274 -400 121330 60 8 la_oen_mprj[22]
port 686 nsew signal input
rlabel metal2 s 121734 -400 121790 60 8 la_oen_mprj[23]
port 687 nsew signal input
rlabel metal2 s 122194 -400 122250 60 8 la_oen_mprj[24]
port 688 nsew signal input
rlabel metal2 s 122562 -400 122618 60 8 la_oen_mprj[25]
port 689 nsew signal input
rlabel metal2 s 123022 -400 123078 60 8 la_oen_mprj[26]
port 690 nsew signal input
rlabel metal2 s 123482 -400 123538 60 8 la_oen_mprj[27]
port 691 nsew signal input
rlabel metal2 s 123942 -400 123998 60 8 la_oen_mprj[28]
port 692 nsew signal input
rlabel metal2 s 124310 -400 124366 60 8 la_oen_mprj[29]
port 693 nsew signal input
rlabel metal2 s 112534 -400 112590 60 8 la_oen_mprj[2]
port 694 nsew signal input
rlabel metal2 s 124770 -400 124826 60 8 la_oen_mprj[30]
port 695 nsew signal input
rlabel metal2 s 125230 -400 125286 60 8 la_oen_mprj[31]
port 696 nsew signal input
rlabel metal2 s 125690 -400 125746 60 8 la_oen_mprj[32]
port 697 nsew signal input
rlabel metal2 s 126058 -400 126114 60 8 la_oen_mprj[33]
port 698 nsew signal input
rlabel metal2 s 126518 -400 126574 60 8 la_oen_mprj[34]
port 699 nsew signal input
rlabel metal2 s 126978 -400 127034 60 8 la_oen_mprj[35]
port 700 nsew signal input
rlabel metal2 s 127438 -400 127494 60 8 la_oen_mprj[36]
port 701 nsew signal input
rlabel metal2 s 127806 -400 127862 60 8 la_oen_mprj[37]
port 702 nsew signal input
rlabel metal2 s 128266 -400 128322 60 8 la_oen_mprj[38]
port 703 nsew signal input
rlabel metal2 s 128726 -400 128782 60 8 la_oen_mprj[39]
port 704 nsew signal input
rlabel metal2 s 112994 -400 113050 60 8 la_oen_mprj[3]
port 705 nsew signal input
rlabel metal2 s 129094 -400 129150 60 8 la_oen_mprj[40]
port 706 nsew signal input
rlabel metal2 s 129554 -400 129610 60 8 la_oen_mprj[41]
port 707 nsew signal input
rlabel metal2 s 130014 -400 130070 60 8 la_oen_mprj[42]
port 708 nsew signal input
rlabel metal2 s 130474 -400 130530 60 8 la_oen_mprj[43]
port 709 nsew signal input
rlabel metal2 s 130842 -400 130898 60 8 la_oen_mprj[44]
port 710 nsew signal input
rlabel metal2 s 131302 -400 131358 60 8 la_oen_mprj[45]
port 711 nsew signal input
rlabel metal2 s 131762 -400 131818 60 8 la_oen_mprj[46]
port 712 nsew signal input
rlabel metal2 s 132222 -400 132278 60 8 la_oen_mprj[47]
port 713 nsew signal input
rlabel metal2 s 132590 -400 132646 60 8 la_oen_mprj[48]
port 714 nsew signal input
rlabel metal2 s 133050 -400 133106 60 8 la_oen_mprj[49]
port 715 nsew signal input
rlabel metal2 s 113454 -400 113510 60 8 la_oen_mprj[4]
port 716 nsew signal input
rlabel metal2 s 133510 -400 133566 60 8 la_oen_mprj[50]
port 717 nsew signal input
rlabel metal2 s 133970 -400 134026 60 8 la_oen_mprj[51]
port 718 nsew signal input
rlabel metal2 s 134338 -400 134394 60 8 la_oen_mprj[52]
port 719 nsew signal input
rlabel metal2 s 134798 -400 134854 60 8 la_oen_mprj[53]
port 720 nsew signal input
rlabel metal2 s 135258 -400 135314 60 8 la_oen_mprj[54]
port 721 nsew signal input
rlabel metal2 s 135718 -400 135774 60 8 la_oen_mprj[55]
port 722 nsew signal input
rlabel metal2 s 136086 -400 136142 60 8 la_oen_mprj[56]
port 723 nsew signal input
rlabel metal2 s 136546 -400 136602 60 8 la_oen_mprj[57]
port 724 nsew signal input
rlabel metal2 s 137006 -400 137062 60 8 la_oen_mprj[58]
port 725 nsew signal input
rlabel metal2 s 137374 -400 137430 60 8 la_oen_mprj[59]
port 726 nsew signal input
rlabel metal2 s 113914 -400 113970 60 8 la_oen_mprj[5]
port 727 nsew signal input
rlabel metal2 s 137834 -400 137890 60 8 la_oen_mprj[60]
port 728 nsew signal input
rlabel metal2 s 138294 -400 138350 60 8 la_oen_mprj[61]
port 729 nsew signal input
rlabel metal2 s 138754 -400 138810 60 8 la_oen_mprj[62]
port 730 nsew signal input
rlabel metal2 s 139122 -400 139178 60 8 la_oen_mprj[63]
port 731 nsew signal input
rlabel metal2 s 139582 -400 139638 60 8 la_oen_mprj[64]
port 732 nsew signal input
rlabel metal2 s 140042 -400 140098 60 8 la_oen_mprj[65]
port 733 nsew signal input
rlabel metal2 s 140502 -400 140558 60 8 la_oen_mprj[66]
port 734 nsew signal input
rlabel metal2 s 140870 -400 140926 60 8 la_oen_mprj[67]
port 735 nsew signal input
rlabel metal2 s 141330 -400 141386 60 8 la_oen_mprj[68]
port 736 nsew signal input
rlabel metal2 s 141790 -400 141846 60 8 la_oen_mprj[69]
port 737 nsew signal input
rlabel metal2 s 114282 -400 114338 60 8 la_oen_mprj[6]
port 738 nsew signal input
rlabel metal2 s 142250 -400 142306 60 8 la_oen_mprj[70]
port 739 nsew signal input
rlabel metal2 s 142618 -400 142674 60 8 la_oen_mprj[71]
port 740 nsew signal input
rlabel metal2 s 143078 -400 143134 60 8 la_oen_mprj[72]
port 741 nsew signal input
rlabel metal2 s 143538 -400 143594 60 8 la_oen_mprj[73]
port 742 nsew signal input
rlabel metal2 s 143998 -400 144054 60 8 la_oen_mprj[74]
port 743 nsew signal input
rlabel metal2 s 144366 -400 144422 60 8 la_oen_mprj[75]
port 744 nsew signal input
rlabel metal2 s 144826 -400 144882 60 8 la_oen_mprj[76]
port 745 nsew signal input
rlabel metal2 s 145286 -400 145342 60 8 la_oen_mprj[77]
port 746 nsew signal input
rlabel metal2 s 145654 -400 145710 60 8 la_oen_mprj[78]
port 747 nsew signal input
rlabel metal2 s 146114 -400 146170 60 8 la_oen_mprj[79]
port 748 nsew signal input
rlabel metal2 s 114742 -400 114798 60 8 la_oen_mprj[7]
port 749 nsew signal input
rlabel metal2 s 146574 -400 146630 60 8 la_oen_mprj[80]
port 750 nsew signal input
rlabel metal2 s 147034 -400 147090 60 8 la_oen_mprj[81]
port 751 nsew signal input
rlabel metal2 s 147402 -400 147458 60 8 la_oen_mprj[82]
port 752 nsew signal input
rlabel metal2 s 147862 -400 147918 60 8 la_oen_mprj[83]
port 753 nsew signal input
rlabel metal2 s 148322 -400 148378 60 8 la_oen_mprj[84]
port 754 nsew signal input
rlabel metal2 s 148782 -400 148838 60 8 la_oen_mprj[85]
port 755 nsew signal input
rlabel metal2 s 149150 -400 149206 60 8 la_oen_mprj[86]
port 756 nsew signal input
rlabel metal2 s 149610 -400 149666 60 8 la_oen_mprj[87]
port 757 nsew signal input
rlabel metal2 s 150070 -400 150126 60 8 la_oen_mprj[88]
port 758 nsew signal input
rlabel metal2 s 150530 -400 150586 60 8 la_oen_mprj[89]
port 759 nsew signal input
rlabel metal2 s 115202 -400 115258 60 8 la_oen_mprj[8]
port 760 nsew signal input
rlabel metal2 s 150898 -400 150954 60 8 la_oen_mprj[90]
port 761 nsew signal input
rlabel metal2 s 151358 -400 151414 60 8 la_oen_mprj[91]
port 762 nsew signal input
rlabel metal2 s 151818 -400 151874 60 8 la_oen_mprj[92]
port 763 nsew signal input
rlabel metal2 s 152186 -400 152242 60 8 la_oen_mprj[93]
port 764 nsew signal input
rlabel metal2 s 152646 -400 152702 60 8 la_oen_mprj[94]
port 765 nsew signal input
rlabel metal2 s 153106 -400 153162 60 8 la_oen_mprj[95]
port 766 nsew signal input
rlabel metal2 s 153566 -400 153622 60 8 la_oen_mprj[96]
port 767 nsew signal input
rlabel metal2 s 153934 -400 153990 60 8 la_oen_mprj[97]
port 768 nsew signal input
rlabel metal2 s 154394 -400 154450 60 8 la_oen_mprj[98]
port 769 nsew signal input
rlabel metal2 s 154854 -400 154910 60 8 la_oen_mprj[99]
port 770 nsew signal input
rlabel metal2 s 115662 -400 115718 60 8 la_oen_mprj[9]
port 771 nsew signal input
rlabel metal2 s 168746 -400 168802 60 8 mprj_adr_o_core[0]
port 772 nsew signal input
rlabel metal2 s 179234 -400 179290 60 8 mprj_adr_o_core[10]
port 773 nsew signal input
rlabel metal2 s 180154 -400 180210 60 8 mprj_adr_o_core[11]
port 774 nsew signal input
rlabel metal2 s 180982 -400 181038 60 8 mprj_adr_o_core[12]
port 775 nsew signal input
rlabel metal2 s 181902 -400 181958 60 8 mprj_adr_o_core[13]
port 776 nsew signal input
rlabel metal2 s 182730 -400 182786 60 8 mprj_adr_o_core[14]
port 777 nsew signal input
rlabel metal2 s 183650 -400 183706 60 8 mprj_adr_o_core[15]
port 778 nsew signal input
rlabel metal2 s 184478 -400 184534 60 8 mprj_adr_o_core[16]
port 779 nsew signal input
rlabel metal2 s 185306 -400 185362 60 8 mprj_adr_o_core[17]
port 780 nsew signal input
rlabel metal2 s 186226 -400 186282 60 8 mprj_adr_o_core[18]
port 781 nsew signal input
rlabel metal2 s 187054 -400 187110 60 8 mprj_adr_o_core[19]
port 782 nsew signal input
rlabel metal2 s 170126 -400 170182 60 8 mprj_adr_o_core[1]
port 783 nsew signal input
rlabel metal2 s 187974 -400 188030 60 8 mprj_adr_o_core[20]
port 784 nsew signal input
rlabel metal2 s 188802 -400 188858 60 8 mprj_adr_o_core[21]
port 785 nsew signal input
rlabel metal2 s 189722 -400 189778 60 8 mprj_adr_o_core[22]
port 786 nsew signal input
rlabel metal2 s 190550 -400 190606 60 8 mprj_adr_o_core[23]
port 787 nsew signal input
rlabel metal2 s 191470 -400 191526 60 8 mprj_adr_o_core[24]
port 788 nsew signal input
rlabel metal2 s 192298 -400 192354 60 8 mprj_adr_o_core[25]
port 789 nsew signal input
rlabel metal2 s 193218 -400 193274 60 8 mprj_adr_o_core[26]
port 790 nsew signal input
rlabel metal2 s 194046 -400 194102 60 8 mprj_adr_o_core[27]
port 791 nsew signal input
rlabel metal2 s 194966 -400 195022 60 8 mprj_adr_o_core[28]
port 792 nsew signal input
rlabel metal2 s 195794 -400 195850 60 8 mprj_adr_o_core[29]
port 793 nsew signal input
rlabel metal2 s 171414 -400 171470 60 8 mprj_adr_o_core[2]
port 794 nsew signal input
rlabel metal2 s 196714 -400 196770 60 8 mprj_adr_o_core[30]
port 795 nsew signal input
rlabel metal2 s 197542 -400 197598 60 8 mprj_adr_o_core[31]
port 796 nsew signal input
rlabel metal2 s 172702 -400 172758 60 8 mprj_adr_o_core[3]
port 797 nsew signal input
rlabel metal2 s 173990 -400 174046 60 8 mprj_adr_o_core[4]
port 798 nsew signal input
rlabel metal2 s 174910 -400 174966 60 8 mprj_adr_o_core[5]
port 799 nsew signal input
rlabel metal2 s 175738 -400 175794 60 8 mprj_adr_o_core[6]
port 800 nsew signal input
rlabel metal2 s 176658 -400 176714 60 8 mprj_adr_o_core[7]
port 801 nsew signal input
rlabel metal2 s 177486 -400 177542 60 8 mprj_adr_o_core[8]
port 802 nsew signal input
rlabel metal2 s 178406 -400 178462 60 8 mprj_adr_o_core[9]
port 803 nsew signal input
rlabel metal2 s 170494 17940 170550 18400 6 mprj_adr_o_user[0]
port 804 nsew signal output
rlabel metal2 s 180982 17940 181038 18400 6 mprj_adr_o_user[10]
port 805 nsew signal output
rlabel metal2 s 181902 17940 181958 18400 6 mprj_adr_o_user[11]
port 806 nsew signal output
rlabel metal2 s 182730 17940 182786 18400 6 mprj_adr_o_user[12]
port 807 nsew signal output
rlabel metal2 s 183650 17940 183706 18400 6 mprj_adr_o_user[13]
port 808 nsew signal output
rlabel metal2 s 184478 17940 184534 18400 6 mprj_adr_o_user[14]
port 809 nsew signal output
rlabel metal2 s 185306 17940 185362 18400 6 mprj_adr_o_user[15]
port 810 nsew signal output
rlabel metal2 s 186226 17940 186282 18400 6 mprj_adr_o_user[16]
port 811 nsew signal output
rlabel metal2 s 187054 17940 187110 18400 6 mprj_adr_o_user[17]
port 812 nsew signal output
rlabel metal2 s 187974 17940 188030 18400 6 mprj_adr_o_user[18]
port 813 nsew signal output
rlabel metal2 s 188802 17940 188858 18400 6 mprj_adr_o_user[19]
port 814 nsew signal output
rlabel metal2 s 171874 17940 171930 18400 6 mprj_adr_o_user[1]
port 815 nsew signal output
rlabel metal2 s 189722 17940 189778 18400 6 mprj_adr_o_user[20]
port 816 nsew signal output
rlabel metal2 s 190550 17940 190606 18400 6 mprj_adr_o_user[21]
port 817 nsew signal output
rlabel metal2 s 191470 17940 191526 18400 6 mprj_adr_o_user[22]
port 818 nsew signal output
rlabel metal2 s 192298 17940 192354 18400 6 mprj_adr_o_user[23]
port 819 nsew signal output
rlabel metal2 s 193218 17940 193274 18400 6 mprj_adr_o_user[24]
port 820 nsew signal output
rlabel metal2 s 194046 17940 194102 18400 6 mprj_adr_o_user[25]
port 821 nsew signal output
rlabel metal2 s 194966 17940 195022 18400 6 mprj_adr_o_user[26]
port 822 nsew signal output
rlabel metal2 s 195794 17940 195850 18400 6 mprj_adr_o_user[27]
port 823 nsew signal output
rlabel metal2 s 196714 17940 196770 18400 6 mprj_adr_o_user[28]
port 824 nsew signal output
rlabel metal2 s 197542 17940 197598 18400 6 mprj_adr_o_user[29]
port 825 nsew signal output
rlabel metal2 s 173162 17940 173218 18400 6 mprj_adr_o_user[2]
port 826 nsew signal output
rlabel metal2 s 198462 17940 198518 18400 6 mprj_adr_o_user[30]
port 827 nsew signal output
rlabel metal2 s 199290 17940 199346 18400 6 mprj_adr_o_user[31]
port 828 nsew signal output
rlabel metal2 s 174450 17940 174506 18400 6 mprj_adr_o_user[3]
port 829 nsew signal output
rlabel metal2 s 175738 17940 175794 18400 6 mprj_adr_o_user[4]
port 830 nsew signal output
rlabel metal2 s 176658 17940 176714 18400 6 mprj_adr_o_user[5]
port 831 nsew signal output
rlabel metal2 s 177486 17940 177542 18400 6 mprj_adr_o_user[6]
port 832 nsew signal output
rlabel metal2 s 178406 17940 178462 18400 6 mprj_adr_o_user[7]
port 833 nsew signal output
rlabel metal2 s 179234 17940 179290 18400 6 mprj_adr_o_user[8]
port 834 nsew signal output
rlabel metal2 s 180154 17940 180210 18400 6 mprj_adr_o_user[9]
port 835 nsew signal output
rlabel metal2 s 167458 -400 167514 60 8 mprj_cyc_o_core
port 836 nsew signal input
rlabel metal2 s 169206 17940 169262 18400 6 mprj_cyc_o_user
port 837 nsew signal output
rlabel metal2 s 169206 -400 169262 60 8 mprj_dat_o_core[0]
port 838 nsew signal input
rlabel metal2 s 179694 -400 179750 60 8 mprj_dat_o_core[10]
port 839 nsew signal input
rlabel metal2 s 180522 -400 180578 60 8 mprj_dat_o_core[11]
port 840 nsew signal input
rlabel metal2 s 181442 -400 181498 60 8 mprj_dat_o_core[12]
port 841 nsew signal input
rlabel metal2 s 182270 -400 182326 60 8 mprj_dat_o_core[13]
port 842 nsew signal input
rlabel metal2 s 183190 -400 183246 60 8 mprj_dat_o_core[14]
port 843 nsew signal input
rlabel metal2 s 184018 -400 184074 60 8 mprj_dat_o_core[15]
port 844 nsew signal input
rlabel metal2 s 184938 -400 184994 60 8 mprj_dat_o_core[16]
port 845 nsew signal input
rlabel metal2 s 185766 -400 185822 60 8 mprj_dat_o_core[17]
port 846 nsew signal input
rlabel metal2 s 186686 -400 186742 60 8 mprj_dat_o_core[18]
port 847 nsew signal input
rlabel metal2 s 187514 -400 187570 60 8 mprj_dat_o_core[19]
port 848 nsew signal input
rlabel metal2 s 170494 -400 170550 60 8 mprj_dat_o_core[1]
port 849 nsew signal input
rlabel metal2 s 188434 -400 188490 60 8 mprj_dat_o_core[20]
port 850 nsew signal input
rlabel metal2 s 189262 -400 189318 60 8 mprj_dat_o_core[21]
port 851 nsew signal input
rlabel metal2 s 190182 -400 190238 60 8 mprj_dat_o_core[22]
port 852 nsew signal input
rlabel metal2 s 191010 -400 191066 60 8 mprj_dat_o_core[23]
port 853 nsew signal input
rlabel metal2 s 191930 -400 191986 60 8 mprj_dat_o_core[24]
port 854 nsew signal input
rlabel metal2 s 192758 -400 192814 60 8 mprj_dat_o_core[25]
port 855 nsew signal input
rlabel metal2 s 193586 -400 193642 60 8 mprj_dat_o_core[26]
port 856 nsew signal input
rlabel metal2 s 194506 -400 194562 60 8 mprj_dat_o_core[27]
port 857 nsew signal input
rlabel metal2 s 195334 -400 195390 60 8 mprj_dat_o_core[28]
port 858 nsew signal input
rlabel metal2 s 196254 -400 196310 60 8 mprj_dat_o_core[29]
port 859 nsew signal input
rlabel metal2 s 171874 -400 171930 60 8 mprj_dat_o_core[2]
port 860 nsew signal input
rlabel metal2 s 197082 -400 197138 60 8 mprj_dat_o_core[30]
port 861 nsew signal input
rlabel metal2 s 198002 -400 198058 60 8 mprj_dat_o_core[31]
port 862 nsew signal input
rlabel metal2 s 173162 -400 173218 60 8 mprj_dat_o_core[3]
port 863 nsew signal input
rlabel metal2 s 174450 -400 174506 60 8 mprj_dat_o_core[4]
port 864 nsew signal input
rlabel metal2 s 175370 -400 175426 60 8 mprj_dat_o_core[5]
port 865 nsew signal input
rlabel metal2 s 176198 -400 176254 60 8 mprj_dat_o_core[6]
port 866 nsew signal input
rlabel metal2 s 177026 -400 177082 60 8 mprj_dat_o_core[7]
port 867 nsew signal input
rlabel metal2 s 177946 -400 178002 60 8 mprj_dat_o_core[8]
port 868 nsew signal input
rlabel metal2 s 178774 -400 178830 60 8 mprj_dat_o_core[9]
port 869 nsew signal input
rlabel metal2 s 170954 17940 171010 18400 6 mprj_dat_o_user[0]
port 870 nsew signal output
rlabel metal2 s 181442 17940 181498 18400 6 mprj_dat_o_user[10]
port 871 nsew signal output
rlabel metal2 s 182270 17940 182326 18400 6 mprj_dat_o_user[11]
port 872 nsew signal output
rlabel metal2 s 183190 17940 183246 18400 6 mprj_dat_o_user[12]
port 873 nsew signal output
rlabel metal2 s 184018 17940 184074 18400 6 mprj_dat_o_user[13]
port 874 nsew signal output
rlabel metal2 s 184938 17940 184994 18400 6 mprj_dat_o_user[14]
port 875 nsew signal output
rlabel metal2 s 185766 17940 185822 18400 6 mprj_dat_o_user[15]
port 876 nsew signal output
rlabel metal2 s 186686 17940 186742 18400 6 mprj_dat_o_user[16]
port 877 nsew signal output
rlabel metal2 s 187514 17940 187570 18400 6 mprj_dat_o_user[17]
port 878 nsew signal output
rlabel metal2 s 188434 17940 188490 18400 6 mprj_dat_o_user[18]
port 879 nsew signal output
rlabel metal2 s 189262 17940 189318 18400 6 mprj_dat_o_user[19]
port 880 nsew signal output
rlabel metal2 s 172242 17940 172298 18400 6 mprj_dat_o_user[1]
port 881 nsew signal output
rlabel metal2 s 190182 17940 190238 18400 6 mprj_dat_o_user[20]
port 882 nsew signal output
rlabel metal2 s 191010 17940 191066 18400 6 mprj_dat_o_user[21]
port 883 nsew signal output
rlabel metal2 s 191930 17940 191986 18400 6 mprj_dat_o_user[22]
port 884 nsew signal output
rlabel metal2 s 192758 17940 192814 18400 6 mprj_dat_o_user[23]
port 885 nsew signal output
rlabel metal2 s 193586 17940 193642 18400 6 mprj_dat_o_user[24]
port 886 nsew signal output
rlabel metal2 s 194506 17940 194562 18400 6 mprj_dat_o_user[25]
port 887 nsew signal output
rlabel metal2 s 195334 17940 195390 18400 6 mprj_dat_o_user[26]
port 888 nsew signal output
rlabel metal2 s 196254 17940 196310 18400 6 mprj_dat_o_user[27]
port 889 nsew signal output
rlabel metal2 s 197082 17940 197138 18400 6 mprj_dat_o_user[28]
port 890 nsew signal output
rlabel metal2 s 198002 17940 198058 18400 6 mprj_dat_o_user[29]
port 891 nsew signal output
rlabel metal2 s 173622 17940 173678 18400 6 mprj_dat_o_user[2]
port 892 nsew signal output
rlabel metal2 s 198830 17940 198886 18400 6 mprj_dat_o_user[30]
port 893 nsew signal output
rlabel metal2 s 199750 17940 199806 18400 6 mprj_dat_o_user[31]
port 894 nsew signal output
rlabel metal2 s 174910 17940 174966 18400 6 mprj_dat_o_user[3]
port 895 nsew signal output
rlabel metal2 s 176198 17940 176254 18400 6 mprj_dat_o_user[4]
port 896 nsew signal output
rlabel metal2 s 177026 17940 177082 18400 6 mprj_dat_o_user[5]
port 897 nsew signal output
rlabel metal2 s 177946 17940 178002 18400 6 mprj_dat_o_user[6]
port 898 nsew signal output
rlabel metal2 s 178774 17940 178830 18400 6 mprj_dat_o_user[7]
port 899 nsew signal output
rlabel metal2 s 179694 17940 179750 18400 6 mprj_dat_o_user[8]
port 900 nsew signal output
rlabel metal2 s 180522 17940 180578 18400 6 mprj_dat_o_user[9]
port 901 nsew signal output
rlabel metal2 s 169666 -400 169722 60 8 mprj_sel_o_core[0]
port 902 nsew signal input
rlabel metal2 s 170954 -400 171010 60 8 mprj_sel_o_core[1]
port 903 nsew signal input
rlabel metal2 s 172242 -400 172298 60 8 mprj_sel_o_core[2]
port 904 nsew signal input
rlabel metal2 s 173622 -400 173678 60 8 mprj_sel_o_core[3]
port 905 nsew signal input
rlabel metal2 s 171414 17940 171470 18400 6 mprj_sel_o_user[0]
port 906 nsew signal output
rlabel metal2 s 172702 17940 172758 18400 6 mprj_sel_o_user[1]
port 907 nsew signal output
rlabel metal2 s 173990 17940 174046 18400 6 mprj_sel_o_user[2]
port 908 nsew signal output
rlabel metal2 s 175370 17940 175426 18400 6 mprj_sel_o_user[3]
port 909 nsew signal output
rlabel metal2 s 167918 -400 167974 60 8 mprj_stb_o_core
port 910 nsew signal input
rlabel metal2 s 169666 17940 169722 18400 6 mprj_stb_o_user
port 911 nsew signal output
rlabel metal2 s 168378 -400 168434 60 8 mprj_we_o_core
port 912 nsew signal input
rlabel metal2 s 170126 17940 170182 18400 6 mprj_we_o_user
port 913 nsew signal output
rlabel metal2 s 198462 -400 198518 60 8 user1_vcc_powergood
port 914 nsew signal output
rlabel metal2 s 198830 -400 198886 60 8 user1_vdd_powergood
port 915 nsew signal output
rlabel metal2 s 199290 -400 199346 60 8 user2_vcc_powergood
port 916 nsew signal output
rlabel metal2 s 199750 -400 199806 60 8 user2_vdd_powergood
port 917 nsew signal output
rlabel metal2 s 202 17940 258 18400 6 user_clock
port 918 nsew signal output
rlabel metal2 s 570 17940 626 18400 6 user_clock2
port 919 nsew signal output
rlabel metal2 s 1030 17940 1086 18400 6 user_reset
port 920 nsew signal output
rlabel metal2 s 1490 17940 1546 18400 6 user_resetn
port 921 nsew signal output
rlabel metal4 s 183984 -482 184224 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 153984 -482 154224 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 123984 -482 124224 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 93984 -482 94224 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 63984 -482 64224 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 33984 -482 34224 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 3984 -482 4224 60 8 vccd
port 922 nsew power bidirectional
rlabel metal4 s 183984 17940 184224 18434 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 153984 17940 154224 18434 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 123984 17940 124224 18434 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 93984 17940 94224 18434 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 63984 17940 64224 18434 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 33984 17940 34224 18434 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 3984 17940 4224 18434 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 184152 -344 184216 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 184072 -344 184136 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 183992 -344 184056 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 154152 -344 154216 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 154072 -344 154136 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 153992 -344 154056 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 124152 -344 124216 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 124072 -344 124136 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 123992 -344 124056 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 94152 -344 94216 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 94072 -344 94136 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 93992 -344 94056 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 64152 -344 64216 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 64072 -344 64136 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 63992 -344 64056 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 34152 -344 34216 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 34072 -344 34136 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 33992 -344 34056 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 4152 -344 4216 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 4072 -344 4136 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 3992 -344 4056 -280 8 vccd
port 922 nsew power bidirectional
rlabel via3 s 184152 18232 184216 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 184072 18232 184136 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 183992 18232 184056 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 154152 18232 154216 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 154072 18232 154136 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 153992 18232 154056 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 124152 18232 124216 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 124072 18232 124136 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 123992 18232 124056 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 94152 18232 94216 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 94072 18232 94136 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 93992 18232 94056 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 64152 18232 64216 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 64072 18232 64136 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 63992 18232 64056 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 34152 18232 34216 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 34072 18232 34136 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 33992 18232 34056 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 4152 18232 4216 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 4072 18232 4136 18296 6 vccd
port 922 nsew power bidirectional
rlabel via3 s 3992 18232 4056 18296 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 183984 -344 184224 -342 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 153984 -344 154224 -342 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 123984 -344 124224 -342 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 93984 -344 94224 -342 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 63984 -344 64224 -342 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 33984 -344 34224 -342 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 3984 -344 4224 -342 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s -326 -342 200242 -282 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 183984 -282 184224 -280 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 153984 -282 154224 -280 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 123984 -282 124224 -280 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 93984 -282 94224 -280 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 63984 -282 64224 -280 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 33984 -282 34224 -280 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 3984 -282 4224 -280 8 vccd
port 922 nsew power bidirectional
rlabel metal3 s 183984 18232 184224 18234 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 153984 18232 154224 18234 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 123984 18232 124224 18234 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 93984 18232 94224 18234 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 63984 18232 64224 18234 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 33984 18232 34224 18234 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 3984 18232 4224 18234 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s -326 18234 200242 18294 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 183984 18294 184224 18296 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 153984 18294 154224 18296 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 123984 18294 124224 18296 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 93984 18294 94224 18296 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 63984 18294 64224 18296 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 33984 18294 34224 18296 6 vccd
port 922 nsew power bidirectional
rlabel metal3 s 3984 18294 4224 18296 6 vccd
port 922 nsew power bidirectional
rlabel metal4 s 200182 -342 200242 18294 6 vccd
port 923 nsew power bidirectional
rlabel metal4 s -326 -342 -266 18294 4 vccd
port 924 nsew power bidirectional
rlabel metal4 s 168984 -485 169224 60 8 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 138984 -485 139224 60 8 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 108984 -485 109224 60 8 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 78984 -485 79224 60 8 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 48984 -485 49224 60 8 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 18984 -485 19224 60 8 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 168984 17940 169224 18437 6 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 138984 17940 139224 18437 6 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 108984 17940 109224 18437 6 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 78984 17940 79224 18437 6 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 48984 17940 49224 18437 6 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 18984 17940 19224 18437 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 169152 -484 169216 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 169072 -484 169136 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 168992 -484 169056 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 139152 -484 139216 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 139072 -484 139136 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 138992 -484 139056 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 109152 -484 109216 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 109072 -484 109136 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 108992 -484 109056 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 79152 -484 79216 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 79072 -484 79136 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 78992 -484 79056 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 49152 -484 49216 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 49072 -484 49136 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 48992 -484 49056 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 19152 -484 19216 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 19072 -484 19136 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 18992 -484 19056 -420 8 vssd
port 925 nsew ground bidirectional
rlabel via3 s 169152 18372 169216 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 169072 18372 169136 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 168992 18372 169056 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 139152 18372 139216 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 139072 18372 139136 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 138992 18372 139056 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 109152 18372 109216 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 109072 18372 109136 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 108992 18372 109056 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 79152 18372 79216 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 79072 18372 79136 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 78992 18372 79056 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 49152 18372 49216 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 49072 18372 49136 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 48992 18372 49056 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 19152 18372 19216 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 19072 18372 19136 18436 6 vssd
port 925 nsew ground bidirectional
rlabel via3 s 18992 18372 19056 18436 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 168984 -484 169224 -482 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 138984 -484 139224 -482 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 108984 -484 109224 -482 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 78984 -484 79224 -482 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 48984 -484 49224 -482 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 18984 -484 19224 -482 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s -466 -482 200382 -422 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 168984 -422 169224 -420 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 138984 -422 139224 -420 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 108984 -422 109224 -420 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 78984 -422 79224 -420 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 48984 -422 49224 -420 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 18984 -422 19224 -420 8 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 168984 18372 169224 18374 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 138984 18372 139224 18374 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 108984 18372 109224 18374 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 78984 18372 79224 18374 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 48984 18372 49224 18374 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 18984 18372 19224 18374 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s -466 18374 200382 18434 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 168984 18434 169224 18436 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 138984 18434 139224 18436 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 108984 18434 109224 18436 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 78984 18434 79224 18436 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 48984 18434 49224 18436 6 vssd
port 925 nsew ground bidirectional
rlabel metal3 s 18984 18434 19224 18436 6 vssd
port 925 nsew ground bidirectional
rlabel metal4 s 200322 -482 200382 18434 6 vssd
port 926 nsew ground bidirectional
rlabel metal4 s -466 -482 -406 18434 4 vssd
port 927 nsew ground bidirectional
rlabel metal4 s 184864 -762 185104 60 8 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 154864 -762 155104 60 8 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 124864 -762 125104 60 8 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 94864 -762 95104 60 8 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 64864 -762 65104 60 8 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 34864 -762 35104 60 8 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 4864 -762 5104 60 8 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 184864 17940 185104 18714 6 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 154864 17940 155104 18714 6 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 124864 17940 125104 18714 6 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 94864 17940 95104 18714 6 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 64864 17940 65104 18714 6 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 34864 17940 35104 18714 6 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 4864 17940 5104 18714 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 185032 -624 185096 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 184952 -624 185016 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 184872 -624 184936 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 155032 -624 155096 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 154952 -624 155016 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 154872 -624 154936 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 125032 -624 125096 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 124952 -624 125016 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 124872 -624 124936 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 95032 -624 95096 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 94952 -624 95016 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 94872 -624 94936 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 65032 -624 65096 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 64952 -624 65016 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 64872 -624 64936 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 35032 -624 35096 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 34952 -624 35016 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 34872 -624 34936 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 5032 -624 5096 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 4952 -624 5016 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 4872 -624 4936 -560 8 vccd1
port 928 nsew power bidirectional
rlabel via3 s 185032 18512 185096 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 184952 18512 185016 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 184872 18512 184936 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 155032 18512 155096 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 154952 18512 155016 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 154872 18512 154936 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 125032 18512 125096 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 124952 18512 125016 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 124872 18512 124936 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 95032 18512 95096 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 94952 18512 95016 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 94872 18512 94936 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 65032 18512 65096 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 64952 18512 65016 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 64872 18512 64936 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 35032 18512 35096 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 34952 18512 35016 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 34872 18512 34936 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 5032 18512 5096 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 4952 18512 5016 18576 6 vccd1
port 928 nsew power bidirectional
rlabel via3 s 4872 18512 4936 18576 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 184864 -624 185104 -622 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 154864 -624 155104 -622 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 124864 -624 125104 -622 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 94864 -624 95104 -622 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 64864 -624 65104 -622 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 34864 -624 35104 -622 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 4864 -624 5104 -622 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s -606 -622 200522 -562 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 184864 -562 185104 -560 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 154864 -562 155104 -560 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 124864 -562 125104 -560 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 94864 -562 95104 -560 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 64864 -562 65104 -560 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 34864 -562 35104 -560 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 4864 -562 5104 -560 8 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 184864 18512 185104 18514 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 154864 18512 155104 18514 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 124864 18512 125104 18514 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 94864 18512 95104 18514 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 64864 18512 65104 18514 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 34864 18512 35104 18514 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 4864 18512 5104 18514 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s -606 18514 200522 18574 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 184864 18574 185104 18576 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 154864 18574 155104 18576 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 124864 18574 125104 18576 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 94864 18574 95104 18576 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 64864 18574 65104 18576 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 34864 18574 35104 18576 6 vccd1
port 928 nsew power bidirectional
rlabel metal3 s 4864 18574 5104 18576 6 vccd1
port 928 nsew power bidirectional
rlabel metal4 s 200462 -622 200522 18574 6 vccd1
port 929 nsew power bidirectional
rlabel metal4 s -606 -622 -546 18574 4 vccd1
port 930 nsew power bidirectional
rlabel metal4 s 169864 -765 170104 60 8 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 139864 -765 140104 60 8 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 109864 -765 110104 60 8 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 79864 -765 80104 60 8 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 49864 -765 50104 60 8 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 19864 -765 20104 60 8 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 169864 17940 170104 18717 6 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 139864 17940 140104 18717 6 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 109864 17940 110104 18717 6 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 79864 17940 80104 18717 6 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 49864 17940 50104 18717 6 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 19864 17940 20104 18717 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 170032 -764 170096 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 169952 -764 170016 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 169872 -764 169936 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 140032 -764 140096 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 139952 -764 140016 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 139872 -764 139936 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 110032 -764 110096 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 109952 -764 110016 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 109872 -764 109936 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 80032 -764 80096 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 79952 -764 80016 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 79872 -764 79936 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 50032 -764 50096 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 49952 -764 50016 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 49872 -764 49936 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 20032 -764 20096 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 19952 -764 20016 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 19872 -764 19936 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 170032 18652 170096 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 169952 18652 170016 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 169872 18652 169936 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 140032 18652 140096 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 139952 18652 140016 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 139872 18652 139936 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 110032 18652 110096 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 109952 18652 110016 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 109872 18652 109936 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 80032 18652 80096 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 79952 18652 80016 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 79872 18652 79936 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 50032 18652 50096 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 49952 18652 50016 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 49872 18652 49936 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 20032 18652 20096 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 19952 18652 20016 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel via3 s 19872 18652 19936 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 169864 -764 170104 -762 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 139864 -764 140104 -762 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 109864 -764 110104 -762 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 79864 -764 80104 -762 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 49864 -764 50104 -762 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 19864 -764 20104 -762 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s -746 -762 200662 -702 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 169864 -702 170104 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 139864 -702 140104 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 109864 -702 110104 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 79864 -702 80104 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 49864 -702 50104 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 19864 -702 20104 -700 8 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 169864 18652 170104 18654 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 139864 18652 140104 18654 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 109864 18652 110104 18654 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 79864 18652 80104 18654 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 49864 18652 50104 18654 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 19864 18652 20104 18654 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s -746 18654 200662 18714 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 169864 18714 170104 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 139864 18714 140104 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 109864 18714 110104 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 79864 18714 80104 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 49864 18714 50104 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel metal3 s 19864 18714 20104 18716 6 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 200602 -762 200662 18714 6 vssd1
port 932 nsew ground bidirectional
rlabel metal4 s -746 -762 -686 18714 4 vssd1
port 933 nsew ground bidirectional
rlabel metal4 s 185744 -1042 185984 60 8 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 155744 -1042 155984 60 8 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 125744 -1042 125984 60 8 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 95744 -1042 95984 60 8 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 65744 -1042 65984 60 8 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 35744 -1042 35984 60 8 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 5744 -1042 5984 60 8 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 185744 17940 185984 18994 6 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 155744 17940 155984 18994 6 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 125744 17940 125984 18994 6 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 95744 17940 95984 18994 6 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 65744 17940 65984 18994 6 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 35744 17940 35984 18994 6 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 5744 17940 5984 18994 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 185912 -904 185976 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 185832 -904 185896 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 185752 -904 185816 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 155912 -904 155976 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 155832 -904 155896 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 155752 -904 155816 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 125912 -904 125976 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 125832 -904 125896 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 125752 -904 125816 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 95912 -904 95976 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 95832 -904 95896 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 95752 -904 95816 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 65912 -904 65976 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 65832 -904 65896 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 65752 -904 65816 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 35912 -904 35976 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 35832 -904 35896 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 35752 -904 35816 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 5912 -904 5976 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 5832 -904 5896 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 5752 -904 5816 -840 8 vccd2
port 934 nsew power bidirectional
rlabel via3 s 185912 18792 185976 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 185832 18792 185896 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 185752 18792 185816 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 155912 18792 155976 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 155832 18792 155896 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 155752 18792 155816 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 125912 18792 125976 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 125832 18792 125896 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 125752 18792 125816 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 95912 18792 95976 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 95832 18792 95896 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 95752 18792 95816 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 65912 18792 65976 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 65832 18792 65896 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 65752 18792 65816 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 35912 18792 35976 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 35832 18792 35896 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 35752 18792 35816 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 5912 18792 5976 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 5832 18792 5896 18856 6 vccd2
port 934 nsew power bidirectional
rlabel via3 s 5752 18792 5816 18856 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 185744 -904 185984 -902 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 155744 -904 155984 -902 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 125744 -904 125984 -902 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 95744 -904 95984 -902 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 65744 -904 65984 -902 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 35744 -904 35984 -902 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 5744 -904 5984 -902 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s -886 -902 200802 -842 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 185744 -842 185984 -840 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 155744 -842 155984 -840 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 125744 -842 125984 -840 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 95744 -842 95984 -840 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 65744 -842 65984 -840 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 35744 -842 35984 -840 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 5744 -842 5984 -840 8 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 185744 18792 185984 18794 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 155744 18792 155984 18794 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 125744 18792 125984 18794 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 95744 18792 95984 18794 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 65744 18792 65984 18794 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 35744 18792 35984 18794 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 5744 18792 5984 18794 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s -886 18794 200802 18854 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 185744 18854 185984 18856 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 155744 18854 155984 18856 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 125744 18854 125984 18856 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 95744 18854 95984 18856 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 65744 18854 65984 18856 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 35744 18854 35984 18856 6 vccd2
port 934 nsew power bidirectional
rlabel metal3 s 5744 18854 5984 18856 6 vccd2
port 934 nsew power bidirectional
rlabel metal4 s 200742 -902 200802 18854 6 vccd2
port 935 nsew power bidirectional
rlabel metal4 s -886 -902 -826 18854 4 vccd2
port 936 nsew power bidirectional
rlabel metal4 s 170744 -1045 170984 60 8 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 140744 -1045 140984 60 8 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 110744 -1045 110984 60 8 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 80744 -1045 80984 60 8 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 50744 -1045 50984 60 8 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 20744 -1045 20984 60 8 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 170744 17940 170984 18997 6 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 140744 17940 140984 18997 6 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 110744 17940 110984 18997 6 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 80744 17940 80984 18997 6 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 50744 17940 50984 18997 6 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 20744 17940 20984 18997 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 170912 -1044 170976 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 170832 -1044 170896 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 170752 -1044 170816 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 140912 -1044 140976 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 140832 -1044 140896 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 140752 -1044 140816 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 110912 -1044 110976 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 110832 -1044 110896 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 110752 -1044 110816 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 80912 -1044 80976 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 80832 -1044 80896 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 80752 -1044 80816 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 50912 -1044 50976 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 50832 -1044 50896 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 50752 -1044 50816 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 20912 -1044 20976 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 20832 -1044 20896 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 20752 -1044 20816 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 170912 18932 170976 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 170832 18932 170896 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 170752 18932 170816 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 140912 18932 140976 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 140832 18932 140896 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 140752 18932 140816 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 110912 18932 110976 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 110832 18932 110896 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 110752 18932 110816 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 80912 18932 80976 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 80832 18932 80896 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 80752 18932 80816 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 50912 18932 50976 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 50832 18932 50896 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 50752 18932 50816 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 20912 18932 20976 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 20832 18932 20896 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel via3 s 20752 18932 20816 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 170744 -1044 170984 -1042 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 140744 -1044 140984 -1042 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 110744 -1044 110984 -1042 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 80744 -1044 80984 -1042 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 50744 -1044 50984 -1042 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 20744 -1044 20984 -1042 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s -1026 -1042 200942 -982 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 170744 -982 170984 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 140744 -982 140984 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 110744 -982 110984 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 80744 -982 80984 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 50744 -982 50984 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 20744 -982 20984 -980 8 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 170744 18932 170984 18934 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 140744 18932 140984 18934 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 110744 18932 110984 18934 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 80744 18932 80984 18934 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 50744 18932 50984 18934 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 20744 18932 20984 18934 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s -1026 18934 200942 18994 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 170744 18994 170984 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 140744 18994 140984 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 110744 18994 110984 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 80744 18994 80984 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 50744 18994 50984 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel metal3 s 20744 18994 20984 18996 6 vssd2
port 937 nsew ground bidirectional
rlabel metal4 s 200882 -1042 200942 18994 6 vssd2
port 938 nsew ground bidirectional
rlabel metal4 s -1026 -1042 -966 18994 4 vssd2
port 939 nsew ground bidirectional
rlabel metal4 s 186624 -1322 186864 60 8 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 156624 -1322 156864 60 8 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 126624 -1322 126864 60 8 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 96624 -1322 96864 60 8 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 66624 -1322 66864 60 8 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 36624 -1322 36864 60 8 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 6624 -1322 6864 60 8 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 186624 17940 186864 19274 6 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 156624 17940 156864 19274 6 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 126624 17940 126864 19274 6 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 96624 17940 96864 19274 6 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 66624 17940 66864 19274 6 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 36624 17940 36864 19274 6 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 6624 17940 6864 19274 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 186792 -1184 186856 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 186712 -1184 186776 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 186632 -1184 186696 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 156792 -1184 156856 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 156712 -1184 156776 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 156632 -1184 156696 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 126792 -1184 126856 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 126712 -1184 126776 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 126632 -1184 126696 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 96792 -1184 96856 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 96712 -1184 96776 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 96632 -1184 96696 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 66792 -1184 66856 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 66712 -1184 66776 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 66632 -1184 66696 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 36792 -1184 36856 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 36712 -1184 36776 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 36632 -1184 36696 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 6792 -1184 6856 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 6712 -1184 6776 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 6632 -1184 6696 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel via3 s 186792 19072 186856 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 186712 19072 186776 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 186632 19072 186696 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 156792 19072 156856 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 156712 19072 156776 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 156632 19072 156696 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 126792 19072 126856 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 126712 19072 126776 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 126632 19072 126696 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 96792 19072 96856 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 96712 19072 96776 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 96632 19072 96696 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 66792 19072 66856 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 66712 19072 66776 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 66632 19072 66696 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 36792 19072 36856 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 36712 19072 36776 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 36632 19072 36696 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 6792 19072 6856 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 6712 19072 6776 19136 6 vdda1
port 940 nsew power bidirectional
rlabel via3 s 6632 19072 6696 19136 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 186624 -1184 186864 -1182 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 156624 -1184 156864 -1182 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 126624 -1184 126864 -1182 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 96624 -1184 96864 -1182 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 66624 -1184 66864 -1182 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 36624 -1184 36864 -1182 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 6624 -1184 6864 -1182 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s -1166 -1182 201082 -1122 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 186624 -1122 186864 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 156624 -1122 156864 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 126624 -1122 126864 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 96624 -1122 96864 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 66624 -1122 66864 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 36624 -1122 36864 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 6624 -1122 6864 -1120 8 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 186624 19072 186864 19074 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 156624 19072 156864 19074 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 126624 19072 126864 19074 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 96624 19072 96864 19074 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 66624 19072 66864 19074 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 36624 19072 36864 19074 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 6624 19072 6864 19074 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s -1166 19074 201082 19134 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 186624 19134 186864 19136 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 156624 19134 156864 19136 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 126624 19134 126864 19136 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 96624 19134 96864 19136 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 66624 19134 66864 19136 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 36624 19134 36864 19136 6 vdda1
port 940 nsew power bidirectional
rlabel metal3 s 6624 19134 6864 19136 6 vdda1
port 940 nsew power bidirectional
rlabel metal4 s 201022 -1182 201082 19134 6 vdda1
port 941 nsew power bidirectional
rlabel metal4 s -1166 -1182 -1106 19134 4 vdda1
port 942 nsew power bidirectional
rlabel metal4 s 171624 -1325 171864 60 8 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 141624 -1325 141864 60 8 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 111624 -1325 111864 60 8 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 81624 -1325 81864 60 8 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 51624 -1325 51864 60 8 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 21624 -1325 21864 60 8 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 171624 17940 171864 19277 6 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 141624 17940 141864 19277 6 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 111624 17940 111864 19277 6 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 81624 17940 81864 19277 6 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 51624 17940 51864 19277 6 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 21624 17940 21864 19277 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 171792 -1324 171856 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 171712 -1324 171776 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 171632 -1324 171696 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 141792 -1324 141856 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 141712 -1324 141776 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 141632 -1324 141696 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 111792 -1324 111856 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 111712 -1324 111776 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 111632 -1324 111696 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 81792 -1324 81856 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 81712 -1324 81776 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 81632 -1324 81696 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 51792 -1324 51856 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 51712 -1324 51776 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 51632 -1324 51696 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 21792 -1324 21856 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 21712 -1324 21776 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 21632 -1324 21696 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 171792 19212 171856 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 171712 19212 171776 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 171632 19212 171696 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 141792 19212 141856 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 141712 19212 141776 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 141632 19212 141696 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 111792 19212 111856 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 111712 19212 111776 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 111632 19212 111696 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 81792 19212 81856 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 81712 19212 81776 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 81632 19212 81696 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 51792 19212 51856 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 51712 19212 51776 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 51632 19212 51696 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 21792 19212 21856 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 21712 19212 21776 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel via3 s 21632 19212 21696 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 171624 -1324 171864 -1322 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 141624 -1324 141864 -1322 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 111624 -1324 111864 -1322 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 81624 -1324 81864 -1322 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 51624 -1324 51864 -1322 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 21624 -1324 21864 -1322 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s -1306 -1322 201222 -1262 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 171624 -1262 171864 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 141624 -1262 141864 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 111624 -1262 111864 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 81624 -1262 81864 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 51624 -1262 51864 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 21624 -1262 21864 -1260 8 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 171624 19212 171864 19214 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 141624 19212 141864 19214 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 111624 19212 111864 19214 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 81624 19212 81864 19214 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 51624 19212 51864 19214 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 21624 19212 21864 19214 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s -1306 19214 201222 19274 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 171624 19274 171864 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 141624 19274 141864 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 111624 19274 111864 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 81624 19274 81864 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 51624 19274 51864 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel metal3 s 21624 19274 21864 19276 6 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 201162 -1322 201222 19274 6 vssa1
port 944 nsew ground bidirectional
rlabel metal4 s -1306 -1322 -1246 19274 4 vssa1
port 945 nsew ground bidirectional
rlabel metal4 s 187504 -1602 187744 60 8 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 157504 -1602 157744 60 8 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 127504 -1602 127744 60 8 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 97504 -1602 97744 60 8 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 67504 -1602 67744 60 8 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 37504 -1602 37744 60 8 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 7504 -1602 7744 60 8 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 187504 17940 187744 19554 6 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 157504 17940 157744 19554 6 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 127504 17940 127744 19554 6 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 97504 17940 97744 19554 6 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 67504 17940 67744 19554 6 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 37504 17940 37744 19554 6 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 7504 17940 7744 19554 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 187672 -1464 187736 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 187592 -1464 187656 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 187512 -1464 187576 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 157672 -1464 157736 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 157592 -1464 157656 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 157512 -1464 157576 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 127672 -1464 127736 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 127592 -1464 127656 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 127512 -1464 127576 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 97672 -1464 97736 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 97592 -1464 97656 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 97512 -1464 97576 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 67672 -1464 67736 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 67592 -1464 67656 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 67512 -1464 67576 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 37672 -1464 37736 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 37592 -1464 37656 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 37512 -1464 37576 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 7672 -1464 7736 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 7592 -1464 7656 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 7512 -1464 7576 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel via3 s 187672 19352 187736 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 187592 19352 187656 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 187512 19352 187576 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 157672 19352 157736 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 157592 19352 157656 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 157512 19352 157576 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 127672 19352 127736 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 127592 19352 127656 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 127512 19352 127576 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 97672 19352 97736 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 97592 19352 97656 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 97512 19352 97576 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 67672 19352 67736 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 67592 19352 67656 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 67512 19352 67576 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 37672 19352 37736 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 37592 19352 37656 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 37512 19352 37576 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 7672 19352 7736 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 7592 19352 7656 19416 6 vdda2
port 946 nsew power bidirectional
rlabel via3 s 7512 19352 7576 19416 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 187504 -1464 187744 -1462 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 157504 -1464 157744 -1462 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 127504 -1464 127744 -1462 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 97504 -1464 97744 -1462 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 67504 -1464 67744 -1462 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 37504 -1464 37744 -1462 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 7504 -1464 7744 -1462 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s -1446 -1462 201362 -1402 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 187504 -1402 187744 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 157504 -1402 157744 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 127504 -1402 127744 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 97504 -1402 97744 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 67504 -1402 67744 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 37504 -1402 37744 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 7504 -1402 7744 -1400 8 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 187504 19352 187744 19354 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 157504 19352 157744 19354 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 127504 19352 127744 19354 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 97504 19352 97744 19354 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 67504 19352 67744 19354 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 37504 19352 37744 19354 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 7504 19352 7744 19354 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s -1446 19354 201362 19414 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 187504 19414 187744 19416 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 157504 19414 157744 19416 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 127504 19414 127744 19416 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 97504 19414 97744 19416 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 67504 19414 67744 19416 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 37504 19414 37744 19416 6 vdda2
port 946 nsew power bidirectional
rlabel metal3 s 7504 19414 7744 19416 6 vdda2
port 946 nsew power bidirectional
rlabel metal4 s 201302 -1462 201362 19414 6 vdda2
port 947 nsew power bidirectional
rlabel metal4 s -1446 -1462 -1386 19414 4 vdda2
port 948 nsew power bidirectional
rlabel metal4 s 172504 -1605 172744 60 8 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 142504 -1605 142744 60 8 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 112504 -1605 112744 60 8 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 82504 -1605 82744 60 8 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 52504 -1605 52744 60 8 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 22504 -1605 22744 60 8 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 172504 17940 172744 19557 6 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 142504 17940 142744 19557 6 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 112504 17940 112744 19557 6 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 82504 17940 82744 19557 6 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 52504 17940 52744 19557 6 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 22504 17940 22744 19557 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 172672 -1604 172736 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 172592 -1604 172656 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 172512 -1604 172576 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 142672 -1604 142736 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 142592 -1604 142656 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 142512 -1604 142576 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 112672 -1604 112736 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 112592 -1604 112656 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 112512 -1604 112576 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 82672 -1604 82736 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 82592 -1604 82656 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 82512 -1604 82576 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 52672 -1604 52736 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 52592 -1604 52656 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 52512 -1604 52576 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 22672 -1604 22736 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 22592 -1604 22656 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 22512 -1604 22576 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 172672 19492 172736 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 172592 19492 172656 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 172512 19492 172576 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 142672 19492 142736 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 142592 19492 142656 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 142512 19492 142576 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 112672 19492 112736 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 112592 19492 112656 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 112512 19492 112576 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 82672 19492 82736 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 82592 19492 82656 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 82512 19492 82576 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 52672 19492 52736 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 52592 19492 52656 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 52512 19492 52576 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 22672 19492 22736 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 22592 19492 22656 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel via3 s 22512 19492 22576 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 172504 -1604 172744 -1602 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 142504 -1604 142744 -1602 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 112504 -1604 112744 -1602 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 82504 -1604 82744 -1602 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 52504 -1604 52744 -1602 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 22504 -1604 22744 -1602 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s -1586 -1602 201502 -1542 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 172504 -1542 172744 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 142504 -1542 142744 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 112504 -1542 112744 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 82504 -1542 82744 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 52504 -1542 52744 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 22504 -1542 22744 -1540 8 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 172504 19492 172744 19494 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 142504 19492 142744 19494 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 112504 19492 112744 19494 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 82504 19492 82744 19494 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 52504 19492 52744 19494 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 22504 19492 22744 19494 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s -1586 19494 201502 19554 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 172504 19554 172744 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 142504 19554 142744 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 112504 19554 112744 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 82504 19554 82744 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 52504 19554 52744 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel metal3 s 22504 19554 22744 19556 6 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 201442 -1602 201502 19554 6 vssa2
port 950 nsew ground bidirectional
rlabel metal4 s -1586 -1602 -1526 19554 4 vssa2
port 951 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 200000 18000
string LEFview TRUE
<< end >>
